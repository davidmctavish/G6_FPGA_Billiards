`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ht+yYNL2dUNWU1Dv1ERgSRMgdP1HiWatsDXZ5YD2FmPaqbvCIESwS21q2Bgw77M+BtZCZy/MZLWU
TOws/DAAyw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k4lNdMlD07BNffPZpUqmwlUKkdrmavSi5N6vi71rrejNcnm/Yiy/dYg3dEgJTJMW2NBzGWeSP8/g
F4V3MGCDAXXxT6LX3akmKYKZTuJIS+4o/XWaoiCzGR9jEv86DTS3Czx/WZ/K5DOgfzhuFVEIh9JO
UrWUQZY/z/WUeW/LHzI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CW7Sy6Bg6Drp7+rdYEGZNHSJJMRAlF68/rTQjhRlKtDv+ATM6NXgh1fhd1UnMTj16ifJ/kdLG2KG
OeFStkpXKxhlDoRNoCeoS9fyj77+QszEdPrBxF/SyNrVAIWAq0V+xqbaK6lk4m6wfwu1HuWDzh2a
GZcT8eAdRtWXLxw+oIolt/HKtyce56jU9CY7wj+rORqGsnloAdJwVj96ZN/1I6jU/g1YhxqkcgDn
GlOlA5rQmPYXWUslebm/NRWnv044arDZdTCn3G46Wfss1upw9ga4NysonBM89HwygV6nXOiVR1ky
JreVphDX25qv8Fy65hnmxkoIWKJlBdXQ8MBdRg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SrC035n16ITCAg6V8YSmmbFyvIBvKC/TfvWCoCuODmxbooOlNXLPqZLkCXchl0dPd9L+la5OgODW
vawUM1gFW6ww3Y91w42RevAS6PKr2U/hTzyK2B0U/fzuhEXc0umetnHnIbKjgE7xM5V77CtA0TuL
NJmELqGq0GwneylbcDo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vgm8m5FExCI2v4hHQEWr+Y1rZL1nj7qMCX0ltzTCV3lkAs6mcYaDZ8Dyr6Vx+Nvu6twpWkI/RS0M
mRQ/z16DaTzP5xfRukLOcwwIMGOrRtXaHS2tp5f/O40TfNAdP3ufN/4fCs1OpDMDAtsmu1ubj00v
iw1tZ3foBdzrttlZxqzZRsHI7wFpOd8NL7MruBQX/7RtRGsmJdEytW/mVVghHzKCJjaeJU57Ergh
1dk+tHkwh/rZpsdfcwuDBACoI1R3cyAv8Z0y7KZh9EMBy7HaAdf2kmUzS++P1peJQhCV1Z596GVd
finUR88DnisN+Wwd1LRi9uzfdp8q+WdM46+GDA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 28960)
`protect data_block
Ek2L90rPggu2HkjGrVP2flzx64DrO6hl1ebj4yvCtwKYkxAzN/bkcKZWBPkiwyD4BTztnnDu4UYw
kAYKGCDzsIMnI3pJ1oZ4HBMoGwbxHIMIayGXP+jNPhQ3E6o8YBfuNeTrIiJ1hjBxM+Qm+SQHSS7l
W5iSIlPF3bCvgJq+OqfeO9kaREbxhJpuCXFoWsZpYRxXiDhvVfAppK8kf4vZ5kbx2T/epUJDV5uk
dbAjloMsphINNnEAWcPAw/r17XkHszf+k37RcYFFexNr57P22cfwdq1F0VWocz8Nl8ihKP58Gm0z
hXstAbhJdN9xVbJtv0l8kUJFIwlriqAkcUB08eDp3bAm9fGWdqw0negUP4LeCSRz+FScHRCEjFxL
7bFRdUYwCgHaLSZ2HqBENL6ShgVNRMQuWp/C3IgqR5O6y6rXz534mfD4KfusfG00tQYU4WdwymOX
Gw1DtDXHJPLEHMbyye4/wEC/DSUCSzDsHE0fFoJtYNTDxyYoPqwqnZcxE7G57CVrZj0TabNyEcei
RrQeh66V4nRqpDlxQJLsIp2BZeAmS0Dar9SOUvqPVULh7tSz0tzGR4y+Xxa5Kdo23ok0X+q2S/9r
ykCpBNa6BcvjpU2vtJSNmn89VX+BQ6I+Gw4MQby+eklV+5g0+nkl1dL1o0TCkMwV5Efb/liKio4v
pl6+y3sQUXN5CfNX/W7tdtKOg9vRAsazwN+yNB9WyqqFKTY1b4JK5Ac0Krx2tHl/YJF3VrzDk3d4
PvRJEj9+GWkPBytAnBlX0annvo0oGx+TfRHdJENfUNm+NE3paHg4pUHA+esGjqpAGnsQTU3dPFOF
pSwWcb6KAeS/mrwDDRDQvbdlO2mMYQYsPHCuLglpDj4ood6DDRwyiOyKG9nyPYYdn3GGj4htzCyh
Ida34eG/0IK70Yb1wlDIXKavTEwwupz41TgXfjlYj7p8JWXA6+zOam2Xa5Gs/T/loTgBd+CmpLHr
ZXEI1ALGnMB1z2ulpXA6cWPt8Qt47j8dm8kw1jkjGLRWzQJ0Q3hPtYUiX3mgjbkQvYQSCH1URAl/
ppvLbK3U9ZFpWGHnv2PmsoULCtHze5tOiycNo+u+Riwsa3KHwq6FxbGvuvGeFZoqxxLl29S0Fguk
gRsNAhXl++ax73S6TThq0NPdctBE+f0YvfKYzj3lVoIApRc3QQJ4gV9PWeGquBcwpWVXiRyUZfGC
lS8f0tXf3RAoDSP0AIQlELOqeZJHjmul5nHe5UN4VQRgtyCr5LaznEa/pdJQshN9bs0tIVXq8ym/
wQyJVfNnvw0QXRnGuyT7ZdmnXJVTrIfHfKHc2XYnoS+tJmjk5bMehx0KNUr02zE2F6fVkQxwgvoL
YUcma0+ZyFibulpQuTqFeZgAJSoajHS/iKUZl3D9JcuD6KA4sX6E7BlIj3+VwZMe97UiDAev/gdM
ZGWz9YhmG2Tdiwo/G3UCUiQ7KGnY7kH0fDHDmnPMn7bDsDTVtzBwwxvfLidSh+MfJZt+Su+UeRHG
RtnwOj+yqPusLqSE2Ewn4K91rHfLrocfhG1g6HurQ9ZEnVzdJrA6CZqEFSPTMp4rVLwy8w4Snh0e
3ClcB2sutAJkBHLoK5B+ZeKetzWEs/VStQ18v+cWMED1kIFMFHty2mgXpdFpXThQwfnUc8xmP9Yd
O4lD6WAIQXZuCd5UAynR4hqxEWZhLZ5xFrx62QQQYBmmqgbPl1AHKZXkC1P6u2k8EA1B5IBpFd4M
nUuT5JXYzpqNZLBqBurvWmEkSU8NCsoNKge72ZypArZRtyyy239RhMFX4OUNxQHEWWT8snCu9JRk
4y9DylvEZvFLfkOaTo725jR0dA3gc8jAZ1l4yJAlpHJ94erGHtVw1SKvLC4zUP/kJqZuZsrTh66I
mMqvwb2hnIhyPbCulidkhtsj8aII1AoACkr8oaAdRHpXzOAevLhENislEpYisyBW8SKOcq/K5Jbv
8GUxW1sP8Jlm6SEq5hamy6oAv/LMQ7gmWSk41AuEfcHIhMgCIy5R1VXvy3VSpvBAQCz/VuODIl2H
siolr+aKgU1C8JI9vdN81cWGv1PqmTvTuX0Ld3tQNLqGNA+UDlEAbqfAiuKniop+EQy+46Mq5DqR
pISbFm5eUQo+PoT2RhswvXJjj2Y+b3AZgo6gXZaBFpY0NYQenXwZWGyf78QfCjiMz5FnjWbTTxK7
7JoF2g2DlzQGZpNLw+SX827u2ZVM5px29S+Pj6TFM+CNSFHQMvXh5hCmf0YH1EqHMrAYoHmgs5tA
5YPpKWd734jtOA6PyqnfnKx9VrMHlaq/dXOcjPzgFdc5yyM1ElaoyZRNNTEGhr79r7nVHiKpvMcJ
gCnfj84qyRlhRr82z9vluiXLFOEIMucut11wx7J5L+f4Lhu045Z7qTIaBGFEWVmOQAcK3rsA4uzu
a1eMXqnlt0To6h5YdBAAfjPb5UQvRrKMcQ5OJ4bVfU+aLb6S1bFqDFcetwqrFbZFabAU5ILU9QDo
neyrIt5kR9Te4IBIrYxpv6RnQRATkaDr6yuci+roBZ3OhHW7nojbyB7fZicB5DUhGka/dQYNb64K
a8vEjHcHdazafm039MC6k05kgcZFBJSIJHSw4H+llIaMCOzkRub0dBjzIk/Vk1OPb9qHnG2bNPJg
Qw53bdM7Fwt7MzqV/M63lWSq2tFLkjoY1EXCBNDE99/UM6hyJXRgTjLgA1JQa1l1s1+2B3xyRUep
4Iesh+Z93HtBZhP34X4Ga15yefv2jSYiLsQJ/w8tqU/Semm3mIIBFn2M4OEKMOd4SAFuSLg3Tp8e
NbupnLUYiAKUYz5hohW4AB+7jxPW4k9Okz80UrpaxyBS1lw8vgT59wiEXSVU8H05bJJm5L1kk1lE
9M5t7uaeujHdQhQrZCVcIeczFluB40cNq1NSJ5a95fPTAOsDJi14Y3sTVXXgO3j6b4pIsuVprOGl
Glcq2uepUVG9bgzWj13RThQyvkmrTSHeFuVjWE6aXnbhvujY0n/ibLnu5AMyMYo48W4uXcFvv1AP
jAQibWspDxFLzGtUNpY1BUDneMSEsgR+O886L8Gyqnw8KXom9rZ9pyMvGfTCsseBsSizG5vFWRnF
AYkjp8b4Y2tRK8BDN5HZ4W6DYhCofbn75vRmOV92c2hPcfx2Mhq6zfKQqAJexlUEd2wrPel1oZgT
zng5D/otI+nVCIjP8E3qQQiSjK7rQLj2uowOuFegNF8W4Dm7zVb/dC4F3kb586IcMl9uCN0UtBNT
dl5q2qbx7VuGGJxKirkYejffLT+Sz1vzzaaqQcHfNJZsPYx1YC/1ytUWGrfi3TQjcha3Vr/RRCoZ
b8unqwqwW3cI764DfcqGXV5Zl0D6tFnQmYIvTen6FGE0M7fyebzdkZscaKNSfpg9f2Pb3xk8edrs
t/wb29Fn6ARfQWAtK5E0l4TMq/ACICIJy+4o7JjaETe/t0A7MluQzBHhyg2REYkSU1BVD4z2Rs5s
URe8faukdtIKtUtq3X7YBgLfgKvwRMKVo23NyskbDIQ+8u6oyya4C2pwAG3/d2DJ3qO1wW8lq/KR
4Peb1sLUh36LQ7ZBlKmO3Ky09v2sdMmYwCQ7xdRuN61pIQ9YKRBjinrMIKv+yzR96/IOavphHfTT
teU7JzLgcSuTi0BPIQyUl50ayPDyDs4WWMdi1sJTQ8987eP4QU17T0UJETZkOmLgNT6XJfsbOfbV
Y6nSlzd5R0fHzFa0yi29C8u5rACohqYaDg3VkwSuKrXX4xPIdJLzvKpWNTOhVzPCx5e/LziZ2upZ
P9T8dihtptmh+xF8Vi8YAbAhDhQQE+jW6qpat39x6hsSrQprNVY1HuFgpScX2kdhEY/Et64eiR+A
qDFdt/X7wFjBTXUqIMZKm+yuoyPdMykvPvt+6gM65du/xsSKMGSk6SrV4MgLYxXOV7NiH6elS/CN
5UgepegTrrFpbv9D8R8nFNyQ6kFuEppFdiNEwyNsmVWHgJZut98v2ckfJSiVEBKwQvWbhUURT8HN
IjJqO+hqPo0aTG/OA9Q907rklsq8N6HZzXqhz7ne5TAcFMvpP5gUAn2E6dkv58eRXv18PNqeWYbL
CzPfFNzHLWN51HUawOaqe0epb2vPlFciSKPi5B2ZgZRlDv/DhNbn3vdQ6Q+OzxIj0VhzrP32Jhys
3YoRX5BCkkaa8DNLhJnhDYWPuOafWVaZBY45IGutzNIRs6Lm37Pf97c83LiDOo2n6vKkAIgVV7Lo
dGk+qhYPuFzKL9aXtp/GdElwfoiWmgJjHSZdNBkz9zkj+Y9ZuNR+ksX/u30pWrCh6l2wrpgq6J1J
uYUJayPOJUTW1eYrekvR3wxjiUO+Um151wNWlzggg3D5/QmZUOipveJLdAuLKEsGNMHGxh5vCJJS
rURGQDGCvMqnxkyBsAyIL5QAIVk6cUnjVh/njlTY1TcqcQy360q0kSljSIF1CsuUGfH239qrq18C
FL3rXW2job/GDf92T7Js0pyUlwkx38xU5pobZziF5hZrgwZjvNu+vtATv1K9fPFTiKFYBGa11GSx
bt5FmWZcgOzF+C0TBvEwHu1VbyQq4Q7EV3o/Z083XWAxZKpMdXOQDehEPEs63peqh1iJNAwnuYNP
LxpiRti3/1vjKYK8rcrRpB0PbJMDdfupLCXvjXQZI5/A1t+TE756ll3gNe3pEudXy5nsYJ67QyuV
QTcQYeV+gn8DeQ0yz5M3a5gBt06q1OVxT+r+gqSF1ClCEd9SCP/MJpV0sMPW0JKQWOpBrgewaQsc
lVBVYbLCLTouk8PMTieAKnz2uVk+oJgIQrjZuuYvAEmgqQSWRHIjoL8woY59U0veEirl4h8xCF43
sPOXAZzCmtZuvwj8w78Dp1KgOsMIwCiCVEDMu7ogKAyB3a0aJliyX8SXe2SpILPtttyNNcp7zwyz
T2bxJ/6rUVnFOZNa5/OYincLmN0+l4E2h2U/rssvb84txoSn5vzS6fcbo+ri4A3z5SP4PlzuyFBw
LW2YgouVKS0oc/e89/aHB/z5fpqhGff7ztIk9wg3YZQIfYymps2OmVmxBjT43I1p30zAZMKkuTKs
N0DHvMUqaQhPVwl+faZOFxGw0dwa4CnUUfJwGlhbPf3wnJmhhqQOpFSmLf9ez0xK18GDPHwlxEgX
+rSWYOpa1G88Z1ty8XS7KsmhfnnmSb53veguNB7bdCwx5sno1O3EPOx1FOm6c4VJLyHIu8EFdQGc
FqcucZDyu0u9pwyG2hk13bn7MGiQbrVGiVSrbil3f36Y59MG9VmciAoKxzVZ171dTgO/I+UqPntI
fTeQ9Z86CfnjMrl/GzbCZiYtUQUJvPT2XWFGkBev3t/99i1O8BGjLLzhhqnE1CrrfPqmbxdcN8VC
FMNcaucJE5GfNYVcDwzg2QMfoAQoAvNQB2yWEeErQe8IYmth+60H5qFrvFLhSF+8goWtFAmdO9fr
8Zx7tV3FERI0ib249qV8Hu9Wv4u+1t4PKgFTkxjbKcV7ITkFRDa/jRBABgKHASdKuaAgvQtyotwb
4HXmkt0rif0Cv5AijbuJUTQikhXN+2WaB01kqaVePCddadlzkl9qfzlR7I14iuyFF12hqOYs+oNL
VF/lGwIUjjLRNgN44wmzyaDafYzEl6iX4veAQjX3BJBVKd72Pyf5kDQAi3xLdN5cjo6XwwMP63cc
kIonM6ks/q6HYj35pWqpC6Pi80y40wnguiYGfJk8vxF/vVfdK2zcC6Odi5AencGLv//EZLApfvPN
Fkwff9naPEybVl534PH4ck6hphhFwwJsbUDuCGj/4/E8C+OBohhoexycKxkrCOoZwZ7T78R9bvfj
RM/Gpe9M7PdQYjlISG9lOfofduKuG9weiJUBFYC4O2MflzXZLQPj4zEDdOWLqbR30mzQJiqnUdk6
YZ/E6hbRYb409UTJa8ejIuThOkKm4pIbKIpFmx61yiDuGyx14BkNWhMTTxo13kDliZEg//e4ggjV
HAoIbUcdQRdsjy3JhRtpLnqQE8lMXQNhU8ZK8IOKxsw7cEwLO618RW2qTgD/Z+aRuVUwlhvD4k6B
T8bQz57xCiWzWCfZktKOD7RdQwfolebIxWHSL1B4KQWmd+BGWJIpkWGKjaQ3KXdu0wbLoi+iot7L
CaTfnwHDlyVoOo/rrgpp2//T+F566/52xHhCb2bFXboJNbLIATI/HEZotniqD51SEfezQ71OyU/j
r/ToWzKGvhjfx1OU71YR3buPLuMG5x1N+AG5C7yCgc8/iIVF6VZW4foOna5nLpsCy2yjRrDgVHM2
aDZLWeXJJ44Jw9l8+YPYSP7wc5UEZq4HYUGpCrEv7d6D7nrNNl4n/jkEYBZHFcjFQHjo8dNtuF8G
Vg+D6vKfwFOtYtlC/nfRupbfdjzR+umoxsZhguUPEet51ROrRMSygYl97QC1RL7iIe3ciRXQo6E9
Ib0ywknLsw/U9DJAhU+rfREiWSNseQ9vw3byfHn9W193toBXW5Lk+f+VMMuvmVCHMApoD2490uj+
NZIuSPwKOjSqfVdtCQoZ4hhwo+/KY34mve9f3uoD2fCMQ/dwQSnNOIav3SFWSGlAxCQWLxuCMRZX
8JjIYGMHuiJy6inzR0XjYDMiWWvVm4njVNr/Vvk8TjrVs0QcNuptB574txWIUGNtmpwgagYyhpIJ
WK8r3tfjQB2kpEc0VG6ntyishl55nzJHa9/bkGAUcNs8xGedkJcPvep+i1pqxJY6uC7/yS2itA6L
5pt4ZLYXOhpdNlahPvKycPR4wR5apC6xLrJm+IRvqLA4NJd09i1B9mIhzoGYXh8tkeULvVp4/utD
u2kUK2J1c53+5gqGyDlhopH9nU7JwN008nciPnBRa/ctVI/BSKuY7uQPLtmiY3aX6ehn9mRQg+fP
Z/mk7s3joJhMBLnKB+ZpnKlZU2vufNNCqwovRJyo9AqMD0RCm70WwTy//3QPkKVjZ0hUqENedBYX
AamVLtj+giUWKnobmAOrci+vDfc5iim1VlxuROZe8xScVo32loWAkoYCPFp/52n7DF7/hvsLdOsU
WVvpcLMJVV6uROipjRvkQIx+VQWcXSdKB39SOsLYUpKWp/b+7dk80Wbmh3qgDqAOmheXrqB4g3GE
3NNw99LiGxkUQZqBNZ9ENvrHXwF3qS5Zz+fqmolSWAj8XQP+xlA3tTYnBZ8YC9+I+s0+a3Y+6kb9
mZjvv+ZIZRaGC9xuCgDDe5sGrD0wkOjDrDA6DiMWp+IR66CfGGW+W7iXEx66/aBJBxNr6GC1hmGK
EW6KMCx0NSSUYqaj2HgA2E3ZvNM+FwMUeev4ORvmZ31U/0obbtw7SM35UmGDoLR9LeXIh1f13ole
MKa9CM9+/0fLcsSBodwisaOSvAmZ50CKyF1CNjDBoTLGExMKJ9+CIidO7xQK4h/aaZ8phUhj3mla
a5UY+kiYOrmiPNn1pDa8b1B9iHqb5trjk1a/HBuj1H1WvxpW0Qbig/qXo75dpZcHF+9kDuUNAgSb
M95cPn7ZvSqOdXHxbjhp4B30smcTBWohCVMBvLW2D+hFzdRDJHcZkEy/JjUWI3xg9nJrgPSjti0y
v4C93jR7TEAUY6HNeDO2xbS6q+ZnNFrWOhL0wf8affDeWIbrHMh6Y8CVotSTXazSA6lw+UCEJvZc
UbE04ThgeZqz/cH13bVZR6v+VxYI/ff6itVbMrc6vM0dQrabyZw34Oew8Bzzs0SzGh0RdQTdJH2F
CsHazSYoSv08DzkR8+Ewx3acsvgHXdwNAS6EkR7vrz5sn3QGuVkTSi2XVpCzB/SPJLoby/5cBuaU
+Ncv+Dvda8/xuR7iR7OjP2qNQBXE53d7VMHBL6zMWAunw/poC5XCGpyJgmBDy3YwkVbP5JczzPkv
6ArcJghkPe+zjbF30jDReXTVMs358MCCS2EMjKsCBixbbDC7gno56jQe6D/Kdju28JCE3O8fwa2R
YhZVxgbiaBVV6J5bhZsVXF5AQBe8yM+6fBGtZHbC7g2FyDAqWS9Kib6GOiyNwKvaVVNR2kbhekAb
fMeIhY5QcdQC/GYYUp9kxoeiGE5Go67uZF3yY+R4uAnMcjcgS2HBwGxxIS1G3HkVbKNWhO6gXpGR
fX5HHBi3ElaIxoF0nkQMHzgYyVn6TiwiKYo+rSJTVx/BjjHgrdlYfT9qZt+DzYzpPCMYNwWsn4xV
DcSx4iKcPiy+22wT2bP0ku1yql2U+e7kpWlO5DRI6GpluAs2/B8sCEvH6+tx7V425h23rPGGIgyi
LCW6VylGWMdWHLSsG5xOnpJxrOnK4YFfCU9DXjbMNyuCiZ6LyNyvBsfx6IajSMNlTlq3RfFGmhVb
rUpKFg4G6USruwio42iEg22y1Syj0dUgK5xon3GbrqyVYaA63Z2yQoOiR9KnChmWuFN9CRxE7M3g
OHpM6fVTXQHNrTc3GdWh2b/hUk04hbPPKtOXDXqYQ3Ic8RXYKP9xWn6Sv1u30U0r902MpNNTunMF
Ax/Ga2JTcdeb8YAgmq393Nn3H3zUb/b9srhq/SdUiCYyAXdPLsG1flzbBiufq3HnSE1Ig2659N1L
Th8cek5J/IN4H5f1kXKtZU67zPOndVSzJni4JL4b/tIaI+4ea7/YYiNH/cBywIZGsrDeijpu0/D/
JoF16BBkZc3UHTCl+eX32CTnKo5eMG7YlNRcEdE0RsUmOVODS2ZH92ikulNBsg8uk5+pkeuDvdtc
oYyXyxK+u++7zKR2uh4MaI/0RXy8nV7Wbyyt41TcFoXrEMk014dzm1i4/wbSg39ReVs7A+hyjAJK
qwcdSbdHx50ooZ1gB6jpeCUGOBMcBBlbWCbTT3k+6GtuUS0LRWrgx1wdykEnOJQIFeSOwWfg42n/
DfL6n9SJtUsXonZ0nsAat6k2IzmGYgGcigibmNRwxs3qkVdJtIV9uJz6bOgWSngDsp/rP73BW2TS
uEICfhYGC5XqbHAyiya2p0rZYi5cxVfth1YzNjXQA94uGEyPizgTQo3AnqI4qzBnQcsY8AW1+Z8Z
q3A8uRRw/q3pNcgxZpaiFNZUNKB2bzCWpqUG4LPlKKYFrKg8uVB4JkA5ZeraOUndIHeYqTqj02MH
swQOmmoHNY4Su16XgC19hh1eXMkMPxaLYGJCYnBjPugFUu2khYDVpOad05nGFC/+Mq/viLIkbNJe
paulqyDjpoZ0J7pIC11olvegbGjH4sd/ZqbKsOKbaJSr36xkAB7iqFuVXT7CkVdlojxlkhomon1e
EatzXKhPiMneZfQVVTzj36VEnKaqhyYd+/yxxFuP+x2KeiP5GH7BFiP8/Xo7gzKCBnGPYo1GGzT1
YY9FxoxoEw5vkjs/MIjD7ioNQC/MWIpMIQsjlQS9fOx4ZYRet2jyAbnFKybyw/TH4G7JvGYXDO1P
GQbG/wvKB54unwdNFJakPhvSwxiDLYqRWvIP2X9EuRg4bNfyGHDTMvsgfeJGkjbApUgoIRc7+e7L
L6NRkOsFF2eHbEn5kaSGsxGBSKSH+EfKBRF/ZNb4ujKtw/qXvUY294m+EG+L46FUaSBq3qjG4Y0H
rDf8o9j+DnXf+WEMeIoSABg5blJ6JDcGOWLsH4K/dsX1I0GaVZ9ox+34xIlUEieR4Pl5VjIoJ9+C
e/MPRDIeON4+OFkCYoQV3/vjBbaOZ3h2wxn0gzAmyBlLyaILAXkZr/tnYgtFM2t2xdsxVn68T4uc
x19rD6CzBaCR6DZcAr6W+ogZ9bbam8QjWEzq32YAeA9yf2lr+nqV6I8eMNxFD4voawCZll9aeHeI
Pk4TBpOvX5xGYUF+o2Kam0JiUnjQRLaViCxduxtB/UZAFag7gotS9YCRHjSVM+ArN/L6LjewbQRl
RjhRU2MU2B+jyGvFGBq6Kyay+VGdEzyx2N9C6vXP5RcEowAF9a0vyMloZvS6fQVLKMijR56GOkUz
59+vSkCKosTx3b1R6wZzmImWuT0vurKpi52OC+JURGushc99zMlUxCfn7H0nf60+T6LV6EZJz/eO
/rsgMAMEP1aSb0X8lnpNVwK2k54dv/IKM4rV4OeJv0i2SVMBQiyeotY37lAJH5Maj15do5JbyP/4
ppBO7OoO8mPQXD0igAOwaB4OSQTFrok4Ifl03i6qRKkFy8aDhVGkPcAB4xe5qBaGj3T86Yjg3NXw
3VBvUnUH4ROMOU6Lo5w9GY03dA4qUG7cwft9nEVHpN9qn+xe4glSdb8ELtas4Eutk8uik6yFHxfI
43Y6tSk5iJurYPeoa7aLbbhJIpUcNFamR2qdDOtJHOhLI2b3DS9LeFHwXmLthCv6TJQPdl9W06zs
PVDoF1epkt3FNW49Cux38KAdlaPNCfJyOFnsfSeyT5ns9eTxTSn1P8f7WS81gzMU7Ivyn7kdWwJz
4/o/10K43k0uSl08CIn0WKNYv7ceuWRwoHaQGhTrwBZ+GLz8VGF1KXiLx6KPCp5b0bLKyaqHS6D8
VGOXMgzq5cuAlFCLiiTsAYCXYgpYQiHU2BN3RGvK5P+PoQfgKlMcJOE58iQc8oQzyNElwTk2XI6o
shH8EmeCQT/MmgGH4+xu9q0jiG0+H1HWQNEKqnlVdSfsjvyn1Qt4YAc5PGZvhAM7f/bOkI4mEmya
rgZl4xYMbVB8fZbr6ktZUclyGvE1yJBfBqvwqY2ucuX5Rg/gePejuXf54KB/KUw94vUYTS/4kQzg
AhdNyLFEzSzxR+Qxlcfrahwga2NdG8mj03SMznYD5WvRg28b4/FLYeuOOyu4MtdGF2XFldOxMjjd
rj6ZiOC22fqwQrsisw1qHxSExkGxc2jpHks2ybLOE8GTIYAaw7rl30M9IeUbd7XoYsfJIs0+L8FS
8M7lpdcePKJXGlZvh8W6cvKR2XFf8vU822SNFmBT+aeT1URuz/sj9+Ngkw77TqcU/nIUzLu5KaAz
GB2btsX9W/J6Juot8RLDLDE7XB5YuUkebn/PKSLSIDMHFxAV4CV65UgKR23NI23Q1xourm1bf+UX
q5hreR2BPgAw2DvpLhRK8tLq1vLgiLOkHGX8J0iyz/nnt3HHS6m09iRfB8yYmEIzlh3F41sZc7bb
hVyT35zTDBNUMtXO4OrnusgKOUXyhOrVTQ2N/DmK4kL9G96qUTIKjU6H5iRUTfHLQ5wSf7IzcgMn
qAVvMznDcdn9a2G8SQ1RwYfwdF28qNM+5k7/GUUyADxJ6pnLZnfsQ64IoS3kGt7jcOpsCDWWw9GW
+RTT77i6lRou4sRzyXp4UDbVQxAmUa1wMLJ501QfiH477oSo6Ft15CC0RCjKIJVllXgGiFlhjHbW
RzbhLU6aDp2DGmvL962CvmIwlDJUuoWZ69pRBeidduP43r0XtpAjXbhLJaX325j3lvGMr4ROGJNc
Po/L2NZhoGe/rhk8+rNC56469PHD/geq6o6YGZbsJfVDH1qzjP3z1O7swkLEB2JQ/qThITBpjHJv
0E+bgdylNIhA5oDkBkiH2ZbOaHYjfXGyodMMv51ElusrtNhoaN8VjvPTMczjhHz5BvqBGAVTFMYm
7YrAewe4xYC2lUII335uDjTs2COHGKpFVvaus8lEv2pp8I7F83Ce5+oHfBdHTvSMxKqYUHioIlqQ
CwVfoOeE7LaaQzCTOcxP9F6/0iNOmP9oafWKr/ToZyqlM6g+T6Sx72In32wVaOzMVM3lDEfTPpAD
rGcl8t7mzDP634DyV6KueG22ZIQLSHBbjjhcxuEJ0pIKTvUtMdmuv3DTPcEK3UX0946esOGi1sWo
KvNpg3fVrMr3mm5FfAf2gvfQ4qL36iWXxyOK6L7XpwbSzSX3iJIZWSZc1SsYfZLeVknIGhr6IjZ6
BqhRXjUvGdx+z8tyjNeITFd6FboveUHzMWMrKfwMEUHUhg/PnoiHQMlSHm5zCsfbvDfWzmCYOPIN
9cCc3EVgigK85fGQ3kbEcqoWFoYWWMCLk1RE1q3aiRsO/lHD+9laKoITYXQuVMQAC0RR9/mDC0Mo
Q6vIWam8ZyN4mXYwYQNsko4bXE25x1pXptOz2EQzIKvqNncLfjDpkblBZ9uPBoHFFvdATST2+NJC
+ozxOBxqqWMIucZNYyA72FVS8Twk/fE9XmHDiraSswnasXfUSlL+QeBnIqwjKnbf/3Vtkl759YQ/
00QMUVsE2bKv9GlIXYlUK5ZngfvO0gdTGZ3z+Mgjl1ninINkNenAvL9c+gMcIIOtTVFXf5V8+e3r
6SkNrWYUnpHQRl54RnMrZzwPKVNEBe3XchlKbvpvSXuM4dkjrC3o4A8yTxxo6aSMP37rwO6WZNqX
I6okXD7SAofnMtUbj8xL7oCwguYGTTOGFPY62WP6qaV1f891SacflNuopcPIn1JJTTbuyAkVFLMr
0roJNN05hZQyUqEdF2BW5FtP0wGfiGQEAo69ibqBHg2PPnPcuFuP62x4fTSsyuf+wCOea2e9W7KR
QJASZ1ns9QZDot1QSkkmqBguwCKvUHUhHLP1VIB6JRFZfPsQcRrl2nXbbtPSxAuhdo0173BJQ1T2
AeDDfRalL1p9k1poGb1NIblBckfNun83d3BgnlsYywBDSN5qnhy+rCAxJ1xQVUiWuCJ+saftBv01
ZToyaL7wP6eWrUOeRGvwHT+i/z1cnk9jcH51qeTywcqB3E19bJm0sODcQmdYNYDB2BgoSyS+yHSZ
FM0EECvLcN0yvRrMvaSgytUQJzUgosdMeyrb6bPc+Vu7hZ0IdArjSHQy+GyVcsUXOnAs3mfFMg55
zm+PhvIErAw2HnAD5A/pd5GRnWphX6YagIZD/AU4ydaFA5oCbKcb3GM7qugh6bxx7NYDNmlqN6Hm
D3tw1ukCsXYX8OYzOtrR3qKqwPQpMGMtPZHg1Qt5Xw+WE2KOg9ZLT9v/UEyDoDQUeDUzzVs9A8SH
IkpA79s2g+Cb7kI6sOYWm7E8Dby0kBKVym8rPKMU6KeSP+ueDC/JNUnnw+3CZZe2ViY8SbScWSn9
IBHrdj66CoW/cb5aZlgSSV6QaAHstFU8U/sEFTUY5VJnBDaGXE0NcaF+KDS4OUeOa6d3iSCPDX3+
v2LCVdOFgMtb3g3DrKAjsSOf19oSQSEZKTn+spcFf+SBMCvVLPcxxaNFNuy+sTwGVt8Z9mv1AOv4
5yWjTzcIygWUHMFDrBQWWTLdOal4jdRR9M/xvcBpsJ4ioleOuMHZRUbrYHxMtbr5KMi52cltt0T8
fdXIlBsEgp90hn7EzcIr5U5z/8HDcEI/d8zUnoyjafnzijYyCTy7A3tCz3wgH1IndYxnFFo1YwzE
zhQpvdNRhvOa+D0CFrrgg+4NyfUn++mSa5QWnTLvSyQO/PqAVeUab/VJyd+ySN9kJ6ZJahNQ9j7+
5nSb1NY8TPlkPvviXkO3vt2sr1SQ353YG7n1LH8Emny03Kdex3+6Py9zs+jDNEeGIyN4uaQDZUuA
lUo9vtkUtvfFbRHOP2PpPRheqbxBFx9/V9u88mS3WGhAfQBZlXyhSaCsGsvT5zA9zI1mhAJAVzeH
zinYE79JJkN52SrT2fh0cIvi7K1MHTSqMbBWwlXT8HNOaMy1Fawiz/aylOLbumDzip03qKBC2f/7
FmwwQjBBfR/hqZQCD6VDTeoMhY0LgNCgAW2C8uH58ZGF9ha+ScRh8ioCQ3rtFbur22PlUmX4cyuD
3UNCwUdVNivrxfOG/B19tndQlfwZGxD5nYJyhuRDMxffSJsKi3T/KGUW27yjajqcZuILZTTMGbJ8
UM+JJNnykBFZntzLBC4ksY/mo3SUs54P6OuaXNeGtV1cde/uaCDfoqXbgiPPsXygCkpDO05vD2oA
+DdRp0MRL1SljG61RaHaKKYreqclb6Ip6+GpZxxgqgndJXjQhHvyUWqUd9OmrB+fnRhSXvk7zVEI
U3cvh2vXTLfhYNhg4x+Cc+3FaNhR9DWU5kjtvCTD7txztR/mwRcZRWxg8VB84QJCR7hllGJFON+6
3llChX7YOdgKT/onntXrKu4moI6BqMkEJLR11pXK41xXOMHBH+RE1TKTpyFwIMt3g1g7qHm6Wnm5
fkHgWt6Hh7N6t0h7zY5705kEeDmNHDYl8AG6FjqCYDqH18nwmZ+dIndQaBWG+spW/mdnHwzbt6lo
Odb1WrfQh4IA1xwanhBZWTvxNRz2Ad8ewWQqgqdisRoJLB2uuxkyRrm6U2QGsxgIlR9QkzFInIHm
O/DCleu7KL329WHeQBBlNjTmq2ntftpwJ/31s9kmQNj+Vi73Io0lwrv0ggrX2K2V/rToCtpXOSs1
xaAKz1BJA4a9LTwprVbgChYxt9hn82J/Rqf4G5rChcSBlx72tHn0xPzq7EG0TyT5UhMjhJ+TbsfV
cQ2RdPnXIrQxjiEO5kC2PVg+hIYIZ6mfKxRzXW1SjGTiSjfRBZ2ujJnOKCz1qRCM27lBv4QZEdZ0
zB30V0ceJKGFD6Zf1rQziPhG9ffNg+6E/B4I2Od0dinu0pLSvxOaNTA8UHy6ltSCZG8Bwd2dIcaU
IWIaKsseSbH5Qu58StLzxMOG+7l7AlkOWLU7OieZ6kQK9V7eyfMbChB8LO7QCYehSio2PAhLlpEx
1BR73acc2DXtCqdN4vsb9rMZbhR5P1bxw7wCMZNS8A+TZW4COddwsxGeAtyTTSrzL49MP9PTZlhJ
azBRIntZPARUnEFCj4JvFfYPxEsl5KCisO+LTx8rWKzOG5HDHgQXOpK+ZD5aLHGvuvkwQB6XiAUT
gwY5+/5ptprHSs4jTN5W1lWs2J16UvqUtvpP6ThwDqjDX0bEF4qyYK9s7KY0VGm1e3+ByCuCbvLS
SYjd2icTIfVHYfdx6cl27UE86HNfwkcGOaSgaB1IcTfn2lDN0hxU8wiv6T7QGOoZ+GePVhcbc5pa
zLt9yy/19nM4ROqRiACXr65I27mrWSHPgbEX/OSI1Mzke4y5gkJ9X85JtolW2KfYa4SPFdBo0Ywo
6N98ZMVm3dynKEAKIalwjLmQ0E3qQ6dI7Co3Ge52QF9q15/c06cunpIyG7iROPqtH2CmMuiPO4/n
udf0wYfzD93kw6ieCaOAI945UqKIMg/w3hoBe0D2qdT/t2CgStIwcnc+WYj8Gag7LECt//36GXTw
UJY49C1TNkNyB9FpyafEaogPzODd16/w9AN+P6tBI0TixqOwiBXLAZUaKQIh6VnlQWzsq+wg45Y1
teH61QO+IbBl74BvUFxiCAiFpLuVbJuI6DW1mbSlF0pxZSpnAQ/O48Jy6fz2C/JiHskX4ZnS8W4Q
NQAzWuzJnoyipvuUzE+1zkEbfo67ntB5+QqsqtUo0x43qHHSKMusv+Ju2h5dYfj1Qi1dbWhUpleA
Bs2Cy9zaM5MIzEyRh9hNNIW2rbo7uVLWQnBR+Izw+7rcJWGn3FNnrkm4lkQAW7oFpNlIvc9vimfl
yy8YR938+P9hM3gT6G3BRG7ZxIg0ZW9+0mDdVALl5zTv7ptICFLUDyDLISt79PkVaqQWSFbGkClT
L7fl6zQ0xBFbD9uKuJw6bSvEnn4giZDQJ4wewlLSueNH/WOp56nRRsFdUNEMsLb+Z+wySRIIOoPB
oavM5VxXtNS1haMA4baYoi5kA1aE5ElCvCDdVYpsCs7385evOrtSnNTm6sPE4lIcbgvQcVt0mMZ4
6JnClxjvUZJbzEyx0zRMWNWCxWKesWDVS1b9IMEhV90qZsa0SLOh5UX6zwEtd8OzBSCuIcS8xXMh
mWBFGKZWQ8dO4u7//QqdLPW9gsmDSZthNKk1HQmOSoRHQAmgpDsaRBAAKpUQjdGSz5gSiKGL8W53
SbGzECiIew6yqkY/Bn7bjL2o4KEJEtlK1NmNwzyPv0+lVlMeZRJG6fSiC+yN8Sukvd7IJUaG0/9F
Ja2dlYfNxi3ckMJJZ0oA4JzThK66GypK+jYm1MzD+mfNtcVpT5lFI/y9Cs6Z2f3Z9pdcFsPPqS5e
SWcnafdyGnu18RuQSFAal1goTktxNzKNsozLZZgmjLEpirqvnvpyCGr/1JGnD8NeftahXwxjpoJu
h/fBjvzy8tNl3TkdX8zgN2F7cghuH4pkuklMNE08HdcbVhMDpwLhaPflU7h0WYz30MhAdKAdB8/Q
F1MMnqz9hL/mpKgEP84JPfZJGJ9vP9/2iyXEwwBWVtPVx0WVDe7y7R8Je6nDq/OoDtQeehnM0XTT
7N9JSSKwsQOjWTfjzKSWcHQAAC4pllkjm+2OrRiI3lvZZ0dvEuRda0T48BbJl2dvSA6QroUd5Q4r
Pg3xk2hNGZyD/qxTnb5UfG/kIMlDjF+B55/9gPcMrlrirNfAGIh5UuN9vgS/Y7dbxsn1VHJuYPZN
W7BBRoYvoDpBEU5UPCiCKSa9JONQm59bi/m5J3p0GuXLwagtckZjORk8e1WfdlV5wn508of9a8NN
k4moXD/cwxdsmd8HoZ25VTEEGSIM4EDxnWLm9Cylb6oDdgzDLIMdu20CtNcBXVRBwV7z6mwFZSJK
ZpvOhp061UpcgqWRQObApiB/cR6rDgLYM/rlYLu+NkLzPcGJVhp7nMIgPWO60OGBZyzaJCHHiOPm
b4yDsTf2cpZ9mKWQwWDKCzPUXDteKj/R/OVjHsxeAaSiZmh4xt77z/jbdGCCVTtcnsvjoae8PMPQ
IzZukDJAkDmONKCWCQD9ueEfBbjg5+m/5G1LZ+wIn9f0Akcc/nXdVj+DEUiHMyy3sZ/J0jsZDDYv
HxCTddViTghOcByRGa2D/5IY6xqIPqSiUelmPJhT54xl1nJtSIpkg4CITDommWJPKuYDHm5Hz/u7
blf56BRAaJRYmjcIP/CJ3dJ5o0LHoqMUE98xzTG9QQ5hyI33USqHmeaM4vwpKbAWGyxhrz/L73A7
zyZdYkKdToSgo1yO8kUVtNX2tig9SOtLcx6aeQLaU8nyDppqKU6Wmtv53Y0et4DXCJM6SDodETnG
uWBz+Fni2ILLeXR27MkpriQqVeNgKQIhiMG94khKvNhm6nLbf7XiGMlrNplMbqNLYTbyva/mCQ8U
TY83TXBFaSor51zZA1sOQR1r8gpQxfj/xnhlQnIQqFaLIT5fCgaW74qQiPKtC/bvvC4NnBr5PLRF
8ZyLXEYNc/fp0B0JnOgWDwBWZXNz/uId/7Yj5uKurN3f7csnmgD2/S+5zIru+9BKGUbSmKsVsdOO
xXB8KLdFMvWbEJFClwkvjWTj/mCigqs5Uk2EwRNmKlh6jro5Gsy2cXhTQI75e04JwCeqAqe0X8xt
S/gcVH+ylRJgJ3slddCHa7OveyNHfSl9j00DlMGBbAoEauA8gY4Z6WRrugGgFAOpCN1DLuzR4CrD
lMCXjjdxgtDQUmV/90OW0rltgpKrWXATIdgPxgfn3zeqniUuxa/tXtx4SvmO/TcrGs/XY+ZmMKkt
OWmwmEkte5LPycflmiUgOHOl7mNg+/YTUM658/0IeEqkr4qhOa9jhUreWO8vmtxExxTcVYqL3Y3Z
vMCy/bEyvTRfYXgMw7sveeHA4F7sstFaZ13XkGYoSWFWhH9uUQujqatGLaTVp7WQ/HSiEjizupQR
RXhLMbXKDdxH1+UqkHrP91JJ1Zr5W0lj0mGqHCxlrnFpm0ZHVC+4DRxiax5KP6MrM2TLzScYkE4z
bJW+JVi8Dn7CDsiyF3vIBtirkzYBLXnwFDN35BJ3+iB/OReYtRbAP24QGq2GV1IBwW3qs2pAmmRl
N10Ob1+tnf2fyN754psXrN9Zyd3VhTuqiBMkSSAONLaHY0NfSLto7xwjy471ZHV0iUXrpYNH5Wnd
ZoEU6VrjkxOyPfhJ/NkjHfgC+C3ohAxV4+OhTCHHPO20C6oZV056U0Fjap8byU7sGt91dm8UYgxg
tt4oJbYX4vhL3cb9gr06/YfQp2Z4MvgEmNFifxAjDjmi8RVjHB8clnhIGU4ZaiiabssPN3aNvzkV
+zKLKfrO599O74VIAVpeh2U6gDR0uTNMKiIJU66tvyUpJcIkwjk44C5FK9DNOY218hZ2lsoN70gy
xAuwEk6uemXcfPE+v/IXy0GTtX93KNNwk1QcvWCcWIsK79vhGe52Sye+EHXwAdEdvLsnx1PJJGZN
Uo8A5PKSJjP//IMmhLPz6exuXEgWVNuguundAkqgGSdGzby/hTbjqhcQGAipaPFwoVQiI/XYCapZ
toS5GrbSC8txGIe0MJK4vZlHYSINRxOlXRDDyAboPYrjFCJ/LQCW1Vb11jYgUT5qmO4MHCUHrPPB
gYUimQcihGpFS0/Fw9dGs7kOepXtHb3T3oanr+nCqMmGaRhKAIq2ylLAUI39w6NRbz2o8JXdNRxe
Uofv3ep5EtCqnTO2LRuC/jJUc/7D+cSdEHApz32zDk4x7rEifncIRQnS/1+sCBoQ/fvPN83WeJ3G
a+JeY6azl1VIaDGGzGfOsVEiu+/eIDAk37FlMrnCfL2t01TB7Sk12EhPWcYONI8yIzS45FIC6CdF
zfSCmSmT5rLPKeaHLP03cuZJKNP4leJfiy6EAGGDJfcFPPb9MA6J1p+y9963E67ln9rrlOkvvsoI
Jzndcj4idqB3l8yOWqEKgCj74PuYlMluE3+wr5zxnmq17CuHBM3L8b3I/+QpMUTaOQUFAeVvpcwc
Y5sO9gtxIr3zS/BQgckyRp9+eJ/SdaUfzcaJtzOCxaY7UZIeiA7MuLMHz5RcADTKmtaAyUcfHda3
GMuADluDxo7TZRmiODVI/Wr2BOWm3vcEY2wXWG2lXKRSu98xsDawE//qf7EFYkEOsINXm7hoqj4p
P+l6wqg20vs0jnEcerUdDKYnjZOwhysngr4BzpOQtXSbRFKBYMKfsiVF+scvXdCt+ZbDcjItT2XM
EAl125p9Hth4DxIB/nz8fcldacsQiA/6FvBcFdiFrwaSsaDVFwWn7ggAs2bDKzjNt/KwQF90dAdB
CG/S2YjFl8M0t+xubEug1w+TQND4OCg5SVC92t6S6eYg6BoUXqgzw+EVqlAo8ve3hlTVDYbqWPUv
f0NNipCGomniL7fxlsRely3nj4XfBRejJDUW8jRsktWIbzibhFD0urBlYqdJ2eNjnx/25gk81lYH
g+J4OTsV/V3v3tsrEMxhp+xwNMMoFC/f45glfIoyS8Dp+ZXNCbO/kj1rdEV9ytwzF7J0QDgGkZJZ
BWNPlHr2ZO8G/9Lwoe4/c9FFbQXJSEvbgRpOYQ3EyxqZESPDZGFnlxmT0/2AbLyuzlhYM3uhCiyD
bUEsh2E2mm3dCxHYoZhurxsmhHuAxa2i0l9O31gOsI4/vm9DrKCbsyqcr5JRAaDqI9Nm8CHzdbti
siXpJ0rix11NjH93y/Or+DJGOq5wu22XGUck8cThfhx5RUozen9ijicFZnwW1N1IeQWJR61ii2AK
5wcwJlvxq0aDUxCpAsxD/tSKpHwjc7QZWqvTl8oi/OjeB3Ozz8y7mYPaeJQ3kwaaYUb4VQkdfez0
5TQ455tzjI89QZ9hPJmdU6noneD6h4N6UC2tmDxWlLEchTeCKOQ3ezA/6QN92iIOGXmAoOEBt1qo
uC+6I7l03pvg9wlG/uWKj/nTCM2xYE+Vl9PtsNrrDLCUirOcM7kakCOSdmFohYq+3eNl9B2525fc
Sl4MTl5RwnyY1gYUDb6mj5sgvIVRJB4RKDxEABJLiH7PNIzEWjlaRF6X3B77u3rrXBVbkSC04R3g
P25JC8nbkl7xGJiPj6eH9CqelTrDJEiYOP3Ks29cxZpqICdpq+VsKNLncRERnD0k4pi2PYKrRQF1
hL81jz6rFxsJmdJ4tYm8qlVQHOPVRaBeKfK8LhKZXmqjd3dpzigk3Idye+YmbJ/9jLHpMnLTDEhA
J0ZEKt4NEopXnu8nvNfshXGKH76Bm85Kbh7uds39kLB3+UUgndj371UHybig02H50a0N4pMt6qMH
GyD1qsXcxoQosLJAj7dEM5ietQEC7bCgHvC0wRF/usrgZ6GtCPmi5EPmpTzQ4NTfQVPIic+NeLvN
+FugH5PCNRIZciDS7UihYNsnP1x6HtX0VUfWqn7ov9XpmsXnrImdVa2wLpoews1RBqx8yYfzuFbG
iyNOyhmlP4tIZ6+r2bUPmjSCR54t4dB4Ox2Tv6vBrq15q1ngPss/p7bMuO6C7uhgQ+XrkIsPM7zH
Cb/1Gt6hojAXzsC8hML6JaMnF1hC00nR7DLORf9UGdxL4mdfPtU7f/KbuzUEbrPs4pexRp3tPSha
wqcYr1MikyeAdoo1GFmqQX1Eg1IcLA9HPjfsgHGF8bRL8584NY06AxjKvbvDQA3sXp3EuwwDZPQt
fekRGXLsspVc1vD8PlzVWSS6ttyjpwn/aD50JaVvz1GRS3NGdZhAkuY8vVzbN4nWI9XeRoFHmIX/
JlsPqoYw0lIIQTO61brBb63shsPOwWTNzhkckCKKJvFoccn1Zb78mN4s9PO/ZZpN2psMTvPo+urR
/xZLoy8xtHkYCsGzGCyakOD0107RjX61y0N6xexXRYOMOkXNxxcYiiDZHtfX4tkR43Hs05gNvnfW
hviNS+ZmJdUTnFubGhfdTYmo4MQ8yAyTSpQw9448OITy+RdWjWsZm2Ec+CITNBAsg887gnhRuExj
uOc14NvvlPHhrDf5FxWNTh87dvE/D8gNh7U8A9pVkix+B47Md6dR/j+lj/MzJXqL8szLzvWMyIV5
4yn2Fv3TGwDrCb0v4w+PoT5WDltIQmh2mFmpKJ6Kx4EJ1v07gVT01pCeZ71xLh7XZY22xJ1ykCGi
IFh3p7Ct6UKNfQiVXET3wipIXCAPUxvJ87Oio9DTYDL/tfSTCKPs3LTXn7huLbp7ADDZvgPERUcW
Mv4DpqRo8rvXOWoURSpNUc78KVi3cub/SL6gTUpEh/ne0hCmKr/eB5csahcIhO9edQiNeenlOoUc
ADRYHw4cW3MqbeT3CfwaYM0UQWVo2O8qx070QzFoJe3sLGGPDYbuap73ggFhBfQjdez2vLfixuI8
+TTgkBVNl7QMRH5nkK0cyv7Vl1GKDsMOFK7KHrYu73gSTt/1MJjktYlXvIrAOo+voYXeAaeX7jDX
6UTPXbDs/cZsZuJesBu8wja00xmglz1bAOOXALcFO68oLeOKszNiHcsLeJCS2myhfxy5L/xPUugC
8tdpNjVSqYYsc0S6HZmABpfUkPCegHGlWVzp8F9IKOnt/bboBjtojh3NEk2NIwupZG6oTfbLRFp0
rekTQhAwMhe1NRdJwc4/mDnoXWJkk0gmw17gqlLqOsGgyQ2odDQxdL3344nE1mMS461MmIsW8d/e
ZQ1NlX5IgXBkWPSXR1/UYRYj4IBJNhuEO/Lv8r8eAAm5TBiqCmU4fkWFDgV2A+V5Uzntc9kRuAYE
w62M62N+Ci6x4ud/yJB7fgQII1fGcCWvFWTG7mkRpvgDKoBduluLWpMg5HHdPv1k2yY17eVRPO6Z
q8xFpqCpw8ltNsIrSCnfGDnqLGY0Ukfkvn1mQTYwneB+4ppuX0j7/PQM7XbzAeazO4XpzawASp4F
bjz/ri60RosF8Z9cWxKgOp8SRsCSPEfRLeuEMa+6yIU1BZmOZg92zkDlhfSkFObTKrWLDmYRlsBi
ZA4GWPgMIBc6t1l3tiqsvaSaaOsgzQ4pNTgaPURLWFQuhqxtaROGmAzpdkLkoK2fJiFhblge7wvA
kJ48nHEHKI76jq3NGNQ2ov8gIov8LFIBGRJUUL3u8sLRQyUvQDwQELGnzPiVaKMEyV+ovdxv+2rU
jhcvq1DxLH5lGUJ0HouIbE8PeJAqD0eaje37125WOzohlhkAzYi2gT0kny5jrGVq3QNbXu0N3CEG
Ly+WrDOkfWzXVMP0pRP4CL0ZbZnLY1oqohBFmnm5tuBUYdGkMwBV/CJKXFynXt8aDejjPki5V636
hu/Mk25uwhM/NPswoEExiOCZDTcdTrf1KnyawS3x9MkyDMGKzLPLo1ImFcQDaBzP7CEbC+zKivTg
12KUVwdRorVXAPLiaDKHa/WeeRIbmULF3cpcbb1Qa0Bf9vPRBKuJqnYpWpp/uhJFDKoAYbGHMJ1h
g3hVVgvaJLKkV1KRJr2hXnu3j+96t0eMxsgwdNJYbC6/VfuVrvS3DCAWpPMWnbzs55QQ5Cy6fQag
KrkztF4wixSNeGJxjgSKE0RhwBQQ2TX9FTa5lfTlV5OSpJEuo4akiL9dm6WnZqRFtsU7ykg+fzm3
/Uk53KtGNQi1mI4IvtdCUmK9h42BGhbAFtNaIFgxlAZyfq109pIJdtz0rit3+XacArxrp7gRWGVn
V/9P130I5/yPx4rw246SkirhGgLScG7m/FyNbybbusHKXdZSxA0ZPqtMfbPfxZcMl3zraV7synaZ
kUynWcT2HlND7qUEyfaKwD7yHyzgIZImu2+TduSharR4DqD2uJRJvIHsQSoxP/9b05LSQZn55Kyp
74atCI7c11wO/RwofrYyiftYal3gIOyab8t8aJvDuNtQwFkFZ1qykqV0DWKJRpeuEkBitS3rCLLA
5gVodzdNnO/mNLT4FHG+IvgyHK5MVwZqLP1FRmkvGcgJ7jengZn2USm8iHs999HeGPFxKzUO8Xl7
+orKe5AN46hVIkkYJY58ZBjhY+NwtTcM2aN8O2B5aau/9pG4MYgC0I+X05EnZK7nwK9L3xsJc+zj
iHMsqs/laiNBJPkJtVkL1ZlOAQyulcPFUCqp2vNLPFw4125OF2i4/l7MSis5M5mwhtf7CkgUT7VQ
KH8EwKUfIQY8S7Wg+24052ey+WIWmzn3Fj+Rh6Y4ZhaXJ5GlYXRO+SzDuLf5Q5x4cNqERkSpnWLP
wCF/zZZA54tn+IwF7lrlwEiaEu/wwVkQnVRBcM68cuK3/2CX/TX+93+U12YyrBhnIoRhwkYZBIO4
2UJX8i+EYJkfBD5K0H2RFtczkE/pL873LtoTPqtrgMtt5pjfnw5Zjuz9DvhDWWi0xiA+/JWStRat
zhL9Wn+Ec9DSFK9+ZMQri6R4PSANI66IZRwJOAsUwGh3doLlHcFlOykgtoTLPVkLjbmt3/w2a+vH
Uge7URjUYG62wQliIpiZatFCrbGJL4ugsbqTjC4WF4ZzqEC9fo9DYX/ozVSkk4h7usdvPiTWvK/k
9gDnYp6gj+THogRcfQWE/UpSPQTFdmXM9o0PaullgsOJ7al/DV2Xj8J781wH2uFbSu9llCzz239j
UrtxyhH9zktgAnAAc2UbekXXebzdfQAqv9PJqYlP9dj4m2cIfhUPikTy24BXFkcHPwFk+80s8I96
uh81Uf4YqEwMkufmJZoKXeGul3FZAuM4GTAR980XjVm4dYHwuF2vagA4eSJPJG+HVHHtCaOyS+ky
1DF7v3dQvzujj8dXsuBBqAw6KUSEG+sGKbeuPSNDbP5yn6LheEQrGMXwtFrucIKL63tM9g4cgk/0
TFZuIPSWgcjHhO8084liGsBSvLvN5pHMN4yQYAU9J5JOFc3grkjTtX2N2BBVotzDwGgMfH/+96mp
6lQZiX2VTXpiaBjge8MaMtjaJdeMV7t9OlTWnC50u0tKwuG3tphtOQuNwPKLNohZxR0mK0jcnUFy
9WbFYpXRLZ/Wk/ELxOXe24YPlKwCxVGk+dpo2GabZhyHEpZVtGZTWY5x5G9x0VxAA4OqyCXdwqlF
920b6XshKJCY22yMZd4u0JbD6n8+j39/hLhBHyV588aJAD4UMmuvk/umYRaHshuDHsQJmwApUlrC
S2pgPpBl79fKEyN8OxrpTrWTLS3nDvmuVLJGYB6y7THjBOADSYfTMat1aHRvrEuUbDEuTuifQTOd
6FZPRb51ryre4VvEbXnI+nsz4b6h7eeDFlQVnm7eg7t996r9CwyvFA1axHgE4nHCm4iPmSX76ap1
uXjUF3v6/5eGP8QFiIbeeCghf+a9YCR2PH9yXxXRuhir63cg4GAYgJZcUFEFr3eyuXDLF3SLYsS5
Hf3XZeQ7aWVFcrSvX/ZYP1wiZHrJ3vQHifZIsYqTDAIFKFT+UwxHoqNpgme9WkolFr4X+oAoYUHA
eyMMDaIc+6PH8G4vAz4snPGZDwLAOVW5/h2PXBZMH28MOV8Gv+7lUIytyr94oMwzrbMpd5m6MzVt
Se4O0shzyq6j/yGjbMKH5VNdO8OB+MUgf/V2TdsgOWeT6mq1DfUOJgBjLkhsZCuS3CoXdM/iJY3r
5+u3mFSui9gg7N+QBYYxT5ShPinWK+cQInRpxUEWPCNiVFUSt7kCXGnhyAUfok8F1XRyHJW1LhJi
XOKrRDGQFeMV9r3gyoohNFdZpzXPueRly8vNzSzvnVV3KklynxnZ5scoV29cnC1VGOto5TmTGJId
J2VETkOPkN9lqiy5SUaURpPQuVCJAAg/XsfO3m89EM6W+96d2suE6PaF3pMZ3IYXvp/IKIu9negU
KV3Dwx+sMAz7zvrvq1McNNNsDHRcboxyRthjZ1vmYFdARRHIPNew2Vfg28emF7uTh9hYsJXudSVe
J0jdQ+c6nmKfdguLQGeB+Cd71/YZzXSBvrWWMEjfGF7WdiyEvnmy9Sjn1jGPEfyd8KK0P7RmMpnH
t/lXzoQJsrMd28clAo32YpRGgHS4d1/7MRdlh9qbsHQlbdPbazUhcU8CPHz6Ah5X5I2g3dzeuG+g
YOBKYdYbwuz2HbbGt4SyDQ66k+TdBapDf9Mp22HjoDJLLxGSO/TOHsgg0iKYd3HChL6U2MlOB0U4
4uHEUPc5J4cvtyzHB6sPXX6yebF/s0GGT8Nl3RC/ExQ9ZgD7veb8VFJ0rlZY34Tts5oly2MndlK5
YZ4VeRM6jObNGDsrWW0zoOTq8mr3PgaOkrxln8ZTBdQrxphHnPJpCfyU/t5zEim2iwzH+uTzYtbf
LzaJeLmlr4PJBMMs/cU9EaOZu+3Vm4i+n1tO48Oo0Aov3HSuFcCBi+WgQc90s6fsUvZggKnGZ1mu
nZ78ahpeGooPOgHBaBbyH2pM1g/K0QfSaXHfAB1Sr5EneOLlsTlX0xrrkSrOdAN/2lc+MLaVjUyC
CCTAdkCGbKb7zWk9jgliwF2r4ILrLLqKcc4d/rQIK/rq+JBGmKPnug5u6B1pZv5cqBlOOJ61goM5
TrwZBSdgU1VWtPtCmKw+mUQ9W09AFgck4WCxv46e+EdFFRJH6oBugAYD8VG/n0l53fzMoBBOCg1O
IfEN+KPNk109rIldfh+X50zk6xrjyjeVhfuouz3rv4t7ym7Osnr6UQEYD+k+dr/v1VESWX1+KUd5
pYX4DmhPOi7ZjxxxR7EY3UkTzOdB5Y0HTXzhpeg/v/nq2V/Zkgl4J11rpnauxgytASk4KTXHD2NK
JOOyo5mM1Rhg8cnh2AEP65VBHRFy+qeumBrbwlq1g0ggnWNypxrXdDy/NHwpmaamy4v1m7CBmKe4
lvP0Mc4LKwFYtlojBSx9Y+qdjMquXZB7YHGlrX+XAJbd7pqMuwqbz4Jr7U2+ZRgYBOLrY1F3GGhH
KjpkfFs3V/KQm2sNcKA4eEdyWBKzljw4TI4wRfLXbuAs/Gu94cqDegUOR6+ctjj3i83G4pNmvCmK
VJmRwkPR6D4efXz5ufIBjlrnk1dSMaXYnl/7NFCsn6zrVbNvDt/PNduUAEWmNTliV5CF++jN3Bqu
qUsSgH5lb4YStWRAxpR1dCw+tjlH6c11bHh6w1XLreygadR/m3egu34HsVMGfKKriNank80ITqmO
da3fxWHc75vFEVTbU5XxU4kAbHINjWAgMptcqE8Z/3Cy5pjW3RkORI4uypsDiZrktd1iJGQgNmBI
0Yf32V1f9hpeOfM0Hbj1Rc09FwoOJC5vxF4lLP6aIFfGgU2WvsdDk3CoJy1nPbS+aJi5VAlquyjN
+liWWU74RPq9dd39cEhxThSgx6BnWvCUeGdIBGpuWfiybdEVTkUx0yDh9ZFxbxaH9GIeZeXmkhSf
tvElDB+0ZLVZe9283qqQYi2wq7AiQIxl/mQf4AKT24D0G2jZG/6Ae60YpvhaA8bJonQ+CIpW+HBQ
OGsjWg2Vdc4qug1WWt9HBKdEI4OyXvZisW3GeVz622C7tGspqUC3y6Fj4Ag8ye0tuicuz+8R3TCv
fWXS2gkf7yoFxC+M4yGdL7xWIP+FeNYE+6TVlxNZ9CNLhPT8Y+9zaslPe7FL1uknXUC+f2YipqES
4MZf2BLLnHq6V+nhqMPAC0RAlqGj/kEwFFSyZK4wVwuNoBcp0rFcw+HncWWyicoLX/qoPJarpIqL
Az63VatesJpWv1CT9p4ct0a9cVOkCYKsS7DrP76eNEQ9vq3DdihmqfGiO03MUl1Ji4zBLg4m9FCB
r+9wznHZFm/o4L12pND0HWoKlhpmthBBJw4rp3ytQPAh5WUHylrQ2HD37v/5AX0wsIvUz+pUnf0x
xJcflGC6RS2Tx1CcZyyBg0FSjW0Vv4ADKuXLuv+OkTG3Db4xhr3U+0cdiSaENominJ0pJSDFZ/IR
+0L96gB9y7QdGICScRpHIq6Jxr2PcZmxStrnNMezM1d52unMNxNCBXx0UUfJtt6OpTVvg/pde/Y5
pVGtlSmZ02NXjz7dvZ/GcN0hyTNNqkH0zlNgWunnLm/F/m/dRCm05F3XgSDlPiKehoBZN81dJyTk
u3ukk5LltlSXwPodid+gS7zNNZ9EuXgO6szKYxo3ZSIEqCrTaSGyH6GlLJgS/SmL178aOCMKtjdi
B+yPY0AcOiZhZMNlZalByt4e2btmBSWXmBsVcgwBF4HXlMv9y9d4vTSjJ+pb2Skb+RgQiZmYY2zX
TACQH9fmXoH394SCQYeRYRUwFA3CP2F2y+6AMRG/67lx22HtcbL2QFex8GdVghk3vupPEc4yL/Fj
Z1PTsWyg/xrqTUJISCP1HRjruafzQBDJxH6n1as5TPxZNddQesV3pLCMXgEsejy0E7JlIS0j3op2
oG2VFZzCOazkYafI5xuUk6OewXLdjH2HcmFN1/jKyUuNLSqZ+GTXapxsYPC/OgcfbWKueye28d6T
7/UwHNHbbGCUfm9axcJFxdfH7D9hwRbprLeMeIjAvyJ6l2CaVGfbf4wbHpwAEhLGN0+vI3qHEhgT
czgc2WzeFeSJqGpyaCI7dZ1Y1IGgrF4gEbXUgDaYiM0pXTXslf0ho7trG4j+9SAyiaUsCVd3Gnqs
34NZJL9gegZnvz+UAKFkqwFT3M1eVB/zMWU+vRNKTrgaE57NyxSOI2xvgNH89bLTH0OnBH82a2U8
+zTg+RfNP8CPJ3FkGUYgofvnGsi7bI5BgUGJTy0Y7SPaZw74oWDUKboV5pZmnr9KgrPfce4xwD+X
Bp75sQsPXvaJi/Lm+mZkbOtep7yCVCqko6qYihVE0yCUgrk9MvxZqfC8e6UEZIr9x8e7jRZZeR+r
8C0JrmNLlrfmxUPX+vmADGQLaCBK0V4Y9EDmP1EomL6X4pWIZz5NV7ar9hGuPKcsyC9YPm/k8vcP
t+lPCtrtGr0iyrJX/ecfEuCVm9f6Iq4P8++4RbtBDS4HdjPrfilD7qgTmtMWq7vtPnErKd4bwonF
sADg76HozQxGHdW4/CaSkoaEVH6LX+3bpSjj5QP3T8FCSqVSDQEQijjXzxirBVnBEnck08eB3QCP
rDHdZgh+XTbo1g5kmg2oXhHtFRvTYHRCttZnGp/YHs6x9iWC1fA2RReKL81WH9ZQXvAzmWsR396u
KN9yP88uc5nhefO3knuSX5dLEqZeyWMy2YLql7zyIC9cc/nvFJblyGlbgY0wnJzXjnN+0CUZ3i0s
aACLKpl/YK+HlFrKOL65Atm7nwCeJdpB92hz4aWZCOgPelnnwghs8tu/iQBNeR2CKzhCQvGADsL5
QThwmANhoEZR7Cel0NDUflhOkBEaNpc8hTIaQHNIRic2hsKzUfk01cYuMfgk5H3j6QcP5RkOtTTR
4e03mtrB7mfBOrwCDYVPZEV/JSl8QDnQDzfi4+w94lmBSBtGBV/T5pg/U0TP7saU3R6TpNC5H8O1
pyRTVVa/RkB3to3Cxl035tc1fIqPUWyS84TAytz7AfkJyWrb7KTPKwYqBWMpg4K6Woeeb0tU9ufE
4d4+A/Z7U3NG/iSdCZBFSooG1pNZAEEjd79XNPaIJ+08b/mCrHhoGIbCYKEWGUel9bSw5/nHawO8
e0/UPLWJJ9oueYfvST4Uxde9ZI6HflEgR3JMBFKBuf0voSvRKSOqKYLIOo2ax/Kl6u821ZxGsst0
VeAGEL9jCIhBvi73bM6BhvDfrs1oRR7NpU0HefVGdzxUtPXhnj0xAazQ0/dkirpMwd1/tL5AxHXE
78qy9Wsuyz8v7zIMUyl276PombqTAcVKvFqDmqqsqyPlSnmhevsmqH9SmIeWLZcWLSQ5OJIruJNc
vR5MF1lADpNRe22kWt+RWjvP3nzP+x7rkvky0rv3o3sdAr5+iZuku9N2aamNkCpZ2yM2bciwn6Zd
5DtTNi1Sz2PY9sftwgzUe+mRlVNbzwAr1Leo8d/Nv8gBxX5lcB6xBa/UaPqs8u49Jms6685ZTvnE
tPkirfVnP0yY4jPAde7S+dBN6HGBg9tjJGen/oQYt7g9y6fAO1jgjmN3GgIvh0RjkzQcasTSQqpW
iFaY4j6ev8XscRYEBdXSe0Lm+RzZHWjGdrLj8T8cNNnRBTlsK948GMNrXA9xS4CJrE4PgiSG02yu
gC8JTmbiVyoq3XiRX4gOo88GwFoN1M6eMQ96Ncajvbd3CMfqOaDD4CycFeVzCTIHsRKXo7t1yl/d
gZm8KQQMrLPMrw4HzOZSjsrF/9nnhDHrmkktJIDZKX8U/oHu39or8uYOovtjNiISa797CuBYJD4V
GBSeqCOqCHv9LgW+8X4PSfK4plcmeY/OY3ekIIhWa+3FAE/JkYw4SToWR16OHcJ0nQIrU1CQDqYC
rPR/Qb12AR7s1njq401lBiGjm5kNSkpbK66wraHU88yERbCTFAVajrPG30l5erQvJp5LBi2zjW8n
k8bRdn2sScgncR7JphVnjZOpyyiqUTPBMnC7o8fI8GDLst+CVsllKF33+FjDbIrXmW46OgNuPYL3
lUpkp77DlEe6eUDE1D25NVVo45O5MpTmLELP9bJk10+FUCMEsTMFYIDezhM2i6Uf8gtchkryyBz8
5uxpt7hgLbTGM+JluBbGoUBtzjkBLWcM0HLXgzGgzka+QqD/BYtdt3pYOgE48qdhuTCZJRezUd/B
Lw/zOuGrPmJCSdWZYC/uDxxxo+RwOafADEXOIH+LMb4tMJNE1bf+noXZ1Cim4MX6RkvTh+Ou0YZi
F64dW1Xg5opKB1fiH/LEDXqseQGdzZewoy0KGMCzKqRK/qY7ubE7/6jEtIfE1dxO+amr+UpI/wBN
J9X5dyvQTL2puSLO7ZcsmG3fCRUbAUXGnuc6QcfRSZImMRbZ1xTrQZqo89iL+orXpXg9ftPccI1G
zoKD5x5G5Y2CE3hD+KKTM8+vxEgIxG8tKgoT/Zr/4nt9eHKxQL/5Ci9UKKiVoetemcrwSMfR6t9v
se3b6mfWcgc1wBjtMk8uq7eBSl9Rn/mouglAf+1H4Z/wE29+x/fr7BYhpMfHWGa45YMZr0/U8DjE
foHK1n+3L64oZokLfMwL5HOBAf94UeHmdlpbiLn18btHD2BpqpTu1CyW0Ga0ArkJQDNMB7gidHYe
9ycEX6upSOHDnR2BO4yvCWXh8ZVKzoQDzQpksqy3gHYupN/B4O8v6iqpqxQkUTqv0K1yyDE59yIV
p0B2jHrgsfon9qHnJYOvemFGQyirRxXz4YOaitIenE4SpFwL4ojBgos3llZbXsMAXGfU7mp+4mRf
UuIshijYW2Vz6EjjwtLLeX/X2KyAae0Yw3quL2dkdN8Zzdef9JA1+qYMgxZPfNqoDSXHPHFZ6+CC
fdDTKCEUDhdBl859ATnZ/XnT5IEAcB/hR61B90EyDB5X00H2W7VB8DagHM/KbgYK3WU30SaUTTn3
e6+Eev3qaGCZgM18YkoNSTtCHDCPm/BnacLxp5HJS/hcL5fEFAvCLL3O/Ie4kZLwHhthwXLCG+Qt
e2zpOtLXD361OIibtrfXcXuh6m9EwjJ5z1rMrA/qWAg3IbBkdyC90ImpuFW26aCnes/IvCWTl8o3
0vI+ECKkMr8fJ84tJSJw+51i0TA2gChO0x9IHmltiTEcBBVMz/v3aCRLzxXOJFj4wWY+7UbLvWdq
84Cf0+TJCLZqGAksHyq729FhvbP7w3MhWtWNk/SfHmt+TJCsm+Txk9ZvCj3YgfBAWplsGhbark35
1e/V5IMuM3JrthUWQmAO7TE5RrrynfICZdCz0YMswuss+XbSRiEjkIOSnB5JEjh/+1Uu8Pf36/X9
SEPo6Mp4qM+Q7+p+G9PkLp/h66gHt473xvY+QIzLd1JJbzcvFsLKwBG13rK2YTPDd65tuTe1rZID
j7kdA0tyVApA+wDIDNxpNrHhG/kUkAj/g9fXp9mfY0XNQbW3fC3Qurq+YgjRmXjwALBfLo4UBpLI
M2mW2MMWnJpp0hXZ/VRVe0P1VaNhY+LI2PpRZxG19n8Sf2v8UzdqHK9GYdDTvw7fcwVP6FoCTtVb
kCoRp4fkmM+A+yUJxhgzjiAlY3FzeIjxzyaThBKIe7PL1cNIhXAhizBYdu0RxSAKHHR0UNS9fTfd
Z5z+C1QBUNh8FnOmhb6fNBQpgs+IQsHJHh+Lah1nfzFJNv89+Vvsk+082miMOfr3+vpkni34SuTx
xSEmaUB4a4jY0UEnZFbujURE+C9n+QuMj+IVPBWRMolLbUVcN6s3KwZfluTuSBxbyi6k+b6JfDKu
KHKjcbTnfQkVr8S1kOAg/+yI8+SR89wPw96EB0wUfKUoIPJvJQ1Skl9QOfyOr2trg69i3id5mfPs
7zJq2Zdc5reWxvAy4+dJGnYJciaR7EE4lfhBzSCJaK3dCbdxppBlnfzIZa5MJkQ82GiJGO0wBfyh
XlPdBXepSRPUIFkTFCHzoSql+LF4iQAj/HMKvVPfXl04NToIrkxAk7L0Z5Z0QCZf3PjRmKpJjlNX
vt7q8muGkvrbV9aaxl7rvptgU8SIgL39blxxzmo6mqT5GUgeWrg2qNVedeQm1Y3MZoV3q3Kw7gNt
j9DC0+9NNE9W1ZHXVxTQ2XkZ/5mAQqPsf/JZi9qzO4+QOF1A+AbBouGPhz5XJlec7HcLnNianbVc
wKKxcRK3dB7l7+Q2pHDLSpiYHLEDmy1cxKqU6d/GeWACtxmevaVuEI9oMc9r7jBRJd9kPX9latFR
pexhN2qaspzRJ9Jqd1C+euGKV6bo5a65cfoNiz3QJGlI5cUkiZtilxnsGKEx/cZb+aa1IBCHj6mT
XwYk9JcnvGrmVxu+MLG46luaTWkp8sQt1WshdD66rIoZHwzQfkR6UtLYfyLsuPCg4fj/ri94qr7L
0MrepSa9IQsDDcU++I4KcChNy1YBnWgydCwe00vKMj11rwvTQyXqSpf9ghARa5pkgtDoaDTPTcOe
D2rudGNsS37NUIsXZ6vKSrDQVGRQ3oV6/GZ178ZRk9E/VikE8+1DzUDnn/1qxG9R8K7/VQs22Y/D
eYaxqYNjbewHIrVUeqLqwusoXQBdJV5r2B6T/aJe6V6lggytPZ9YNJ5o0z/4kEK8dmfhGbjXRpMk
2PdalzayjN1EvVkNxCErMUzYb5UZGCpG0eduVFTgd8g4TilGk94w6OkNISrJJrvL1/jqGAxqLTP5
/BsuIQCLgyXNfRlwjSlGYnVqv9X3Tee14xiUMU4CAmoe9U1SihCN3Hu/7vXDLSDpHLLUbd7mb8nG
TczFKLNsGmkmccBFNevDB3/wqbrCaI3hJ15ekhV2yznJVCCIcvd5f6iCauCJwk8c9kPKYCL/4stR
WZUd+4liNSeaW7kQEi6Mbhn/YJE+Rc9t8AtRh07lZIaw+uTxvC6kqdI2vw9+5ndITKxrvBrc/7iw
MgiZ9AssqRMYp12l1YjIGyxoTMa1rDNFxwhef3oZKcDyv+S8X99J3sBsrQxd2YNavvqNSDeUTEQG
wtcB0wTCjRmPb3WKgOcc0J70jH9kqJ2g6RcK+8MSgQmrzfmavLK0bDNKcE18X67vJL+aLZUTzvsl
2rR+m4zSI+kT6vALIKBNF10oiTfCRCKHcvQlmfkb/bXlytfGUfmxts2M4WUIyHbymCvL45EYPMj6
cwl2KYVKD9/FZfojCmPuZbmiM3OufHG3GKEZvLzLgQr0Y4g8yrgvixpXEueEkkSs/VufJinTiEa8
eKtbEbXVG+M8u8dmSWMvd/msl424SEu/5CbL10clZO76L8xfT2uV+V3jxCII002/3cJwLi36ZC3a
Tlee67f4U4Swo4eCt9vrsZ0nfWY9dGdqYU/X+5QxFloyRbytV2qCH0nretCNkO+QpakrE2FSTBqj
lV1xfneeSjGvzMGClu+Boi915v6dM0bp9/OuDmGAnw9dZxW2PW2r/kHmGFKh95v3MyGRIIYOi+3M
075QsqIR6I+fMj4C+uX/dnn8xSWjedPdKXb8y/VmdnPvo03SGrWzP7BP1qyiox541hOH2vLc9sXs
wf5vbHqlfH7+J4NTMjb5/+/w3qeQ3JqSJaHBrqmgdeReJSn/STO9JsReWlc7x5QRNf+yeuqX/Usn
SBA6dT/z4Gu12R1xACcZuOxrXruTBn+hApFUstjJi5q/GkPYAunlO+j+1Qt7LiyjwjBVaFQZxb++
e9p1fFdUTzX5BBs1iGTWdmzP+NA/k2SfgYjfqYlzUVjuHfDQtXy0wbdKn2UXQl5/4Gc/BLfnz1+r
9dw/QvNIKG/wglPbobq2Zz/CXnljDfKB3wpW8FbTLD3dJk8AfDFEvMNaXQcMFEAlf6GK98Wm7yEd
P0rRBy5fgfyjHxVNKRHWG/F9ax7NBxJlpeyBGU/YPCuS+iVRiV+u8dtdgN38jiZajEhT7gKLXy4x
e5c9MLUszUU0WG42utDBl+J5ki3Mt0tAVmirbtBBttnWLLvW2chmRLHQpxQ9k4BcAdsra9gOOT/J
S/JCShrh+WVYTKAwkaVk7W7W14yT0CIGgWv/Je4Ovm6lskMvpIN5HmyEr9aROxvgxvMQUiu8CfNn
H+BrQlKjUUdnclGP+qdNNwKK39bqjXARXWVxW3q8vya37Ce/4DgzvwDyaxOsA15IeFNIxuzxxebn
bQ0UmuPRXEpZhXCYoozR6cCkwBTwka0KUc4c8EeLFqVP3D5qtrNXGtdTrBYsJg7YxTWX5SoUKqQ7
alHgq4iLhvbx4KxVSfXOjOLVjTfRj9wYa62JaImRA5aNvAVVc6JvRyNAmnFOzPMZbMbSGsde5ub6
b6znGeU7SGIa/azifdqxs83xn1r88ouxEjfoK2Ot4G/YiI0VINjDQnpWi4cG8oPrz/WULa4gWSiL
qZCs7R7I/z7hVuHdflZB0XQy/3I5UHhb+2KGdjIdeoInKga3JbB8E4HODORSpnbnmeKqK8Pb5vLE
cOnam7JqMdpEOETmc4/64KPHpV0eS9E0mQth+sRKMqnSQx6t6xCqPp0yGhegutWJkC9XwNZuogxL
MHo6atPEwQGbfl3+zG2WFlNK7clmds5R+Ayf5Jy6TKnEHcQgTYlWqdv0aRN4EKgweeLYSlRIBcN/
PzeHFERhlX2C5IDeZ+tlHzPLwt+oAjtZ/6LCSyBpsuEu8y6ruiXqh3vL4MsgxgjE2ldhzM6v7Kwb
U1/ZeBP5qfyVEz3OTn1wNA2DcMZJADD6z4PQU4aFJ+w+mPEq6lyq5xY4ztzBLU97V3pCzXKfFyRg
BOM95cBT0oj6tTxOGiknFvkxufgUs602GbcJ39aTadWRUnweb9MgbQ9xtpnLijaqIWRClrhBTimW
UWmN+eOOQ6UJmQ/2c2axpo334utcxm1hF0XjwnE+kKDG8wLN+RCR5G4vtbxZvXSNmoCrVFXKIhJP
EvdmgZ6mmRQcOhkm0ArZ0bqRy7KrjZofQNTV2eMohaUBzI5OBsskPtS2Fw6poXgk9UX1NDHJ/Ey8
v1scq1WDtqYHknlEA3S1KwjTfkmJ5j70VvnPtcYNl7Dji+rrKuHlUdQr+fPvQzqifnd0KfY3lvUl
PTe9oCXvstmUq4QHgi9kn8flW5RD/HI1c3GiXkjy5TPuV55ocDu2X+1vTRqN8FXgD+Dn8Xq8uHEK
paO1xDWZ91GypAc3KK+1Sjnpw1Y0sYO0cXbeDc9vKqCmc1BdWt+pzr3H8hpB+wVz+Mdzx7a5rZbI
UQ1IZfq1DA+/9aQ69ZsYHfrbTUcARNiGSOMhp9snnH5398mPmYJ19KW5WsZqlKfxHLf6XdQP8WR2
2+Xbpz1I+WhfGZDR+RqHMh1X3xDR5FXTy71TqPjU+e/t4oK1ZAmKl0vzheFm/ZrLInkKLEwhQEpl
gSzVlRNLHi9NObbNxrebJbm3Z+90Ka4Sxi/Rc2PKTaQ/7TrczVN6k6vNe+REBeqlNkkT9ZP/5ILk
aWzxyIXmcrz3pzH7Nn2+u2bmULH9nlbZDKUcmWemLsnc2Q8s/Dc5zHkdgmqlHSe7RiIzOIS9Qzxn
EyqPiI4DKWuEul1+tEb0TzEGUdn5i/TzEpOmrNwdWunOiyju8jWuWPUjEYC4G6oiu1vjZ3I93vIq
w6ZYI/9kEC1RWikBQLrIPfiCgVSJLfpjBSYrQAZxA8m0n2xZ0Qo8K0/L4CMOQ97sB560Px+E7DLY
B+nbPXohQkFor2TRP/cgf3H3Z5u7bituhW4mo9wEqBMvrGRYRweeIfLVssUDo6jMtSw2ZDwVItY2
VFg8y7L79ICallHmqQ7ajRA91LGewY3zAxKZUtjyOdmn3IOiNeB0oz5HATLybSlApsG61AiDCBGw
HiPcWNNUB+Srsklnb/xc5hAECyoI0PJxqXa3CXCvF+Cns1zp3bz6YGH8X0QIBLTPzZ44Xi0uyTNB
LuoyTSW4gvV6zPBDJcO5jXFOVMXjiiqGej3V0VxRRcmH/s7gILrowLjTgOFec3L2Q6jFUN/vgOo6
Iq3FFjwtUbVS4RVGmngkE0bUPhVPqNxSo6eg9unUhhhQq6wlCCqDuPqXrmb9aOKG68TA37zQPpC8
826lCtfs9V0yIYsD6oIuI+r1P9XywGEgfzKHoYs7tSqj0u1NylRjrbsRLiaIfE/F8iXqnZIA9jAV
Mom1elRGc1R/DyvYAOvTRY7zkKf4PUWJxD7F1l+8DOdk6ArYwSJw3WP0GrubW6SJJtzaLvH/hlXF
Z58vvqG+YX6byEcjydI8DgNnrIVFbA6hLJAzA5McSZhaRgBGeSVMPQOhPCt9F71RPvuI5rt9e1BA
2CFoGD/FZI2sa9SNuj2JH3yKqWKPL+eqoCl3wpYyWmv4vOQvXMnpIyifBNFxaRsblplcwzpF4uxX
/M9+JT9drdhA/FfrAP1bg/NvuWwCR/fKfS5pNsMQcicuofSBTG3VAEIczeyAIh75gZUtJaXKcjMw
LgssV9BTUDrP2RB1GS0S6KlYPa8j5GRvmnN4/p5j9u0Z2iZdckY9cBYM0uBdQqcC+2K6mnJfeKRF
SGoV0lXjg8V3ZJODp4dDn8x2VAzzlXyEL3ZWXaW0MgEKGZ/2sXZm9ojfRErRXpAf0AtgrbK3mz/y
i02AOt/WVounm0jPXjOonSnGUdXnr4zSh4BstpbWszhb6JHJYhs+Phpx+RbRC83408EBibqJupQk
ftNEJvGtxYTDXNfbg+thWvHSb6HhZjlRoYPWpuNaxJH+p7BM9koHLl5P6DQ1S7qLC0/hV88YI82S
kb7pFAluyRUkdMDJWyizjGUpdYcLcf6gtR7ZRDwEb5LU1yw5M4KEFhcmUV+Hb1q8kV/OU7fPidjB
hAiRVVxoYkqEw7vrAY+0QXevwhu/KFPQpHZ2EcwQlDdJ9XHVfit0XSc/UAeWhYwgM0fHeReRg0bF
zYeAcbVs/2Nzqhp6sEY39h2tiLnBsfbEBt3gHgY3HRJgjKwfsvRZaYn5hoPZsZAGsNrCjhN4XjTu
JYbZ5jbDyfAqiBdn+Pg+yBr3okf6UhdM1suVqOsPqD8byCJ3IU5Cxd7P33jaDSBqw/oerSjNH6jo
o3s+Gd2Ha72DiUuk+LCpRBGCAnEYpG7bVI3GdINe9JlxU0tA2aKeFqh+V9VKORijQK3tFF5PY5b3
8A0nPlKB2nJoCymHYMXzE+CxbvVaQK2M1Ii5zmMO4ojVO3MhDQvaBbyoUdIv5zPTlUYw9pURaybt
A2XhT45ofOzjreVWwKOF61OPQa1zDbY/xdBrzwsMod32RLxWis96P7TvTulrmS8RvJPL4bVRflaf
c4tiDV0tfz4bJXmKJBhZEjVgvOtyd0jBof6+CStFo0xEZQUvT1yp9spV2Vck+5G31DXZHXjgfsIp
U11ZBQ7M3wFUHh6rFZQPjWqk78F7lkyyCfVC+o9Zjn5/BiAiEdmfVRxHV8Fe7NHm/qrBn1VSd+g8
a3UVqGs9znkgt9i7fQF6rFhD7j1FNOv4p5rTdSt5cLLtoi+lbSfz5vFGyV/1hkxhFMURF0z2pIhQ
+5J8Wjq7K735RrygG1gGthKNpDvlJDY1fL+HfuPWOc8lKuY5d7WA9jRIwC/8iQ+/37QXec8fPaUv
MDYwXEZiiRjlL97AONtTmu9HG4xwXS+mOmfYJtEAJiowyGg1m9N3Lg1JVPNdGR0nnUsfLaykw7I8
CsZ6XQpGIEx3dG8ERAvJDYyoWYzK6IYLeO8pxnTUGgvKM3gd7aWN6kiAYYmgagfbEELQgLxg4BP/
SiLL11D+K40PWqlpi+dqevGAf8OmNLsRIWWDhkKPy3Cph+B22mNmI9LqvObGyiuAf6ZfDBOprTgC
Ttlqp/M8pb2J8invoJKXrBolt6kSmXry+Ml7ymrOK1DNRPfvQrhR+aP4Dsv+X89kiQIDhPZTavhZ
z8hrWrh9uF1qDFCGHmXBHbIJ84G2Zr4B9mxXRUSWbj0OnrWK1otnTFwPjtzrAmPABhZ2eFaCrjji
pk9Wh74kdyJqJSlXAaeYvAjR7IiL3i6Lfzr1fl5btHQ02Mdo/cvN0Sd5yyxraFOW8jrz8oGTA6Z8
yvGMK55RS7Up5mRuZwQuohqL0++buryS2rRXrONg/w6YyUcQRtIe19SAkfaIuiyqvt+288OXICD/
Y5OkDsLzdCrk6WGmDh1/NJRGV/IR8MC7nCrY2umFJ5+H1+unCAhxFgRHZM+Y0Ikpm4TmS67RcCf+
eBWV0eB7sNUiYEhcpS4Cde2HJTz3fYITFZ9w6whtE286/Ai6Dil867Qw/8HRc7lXETWCEblgfNki
BMxRcDJV7F1xU+dbo7JB32gDT2SNK5c1DE+aEAc/tXaGgN9CrElVYyToDbTFAVcSt6B/s/n4F0Ml
Lx80drm1aQ2KNu+Iwm7td3kaWRIN/0cl7Eo6+KFQc7vdBq3ebFCSY8yw9+xheeDIMVsuCBIuBwKw
rAdeiApcsJHtrC2AkXl6eIKbAnB/ZBRC4Ezz+R9MTOei+iAx1+yZUXHljtGE3q9AsLH+i18KYCpF
GGPMU9sA8vkiAbMS4VAoULrLAK9+5NbUsZ5UkHaw8/fV00grNZ6kTKu12oQLaPmPUTJry/+1SsOG
6+E/4bIl1rCTr6U+mFZ3hNCkPF2BwPjNeAvrVEq18BTpzLRoRWghjfx3wQsZCuLqBiofwbx3DoDG
wPxTfeU6riTUzX2BDLW14ePE/WI7F9uug8MP9W4tk+ptufogBUKrH56gkrE89ih52tKfY/+KFJXL
S3maD1T1xXQQkxiJe0E31yRQYD2D0ugYNuqcSrvIhvIWWQ7RbYpRxfiJ5bsDvIj81apd3j2RcGGW
7ceFb591rhHb/OBJIq0waPUhIoMgna8Q6QTYiP/+WQybXIeCd0K4o10vu3yYbnl3JCvzMf/s8IXZ
HgtnfkKzbax5J18yT0eEnq827GZC34jangayBw2Vrv8BZ1lT5JjIV514cE+xWH/UICp2IgaJHV85
s7Z2FOSKpVhn2QUzPr+HE2kXzCsylmNqPmg7vuBwqwv73ZaaL6UCdoDzeAxoUV1JAIRHfSOUtTq4
uahFShMY74D9en9FPXgg1lyIJ14BN89tk3cQJFbMn93eHC7M6+tq8MSD1xiMx0JOUtWVLBkM21aO
rrJye/+juKS3KajhFYl9aoNaHme5b8oeH5nBO0rnAVMLQUv6RwY0it9XbrFv1rBdxOvxsy4BzC2A
NS8CTko3hZinPtgDOscMfo2bwyXHs4XfgCYlTsyLTh38VaIFuyXK7fA9p6MBcMFKlRBNUsoVo0rp
zPeaqUjhUlzqoPDRpZvtpNzOGgcC6OO5SXfEeiPRCxzH+TJwCyswa5V8ongGUkE9fZaTCK5xTgJk
rp2PzEu63zLfzKwauSszSDQ9GjnIDX3KcBHrQDFDN7ioWYzTaWp6iie+sHeK4uR5JgZQyj7mVi/v
dE3TKc1k/UywjoJjSAE2hr6nTAjdYkdwUNZ0qevqFN1UBOE5ru9b8V/Ux7/JueSlYncC3lcAkFaR
o3ohGL+H45XWu2+FpLrhil0N2cSab8fAXM8+Fvp/dLlwH6JFRDr9xLRL3bdQO+OVJgd92TcBN9L8
lF0MrIStpjsO7i3aawlQzdXbMEm5fjgsy3J+uDVZFi57F6rO4Yhg/m1k54MqaCiDFE6PzYJUSagV
elhTBQ==
`protect end_protected
