`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xbx7xIwGr9qXZQ31E+UmA9C3h+YfZtr2P8H27IAFCW3y4CBtm8Zjq4slmC66fPki1Wrkbxv5nSOG
c191mj3oAQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cngxHIRmPnvD76UDYC8i1mLoI09H0Rd/jxtVnGmOQjmm0yFs2TZ1DyXI0PTya48QphNacLXxVUWl
4M9FTFPiGI+Gop5X/Y7wffM9Vty7QS1QY7iu6XYVg/WS/DZrSD6glAhLjXl7DWCCyH+LErWR/C3h
mcG0DA3NCT0SpFK5TkE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X3AO1+Or3X1oPf5JAwOFRMc3APjsxbAlM69ln0GDlwTkdzT6TmmF9nm/TICkJc5QMBYjEkDvAvcV
l/uBda6CuCHkSDPUJZLYiy5DLYJe4QtxUqRiMAuDUDPyeAEb992OusP69lvY+w/jwVu/NleXo2st
ICklxkq+4GpQmLO4cAGFFWadUSHJrtuysgXlfbrN0T0Qj98+yn4MSxwajusFVzDnG+lIBKBUlTFX
K5FrPWmoKcVyToz8KhUGOSpxDiekdw9WAmJm+LcMpwRRW/MP8W4wqJXrGQhk7o7smjrBHXxSOilu
GkG6dVnadCpB7ZYudf5iJfN3HHUhGy52Nhdx+Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PHVGkZ0eplvhR/eVfIDv3aQNkNcNXSy6MqtGCVAGrYH/wKDnV0dNBPO8CTFTCD+okrabp6s17DWx
fAHODnyrG0JxGwYvmvDhiq04fa+XVmbSYYnfv4RasttVHGbP7KR6fWqawGabpYMQvrJDKcY6Gomw
/UOWsyM1QyZ+5zQzpfo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YNW/V0DhpbLywMjDrIfltjuD7H/e/cgieSHanRrC9Q09NW1viD6qoupmzQ/u5vHvfz7oC0avz8do
u+vj3Bdy0S2AA/hWGDSEbc7VNZuTb0KtJBLRrHsF9yp0GOPHuRjGv+bj+vZXtWhE+Fu8M8/tUix0
EyHPN2zxZATRcDMXquMegViaV4kvga3EeaGYX/TynTrq2L0t5zpt+TqQrA48t9y9vyNELnEsJyDt
YxIufI4G9hi8oWxLWSfcxVT43jgkpD4L9Qptxnjj0DIpk8TmpKEZa2nmDN3TINPrk6xC+73HrhKf
4AFsXnDZwPfQUHPSJiaPC6tn369OZxrPl7Q08Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
p0oeFt7PwGXPFOVihZOUF+GzngUD+srjWXn3eYn9R+w9JopMdB9FrA+zWpIzpIvK42EahO/Gmotv
T6u90aiEfR/5Ccx1XGQohBoW1f5RPOqbXVIUyNj1PbmytmQ/6oCCv+Gi4/Nsrr5l+Hi81OaLmVLf
k911QG++1CBDyzhH5CCK+6l6+eC2aRMPbJk1Yo7Zpw3ufXXLY9ylWfbob6kLlDaEHo5h3r3nO/k9
XwPUbjvNhiYgKBAMRLu0kqkfREx7IZiUY5IEWoK7y7JvYx81hzCPX8KH6Ko3nmHbIHZnajAmbRSX
jM2LwEjrs6o7yaGW1/gWyxTO8b236Q/UNGlt1wT1K0KYlOP1+upOkwosngDPzV2dEfeNAAPgyRD2
bV8sZvg1FdUvXbspbfkqhQaHO3chPp6EkUCoY2OUbnzG2UHL2oPkWqL9j8mtkXYgMy5l8J7jSWAu
TgXUJ4jgm40OMh+svn2vZu4UAxzr478iqH7op0C7nv7YmSfCsOL0LM3ycwel9WwdVPk7qAN613EZ
PBRg5tZXczp9VnbI/BVzp9BioGOFNoihJ7dbH0kf9GDfpxcUEoqXv3w5xFMYl+2sBVqcLCaohZvM
sKpWEp3klWR7s9eG8Gh5gEFjwSe6m9ARFRUj23dEgVcSbYV+YhOVybY/Qir8nuBxKEz3zAm6u9/G
08HSPT390FScxa7CiuRCib6cSFag1B6rEAbI1PArQN3iC+TxnXMjLk5aZqVg3As4UN0vw0J35cRT
KHnNVqg4iuDd0FAlhaFxgk6dEtMiEfh2Iangz4SsjIA8kCYEkRo1ReDv0fHpKO7meF5TzfK49Yla
3F7PYLQEd8fqUCiZl6SGS3rFtpBCYaifWJCPCGXqXAqCRfutkSnGXFGN3i5yNAXl+usYAkOkam1L
jC7Qc/eaFxA7YKIGG7sdsx/gcgMZ3Y2NO97Hty5OcSEPryJIUPEMiPKhO+HUPAliofSouQRhzYHZ
8Irk8yKimOEslqaPfq6SUNb5jTNJ8Ww4L73LdzD+qNm16kFA97jpRj2LMCAzledNNyS8rnZhuz4R
mSsUUKaMkOe0Vcy+cnKhEGuZCRHcOX0oX8/yElpNGt/odyRLyW+7EbmYbnRro3ZOeGjjWrC4B6od
QqQu70QmItrhm2971AdwNdH2ZVqVlQ9GKUq4B3K1cb4mhkOx4ZXZEYMV8kg+TF2Tni1whhW5Fna3
jqD5B/8nJ/B1O+XgSOAxVfrPIY9o9q8MZqLSqya/CfwlW034UmkkFt3xjmZ6vgHrMtbbQcBCrJcw
EPNOsOEsbcQTgzpwWrvsh3zDRC6ZDF++vKQRi/LQdXdYENj2RP5qv0zBhqzrVfManklsUDMNmFfS
nD8OywIce0Dxf4DR8uhRoRbOELNsWWDfPO/X3KOwcMoGf+1Pb0Ic9fTXnBm1BBDcY0on96s1bn5T
B2TZvtO9upeOECyA1Tf+VI0c9qG/oDI0ADC5AG5d1oLvvAsHNv5wK2ElALS3EzTT1EoqLhhEJIbX
4K2m7wP43Sp2JWWXDycgBIPS/i72KEgli+Hmck7cQTbHj8gKX/1ZgSGrNEMEbmw3ROnv3ViGxpMS
YHk8S2TkJG5GGXmu+nMsKkVtKmg9cHR+WEK+/gK254hocuBD3I5gDmly4Jfe8Kbwx4eGZKbT3SnI
2+DeEfUfZ/swwgZDYAJ0eZ2W/mHf5Sin25303aiNGA3MN30g/OOiFZQTWOh2IhY3syRby+l/p4hS
NH3MHENPYaE1KGTcWyttZbO9JJTre00Cc1Sjgb/Q5K2bTKz3GeWhFRN/oxa+Qz+kia5Z9L17tPoe
e8vdrEax51uBSu5ppXpXXxMNVlsm88U8R+8wPaiwtdnKp1elNCluYfwPSUi00jHY4wNqRjiUCwfQ
leQuS3KwLehlJ2Ymo2LxNxrczVF5/dOUBsWZncD88fQioeTMhDZUZLkO20wQ2q8HCEC5rUyNy96V
JG63/1+Mp24cWaolXRw9jM62wC/LGgUIKNFmjXvuEPhFXg7ImMhJtxd5VmPbEXDbZiNlFu6Z3KU0
0KKJ+xSNzbo1Atbvs3z9JjpMBaZsAAZwv0Rz/DZx8eRYbUvQ8OQJBD4hcdiZSYxr6ZkbbTyreT3o
SDgpCSmAWQwb1kg/fIqphKgPbS+UTsxofQ0gspuV4GmtWlnlKaBzrS5PP2avuDzqDMaiZCt4e3qA
CB1QGSPiRmX04baqzY4L/Lb/SXS6UMMNJTKNPCz/FnSUQFysqrZY1HnY1N5VxSV5CieJfgGCRmmE
0pSr84s7Av48+lzuep6TwPp1j6OMtFMiHUHO2GDktJYiZv2sEcHvo0vJSbv5J+DtRujQpuMku1x2
Fnu9ZGDW/sw08ynVLM1y00vdmEc2NEs8avKdezTUTW2xBxLAKojkxDD8p+7yFvuREXzISd2B+SeU
8+/SAhIdXmX3jrUf9kHxz6PkE7ZOYBHyw18K1BkSP9d8J4ffbbswHMawu1JQmxIDMcJfhXn/k1WK
KTRaP3hIFgoULbNAgo92J1ZWWRlkhqgMRbQ+QBdwuN2HAZgz5DJm+bqHu6CYu0ac+5RH7Z1w8il9
9BQswrenp3kKrV0VdLbCMgvdl4bV4JD+Hkaw8U+9a4A85MtXtSdzvqy/BSl6Qj+V1I3VCjqWIGLJ
5D8sIlmXS4Fb33WwD59m6hZch7P69h+VV3prImGXXA+xzgWMvWB3Z2w/1o8owsICCvqF8oelCL8l
h0o4P1C/bR+sUVn5VK4voCmYfViHc+Dv64p2yiGzS0xPoxISDsnVJZQg9tThPs5CSbZy7D/kQlTk
0uJhyh9ANptb6aJrdvfJ/SvVZYAJkFHozFlav8c8d/Le69l0u8wLKYmslK910ZjUVGIqV2oeMQjG
S5zn/mwYXShRMT93u9tiNMsjhycqXGwaSk2qdJCvhGPwNyS6MBpgr7eH8l3skE3S9RJEFNczEQx7
+kTgaZwxOwNWc7TB/dbgCXqRKUe1nFqWGD9NBc1wneyLOnTSpR5GrRvdVdUodrugFssXbVoMXuyw
QcuEfqfpfEpGZz/5syTPPh5upznxz1NbS2/cfIZ1EwmoxIG8wd+Rj7oPRKV77IT3aY7mFcZLhfA2
piZMq8jKlBmCDkbDfCAD0iNtUWaPHHfPh851LetotCrU+XppTOP77xbnyap1SUldodlwK03mGeF2
Uqty2VAqURSN0twQM5dnpTJKw1oakjTh3r/PZjRl1HFoOZ7bNjQWXQegRMAzROyLr43KESeFam9P
LzwrJ9F2cWNKZbmx4inV69+m8b7/7YH8T04tfEtUjR9uXXftypte7K5r2M2BI+wlltMUQ4ujdNpp
Hw1xvq/0JpUIFpBrcoBNVZeu2Q6g4N4wTmFD5g/Ar+B/2zsFHr1EhddsMqEVkAkuuIk9Y94aFMGm
wZcySvy5kOAwjyYX0kDA90LzR60IUu3cKuIA54SkI7MkQ+M/EP5sUBP277gpBVQgiB/scBtGgluE
pH2I+FAgpH/UBDFexwMO7VfnxWPtF/MDTq4eWMPHldW/g4a+aMYiKAWn9koVpdds++dfcaZjnXOB
tvysFCoNiMNDgLJ5h70DoGCgERg/szF9wKA2r7I0gV9Gq/uvbXJ+ZyA/FQ2YE95HHxtZQ3+6SiM6
WJxiB2MqpiPB+Tm2akLyXDxJNsYRz3c6sYnqvc5wfxTK3MmDBWcC0EPlZoa0LOpu4AdeCb9pIqy+
OiqNZerO6UbHzeR0ScakY9D21g8fQdJmafkzYtjV2Qh71OyEOKLqztDdBiWU6XsWzFrsrWHMaH18
NYRwisufhISg35LKR1RVXf9aRvVVecGZeBowSQJm4kPZYPCm598Cq75R71Mtx3s31UEZO5lS1WQH
7PPUARUU2DvGRTMOjLA+Y1Mjjov2myId8An2n2rAygDWLFt+f3CZJcd+lrbKHXcmjlH88AUpgHHm
V5tJQc1uCra3hTb+GLUEa55itbaBny2qyhHvQGEE0EmlgjKpoOk/i+0CTF45G1cRpAOOIwYgOH5I
D/PKaZ5tjgjQmnb2ewlEply86FvqQPkLM7hzXWB7Pj5WwXgJtVTtXF/KoNmJ7CLamOAmqkwFcVwt
tkiwJFdmL9h8SgQ8mVZcg2Ha5TfPTgST4fvWdcQH4RAbirtNnFFEDAXxd80FZsw2FxO6ocyg8DsW
/BbYwZZ81V3CPGYw+FLo7yc2DY4xPOYXup2wCbL5MF80ojW9L2c9yNJuy2MP1SZGZYY4DEIjD5Tx
pv9+OyF94BqZ85uJQEDjvn2JtACws9+Dhu3P0O/0CJ0tnZtMiIXiZVHx2QQEjSF8FU37DLgVbbdV
fB61zzRaHZSpKQluIXXQ4poNDE1JYpn8K8IMPjrgH498fXGXr9yZ11uVAkAtImJBWq6MmgQNzSsS
kh/evwNC0mpdi3IYA76NaNI5Of/F8bVM7AlEx36fOub2QQFPOOsp0VS/ijXNJzxm9yv1ys8sA9TK
zEk4S66GEyu6zCRw3coYcMQG7kM+OfpRJ07QZZA1318rsxn8J976tMKWe4fZSl+GFlfv+A9V1oXR
dvGZTN6MJmGRM/nhCoSq4xJqRrb3afQA6a3yaZpWeLzJMZnVe+KlK/UNS0YihO4ggWPzr+yh5LiB
3X4Qwsqhjx7SrzUyuDQrDisUczsa/WyL+S3sA/StZ2IAqD1e3v1m9BAJUI08VUm5C+HtEJDv1oWD
AkY0Kwqn35fdV28uTYTN+rq7GvkXBbA4OvwxwtdDyXMW/V3p6/FqqMhKMl0pj+eBbuLn3ClFy/uz
QBJTyHnOhXEstowPGt2hV40IKAKb5jvNPJcOWbkmsBaDx6V/cG3WAXv7XEsuXtXxDUVmnOIiozT0
osws+HMUXNfKf1LdAWyBnVpeWAtSK3GHkdxQwXbm4R7Ec7GwH5BCh/oVDYHsN81rGB6I1zr89sUs
U9OYnRaF2+/pXaZ7YSdXGSkKoQL1Td4VS1OcdPJBn/r542WI2Evo9MDbb/OgHYy9Tp8d/kY63b5m
inQPtHYZVNIh3LGsJ1R0XsndHB7TJKCUSY4rotbFQmgHBIZkZUn8xipaowuyTSrbp8i6RJqLI1+k
u+kNc9WzKjksbiXFuMt7DQZzybtCABUCkKDfgtyguf9vLTeGYye6YfeaqG4TQ1IWKgsPrB9Jebtq
unC0gFFXBG7FECdN06DbyrmK1b+Ewan0XjH1gZ8/fv4yRTeGYk0vVJB9SW9Z0h2uNkYh60+6It0W
Xnlt85N/fvt2ixVTN51Oj64nRTdmc62L1iVHx4ibD+vJIUpxgAu0++027uARXesWHWdbedzAsPUE
N/oniAQHUimfw9gmldL3qj4oTz5hTKuLOIlMKnEP7D7eHYl1QebGK8MAQoSGA7mO7He+0VdROX2+
eXlolHxy1V5AagJIwVMINA+SiL/HjDX8Ot7sUgYD76rggG1DdaNEf7m6OAVA2yWYzKv6ba2gSPNn
Vt4Z6SJ8qchWKl0T6eamtSSArrBM+X8akE7U0kc2wuuZ35KNXPXnGHsd/bL3Yi4eOxGmMHVdHWZs
Fy2MoCnnIRN1FCuXuzunfH5gc+TaVMOONmvX6Ak7owN4EedrJ/koc8A3DDcLXKy9VZHlZxVNN4XQ
yDj6RvDICAsG9Ubg0EjVfn3q+Exd/s3WnSGm0XUCBx30aB0Vb7qDfGbs6ZYbQy3227cYHLdfJlVW
ZIWXDTDg2f7/2e4HdyoqclGNmIlN+GAekPpHzCFdwhDIjwK1htBwhxVX4flKyeE5BPXbQlMTg9Yt
7wXun78xRCkv1VPYWhFCTgvbU7EbfraGJ4ZWEEDQ5NjQRtW6YEpDqkd37RS2qr6l9Ad6C9Abhm3s
M7xv6G5BPplCuC56evxIrrbnGLjjwb2JkPzM/0pm3HgpKR4OZYSPI7cassxH4p7YAICDTBgc/fjs
FZiBSAya7b6bEqCO2cse3Rb9Epi2tFnuenRgFg4GXzbe+AEUTso2/iYqrme4cCCTnM1Z7MAOlQqI
Xhq1hoyYiaLXpJyVRX/oh7gedv73pUCF4uuBEUywXXKB/MHvNQ4hw3S38A54WcMzamIjRe3QKN4N
HhLFAVO4qHd3eqIl/onohMzdO3A5c6a1YVl28rI0G27kBe2pqiQ2idp5FAFhbv+WUUrUEG2qESKG
CydPcOnsKm7GyuMAWz1jyxchO5rb/Gx8IPlFyldit9dfyUacFD5Swkd5r+lI+vrOVRLhAfubcatL
kMBMURRSlqY0AoijrRVC5Ypo8bQHO2q0m0zqoHL+uRJe7FDpjye3aBHbVD34VphPWi1sgAP/BCar
NqES5EmU78FhWSoZdv5y51xSUdu7yMqVp7kNZ1qQnkTd+qO2GohTIuWHr5kGB79IFszRXNQn0XZD
BZ2nT3sGh8rI/aHae1KWikE84pCzwJolblGNlqx7Ig3g10vcwyqv/joMdYo5Tpe0OOwPwOal7yQg
j3/a9Ci//ONrYCRjwhrBp2E5i5F4ID5+6EB+2GmGbda976N2jeF88Ejh2Rs6P3uBdwRw/j4bBCd8
U7bQtB3sLnszRmCEJJXQ6CMCV+LuzXd90/TXBM6F6IyjJxjXwcoZ+dwwWTqxkZXSOM5aWXjp0oYu
MgwMDHz+N0LPmbK3hGhFKTB2s2bZb7kBDmeJDfokPgdye3pok8rPV0UrIc8LtAcIVw+44uDDzMaW
wBur1eaUnK3Y1zuT9+mtKpwiquZ3p3dlNRQCoP9qjYyTEh7/3DFo5gacbBgv0Z4O3jQLDgm1Nyu3
PH3p06Iol95BAeBHV9kj0JxK1EYw22zly7zGdtk9HC4QzdpTKCNq2zQb7SeZtsvA0HDQSB6hlTt1
Jf0qb50aenaSRDnzA0/HGLygS0QEJchykjyyk/bnO7WRz93FoiP1AI+5mfkTBtbb8Nh/ya6l6hsg
wBYs+qg/Wu3KGrxM7+hIJEjBr9HVSBeTaixSSNNd6OXhygWCLOX+qtpSFJ3rmSqP8ZeuwtF+4ou3
vmVUrKnge0l6AWDZHTjgOtJrgo6e+1fMbLehc4Xsvg9FfcB0hm/SUwmAshMknztda0GVR0ThqjaY
lIXr/nqQVuAVsKPQxG4wz2DI3aBQMBm+K/sPgdWLNxmzDSYchbWhANWsot+hDSTr44lJPcjcD6EX
xflpm9YXbAAdqQOVKncILL+CxkOfqfQ+PGSzW+HUmCcnf5V/+iBCAxpKXP2l0OPl6Xlvq7tNOQYa
XK5GLi45f/fHl3iq/d48iXfZQyw0uUbzBUSqW7mOpivWKemMjjGRivkJDJn8ss8s4IuJAsKjZznh
gGuLLDWy6msxKPGSXHKdP/O2zU2lSd0zIUXG1ZULSwxnnA2SscYrdGLiZ5gFB4i3CvDNOzHx53Vk
9nKc3Jfw5fRbgvuq56UkFDmlhI1OATWh1fGJbQbccinMj6yEqlIfX3qGs8hMYkQqgCZiHZxHpnU5
RbfjW3lD+HN5XtxmudzIftYcySN8GxMDCz8QyUUCTwKsEUEKOEBeuiUuKDUZvjv8RRhoOFm2ly2k
rXK1Shr54HlDywK6e4JXP0fJj/Op2BvmUTLFCAm1KxIrQlkCCb3cjVbOm5lfYhVyCO7Av1P/Rhup
OJWsOx/wIwClBW8SWsC9hTM4xFNpancJrtOfWvJOpABeWKXV/K+XAT8FDasfPp4Nagfv/TU4FJyQ
RMx/cZMfzbKKpcE1b7FttXjhMKUE4Zk4BXyl2vEGuXKJhlwdLyzteNyDSqOlziUKqBCRYWZn2gOC
lxZ27ATWXeAUiVkZMhC+rdB1eX2fnHW61ywZI0g/RgbwLNx5pecU1pJKlJEO6IN7KxjEsqx+F8DE
lqK6XPNOrx3bnj/Cz5TryxEndXEEw9QZRfTKe/iRqjB70Hl3vX3fkQuJtXFW4xuCXiKgGXhqJc/m
MLXxwWkNoMe8iq9tLqgLvqnlJ/RnHth+4LMgebupiIYHWXwIOBR2eYYaLQ+axo/6rbp5ISDgdya1
uUbILJ6d16pAyc6eOAu+L4ZM3z+G54SHQ/6+ruOCsvL3MSPotZcoHH66WTaVN57YMzmSbjVLhwB1
kIIPl/JmBYUy/tjV3cP3aIMCs3l2oDI3xujnHwC9ZV+XbQOZDo8SCrQa8/5J60JYqyh5o3yJAIY0
c6BLnWv++4zLHQ0E9rl9Qh4xl3SEp5+gEy9hyfq/Moibb+obO54SKgfioHnm18NUe6MiYqAUwsgi
SpVxiwbB2AxFu0W16xdcDzuiuVmYPU5VVjaZB+VzWEA9N2orvKCONpCJo3FmSKkFXp7nWm1JtPok
qrPpQXIRGlZjpDeOfxS+ya3LRVYt2ZWaRVN4eym8A97w4Qeg4uehTmilhgBrGQqgfsCYu4rl+bpG
GN1U7ZSHjYvKi4EsZ0hMNbKblIwpZY9G4V0L5ocQziOAdk2Fjlq9t4gKikEUl0vNtna7Lh+w1tSu
CQ9qcoSo6o4RIWTLsVzjnHBc5Y5H9SXMvM44cge1Dx8iG9V3GAzEv4hqKto8qHkXhjq7vuNsIyXe
q774HrCXs+QclTXIb+z6S+8SeoIC7l78A2kDej6qle1j1fLZEl+nKtDwMuhWIWNIMvN17eH2g23C
gQPTGRr+dZy3gr8jEK2wEUJXzdeNHrcswm9/aNfrIxpOFhSRteF9KJki0AdKmEhBMkicOtpG4HaA
vJiSY8xgfV6u5NjFACxdtB47XyHLZoiAUxZHEpASXWjo6VSuGbWmbCiQnzTviayTlEGZGMlfOJtN
2m5fDLNF0XhI1uVJ271hkJ05qdOo/Z7uqvgG48+tugaDd1KRyivC5SuQteW7ZMSsurhQO/w4JoVu
hNm1IEpz6v8ZQeKEU1CWns6rjwhuFjSYj2yI0la27wPiuAHg8yA695Vht1Lc3a0WsCPjaMPZ7lKt
RP0fOaY4nQApHWPF+L5ppnKcmf8dxxDMRMCbD+xvk60uZyey1ZHG3esqjSmEL+EPz7ca09fmGkQT
g88HUvvBAW5BITcT9egarhLFV8t/Gh27kgBiHFTQJxTo0IKo2qPiDqDKcVOHvnZGaERfwO7/7Qey
1NrqzvZonVOsGHa5u2al7MZPvpqBepJZu04O5aDIkPXioOFgjBH8ZZXb7yBPBoSongY878YDnK2g
Fdd1OBhlBQADN14fds817T2sRoqmjE3gdTmcbOwmb42oUyVhveHy4lhd9/o7kTuWknCKdYXpPD08
knpy93gC9oD/21jnxQ6EVYropZu/bvOuJoHkZn0uREE1UBNV6xPumRkheJCg6x+p1TaClp3ntIN2
att9rCCUfyGG9SGXY9F2dtFSFfam3AZB0HnFmlgxrkV4bGR24nYvL5YHc/voEbXKxrB6S5wCrgn1
AKZWXdq4NaY+pUCNpR0+S2/FRY66YxrGIXmTLSIls58X4JWWZQQHG54sHR60CmHk8HS4/VNdIgWV
Rp80GR58xd4WSkKYhCjGaj0fGZgE0a8qJjkV2bE/R+mD4Fo7hT/N/w6qOqoNeOk6504cqv1r+lSy
8keb+OrnzpvEBilfcCIzACGFrBk7aLuMTNC4OfwwiwLePpLL7lmSR0UfYy8OsR9XeijCnvAJQbKT
PBgDtMiQ1zzbpRq7myreFi7TJelWOgfBTwZiadvM+ubvFww9HuTAKIM04pkrvgOhOOCy1VZRtywf
9cLj4I9AlHp7Rs1pgW/Sgc7a3b5cJ5GuWRTrimgphoSA4gqOtpnaIFSXS10xlPjguDwHr/27uPcB
VSHkErfMVmuoyRAcLIEp+zq5PhoD/Jx0r3H7Me5/v0ztLj9HXWNiZ2aRRXa70LQgDuHxMTG3+R2m
sGF3re+nqAjNGZcrbjEXWQsqjp30aVG5XoAXwoP4BcIQVbN6THe39vhAKd/j4qfwxonXDxylR9Wq
BQccjcRdJFIH5Djy18asrix/dDXSpFH92oS/CdHKNXhgrqjfzutJWCvYjbiko/nIKQHjE2J48js9
QMRVamXa3ynbm539nR0oOIUOPJXDlAumHDh5nHV+WqIJ7Bvx11NAN2P3/KWs+ZFhy9VHxgcUtMTB
gOlV/p0gTHzWafN59h1l1plaJlGkF3NclBd/XUZVNhBWZN5uv7HPjzAuU4nYajnqmLKU+belD5Sd
I5MqLWp7GZ7yH59wQPWf3vAsJEm36RvjvcnZMoAV6TlR8ueGOURt1cgHL15ie+SueW6j6Yr4LXaW
mfmj50wS6rj1ByCRadLM3gdS8qoRVDNp6BhV6Lykbyh4gogLGqsalWyBSbD96OPIeixHBdWuY/Kz
+uFeukJTa/bd1KPnY7IjQqW76vmm/933/qbr3D7filVPW6T26pfU4luCWOVI0yB18HPrGe5Blm37
f9VMbwVCaL92JgSREd8TUkbV3DUzKrLYtrF0t9rlTaQYnjtLvAt/ChUkBBBs4J46R0xK1eykrb4y
O3GXTMIh9M+2QYuJ5DxW46+InOaflZx0u4Zpgz9YypDuUgVEtwB1DMuIOjRloLHPVjd6GeEimA/J
VywA+4pvX8MNsuuU+eAeVUOELZDRfQNaJtniJ40hGAVd/azLtE7NIuVvmlE1eOH9kNO0Q9kXS7MX
f4RLQ9yypYIqo0I6VLbf1XC63YQ9SUwobc1oYii1X2Epmn0AY0pp1KcjguhUWzNCQFi0enFA4Da4
ZuY8ucxZXDcwbzGvyimxnzXF7fW5w+P9Jby/8eVpHD3mB+TQB6/dZKvTyFtnyQYdlDyR2Vx4v4+9
nek5/jvRyakeb4umLa5Ud43MuPfJCwzPxMcJfobXr2RnwlsLYK3m1Nazffc7we1UQ96W03mn3gki
BpUY1FnAjakofRHCmZ4ziu5d/m8Xh5Ern4I6rMDWKv8s+pZlxbfNezQiQLuEk368WsUatxxmrgK8
N2l9mZS/HLKxpJsqVSNVyPshGQOsPPMyR5q9kk+ZyocewjT5NpcwwYAI4GhfCMB4D2PB0UfQQ7+s
wn90lGWD2cWbs5x+mLmwoKhxzuPhGB+L3/GMVtC3kiZ5B5XaxU2Eyb97BNOKRyhtRIKyjhmB2Pqr
+pLUIvzfTmH1c+R9HoPKc4aM9T8XyKO/sXTEjI8D6g8Esrtpa/Ap7PIJ4l33mzlpwM1lCKF1JZvL
utjOQU1avidfb40vxwDHo4YFxAPD8AN14uYDZzbgpyYXBCYQrQJQ1d5AvDaixKQvXMDBIcqbmCYx
tH5SJ9Tuoc7pLV6E6T7Y3sippHPY
`protect end_protected
