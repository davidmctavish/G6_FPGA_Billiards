`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
peElgUBnFYE95eKYTfZrpnIvdxmsESRHI8KsUslKl3wxGUHo4Q350QpQ5Daeisknn0jkGzHu55GX
rcWj5kY+nA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
foXL846WnMuQyS+KnySX+Um8/BzYDJh1L/Vkuxz872SKIxAGcCGxqYVxF57yWDQolsPqtbmbTxiD
2XI0fyevzAuClOgGeMP5ZM88Vm9zUmlH4Rixwqs38I9V1l2L8Gvg+NRN95ddYuuiy10Q/Pt4UEEs
qCjQhrRbXX1UTL3tnew=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S7LVSqsd7mNTg02/lZZbRNeWCeanJptVPdmW2TYWEaUfEG0f3QgDXN6cw/ZtDCxyH7QM4o1eCLDV
RxW6Rj+XGbob/LSYNDUSrRqgqf3cilsMzV16ouyMdQzKDi+/yGo5EbTxg3o3GyQMx7rclF1gU476
Kqle5cy0G5goKQaLHYAtAcuu5IyFw62vJJCwLKeyLk89phhJigrHhEAfHWqibymGa90qdDo172bZ
wzci461C/JZoOjYiTJSPfBMtWF+CQn60xf/t2CPjlSGdrCt+lEUMkQNtZUjOFas7Z2ND5N0JOffg
Oby33ERGSw64g78gh717FBsgC3DWgp1tEQ+Pcw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DE4yvRnHc7oO0HWP5V28l9C8UDq2AHTE+Xd/v7COjBqDFLp+G8yc4rfOTqjOcSMNsttRrOwsbcba
7YcOCAiaOLriUv1Gry3a7kcYiqvBODr6cEj4nGbLinNtjT5raCIA9alFqfNOgSGkheyTfqzDuGa0
z/F1Lzh+WG6J9HzTI58=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
reCKS58wk9DvCHzX2jTuq4IGql4vvQcZraOqLFE0gj+VqiVbOC7zHTOkYlRpG5HtC3W3yZbAF4YB
CbsiltQhm3AfPuNR3vYI2FGLfud7FKeiL++y6CbzGTaysnARY7/FTuNDhCX5jAVm3MFsFVB0Fn6h
m/iRfUJGvHOI4Maw+HD9o9rbNphlJF5aOxGMoI+JxKNMsk7o7W1F5Ce7gh/sReh39pbvT1zX2rjZ
sSrRI1kvWPBRd5pNUI0fINF9C/+wgu+qPRNx6NKuNsUKzV9LjYwEHd2rmNuPVZ2NADQdFTsgp0aa
4oOnxY0X3MMLNsSk5palQw8GZMQRc0Ls0J4dUg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103856)
`protect data_block
2SL1HOB6XgboWv1VFRDStWRlAKGMbHbk/5iiClYFox0GSbSNI8E0Jga6Tlg+4qTcb72LHcmGwBeh
JjchL4v2t3NVuLhIphCefaiVM9oDO12qHvILHf5GetQBzARStpUIofQECvmlP9f9MSBqVu5/OhlO
56BWK3hRl0iFR3ognZk5M+Wd+GYAlF6f7PIr7DgjzySCoWSzW/tQ0Cp2/ChUu+OYQkPTP6jMNglq
k9u+4WBRv2dqeT8H7cOHE/tvYdKlo02jxzlULC3tlLEQZOyf5zF1XmekoqliMM7qjWagZmUBoLjW
0zbnZYzXksX22Mt7iAqEqO0Cf/v5bC3Q8+KyMNzyt8lIHeKcMheuO7eL5rl8G1iX+OcV27R8qxqT
BM5JIixUKCwcdezToqAdTibJgZxrwdNpZloV+oTm0dC6cYWKCqi0wPJSSzJB0/+1xMZpHQzlbDdz
nxOdVJir/WoBRH5JOOeH+kam2R6NDWDSPb6nmn5DDJkGHtfSZQ3KdA3HtnNORuC/Q33L2owJq6FO
ZDK6idZczP+Zj25OCG2Zh+fgkjf8KzzCQK/qOLHSMcpDU0GGbkRC8IpiiOcxd1yWFGzGNgja3Am6
VnbU5PBbiocQpQuuLGnYCTFsIgQS+HVfQ1/RpkIippBzGLyMfNO9izIlHf5Wm6V9duc/KaFix2UM
b8K76hback4pl62qCgNJGUCL9kwMddkSdl2natCVQk1IlEJ8nw1w8NiJIYXv4wmwiQq7T+VclC2r
G49rp1Rv3CZphS6ZH8DKcXQQyzHy0hWI/X/VuefOx252EJFhOA9bvLzqanezBO+7QzHA6bYGr/Do
MnAHUR/bkma7ymXpdRry7SZsyss4VKTbPbpv8XQz30AIGE5tjw0KrHOyF+n+X4BHNcXetRELCWY7
Pi7fthaCDfqq35RcXqY6f4rEO2rEVQUUOmZ8TQxd4TpdcCBcGLEQNoxBf6cN3CsmsDljoNDzFmx1
NPHFcVn+R26x+BDjpa4pe8lnODsblABxI+zXqpKn31mdmvMib0hziViraOCEC6GGw1eOWmnnnMVo
WRoRA99OmlMZBRZwG+VZVOg0NR3zZc4nfHhuGxpPw4jEjfxAXkUSaHS4vmzHg5K/Qp910BMD6OSB
lhhCcMIBWLG6g0Q4Y4g0lDrU7qBFAOfp0zKvypledlCwqq716epeF4bRc0DXimEpVQs8DH6Mnuuv
Ze/RiWS/TZfMHWmUqtCAQ/Hq5u3KklXyo8+FB1GpmowggB8ZuZgZ/t7OngOCkBFo1azSa+6uiTa/
HSKzL7l8WuyuCiVKfew4k/naNo7XQJEAe4q2tNlztC/1ue4sdcSDP0xbo8piQagcrn24QYxxC/Ir
bqM27PN/vECTvArF0Ryfv855u5aSb5d4S67F4f3m8QWGB2W4CW+Hy/Cz3THB9T+5UeGSk90+WC1U
z92+iCa0tcpttptGYOH7FXIyms7kfxJYXcAC0BDaHnYTgWJYoj4kaAw26Hs4d+lN9VIJqqreHEhs
iuafwwJ5bAy06JhH+0NWg72QFJ+RlABivF59xGmogU42v8homq2q0Tld0Z8o+sxn5DsMWAjJXpm9
eM986HllQK+BxUVduue5Z4atP0zt36/NAGfSl0Sc27RnQVg84KQY1VZC0SNj6vJqubIWtu+kP8rW
w9ROVvZf86SIq4qjg1D8QZMY+nOo7jNL6djac9Ei/6jZG5TYBtwRVZfxyO1ZyI97xAkKxq5UWtVZ
uzOOL+AqODR4/Ze8cmhigF1r1+FPEq9jOT1/94MD9RyUg7yt91R10QYDqma+ZpW70nFoR5C/h1Tn
rmoj1ABlD0nywt46GtC9jUxPU1HJPx5aylkKs0ULF0AdF98vYwWiJwXCjDijzW9ESDHgh+bZ6CZU
mOyYCHzAG2JvWsT9/zk65yKZNI8KREC6JQeRFA6c3SlpJTZ59Faoj7VQ1gXjwvnGmzgY4Q0rAY+f
IyK53fCqhB7vp4B+F9I4UkCZxiYIJlPyJq+rse/8C9KypCWSnKdtZZgJCutdfBljjr+aSoBvdM6c
FaNX4zLKgram8WwOyoNTJl9An7bFMAyfr9xvkBYdw76y2tq3okbxhUPOoSRLscWUu3st94SOsafF
9mGppX+4mETM9wNjz8UwfOFnR5uP0A8M8iBj8+14bDy6D2KZ5eGNesALtnfO1jZbwJBuGHBCE/jo
ystyQRAwSCRAYAi0+uVsRtQdEP9IQFlsdyvSaAEn9QTm5NsuKzAhgN8D5v7kQCFbEN2XwqZxL68g
9Po6rkYpBh9LCrpBH06J/Ucde/HLn3kB7JWNBhpkK5S+loHZqT+80KH3/9iHaBbYeqvxgjRfsRMG
a01ZNEuTzWsjeONgD/CYBjg/SOer8/dCqs51wa2nFRGYVTU2v47Rjj8assV7HLOEZNoeGXb3/aqr
+O42VFxnDG9CYay1KU8Tb8PjfKfbngciVKk3grnpbBZ7lzZ2hofrauUpWmwShIkYPgCWvC3JRksr
C4njak62b+MqF2l+SxUFfkh5EbR+Ijs5fd2vZy4d1HCAqMkCXwxfwsGeXVMfuyrmS/yoZy+OO7C5
fndTnCZv1MpfsHESPP++BYrGL7MLEx7EtEfomq6w51CB/+mKwJgI2S6nCmwB9bsjkLPNaNd5MzE+
ikIn+JOSa5/BNi+B2jOwZT/TFgZvKXtLoNdOJklS4lJ7/++38vejSSwKqz2LATlEjLWJuTxVCffQ
bkU8VILwM9UxKlHB1zi4Lmx8F6kAx5gG+Og615wAxI7800GF3pzZZIdJDloJOa9apHtkV/7WKjbE
rsF2i9CMeO9wGsG6sCfV8HYOUh0a1LHve/dMvp2DMt4dG4jQ/QsuAY+g83nmMEkyCdpVpq1QUc2e
dNS6OqvU2ePMwbP9ItvfkBvWuJOKlJcu+uZ6vBNEJAnw8d/8Kb3VbCwv9WOe8tbdnbFUe7flB0bm
mRyl8r/+5EnvYGlsDi9GWcjsezdpLmsMNAKkKQpxzvqwddLT/9obcHV3Bfex6pTNBgMPv5o6APiA
rU+XuzImof6FMMN4VaXNwLjN/ZIBYEIht5U5vqXuSoT4YD5MswSN7ngrsTWXVZ0Yma3+io71YSl5
q8Tm0arLBoN7kmp9QmYNW2OllaFAOgpYK+aHcbCdlcDEVvjr+1ApCY8NY9OVRsXMpSfg6l0ZO6I3
WBU1js4WYirweNO0i6VjTde2VOPOOcxUeaPqIeTxwiXImQ2WSUoPDDvOB8Kbrvm1SLkFIZ1Tflrb
678+UTaSTS8t8Y0w50wIBgHahdqeJqsmXWpKtcH5L3yOSSb17DXJdnotQLy8maxgvHGDqpEZvICj
YRVQCEsfWl2j738RJfMkUQsR2Gg4VDDnzgUP1PQR2xneGmD7eFUeV77+IhSOKIEWRe2v5toMWhZB
E3uU+U/gu/xuYlWjiYJlD1HL7dgmi/4kkborBMwwgnVggOVkUmTe5lAjxdFDErqAGNtMl5VTNia7
sWIdrrWFZFYvOK63rtf0Ieq8MHIYm5rs+ncFA6vzD0b+l5dGDpzfU7cewSCWBMXoJFxxlBrJ8w0q
w1K+SDTDRh+nQD73iin4rzqsoWDNoxAdDDwa7pfwmlDYRRRScphxaSUZ0oXTC8poWmK+ZRYDw7wj
51m5kCZbnejns4J/vMtn5X502dTE6MhBLL7+imi9+GfijGe4ZqmreveBliDym4udl0ra+BT8s4Lz
srpFGbWMLXoOSntq+Vrjzq2dJly61YlBL5Xoj7EJb+NBd+p/4RvuZwi4NAZ4974ND/fPI4Vdgdbv
6DfY44noqCMiuw8SLOkFIggxofA5nycK5nt3I0CyodMPeCC0uhIaZnMxOL6Y+1YAzRLeoOk0Q30m
D+GgPWj2K0zMtUmmkwXXaAA1azfWbmn4fYdHw6XF1UCIEW9dtZw08Cb/3AW00Rm+xY/Y66p1RCeI
2oh9x/nbppzP62FUVlguqx8A7jXOC6Lr2GMlQ6imVwuYtm1nx1WRHX3uxWbWF5soT73lzGjrST1J
REnH/Qy9GL+e/WnWZWAwaeuUqcZL+jgFWfDmZIvzdtRfjvIhFCf6gzLuy+r1DdJ3cB68P8unI37i
0icX/MPtkVzqxyVrCPXvpyhQhWeST58z1TE1sbnj/H/tkvpyf3uF2PVCP2QoCUIi8BKrbfJhF695
vE9nBtzxigbgm/ApG/tSv7CtnSaxUj7KVXe1w7NBUXT15igqjjIHgxdeNSXTzDaEz4bNSc5tabpO
zDImICW9A9lAxlxtyNhVrY7O8ipR+TRemFQi22oRj6S463XpH83K/gvJULb6HGCBHLgh5k4T5z1l
g7yAxC4gYwsltNoS15D6NB9ltk+9Ho1jvJxzfmRjFm/56lv8fYgl5Z+jORsI9kvfICjBnVrGpbxo
BQeNigs/oNAs8EigF+iwKvW1WmJEASd3HefmAMbG7Y14RXkdkIzePBQv0+0dS112pE52O+9QFMNs
/OhH+JiLolomShrfE+JT/ahPdTnMNxz+ajWpLJcoG4WTnUV2uW0ezss5obHxxud5zAwbrEJQAUXr
KBd1GCNCWjv6JefxxwP0kj+lus1gLy3aQJmoBTc/5NJ+n76DWm95Ahbv8fwDlE4VS4Fs4oSofWrL
T0rdJTF09+4eUv1j/FWKjPjGmh/iai0Ad18PgDPaabIkVXxxozNIMqqKMQHInJFKiHWk0aCn5Isw
TSXifCPz/2CH2o27jy/x42IxcEu7V4rMuwSrIqHe02tO9ZWDu3OmxR5uzKMNwkKuNYncUmG/BmQg
F7Gebva5Y0olVjglYPW+IsCf/CPS6HIrZGVGBffG6ATjkuWfSh2dkpEBPc4wAlMpiZXqge6TRioL
dQCtbdrLWipC4exBejBWFvr8pNDHoELDW2ld5WvgpYns1kKnoXg7Ub+T12lfXogc6mBkOje0dQUJ
N1ISUM2fBXB4sarnPxhpJQlEWvm/3tezCUIVYauNuIot8U30xhhgGPD37L90MHvEy1i+KE22iU+U
O7igciA/m97DIGJ9Q1WsMOamSZOVEMn90NuTUayvJHYLLrh0SvurvxkXlAcewAQNuDaw3usAlb0o
6pMT50dnEKOpOWLFhxXaP2ZozZgu/GAqMo5wVIMHPTd3E27AIdkyD2UVqMIt0bZbB4Bim4SkNSwj
2a2ziyjqPginkN/80pdd+SFzMzsKTFxK8H5V8RnDKNMtXhCyXecThpXdwP5IgA+0BfwoYq/LGMrf
5WYExboH5zF0b4XHg1lJ7PRVmCSBTzxX+r4mbJJsib3+DOpB/ntpKp8I1+n0IYGLPZvLcj8BON0z
N4HHai2fmzh73MskUOphZcedXRe5wTeQ29T7s2sAdbliLUOu5GE4yaPvQAWgXEbBKk7U/pvTlJMe
cZms2exIrp0MD/t/BBuGNhUPJ1wp9pI6d/l/BIb9FCe54jjoyw8N1C0PvXbwjwrdDCOprHwcUVDz
Xar/v7HJRG1Dvv3DC/n5eBdUzfo7AO0+jNx5U53dmf+aUWniG/z7nL3cZ8atIO9sueHPS4ghTdGl
E2iQV9NYcBb5iqgrYwypDQLp8OMN4JmU/eM59ElfrOclFDBfkKScvqO1biQhXo6FgnUJNL6GKlHL
60OffyLYUIS3xPHN29lm8irFiA9wLTjSjNW+jBJHe0Lh3SG3FQX5XHzUNE/p3as7oMZewToR/Kbe
uJNGqOgFZT4zvFnGT06Qjw3TYLTciXe7LClXGRQ7J9Zzbb83c6MUMQQRRhWiSYyHrvdHepuPPuIu
oi7DVHU3tqnYQOuhLiXdivMwTIkuYIOhfjzhzAvpeqm9BeR5zDXUEK3Cgeqjt+/5/7rYNPsxU+/J
78bqz71nI1uYTEoe6PKLT4sv3nCi8HakObPXi7JDU8mvzQseBB2nK0upFi5V4nrMQBVvwyMMOpQS
VeGFjfTHD9cGtcO7/js6psKNR/GQActxAaaop5ERWUKsYtp3OQ9pwlHTtvkOMxC6sf5FU2JClFfs
IpNSylox9h9AzFCi2GmsLAJGWjqLntdHfCRULt7gacitMeqUnzZMo4j31wO4slv+BfQxlyNN7QeC
xKcE+0nv5E41gr+ZxRyoOMmIoqDPuRaxnb/l6Z0PZJzJA9/74bdA/Kvw00h8hmuyQZjuzjPtaClA
AF3wfHXYE4PPEk6Nhu679mDj0kBvsJlu3SCCuUAbxHvgWsXMzKy1Db7gkaJeMA7YjBOv3V6JmwRu
uRXrpWXED8b5Ho+DuoM2XuYgXyg2dTs8ZjTB3OsDkur/T8Lo1d3PneyNyl1CIGVCqjwQ0S/gu5fO
IberFSJN3EB0DPHdt0n4Qfm52roGIo3t1MYBMH0ArZHQT2f9vpeDsZM52s9w9vI9gyc9MAVsDad1
YF6kLZmzSojb+k1gyPu0VBAWHTComVCXFSJJFhH0mb/T07sLfRSkEcKLxwwY8bi+qhNWh10OUoz6
BYG7x5uneJNVE2zSBqP/M7n0434NqF7A1HvjCnuyiHUGI4zqt3UXIPZzzczKaIqAz4m36dSoJqoP
sVRmn0eFddudpSU4eA40lRouhSNpvOo+3cupkUJ6YE2hj+phRPsGTmHDyhlPj8exw8pzBVvw1wU2
kMCvSlSQe/NSbZODdNYN/WPEg0TAHNvSh1RTLcOZOCZ9K7+pDD0B1HE4JHk8iOyv325cyNLch3lY
yv6mJMZ+eCn+t/Byi3fIEy3Cl6MUAcDvpaxoDSatb9/hrJX9oOp7WXvd3zIWXLdxJjZR11sWHMXm
qbtQCubQ1csCPZe3Bq3nzlp3w/r/vQHKubMKtufBPumjR5//Vm0lnVMTbn1hErRMYGySJJjIh1am
aqOkhS1ZqnEuZwW7lp8wx8wHUW6XQi87R3uNhb5Ljvd0+yehczVurBZBqC3n+3JLnhIy+cQSK5ks
FjAS3u+V33nmBn3uPEVG+llzO0Ig1blpv9i5A8iScnamPNef19N5qT78HbYeq7y5xJtl9QtO1mfD
do8eXyJXas6xmh6UQYlP5n6tC1WO9kDp+tjypVVu/prZ1K5XxodiiWTfIuiXPD6+m+hobt4bTmya
hs5p2RVIA7e+NNCuQQ/301QaDGfHWngdkReuhe9vRsMSFtuRnTwJvssXpqlehRBinc2YtNrXdsY6
InBNjH07gV8HdBUr5dAyUBROvsWoClqtelojCpdjU//6X4mxsF9dh6/7zHVIRaWtDqCyy15GjAbM
g0YlIn1qAhiUZGGJrptXU2OvIHRcogW3lad10ggYFMhAcedyFMShYhOt7klU4zdeFPSwK03dVi53
HEFAzrqZPs/W4STois/5hN//CzM2M9RVEUO3Rve2U1MQtnYgGgJ2mOXtoedSrzhxPkcZgk+jt4EN
nFHWKF9UcxoDpikeQqgnSglr8PD10RAuYQsFiWq34KWVHU+w3Gsh8tHSWWTdhajh7MMUpPDm+k92
MKDMYXGonZwHgmKScZQXebVKg+d8mo2gZQZxDKQIB55xKqX19bCpXvXPglj8NHUcZ+4/0Waexm+8
RUf7XOzyIKZH+7ELNzHWKaoe48FHnRU0ti04iiauQLflinGkOay4bYdJhcpkDj+sr5FWKAXiuTsz
5GpZTqJBq+Obzagfzkl3dZ6qf2MYQg1q3BJi9CwnXUDObC75VL7Xr7LYJuiK57xGsuRDCopJHUjv
+SaRe890tW7YbrNouG93WtcM3xbzKgqFrusfJIUZ8y4QN3LK3SW496JfS3R3UqgHbqQVz9YvFZiH
LEMIVRDepezAPosNTT6/4IuNwlGpBeBpSuNeggEViIStFZFB1EfrL93AkHqYQrmh2wFVyijAy8zg
qb56iUMIydLPwP2PXpQXAxNzahDOcahOuDa//cjeVGHfaf5ANQEiF6ABOfQ9f3OjFwRdYVFv9PUn
Mz7uRgVEDGv8l3dR8ZRiKGeoO+54Bsr6M/7FC1/bAV/MI6axYnnu8Qp9bBQMAZyZ66NME6pu6j67
dSEUKt19QsizYGwCAi5ri+VMy/CYHGzcV6b0QOUpvPbA6PUoihZKu0ck4lIzVPJHzrKJSWo95lfU
YCGMyZuFYlDmiCVgad9tjo9uhxJlGcUpWrOlBvYDTZLYjTERDudeGYn/tMDlw05HGZNemds/qwr5
Zov/gAamrIZh1ThoQ6InK0+4nMR5edExFlOPuBn/jNsBk2bGmEKzB9uxhfRP1Dq9pnOxjjFTZ8pu
4X3U4bCIE0VgIdl+VhA2cVXaJ83a63UKHO/Jqt98uMv1MOE4IlWH7UuXCO4JLWqHI6eZoA7cFFN6
tOQzKSsHEY+t+OcVZwbYOax1KJrsuFQ4XilW6k4I9SHnzchEkk8WBZzkiw1Qg2eoWOqu1af72Aey
DLxB/zounKqEZxAPmaJbRN8PW5CE3A/8InZt630+Xx3/jdt+x0j9UPEf0ISi/ChedN/5qr2oKzVL
DlPKkviZEYPci5VXaJO7OzYDtl6Ku8m7RQ9+elsKDdvQbF3zs5ceBclr8fmJm5oYxshw597Q174D
y39LxgFseYnZyZfvvZ2eQubblzktPpc1l5E3SaXgl4BTY9KGtn4SmWUgVPvrMlyRFDPVbQSG7dY1
7RfH9+BtHmV/Xrru/BtpLAfmTchvwcvuo9jRFtMBRSqDuUXvqnvVQZWE6teDKfwg6lao+tifYaUh
hqNC+e3l/d8NwMbfolBb5Ds/xrtei64FWxGD/IdJbyAdQloyxbDTA4Od9wfn2nrdEugqTv4BctRZ
lBieNOMIrIbcJPX/UC6KBaD1qg9sjPKo+4U1+45uJhmC6I0xOWqok5EeTOFlSaUZ/0vJP5gUV0Jq
Kch6cQiUPqiL2BZD0GEuRlKmLZjmXhCcqJ+qrV32BioexgN8Zw6jjCHH3vZgd8qkHHSrU+6iqLKw
ea1xTIMYvM9mBWG02PTM+1Igj131dVxUGC1hI+oUrc88eE9M8k/nZQuZ6HlemyF320L12jqXe0Df
oDHhpK5Hs1ctPSPtCXzWIFQJkU7HVfpcKL5mBr4cfL460vdWgwZ5MqAuiZeBCDvtZQB3AdJ2ytke
Ge2c0jaabuCUD0MrFq5IfGPhSchBcYNJUVYJsyL165/I/rciCCsF9md030RFxQuBKfJSJs8Yis9c
mRpnTB7SRohCqHqWVvU7KptR1S4mlZfnzMbArpduvcvPHcNutvysc2cDPkTkvW3SPOlgQCr7fxsA
Q89IZPI/9XLyTFmrlTGagMHM2Tos5zWAjfLi+0VjYO4f7taQC6KgpNSDC6sNpaDb2ttDE8u/kw8L
Tpfj1B6sGvxasEpcUGVsxjxOEG5ytk9s/a8iyZliViGXKqbY44tyhv21CU++TBFBS/5PW9iMneqw
Gz+smzlKgR0Rly/Q0GVfSIvEPm83TtU+5QdJsmwMAxHcD3hEDzvhw+alr/6zDcgG0xqxOpLNFx1P
ANwdUVIfnhkA3E6+D6iyxZKGpD4FFXs/++2D7M16ex0ZXlqpZ7VoRvb9o7fkUtf68L+o2cyIkKF3
dPEmqt8nZXJ0NDzJtZlbPI+3zMi/QhnTTd4rdLhixCiO990MiTmdRvD+FtNhqAGzQ76uK4XIBefi
K3X5qD/GEt0QPPgYgXeQrBzgGmN1XFhornqH4vJoqzqMlVWKrwS6vWa/Y9JfYN3RNwG+t+J4eUkz
j62NW03nX/P2ro0B2Q3pvYCHglTyO5wcwLAyGCGnUbDNJQPd8dvgnHiAe6m1ZDNpJR9YUPVUEU1E
MzPm1BKfZUsRDxrmmZ90CKyvvkdWP1XkeIJnj1qKA3k0tRQrYiM9BRdYMbeuX3gz3sNcPTbUxG2U
LXzvZ4LOVo2TGafxRwtwaRStgW2q3WH+7HBx4WIcaY2Uwb/ybGCO6P3WombKC+8jPOYCp6m75NLR
tEgx0EXMsgNfnFhli+fRfJn+Pt/ovS8vYvwUwLOjr5W8jxsTXltFqXVJ3YdfBYMN6MddqwLCVvZP
2YB826NhGMQz4BNkKPC3yXnIGCLhc1gpoE7NGdIpAjpEyC6uJ2Cqg6clmqO32KHojTpCJWbF4Oqw
UWCejt6nFacPdRuMO2/5CEthN5PRKowQA6BVAN/H2B6SnT9ggWa1Z8ER0fEkYXCn5O4zyWBjPCKQ
TWx3VjgTBpWXaNGAcMUWNDzEkz1W0K4+fGG46eMHVAa91RAjxTLFp5CLoIH41XyXfXxHIphlFuSD
mSJDeh0dKPYGcyf0Cuf3Gka9muJIgzJbn4jhL1wKJcr7H/YOp1zWALM6b9hSUaluBhDafYmZHhXn
WJgOHVlF04M+c6OeTuMDhpiFNpkBozcAwMxfCVeDG+ObEC3w2a+P2x2uAS8cPx5zkJ7bcoIvAM38
bEJMzQBwCcR/pg0VDrVNf/xWF5ptxlbUxFioORKsS5LdjDmrWScT9Q+KVxtHa3OMoOLHYSO/DQf5
gwMCWjZace8P158dRbF7UScfVd+ovJ2rOQWyfxvfKdbXGyReh8E1sKiAQaUVVYWEsLX8+PZfugoM
DBvCHwXNFaFlsEWy/Sw+/wXELi9fl+3n8DT0YwYHUKXbaqSA3B8YkgqmACzfuOTQ0k+BPetVYkdX
iQfdET4wLH3hmu85St8TuhgZFejs0klPUeVDaKVLWM6jC9q67RVbyoz5KA83aR4VAVRZhgXAixvS
Vay1mCQT0cxUeE4rmNgY8Dtf6pWu8WoTI1O/4uQuVVdBmrZ/FMEHai8eRW/IrVy0vI0fsQCtOQQ7
+EBdC9eR+nSJcjRrfNBoHKLWc5gi8/1zyqyfAUW9+OYNr62Em/24IFPD2f3edMnZgqH7A1U2MI5r
QXYUegP4d4vkYrPMjJyntF4AFVCmpvkxeWWWbgxQ7zMjkiT2m0AptOgz3jt0h/HERLgLZGJDLNk6
e8i2HNmm00loHoXOlAmMsSGVLcIOXYbgF5/aXwQoRWte09Mqjj6GvQzwAN6OMAV18uBlKElm1G3L
KtBphYGgnB+Z423gC3PvqEebDFxvcVlHgjOKQqCqOSTwrxE1NZZw/vKmHt+bCUlBeRjXeXFYVNf5
QG7HBRXbj9k/BicMMHYg5FwxuFcKvJxU1HlyXGxuAgV15BPwta1MK0Y2q+E2G6zfk5Yz3oW/ukg5
wzTlcGSTcSiwjYD+c1cTO3i+Rhay7onbRdLO7ItPHvOOxHWejOBJFoV8Rf0HWZE9XE8VCgR+LhXw
DqhLalR7ViLWMenSjfM17VepfM8e5agcFc+Ocnb7fLJM5EKfMd7B2caTX6DLGovz3jSHTSXtMt+P
RxALRjuQ+ZnnWhtt2PEf3kESH2wQTlcd8tHgYQU6XCfjf04rVqXWOO75DZv3e29AJoKtt7eyQil0
k4Rk9Z1hHbdf9twfDp/FqrURfoSw/5DG4u1XLmiFf9M6ccG9j7c+fACzi9W2dfoS+ESYF4cyfXBz
kyWv/1BSh0HWYFGq6cjjQX3p50k5EclaewRvdOSe295g6K/ZoH6xXlwPSpcAxFJ2cq4umq02CBm8
9PT9K5V+xYsKUvFY1iqxm57ESsiYzDjWXUic4OIgQP7YPYPq9bKIN+yBxHAccEVbr5kFr/EQTD7g
yaohQOlI6r3LdmPtqEO91KoGM6k9XyOVhiKKvBJC8gOlxK1+QydI0c4fF3eyKB6LE9upszqYBlbM
Ld7/smjAs3ZHBqO6Oj6LNjMcorfhNifWPXBj891BsoE9+MlhR8YRz9Qinca9jQlic2zEBzuWKuHi
m+mYTeMEwMUWC1ftybQob1Tcv32S9a+bbeMoaY0DSY7ogXIhD+pdV+omQX5tck+RKcJO8xrCBUF7
EljzlJfUPaxcoJUbCuLxWBubh/geIeWCQcbF3CHug7YcQUE4TiKoCReJbaVBSxpAD0p3+o1poHz2
WrcnDIXTQ8EQ7bssIUpBQZtWaHiCu9daqW3muL1pbihUY/7V6m7gIGhuewqD1mjHh7gHz2B3oPVo
72tqI+Sw5sFku+DK/3A/Ds+aFhRvtSjUokd/llb0R0jdGmvqocxtx0c0kzFWb4mKaAolhe1kW2WG
lLM87VkLTgMebK/jDpZMaDYCjll4AKvIi9u7IwpQAzRk2WiRf2jmpmK/e8N7+IDdaTN+4rqmChZl
anD/WBqwPZq3MeBUpeArK3J/IFFNGLEW/346uX6/FyOJCqDoVK65a4xmMjcjudVsL7O6JG1qnUYf
7hg7990c1WkOKSYFs2Z0wtxgvBdpKZJ4g7M5LFkoyFIlnXsD4ugx5MzgCLHyAZkE9FRV7ObK5Ib+
+cZZ7v/sungt3fHtJ6OM21XW3tRpfj9chC41PIHDAhZS0+NUQ/da4AGAudv7vw0z3vXLmcyL/inl
wLSDBseri2EwyEictzcGZ0abw7z9bNKyV4nyk/pBusp2eYR3qFgn6jyWrLEou79M+h/dhwbY0bdt
XPghaiXVxC1fbQn87JFFz6ATM9HfQiUMb2V7lk8JdFFr4c+lR9u1I7fHijxbQPOWA+IHPaZZqEgT
3XE9zDErio4YASIofcSVfEF9rWx3vUs344vblIasoOWraMcYGAaCGt5sBAlhGEqEBDbg8JKR+h6n
QmSF59Ejm7K6A7TEwrLQQFLFKyxa3KnsTVRQhqnnLxE5uV8+W3ro/1nY8DKkcm3a2d7qRGWowuQ5
+tGyWHbjoVGlYwrJhuKiinS2/19V9AZwfXyUU5lIKUSlftaOJDVM6YwwYidcU1in1NYYaZm6N1f9
lA3+AVf65dbew8RY4Dn4+h7uicP87VUBojll34Pp9Tm78uUQLM5Ps0A8d1E6e4HMaHOM05zgd91/
/kQVJW2PSgyS8++Hf5ykEzucFOqGHKoXX51sjb5bgJj5jMYBicqR0M5noe9dy6KuIHAasBVE9o2V
QLasms4eejnESE8oiah3UjYUCPlFE0WBKQcrVkbMoa21BEsGCDMrEcImSB7GJCkIgiSxi6GHPXv9
/1FPWauACTTE2+ru84wMeQZqWpcZuQLsa34RF6VWFaAFXUQdjw0ywg0zJ5YQJeuduh1/pZK4j4qk
KAQl0AOVuWQUImDNeDrhKXMkTF1x3B40GfQegYS+HIT4aZ30Yi0tTeTv1wTarrwZ+WKskTZCymz7
QkZB2pblKFLmyHhPZnSlX5sV+TGymcqcuGEbOSIhqzjfg2AA4v5AmTdHa4j41VAbasOZOz+M0kbU
xG96vY4slJoghwJvKJPBsvFnyD9LSB5pWifWxT14Xd3ouunwoxCzUmDZysWkddpcWQgZ9zQBCUKN
2cnY/eVpwaHNYbgKqtYh2zf6AZ5+F3TLRToHxjMQFttq/JioC1EtiemapZnMfHdrwYCdEur3kVGS
yytuXqGVS2IeWlLa3aC1u2/kd0CkbUTmi1wao81zL+gT00mxod2Z0rChxAiAnPeQDEo20By5+Fik
iiZf7BMlyyx7o/oRcPj3VdwzjHyXrBiHJKChO0lA29hrpYHk7ZXqwRWyt3+YiqXjsrbvRR3eZXG6
vaVo1Y7kmSLdY4R++220r0hoHljsfGiO0bdaXaB0a5zaGV28do5fG7m9PpugtvddPSN+IVJi96mh
hmM5hGhJQcfRZ+PiQ+u8l3dVbgRUck/xbp+X9dWdLOpVz36AemyKUumASP2g6fR9s0vWqQZF8uFI
tMiKNpsy6/yX0BqWgc7lQoF4UvFXy8RH3NfsOkqtBLPJpUaZnB9GF3aj+xKbwUKgM29k7l4LDSpf
uvai86DSbJDj794h1V6+BqeoC+03JzAzOzOGEW7pl/9djFLq635i6q/WDQWP3QbSW4bwajcGLfhu
LppN6y3iNg8OvZnMvx+/ngMC5a9yA/pyYBJ7DRwatng7VIRW5t/E9HlwlzNprVmzYMlFlCm90/0z
6hMB9F5jXxTRt1n10AVwaBcWUvm9Es3V80XoH09hHBf0BRSpTq2M7DCijuOxjM1j5M6OJSzgsICv
2ac2RgsD0/0IXuGSDDF66zL8Fqt3ms6p20Tb8To6+jh1wVUG0RYBSNbJ+1sb9SLVtroEz6Iv9A28
La+FEfWiULwiWkBItLgwNhJxzuGEXh0ajoTYdp9jvHT+sXfWqahD1ZoIjljYt8xvjshQmu8yQuwL
/F+Fat2HbHP0RXGkv4Rtt7QOM4D1UQpcmff/8tc2Ig0QKO6UF19FpCCbCYr/BjL2ubkkRLIYYt2D
agbWlWR/miuXKZyr0Ho5udBj83oRLCkrSVIjWAs7PEPkn7QFf2mYjV8B/TmJFZQhgy/SGcjUN9va
F/0wYrjFwVouXgKkCal0Hw0m3KSHHlhM35ESwaLqPbQhGDJP3Hi6I+wTboUKeqFn14Cs+16QH8PN
YFbSvErS5W1nm/g6hrbv5bvv7vwIcpWCkjDppbImKjAkoE3NcBHcsJgltTFqMqWLbWGRqiUmShEO
sWBJ5719Gbr4IUc03rJaq3rFbqc+xOGW49ZdCIHF5nhj8pruaoFXqWliZ/h12ZogIuJdM5yMMELe
jHwnbO+iS9FsY3f1pz7pWll40vVtC1yK8OHLBnDOJ8Y29g5CFTJ8NgyYW+aNUYU1D3xBfbOU0Yji
RAWDY2/yE80ClvgfT6M6ONn3yjaocEVEyY/ARVYKJ0xEOIzE6vf0d883TGE/QSnOOAbnUaSScSHF
MwIgvm2fa2r/DQSDTuXpchb4qKeiWqMHw5hMfm6BUnYjBZFRvMrs9zWJLFBGvtN1vHRZYzTHrlGF
l4yeEEX8uYKY6KABxGovo8EKa3M0n+Rma/FTvq4Ro/4I9mRYCxWX1FeGBhhp3fimFZL3Bx8MwCbp
V8Y2asg+Sv5lhSSW8GXspTniYUAEaQUwJgdE7ODyR5KANaSAP9IjL+PardpSw3hJwGav/95LtLzn
ffl04ukOVCSXzbotJBt8Ypqy8SPg1ZSxKHqWo+OAf/TrRGRLq2Who0AzkGFRAjeUs/7/6oocqbji
9gJJaOltIArSEcFOsbVp5wiGBQ3xO3lOwDTRsmA8cPMkadnMARkSiW/xN2H9zU325R4sZfgztDNR
zPpq0XLoqutsnb3KRPKUq5FoyIfjnhDo9ifdoKRkVThE6MnCG0XVOvuBPOYJAgBpy7NpQrrkbDMm
qmnwcl95GXPnAK5H3gKcW9q40dQdLcIBWtXNaKaJtQ7vdqi7tAdGEWewQE+sqnJwVc/c1koTsgKe
6psXNe3rpRMeub8GlbFiO0ZOOHjRkTcnFf6ppbzgNMb9tEy+0tFjkSjWdezV4E0maPRyo6v40/7X
dLpZhR9pmc2o/1ZWhf0cKFmw2EzOlKQzR9hD3uMFJ99WWwgLQTWsNAdRKVmgwc7Jpb6HmWzy7Mww
4krG/cTlot7d5yz/Hzen47wPt3VxMfA/fBRo8DOwcwYAWaDvQRRY9ep8Pc9VkQL88L/G+kcMNJcP
vQdS8umpO8bI4rRWKEIzj+JLcJTY270Br1iFOrO3G44AuXnwYnBDeX9lk0cEOiN5DQQ/P9mrK7ig
/n71GwG0nius05M6gc8HWeANx/vHB5hzG4YFPHh8CPPNCv7mqABLYzY8AZtztq6IX/Z7VwnIWbMG
AvmgQpysIDUyOetOgO2IBxPq7LTnkaSF7MhGqjDo3k/eJuFtklGNXTFZltTITUGovWpaMIRMegKv
hme9IAFzrGYbCEJNez/wZBHu640l/eOQzkdDfFknN3GWQMepk1rtnkwrE8cP0N0psMIKahEKbZVa
/FMBIsahrz7F5UyuPu48z9hjsVXQuajS9t92WI3XoBfcPmSggNA1Ril5B4+6fN477gK5KFd8OBOk
5sEo5FceP4A2PlJ5GpmOFU0CK6/4FU3ZWiuWkZd83aBcatJGcALlsjhe8D/93ZX4jMqUHg+dQg/a
CULlsf1lCX2KORAIGWEQyp/5h3Gzk3kCS0+jCmXRCbvgTc38QHyjFBwumj5y9o0vj+xJNB4j2lCn
8SX8tp6HJnUNkvyXv1l7r2yb3wHyrhGDkoJq6ttPBuNVFlTFkbLPPOlC+NXvj+d7udv/dz+2U8tQ
UIzwHGodZv60QneSfMlX+GCKjuZt8dyKWLGwzpyL1y0giY3jXoG84BNLALryjSJ5zLYm3jsRSOpZ
LF1UCXVEE2V9B3mcEK4P3o1xF95WOJzD6TxkeHLssskFuR12+b17Gt3/8wlSY+FZ7SRFICXYnYHK
u3BnZYA3kzGvvrnomxO+G/YLBDDRLK4AgMYi6pNXOkaBljoK6epsOf2708AYV0MWDBLe03TehKWb
OKYkopFexxCLYpdE2U+hrLbW+Xvdo++ZBofZQxbYOmaz3yaIuBMXJYHG3qIPlgYAxlCT/ipxLnlU
luHHWGcaZN8woCE2Cpc7Oa3iDt6eDz6P102qO05n2a7WBvldHPiDIwDy8jZwskZlTr/XzLgSMzzf
R0NaNqLY5nnNOa7mHuMPxsnQXIw3pzgkn1T96xzBtTkBFUQEQPvpBK+blNVfYZ0lTGHRHbbhQXhe
DmyjCVsxHNllPJpDCaRx/gTaV03y1vtA/OjxMQW+JAsy5UVG2OxlQgr9SKHkFTzLFnCkBgzedaCk
+3cN6FVEuBhVTbTa5Rv5HxoJUiurB9b6YVqb1hKhh7POEKUL57ylNiByNirXE5DqB7qpp6SSinn6
TbNw7wGiw9qOrcNx9VRvecOw+bO/GWWzSdaT6jZPDqCH5iwEHDV8nl3DTiXynkDynXyTCSfIIbpm
kNwM6qXMi8flVA0IMmBarSMM0yKjJuykK01o/7BObkN4Q0A77lRmhWrBc7ptbO+2l5jGVu/qAvrt
Noe7wF5py7r91dZD2/DQ3pAXnRVs9e1+a2Xdy5hiNIuAgaWrrY97a4Vjcjk6Vh163eTFHWXOsI9y
s62hsmE8CH4s42JlYJRERqyHbkIxv67k2W5d3KZcsFPkO52WSkKHL/rG5iR03I2zmaXFZwHLvyQl
45tU0w+kPRjG/G0zB3zvs4sDYm5y5gviP5w/XQzyl+Dp2lqF8OoEoKRqGHa8JSFVxx2uQ6N5wJyj
1kLLKz1jRQAIEOdyUHSvnjMuioUDp/bgTPNs0D3Wxonq52r+clgMhFHffx7D6Aph/elUcj3mGy82
73fFgTkfWQb0LiGxo+HqR9XckvUt1lfZPVasxL9JvfYYdW0u2yvBufdYxqh6hORngbBkNczw6ESN
bXYS8IAGdjn7yLYGs7JfL9+Y/l3ZYnB95DSUUkeEYfcK1pZ8TgtZN97YwR+40WoZ6tSNhHuQUp4g
ZDzwoebpXymVaqyH2p5hIO5iHUENwHGlOufJJ9gCDoF9WTGPbIpPMmAStVrx6SovDR0lSeKuqlt6
Y4mY6aXhd5iOYSj25etTu7gDTwP7ur4T6Q4Io/Aj+jp8WHt5Q3QU1e83aYk0M5mp4vFi5xbSAify
MYjIf1kM8GDO97J9HMw0lvxeGzCiuPx6QhjqBth/JVIJtp+pdhcGHmtX2oIO5H94CSnGVsXc8NSE
Nc4lsleqpkduRbD+hSEfrHspthcPha3VGJnIE4coRDwddsaIIPVbyaQWF+Nndqmdb0xaua7Ur/h1
/V99iQr9O9q8ty39QPNcQhgsG7BfoBK0eHu5cEhaUj42CQmCTeUNW9qoW8hQYJxM4ZbOeq/CC8rJ
rw5NxidsJY0s8eRXmlvSLvNBPDG+wCc/x8glSlUOTiWaRlhWb73DtlSRZmh77vlU+Qvp7wlJF2yw
+2dQM/bII2Q3YpSGs3YujQIEXeqI8ZfcqqIp2UCHgdt3028i4dZrEp4VMUZs8KEQsft47O881/3G
hZEuQrBo0JxvKqG+Y4LnG1SwhLnzm/mZrF/APtIr2yiC/9OXrJdWXdcamKwSopHJc7D15zXwUwxk
zIGVuVHNNymymbEh8OcLLS4X7aBHhHTkQVEPi+zU3l5hhukz++WU8zcOIPmLGSCaIvu86wsFCnh7
GFvzncjAO9pczL/oWEHQAhe5xgM4zW6vxy5A5ObW3HRc8ZUGmNBCYcC22NvzcPJQrjLcb4mBxumL
m9tc95Hl9+eUeUTrp5YUGVMDolKsTkNHM1F1WxpX6XNYlywhD7KxZByYn2sFwDpcXWsBuNW5leDD
odGCt4RDomTUARFg3yNtmUqmVwOvu5Vy2atJK2pwbCdaHMhWdpy3a8gM5aWI2Zp5rRxk9+17evCP
DvlIoEqVqg60c4ODDijClDQhiW31PoiYsMUJTWpDITrFH4S6FhwdgQJ8SnMaY1YCrYT+JJVI6ufY
YX5chOpGJB6Yw6VnUU91Msmvpv0Ahlt4TB9CRavGwJv06YQ0mkFFiXREmFRr9r/80A6cO/B4Sk4P
yS3k/mOyAjOAjEVOz96uI11RrriqRuiB0KqM5nkcrb+Mus+qXI3YaH+4N4y1swzxWivLHAx/th1u
hsoii8QMBC4L/Sed0is9YVP2/lVoFLdA0CXgPi2o09p6B65KCNdFdTLw8/2fxDreuJP/ZXZpofqw
vQ2/8aveYOLdn293t3JHF2z/BH0ro1qguJDj2Tz1N7T5nFa2PUcAzEQ12aj+fpdZMa/fv/FCJ4HD
JIoeywSoE5j+g1Hjw5XqKyZYsvSb7Lk4HlSZyVEC+uLuLbDSWu9/l0BQxnrYlw+gQA5EmziOL7Cr
gUkLHZTX3b8WJNNNMdzdS0BBKk4l3VtmPwY2ezVYJwaC9aIWNPS92m4BZgGsUiV3HDbVKzSuzLBW
QQBbZ1xOYTiuPK8aB6VK229/jYXybmG+wDesYOt4pQDm8gQTOLhItGeAhP5MdGcqwMqpAcL0YwES
HfaP2ooePuBFmrbfL+67a3sYEaB02coQ3ht3o/W3qsRsafZBKOkV2iV1WXy+cjhKU3owfJ9/VWij
jzpcsp2c5Arvn35EjQo3iOdZmjX70qS3pyzni6xMEV52TSPwq8YMJqaXLSmxEcaarKOT/sP63OLu
7sXuLMsCzhJeRag5KLCq6BHJ2Ltp23bAaJLLeEJ9vqXi2kQgMq+mCElysoEFIIleFclJJFuBF0zh
i8YxXAc7a4I+KWyE2RfHmZaZ8qenTseAHcgvwQ6O0d4mB4aFcvB53qFid+0nb7Z5XKdzDQbCM2Dq
0K6w5LSCa+at/uzPe8mVXMoJRZh1fS70rLAXYrTosF+lQILrGXRNO1BJZe+htDwdIKa9AAiO7r0X
S9ughyULmAV2rCs5kOLpfYCBW/EOvMB0lEwKvElClfLMNwyYqIM8mfFh1jABmzYtZg4AHWVsEMF9
DOns9+p/7FuHkv3xsmRvP4R/7e9yev2e6jL3IqJ2aj2AhVZvAjFMGQtFrKCyP7ofTu0xO352CmHW
6OsTxjaVZV9AqeRrXqJ6YKoRE7kxyzc2B37p7ZkoB38IcVKSiWCzeG+uFtbg5j2+GEl3D1W0K+eT
dhFxqfarmm2yMt4bnq5uzJ1WFP8WG0jCGm5h/mx8jZxooDtdM9nUjRqgn8hzJoq2ZzubXnd4betB
vd0y7Jy2RzisLQCZ9i2h67RJicaYsJOE/9doqW+9HRyGrv63AUwJEtGEAVcM486up/VJV0Rcfifb
6RGpGkrplvmAHuiUVSwMibOH2fTyUNtnGFJIuZKFTesPiCtS6yn8jRxUehOq0oG7KiBjq3fiQHWn
0K1QnpQp9qD6JVMvCE37LDeODvWZD1lLQv3nrq5Qyee51h46Tj/vG2P5tBssdTeHydi7zgcgu3vm
PSfR1PcGAH3gpnFOQQwV5YgvQ05UhSrkL/XEpKHZJTNCS9JSqWLQSMSRuUA7RpAVNXyOGM3e0mUE
XFTr+Foh10UgQ+AywwNWN5jRin3bE4o2lmG0zPTPsU49JOJ6zAs2WP0tP0+uetAKnh8KiRMYHzjr
1+D0Kj3rG3cw4KM8GastqNYcibjh0O65rz7WcWLaZaCMiDUA7XXhuHlvaNkDeZ5+ZKmgsMVxP7L0
+UPA+DlWdzj6dmFU/08kzxyyRmvclpfkT7K83PsFhHZUzCnIH/C8+cd6x8NkeVpN/O+vLQLh62hr
/eq8zHmXGge1vN/0T9B74XXpALPjRzyxYQg/1iHMoWlfAR8kGH9vh7W5CG74Xqkr5SBOfukZgp0+
MiBNdpqbVWzQzO8YDHyi086lY1owi3VUSZBThbn7wabCb76TR5QHQ1N0afTTXB6Qj3Fn7PlIjQTP
EEt0Uva1SPw+sV9LRZCguL0zRD59rTJ3rPJrVMgQhE/HiQm1ZwJEtNQESaJjy53SOZePAnFajKe1
td7EP32/q7aYI8xbrbbxn1jnGe8JHJpwIDF3rNc8cKOsoOkcsT6FuHwrvQBs1TXPHbDL7RfMziUN
t3PBOiJgRlSrve7LsEdmiC0uhUqEqHa0AKMzr7t9MwvxqUYmT2kCCEhz9Ozv9Vw1EMIwYH5rYWkm
uTMgr6VQQ2MaT9emxMBN1leftqnSKsIEF6l+o/E6BsTSUoo4HvEBb4x68g4c9a4wtFDq493IJ+XN
13Q5skRsMctICSljvMVM10fcVELtHYJIzUT7woMSwWbth/KvPeUEE+nNs69bw7NDK30+ngTbM95q
w4b+VZZhgMNz/bYbwpWee6Eh4tF7jKJY1lVq6IDusHuxymFK4lDncbDY73Xl7Jxr4sN4FlpfYQ+1
2Tiz6yT2VEbt9z83g6TzOY7DStcVOPDSTp8PGA2o384/1vmTkjIXhfYhPpiAlh5z+m5ZaH6tsiY6
MWLbB5U5DhBJTE1yExeafhM4+Y/y6gZkyeRqTJeFYsTMTqqG93BUm9BxJqhTdXfA8cLIWgUCnfls
zQr6lsNFfvBjxH+e2agq3BPcLBX7Xvv5QoxzymRIBD/ayTAvCbmd8e6sf8PTYXx420nLhhddUPTV
2MA0NVaOLoAyEllbeUA0etaCEfjceKJ7f31eux/lN1WhNFKoXIiDL8FsSzB30ZISq8vG+LBOHFJ+
pS+qtAZHBZw/AIRfoiHyZzFfNFBpzNe1fqaZ2U8x9XrQGYXGqpwwJ08OjJT47WBSVcU+ob3xJ4vy
r5R8mzW5MM1qXMuJ1zA69hZDaqX8O2VMliOwePySN6vveqFOSUv8Eiw8AjWM0beLH3q4NsOD3dhM
ONGyqT5QQ1qqai8/Hm2mJIhagTJpbjRtlrz5auMUwcnUv5WrAwpCzFIyFremyHdJbzxMhPn3vhkV
wuXiraBTQY8YfmcIUyfkzrt5sjr+NftCwSV41Apf9TYxUBHt9RC/f7okVEwSqP/vFqnXm74hnk6a
LiL2I2criUYAFOFfPUtDy9eZXXVPAjqxL31O9ZyYQtLSvt26KJdZzzlRwAqXoobZr0a4hYs/YUal
mmH51MuNQnyvsReoepcOYrufM12rsxAuRt0TWoizPD/o6z7MMaVx1WxmsyR97OxewkjGxCfE5Od9
Dq8ReWrRS66nJodTxvSeBFlCPVTL20QIRFHnGiqf/yUopJPy6xVJ8hF/SE6+B47jN1q/TWB4Ferp
Uj8OyxCNg6NJYwiMD/GWpfGNdUWNVx0NKtvEFl+Y4gssaQn2kEN9Icpar5RJ+F7yrAXaIRu2Xmoj
XH8yT7qIOK29tAHp5SyBzhq2Dkc6WmCEp2kTTMnV7hTAEPQrf8QhZKcoIlFqhkqAB01EA2xfopyt
oQn+e6NDe14S6aII38uCRShcQNVjMoivVQfABtAv9gk3cVIUZeM6MbXj/h0IJ2HnOQNcBGU1J1At
4wPbdmeocDihPIiQQa1NoFOgRDZUZKYwinSr+2AHKe/N3+3jTrF/n4dxeV/8ksoGC4WBERV05ywv
8m6UhTnfMuq2FneEgl9GqK05yDZvoNEQoQMdsKY3wZcd6BaZTtHahTmISHc/SP1CTYl836ddEYhK
f2d17HqXW0irDCjj6hTIS1CtMjKiCKkgNhKK2tuFxzJew/rnAra7EE885jQnxFQU5qz3Q9ocuLIg
zZFbocveOjy/dfgysLBAlQ0O3iQv0NO+i+F2pLtKtS6oy68/VqjIkFu78Q7/XHjBo5Ho+0LO+6hl
EZOlSuWa76epXbNqyCiMCyHFvhpZpUDaUd2P40pAsAdryd9xLP7EcdJ0dQvXprdHcdQPWkw8PkJX
d4VD6pIRbvgPtrxZt//ijwF4F1iYJ8wSXqwHkb7cW2ks/G3N/IWXoUwKTVOHTI44XbSrnEI+Mvoh
EFw49TlezOFGI/mQIxpF4Ju7D9OBEyZYKMuO7FdsTrGsKRBv5kRQgysC6zl9ClTXAqamKSScAgPm
3X5I0DbilJ/V1EfuSqozesgTmgWoBuVeYoUAtLHxjPM7siOZExsf927Vp79E+O4iCLzXV+CI0J4I
7TU9Ir2dBLEprmAP7bKJafoD00yrS7lrNfcRnkeOw/pDyzrgEH2nMcikZWmiAzQqC1EzbDWcqPsA
XqLtzLy9xnyYdToScMKiZpWls08lY7Y3Wjmy7FcLM/eHzTeVQgfXEP4bcul9qVplcIOQqbReV6d9
qYYR9HHwNSiPnkFWhR+6AwKx9tcbaCh7j20il/fJEwI2jMk5yAI/sT73Q9x8MaSzcPN/ovRLMRY7
cX/EmUoTyGs97A+xLW2ytkW2TbSYfu/nD0wllDGEv9JHFzsyvCP8jFnLCzMGOxBuG9o3XQPzDe0g
2ihPeYLW7wDPMYqSUA2KqULKizPuTpuEhfOefTowoGss5MOj2FNDgJfIceZVOiOQrKv7oy/5ra1m
hfmeMb5clN5Ep/JVhxj1jaG1miBzOZaTsErrOGq2Gq01TkxfprP6CPzZS/9u9Lxirqjxcz4run3W
eX3y2YNt0M+a/dcU996pTHLQBsSBz44Pgxl7uKBp2/pVUcewPYOAtSNwuQUn8RquhFyZPghB0y9v
pj1VykBZ346hmmWeHkDKhIT/DlnXeGKSTPtHwTpkWA6eAWzltIpF+8znRGNGlzu8u+vGjgWYRYzG
iZFlKftQhjFhwq2KzynXVMk4x7S43xoh8KTQOWhIOYXuKGMgYcRXQYaY5x3J7mdjQg8p2t2vMb4g
2V5V0Wq67DMmhdoWasgU9/R3n+7bUD1eUai0E4viHBtj1c44pQ4JIgRS9o9JcF9gUr60++sQ8Alq
xr8QFKsBadClYkizD76wMNVpsTt2LkP3adW9P2Qztb96GGiLTYtjPW4x5XQp7gJkGU9odz+z+Op0
a/vWauPXnnf1zMG51jfW6DQgO/ZdKb8sq4e15r9o8/w3WEI7u+tEaxICb6Dsdi/4ytqTfsDSfLJZ
LK2fRd0DVIV9goRGAOBOJfCyPbKh2h8UIfdNTw9mH8vqzOoznNO5CUkUoWPpM6PNcaVgnHwgEoRu
6nPNE3KLYb8KDmDhq3zPP5feGA8NT5KIfFwg4FCko9Vz6wBbO8zIwO8p/ZB48RlV7MCSThd6jqca
MxmN15eqDactn+9baLC4qfyES/QlPUoWuQGzY2Ye+rMi0dL+1Lr1b5M6CPmGwZdXDCJlVNXCal3o
c9pVvOAkOZ1f5/ZE1qSCJcbVPobzb5FasXp6NlydAgBVc1xUfwDMOxV9faiuJK62oLWVzu16lmMW
z6bI8ve7zpoRSfOGFzUqUx6DhPNMs5IMkwaqV+KdPridpSh7BaN/cg9Ff3pHdfriPe9B4hn8di5z
2CGUkA/AeNgwg+RB4NgDAh5dQTdvNR3szAP6eTWO93GSCaGgzQuE62VQKh4BRMMOe4d9MlocUc/s
50e0rahrcRCqOk7D+qDOuPfOOcHq0HVH83UjR0IIhg1HGqzRNn4Lj7Hj0R4P48x7wnuKFG/HONqT
cEaLMJmhsIWQkHD5qeOX+aAx842e83lcLVa2V8b5rf9z6YfmMQOoK+jTrRZdHqDVMOKbW9zdSDh6
q1TjIoIwUbT+wJqMWWmVqDsSVTKxBRyLNb0LDsKdtxRkMrzuTpzP8bNKK6oiHB/xE44Ew0IeibpN
lA+OR5j7mI2D+vFE+m6cJ5Pagy7w0gt1ss+VKqWzrcFiJKaTfeF6r0UCiaBPjX3xmtZgw0SVVwZU
jJxFIw3baTSp8vVKL5jLoiTBjYIT1e/Dc1Lr3A8y94JgsBLp2Ms9WrEu0UuOxcQYD23NnMETmq+N
BcE8knCq1XIZR514FtCNd8XF3PWgB5gfvMqDcB9svGECM96Ls+FW/vXdOIxSu0uYl0KDRRnc1kZi
GSbPfU1i7iCs3gIvqhlIq7n4u18XoauEC8X3Kp0LcbtBPrpx1FFQD7LCGcu+IkhDYukoAuyjymxV
1PE91GpF2pd8E6zK6pfvVZWGuzw4GnQbPA8h7BTrAXRdCQZjILd68KYD3PR3p82hGtbU3dkimUFc
SRZ0Vlf3b6dKwsvof5wEH3vyq2RDvoUrBgfxnZxNROmHEza2rPQDCXrpMF6QPn2A1c3sX2ZjX7oq
BVY5v5vTnNIgnke0VTcR+xhtSjMId5FVw0ymZgYEpImKFsOJGVa81qStc3uqlMfDIBKhYn04DuLb
MpOf0uvGYQgn99/eb1/x8k8A2Pb/3uGKk9kXw84W35FYAgah0awPj+zWTlMBVn92ONukQI0bBxXk
UjpHzX+RjPGYSXv1Am3DivHGDvmMeZfvA1irZ3Y47dqzG3y+q8QRxfT2vlPyoQI/Pdus0o6HqG7u
jhXN6AiNEQ8qWaYUf7OsA3raVYRIvPd9F9jOb7y3Q7T8rRb/3Fevm7NQskiCRiEBzPMUtIZF0NWj
svQdVHWG4eWLDuOrGhTo6o/20I7XO6b+K3PHft6aFopIl1vv1dsyMyAaq4AT/FEL1m3k4VThay+2
GqOJ2noZXIFXtkEOZA4P7x7ukA2juY0mOELL0yeRrnlrI5x+w2pVPPwBjtcSyp98AQOoMjNhGlCQ
DoT5JG1bzjYXhLMyQdwyzbjuzLmn4duDYwzsqBM9wN0xUi916cfrgptNhrmTyM08X6UWhefFpc1I
hR/Nvbk9O/5URH14Ew1uEJKqoQb1JjJaAA/OCN8M1gkQcTRC9goCX6lG3ezkv4/PASNGSRQVt8xR
3jtu98bi6QPDp2uBKT47epIxiqZ1c2BWNaq6ROu/slpEr4t+XAaC3oiVlrCxAu6Im4UaA4ucPeHn
Wq+4XmTzSEa2c4hupAn+I+HdqHWgae8MOV/jTfzTm85TTSndOaRkLHFacDqo5vxV/ynQ/wDScZ5d
mUGT5zzTYFPrRuRf1DQcB1bC5ofVccBn1+KnI2m2o3UODzqhxUz6VgA2vk1v7ECa+UKRcl0QDU3+
stI12/qYWqJoSfcynXt6v2DjKX1wkgjz+bEs0e1nZpVWiSXsVLoA9xsRbDGAIm7wX60LQJDkMFZ3
weIsN1EQvaIFK8/Rl94iB+WRIFdiC5LENiBMZ4HYGOyPF6KBIU/SGoJKS4jdfOi6pDhrZy/rPgNt
yiQUwmA+NLnE7rtJQhmtVHjSfolu37DIgU36rTA5tOVxnrchTuq8NiMjeDIDqXp4/O8gQXsdYrSt
RFcx23qAN6hafgGAXTVg5BFQ4b4n2aBWiQW+LSsPL7FSMeaz8XzJLmjuREkFStnduu9wKPpw8fIb
NjK7yOWCEeb1/eA6Y6tqM1m8VRvsJBmFJhlX7JVI/Ph6AecxwN98WmzA2tPZpM+fVHEs8vGAr2pI
03s9LJk916kpyjBjW+LJdxWhEAnHiGRvSYodWeoYqQ9hgQt3pLf4r6qE82AW7UTiCLvsZQUIDk5m
54U6QC3VqDreWZlRAlgVlHPBZ0bNCoZp1cjWgr0qcMStYKqCAx1rG+LJzsFRp5Z7fGCEEanMuXRy
1p+VSil3bfo9BQvi3TeE/BDoCgycLo9j59cCFYIH9AKKJivHi37WvCjbaLL0lURnPVYD2HxOy0t3
hE2cegyy+SWyYH8kcF4FTKsGbGU3AfUKeyRWOSlyMHQrKVWiixb0ngZqQgdhOac2vlhiWkpZWtMJ
ZM/E8zurIAev3BNWDV4xobA8B2LPWP2gDo1Itv//BvE28YRrh8NuuQkn/FHgMwVZLDJJL8CViZlX
D9i94f5YaPj/5eQYDSEjlX8SNr2eYbfBui2RHTkXpGPfX9CGCzj4PmiuQaWpV9LYu6iMOEGQNEr/
SthCRZAIF7aHF+iQJKJnR3fs36PcOy8RgTu27/8JjNfr4ZNEFI32kjYvQ2y8YS7+3gAutrHHzrY1
Sqg3nM1nh/7L8UNhwQUVLNAgo3Y5Su6ir1gnf+2yEGOHjXskE4YceU6tbZ+1glUPNYKN9sopS7D9
QAngvSzn66cYNLX9FRBY8Nt3wsXMkL0cx/HVLsFFU12SCgXPl5uFmLEpB6PYHiaEhzrq3JdOXp8+
ggzC16zCuiSPYfWDtV1PzDUCdmHS+feY2SP7OUC0JNeySPQV/D+dlWxYKxuQJ6uToKLb/KsdmMnH
1EqqXQOpgCSam68WbFegq/xLNOaHS8/XcUXNh3zJSO9UPmXiM2hIeJgtjsVCz+FGD1eoNTIJ4VCT
5rcSgAS1FKoXTn7C2EG2p0bvr7sM+ptolgvumMNHu5DTeNy7xV1/5MDAQBX4RwsDsxok9QCY66lo
XyPL/G7UAnf/4Zu6pOyjGalIMNggiinxL/i97ochUAPhtZFG9hjagBRFHgpKIfDAd8RIpqtatcI6
xOX4HHoaiO9sY+lJ4pkqz9MUuHn4gHgklrvzi6XRx5C8PFZWBMUWTCSmDDfx0zoRNO7nTh+PUaeh
ck2rF5QPT7DFV1d8nPd1GcgEcBpsjTCeb23JZ1zZxmABWKyxXcluCc5oYVrdBotsLOsMMp/7Ifuf
g4L3EN8dGcSLD3M/i1B0sLI65i1vAj6asIwQrMDC0v1G0Bo+vd9JnqmLpWjO7qah6ZAQUNZH+P8F
lcGtjFyPXMXcHgD6f5RkhW2AHqQGkHae1NEYQJyS7B51PIUYPKPpHFVgygiPlar3fDVyAzR7fcZ6
1kRsCmuyZoNni9VUlhilZKmdZ/saZiqIrOym5+SNlupcdeN8HZolQODHxrRl53QpgBWo0brB/BzO
Rr62xC7KjMKg21Qfj8QJRcR4sfj9x4BFXu05sIyW6NjpV9bY9t64T2aRwIzWaznNeCjkWBmh0qLy
idPHxjphVX8ZPe+VK1WxVnNBxgetIwH36lh/E1gpGGTPyuaT7WlyOW+JZbI751hh/fy2rordsOh7
8IezUF7lzaEHDAh4HAtNCQ8QEWU9Qac6zc4lZ/cjh6qGz7qa/3O7FSsKbz6w/+BQarhY+gYsy/DK
HLiGw3/WnBUmwpXvyI1ELLmDuaoegLv/17ZktDDv/aCFpAm0WdNgF2PVLHcO5DVO6wnUcGNBB5B6
2haADHiyG5w16oPePUKrzBa7zQKMI3oJifsezreNO6blTZDa1rk+NZ6LGAFOQ/KxDoS2K4DD95eK
WX+wVQl5pIXuNcFKvCYyEsudThCenYNLdq9i8mWlgFhSuYA/Bhw3Y21UgJu9UthKdKIfxPDwoKOA
oxKgHMou5zGQSZszuy/D7awBYVtWHLIYqYyYmFEz9OZOCOSlOz/4WNYZA0AKHOEzRgc+Ea7XNRgZ
BSsKlA80T6H6kqUZ90L6AUXt//8T4QGNYnEm5dAyK4/u2DSXzVH8Ngcfb+GOsrubMYGu0NsU8UMT
FCBFLYxExGyWcu73CL2eVHQGi5qZkO0Z/0nQd4lCebGoQOPe/ApPvVHob6d3Iszy2tU/M1xwO/Jv
JDonUIAuIovExV/DUJ4qZtUmyVLPk1mGI2EkjXzA1Dtfsb/zb3YkBJsDlMudSTnLN3IRbMVf5XTR
ecVJzlAcyzq9qc772L7IjXD9QbPB072dAT7ABfMxwh7entK2OFb70JcDtzJYzKKV872K/FCRCbeH
6Ho+uOI3RvUB7YXW40P2JX6FxbHGqXrYSaAuQN4E9Z2HbcgRScIarKMiTL02swXXIYKV/7WhnOt5
oRk+KZ8TF9R1qOp6poHo0TOomU/ccmBKk/8OtvE7MTsRYcfYGPjEy8edBsjmOlS9d1LF4TEPc+CH
LOed4z6v5nhNgghejAyTPYP5KxV42ot5BerF/JUxMEq9BPw5/2KlLa7RYnP3D4StOIqbIdXjdj3M
2cPviAd42Ed0okistiWzS/Ou8pMi3MTARVOmErD212377ocVS0o1lKfLRJkSvZu4AEUjvsuo6EWP
zWmNm4rdeNo9HBBUQq6tHRZXXlMx/QIoRXoDA3UliG25x9RC1XA+DDnwhl7jtrYntTFD4Ro013ZZ
mpF/jJRweU+O/xD7SwHarezqqIKDUUPNPpJlrEkltE/lNuJlkjA2ps1IHe/qxI5b/wKoD9YMLIwA
TqZsKv610GWiUrTou1UHIRtr+gqDfCODeum6KxcevbdDJ03neu8GdQRx3jfW2QGSPeV9m/Ttc7Jn
lTbGo9xJYKFbHnBu0uYwsKOKOMWc67MO7iVbbKAgnph9VB3KWO6ChI0hpMIAd5gKZxovzhkVXkAk
8xpfFyoUHOt51v7DM2Fw+C2uCser7gjNNJeSc3XnasJqvBTensl7t7z88/q+Kv2N4dXiPMuuuVqR
7X4sbDn2NrTyMND3fLPWfxlOcR+znE0yWFXY5HD44daqhZF9GFG249MdWqtKd5bQWEHSss93YPi3
18FiDVIWtB28XSYvsleSYpdSTMC8oQUsl0TlVXNEiAUqPTpRuld2Mmzk2xKGRdWVFGuSn8rSMR5Q
Oaf5BstcTjEZ5ePMtfCRUncFrgiQc6H6c9mJfFpsitHpiBcj2ZI+eVkCN4/erXggNmOgE36/zaw9
dNJjuwXY1/zfftTqLL6oNYYNqWJ0NtUjwEm+CrrV6BTW8gk9asKGnHxUPrR//hn5NqqacqRECTZD
0SqpOKkI++50ZetqWsLDfxXTOFJPiySzx6CNhZtWQbfjp7D/UBgq9jWiwbiC+mIMN3u6rSe1iyUh
SBoTf/lY+pCjpcUL82W2C6yqwHoIQIl+T4TozlUEtmh4yWuZbF+5ZgNWsgn6CqLTU9KLjgbHczMj
BbkRs1v9w06f3z899xGjhthp20nuCRVTUDo0seO4pKaqUR6032xI9Icff4DlUUnwH8a/7zt+6J4P
vPCldkWudfna9L7MpsaYso8EV0iKAaMABeWQMCAT4iXnNFC8Lp+K7ofOFUYzkRNQYdUKMoTNLlKB
++2b+iEKsddbumuCgua5Gol+6SMs1DbslIeTM8VYshH8BN/mpCF5V7wKjV4eQdlpJqGy7GC5Ok1w
ct/rPzRQ/O86pve4ob5gQ9ZLLf/x/Jo5RioLbocCYnSuS8LYTJ6aOPxftEgM1Rxsx5utVZtGrnhF
UmlCnHN4fm1zWvTRzOMFz9dw0MaI5mC1vdwMTgslKR2vMi7fLfeI1rg/VlsrrG1RfoXQM28LldF3
IXyKMKZN+F1hrkuZxStaJCoJC2ZIEtNQhU544GQ40qdhfFmZWtVnt8KylQjnYskBJ99eAy0UD2Sc
79HhIXmg9mMJAYjrDT03LhNLKcQL/TOYFsmnGOsAUGEjebSS6U2KXJ36iDfy45HcEVf5gMc/vGgW
Zehue8EN95hk7ttkgrrTmabx4ydWmI97FEgdVecqaZaF0B0ENYpCRGVSAtyLNLTdRcI8AiXpOloW
CZTUcHVsw/T1LNUGBjomkzyDomgMZv/sjC7ydkNW11zMU0ZfZe7MJC4tXjI6DHwxAm5odmjp+bV0
Jss0js+9xRgPaVdtmR+ej8vkjJR/nAiyqkCh7SU4lvE01+nVIVTbTIJ2pqYJZ19U4YphecNmDLC6
ZXPeW/mxkaHWzfoU7Y23wczTsmKE9QQ5ztZyrEOP69ugUNJkRrM4aEQHgcmMZBiaypJONmutEu7f
GujisbYubkVal7OZxe5A8wnxvaH14ZbR3RhP1rbk1zO618u4B6MkZTU30BeBxzDiKGGs5U9O9QDo
M6UNsIrDQtjjhTibrMr+ls6Z+u/5Z/4txLOfSIWbL8X68G/Y4qMubAUgwM9V9RkABgDv6qiuF3uF
lTAGDKdfZqKZSvkcDDuSY9FgeV1Gd3EMc+3E+XLKf88x5cpQX4avAQKF8siWa1+F24KuxK2ebPW+
3z4pY64bsquoTNquDXave0RRDLrgUpw9xs/NiP7xt4kuGLekbf1xRzRqDiAK/v1HwCLgwXEqrk7w
XHXKZOemKtQ5Pgh9uvtLKGEepTPwjv0LI0pwkh4CfaoVgT9WoXwSImLLAp+U+AB7nmMstxCzQrNP
ZVQ9yTVFWxSDRS0TkeHkig9faswturTShGSiRnIf1chgm+7OrWlgrODFma7tzjcdWZ1Ee5mHqokX
NHMZxCg2JjVQooTp6Qx+3e0/yiWt+qlJsUl6r2JUnQdq6lXQR6D4ZRGScs+iwoqwXm5CvTf4btMZ
1P6oos+Y3egrPgjGonZ6IbQeNE5R6vdLCM4g1WO06dlv1nqgCbzJr2prUDyzpGuA1dT9J8x5udwW
W1pgENV5DgFIhbAuaSldRix6dXnspXGTPzAz4BvfwDU2TAA+WSnxu3b/md6Bep68glVT1im9Ph3T
cdvHRcof3leBsDi7OYACwYIA79vCz4KMHQ1Wm4vHJc+mo5F61dYPBtQrDKNUSDa0+sJ9tUPUKOUa
kpBzf7HAiSSMTMdj/23QIZ5zfnWJuAZ3mU9QEhCik1MpsID3eRFtZIWXrWCRsyrsUOOmCtpmITOz
Ip28tmgaic2BkfgQtZNaUS4KtNd1bNalb0TrNbJD8ABL93XtTKl4qM9GMoAHSWSVPtXXNwiKsdec
hpvsDdIi8KuypPlxOjl6Qyt/SPYZOajGz/CIPe3IatrIy1p+yj1oKZvVXzfVeUh808CLk4EoTCNo
r04ZQNWQBKRXtYzB8UoJXbv1nSS/Td3Cev0ohQQiyRUA+1C/KZhWsuQF3hrq3U5RKlsPUKpeMSyj
rQWMoVhTClTHgudqu+YJJsix1bEit5ytFAR4lkZ7QcEHUFFBCoPPUKknMAdoKZ2A6VvJliLnJY61
NYcMPyuwfjtM2ArRJtxe9pSMY6uSDjZXrUXh78xbTctlXHzTg4nhv4FHIAGg1zhwhNJRiNPsketm
Mg2iuj+7L77gkgQJclcHA41kJXk5qoW/aeRvf81IB2gb/64XpCjrzOCCKLxY4BFKTqszYcXRiVfU
SQaLOF0Jw5UPct/20XeW9AS5PpSwF50Yyr9GtfTFq8TM/FcbWwfw56J0Qilah0DHsJpOm5cEfcMY
R/k9oz5fxjVbBX3q2petNnUdkA11AEVcluP6KIQlAvmGaZPCafAYvL8+7Q855SIpdr8wXjdi2oCW
r5U1JCQNCL7Dt/4K8GNtYrnWRrA35Wc3v7P+WkBCqAvVSCao/6qKqF8oG7bq6VMYh8Kpj6NjodZo
Y8CWxam8BURdKk4ep25wwroFeiUq3U0PzN3oBQyImVmr1EOHViWSXhkGTNnqsQ29z2KdQEM5qLwO
zSsGlQg2AyBAyUsWAoVZvyZgPco6Kwh5vms/xM/kqf760sJWPxQlTiqXBqw6ZpZduSm4FqkuXbAw
4+X/L8JmbyGCSl1w1i6LS34JYGgWtC56NF/frf7QFWlwixvqxSCgkxgi1Wtv8RggTGiGpZIPp7UX
dWZmHFtBMsli7azy/+V8oWU7qSwrodFdzyxr5fzAthIf6zZpk7ZTGZqN1jCh+YKmc40+JNUdnKcQ
UQ4cLYcYccC6GK7RAwlbjQpsJg3NMGBk+kB5bIyA/hUfiJC2I/pIcxKF5aIeiLLmPocmzpMDldSv
K2DSpjQkPlP+OMxXzlQ5pcTS9DF0cpMFt839PCTAIskzfpqK19J5R7jChK/0kpg2uo7Zjd+ssi2p
0UZpt2IgZJOu9hWwPBGhCTgllkN6xEU9gc3vjahOlatoWiIf72hoJ9Gjq3elkDSYA32IsCzLaAPk
jkKpvGeJ7YYiQOQojFrMxcOPsCUS32EwNWNIfuytOezZXrWoQWnC/0t6ddOOp/eEQo3iN16k06Em
LUD22lq0Z80AmvlBvQkUOSiKBygUJ5txxLk/CoBMv+pMNNHGnC86AA+nax+OReL/SDbtmQX0VojR
vAuXf7ttj8GMZIp3EIAb6WvDoiyclegvgfo7yLCCWZe97TXBO759UD8XmmA2BnV1ekIVR0AJA0R2
ck4fTCJgdgT9xStxtxHkS5n8I8GJwSjIWZ0/qu3K8uZ5zYFgwphMqKnsfT2vzXsEF+CprwmQ1JF0
vro0WjA5SvoTPaqzgeGx1NEUx/e9mBxm7XWGoMWEVWVqznvnT/GesnMyFXvFA6adCt9jAICsUAfL
9Su0lQhqDylEfrax+phiOo3FQNYGVhow94nqAljq8bMhnyELYVOlxtkOmnl+QAknHFYgM4x9XAvw
Ypph3C9cEeEYSY3t4DLq+qUSMCltS5M90jESaHGMgC/6d8baDsZwuoJkXLFSA9/77vCz8t/lnX1+
etjbwjgkYinNsqmMC56kWcQjvqYlqb3FYPN9WzNiLDkBRa8d5FCV3jEv1c1B2DSO2Q6iW9Eo/lqt
ArMr0uCT+b0z1CPt+UTNktBc3DS/QowvxWdSV+lrBE09Zo+aiKQIE6I942tm6+QVrO1vIhHoAzvp
k1ZbOJDn4htRZu7ShFUHx1lJZMA1+c29XCvo07mGYRH23COaDFN/ZfQVWVAJlvXMrnr/aTMhiksA
YkBWv7P+m3cvvKG07/7KMgQ4pppF6YrHSb4VfIYAF6cDptRPQ1C86QzKOTAwYs5SCQk7vXbUPVLa
ay2MDjyNCMy9UqRDchgadeJ+wT1UcSGqri6rrfb2ZpVljcqpuOugT050XvAUbSeHZzcxo/dzWmm4
5Pu9/CyRER+zGoJZIRUOOZXDtvlOl4Lyvo+gyFmE7vOvGbeWWbYkNCLEg19JLP8T2RZ71HHLX6SY
v/wu+JA4aJtwAMm7eqfT514DJd9df93noEGz4QbVOoOu6Etlu0FDV3heYnz3wCba6cmVWEyhte4l
6RhHtwJdRBHNo4qblW+shCJKt2h4WAP5pjToC9ILLX+3a5epw3QYMstICjBJ4BTdkNuBJXZ00P3r
ca8l+Ku9RNnqkwrP0NZK1WftyTjaxj+zi510l7a2Dqw408FKqBggi7/wx/ESlheFQ3qbLjmFqz0t
h+KPIKrqa2R2A6WitVrW8TveqKAPpysVoivt0EchtTmVdck4FPPKtQ9y6vfAkviEl6OBOViNlY7A
P+/ZyjpUgWGp8935Y5TUDqXM0fPJYV+Mh0QEHAYjiLu7ba5c3uCXGCQKLued5Yn9Z5JrDw72fDjc
MmffQWjwxRKOmw5E1ktRbfsFCkF0dVwMWTbJQn8GwTOK1IE50L5cdSyHaoFqpBVocZutK59c0fJw
y0OF21ycS0BEOcudukaNjB6701TOH1d5FjcPTOgAxEurOJex+B4QBEP9VKgKRszawO+1x9EOUWJm
iN9EavyujgBCMMlsQxsq0z7TVElVaEBbJe3JCZMNZmrL8wzX7VVp5N3ji5Jf/niBrC6Z2MAljAwx
UyGBM8l/ABJqWrOrinanPaCom5qKMREORHQf+3FzQwnZe/ReTFMwsLa7sZC2soBCzToqekpX5u+5
edi26aGee1r+Yt9rsxr+yI/dWk21I4dE7bw0ALSkUGscWDTlFj3Gp9VmSizJ8Qt6Y9mTitzb9meT
jw/bRdowdsRW5RbcxilKWOBosfZye77Q8SN8fxkRCnxYXmd84aFM5346p7Jwioj6vk/1RhyUDWoB
Zgh7GDVODOY09jCGc0u2lpR4s4O4sS/KprwUVa9B1sAhm7QuTXavPWlHmfX3Gxc3lljyBwl5Hm27
Z8I12xHNlmOijHIQ3ye48DZkxLbsusha/1yTaeXm+zQCreT6oyKGQvXYIGyt49I2D9RKei1AfUGO
M/EOfyO+X5n6yoANzw0n51UhpbM+GE6wyug8l/cbE+F1Vr1UMeYD4MyU+KniFPuEJiY5FDHXzs/6
3xEXa1xLWU3YB9jIzQW6f5vlKo914ZzSjYbdZNEaAZkXwm95n3+q7/93piNYOsoK2QomLMaKwgmO
B3b42RGSaNkZrIL6iioyMrd1S4OWcpX7D3aj1UMgcyN2W1Ul8j41Cr+ggOeTHBc3gBronTmBBi1/
MeQ6yGie4Kc+Oj8iiRF8eECc42jhctxnbJgCf9GGS26LIuPWo5MwbCffB+e3wiydvtotjViKifvu
/ePW+dJ7CU2puqF17OVeJQe9C857DJ9doYo8U9fXdfvb5uIehgoeqXUWiXXV8Bbk8TKBMUUX2Epj
biMw3y9vvq2F2IMxjzm0DWTl6LurdHmij3vDpDJog9yCLZ5AzXr7EvApq39X0ByNAOv31q2PdMTO
3xcg04u3NNkIY9C0YWm/6ZxBDkCqgGWvzDQ5yMJWZJyM2lGURTVEYjgo/ONQvKyTrv0eosRKhPTe
8QoSnnFnylrqpWcvVI6oibIQhRZXl/uCWqRGlOUokwX9xlu38kl4ECwSeuArJ4oy6qqqhnsBwbWl
kHNfomk3dCOiMUMReoGp/MTlxg4u4EHyGh35hbRwv6AwYABYpq4xIqIR55lkWlHqqCC6ICTvsRL8
JREHcOuQgJV/AwnEfXacb0yji62+Fqr/gPn/yt86aCnasi+VndXEv6FRVAJCBi7K2kKuWQ5v8VSG
aYokduknnGJh9EmoampzkTI+Z1nSSEtVVFu4HsyeDmb396AYGm4zRQQk5WadhJIdYmyydVWCzuHb
HfE+3/RgRkOh/GG+7k/uuVrjP6vFdTUp4+lcowsmZ8xehvsaO5cQs51Mp2201RNYfU6CVshpoQw6
xPtVF3dmj6SzweLRbx4C+39DUnh+lRGAHzlRVgEyKXSCKj76FXW65AEudjp9f5vkLYkApHgEW+4+
6DgpPSdwu38C9jHf2EFuKiQD0aZfZNtU8rD7Tr8porrYt9EHwAxU6HUSzcvK2CiSkE9ERc5mR93o
n7onK4SJ00SNz4AQRVQXediOMeB/NXg1VP1BTdTGaqCsBTFtm+tVPVjwRBGGxbMuQK8jxnGtfDnq
5YyG95QplU/W5brrebetge5SdonTInX0Co8AnR8xvURoTGbtz0n8352GUXxTRAB4WXQlk0noqyxh
hyGIN2hzrWjnltHR22yqJWI0xuPUHfGNXSsCrIwvEsXcxHJUe5uIgv/bgtGCb5SD0KoGQLUe/EX7
3QmU3m62W+YaRLJfJ4c3GjxCUHWxsyvTaUH6SLJd02lZFUooXPQG/OuDCpynpFK8xinpnvGIYDvJ
SQKY8DV3fDpMXBbHU+HLLWoZVtPFnIIwuJZdbFo2vT/sbK1vS+qBX4zoVsCmS0aGnX+0FF++QAp/
ONkSWNl2K5sL2FKjF2+mBNHPX7MvX4Q4L21SyDdkQDkwOujl3F/nG8ikAENJAQkTUxxfbiADmMlz
KB3wLvHsAUlT1m5ZcJxDC2aVPA0zD25s1jw6cVMjJRVsC/NBx42nfgSxfXalU4LSBFX2WMQ82wdx
ruqvh86bHlmLmVIuCP0AEzW5b1wAutTniKUw4sFOn0tftPLZlGVqGaTvQbLfLVpjsGtW7V8R+Kis
s19eDMhKrouk7qsVngBAbAUZt9L0GYyw0zmPQmh+uWmHn90rSuU7oKpwZI4IaghrtS0XcobH1Chs
sBASjApXy41haPuLhbgR3MGT3QsOwCf5YkfZgKdictbDNHPbkCZ3u5k58I6SJUxCghMqS1mnR3FZ
ag2ZuV9CQRSuGKw5d62n7D7icuN7N33Yu1/E2hLGo5XzilHoW/C0oN3y8tJz/VzwYQunjPvOlR1+
5Uatw59v95mZ/qKNZt5hQc6hU8JTLtM1Tr8gHepa4cgfznGFMas6vOeTU/YZSpQzCzevqjWCZX6m
p1mvjG755vzM0k4PAuSp4qavoI4P/PrT8xMLZJqhfVjmPKmcfgEKr8O2GxM24af0MT690f3drFtE
x11Eh/jUOMhYGSdtFw4viC39GX3oAXwbxxbKueYThmo0TOXaJROjouCMtbnja4FMUKdODLa6hZzM
iwWoIEePDmZ4mvtRZPGK43EZDwHBOEyTZbiPxmUYLZVhb6PWB9q02SoN7ffPe2lnMqCTYKqutqTD
UQgR9uLyvOQhagBqhhcpSmUzYAWnJy2yMHANBIjcuTn/pZuBhboMBEn6sJTjMZfIBQVXk7LDd9fu
iJQBGaC5nddpt6quQYjFUM3Jg5EEJ4VHRY+Cofc98ZizxZ9rGyfPpxMWFATIuoRzNHhhQGwUUu0h
TZBB0J+J6Gxfzed7g840IBaNy/6LuixysSswBc5uo9D83acYjh8LkXBTgIQyal0fxGK1DhvJo6+u
opg4Cgc3DWnw+UMSr4qkZLK2ik4z4Bpg+DwzU9WbwDiN5CftXe+Us/vhDy+VHKbIHrR6UFpsm5C2
/0NB4F2dt9Gh5ayToaDb64uPetvA8bZQnCGDsJ2KJQ1QqaeSJHnywJcaIxm82Pudv/zPY6tOcrmw
XeTYz6YewrEVL54w3bD+TKYiSuz0YaF/OKUwgE3F+21xUkNixodFDWLMMR/sTDrWX3tw+s7jXPNH
PNJx86EJRV+SNA0laJFoVighw1IuaEf3mj0aM9Bc8a+dbRom40IT+llQ/S849z5+UwQ0hF59ZaVL
MXsXV3Tv3zGYXIah8StTalDaGUFuMuRf5yCb8T90DBLzBy/qJxUqBDIjI5SrunTPtVMp+y8jo2XJ
4E9PnDovrUetg2vjgdpPmrlikvIinC5Zc0Nbd+yOAqPECc2+GaJy9Cg5Z+7mkm1/XgfS6PVs+Li4
DGnS3okHR4+6PBkewKLClW2ZmFRJeQa6i3UtxK/VhRiCOapIRFrhK6A/9NiqZEHxDUW7jiWY407a
E6cTM7CY5IJKaH0VEMn2d/N91q6hotVx4VyLda70Drw2ywEt/Qd5VYG6SRChp2Ux3gGL6vjR5/aO
tZXWDBbAZ4amKzIPv5Rc7jlxGBfX0I20dV8vT5Pz7r0MLpq1Z4EjaO3Ecg4QpM89Z++/kAulQh83
WRyDx3EdLpw3ZHlHKftmSy5fziYbZ6VYkOZUdiS5oXg8EtksEVpZpxkQS2x/gmDT5LZIEVtbwUdn
xtnf6aQieDAM3BN9H3HghWs40pcLI48ma9SIG6yqYZAi46UbnpvfVeU7SaAypV7ic7Bz5TTzYQFo
9vJVqmPPJPRizAWqFCa9usMNpu6nIDFVkr0Ad2c8JDSSmki/YrH7dJ+HqZCvgcWnv6CWCvHMkHTA
KV0hjXLhxwpzT8JusiKoWsNWtNQbuGkholaQNrBKtO5utY5oHr8Mvx9Hf8EbldF1XTU9DMA0lB4T
2RDk9OBERBhDIefB7UegbSIHFZo27mjDo7zaXsNYWCBeMEYiZ8PLKa9egVsJsXQOcWGA0ZXExoJU
qKIsuwCRZ2Fs2KA1CrsjoCuuaFLUe8F9/44dDhncdJoErsunBfgNvwEkF8YZv7nEL65U92OTw5+P
ZSsh1/aVve0DJL0xCwY1RsciMYPmC5PzopR84QJnSj4El2zqQvcWvDFZ2xO0w6nH4Nf3PSwrYjza
LxGRgv5XYNl1OrWWyMIrQeemGMYdeyqyHgyGmojBSGSvouTpqkyRkg3HTf9Uzmoi2EkAd0Swi13x
36lscNB/1WobIH6RU/ELFW+U5hBYr9vb8w0SS9YN38pBpdSQy1opb7BlAyNa3Y82kjwSWSdYAAF+
f0eRL7uhJJr8xayhSYVbstYd+xrowT4nCmqrYczyWv4zUjxjuh9r80B0pzw5hxVVI1QTmlHVbLp0
A+SMWatPBWdEJf5t0WlTg8ZDhGaUwYxDT6kzsuxlsCbK3KVL+TyuIj9eBaemd542810leab6bhR7
Z7sHII7Ay2Kg7CiVqjUK33NevaTi0Gho3dN+qjrkTBc1OxeggCq+xDTOJ5Ukcuhw61FriwOGeuj8
d6gUnJduiUuJMg/gLeDUfMMuC2mCHAZlGG2Az/GgpuTV7aekFFnsYSPyO2QUqDo9jYfoTVuLj7l4
F7Kpn5N9wtyY2o9/0JZxe1q1rrecH0a1B9NmSYPlAxYIgg8w+0bK9Db5CzN3mbNpzgGyv93rv3Rt
z/dxZ5ML7BBJlNHohJyS5ILxYfR1t1g/Ht2h7Y64Fs1xjS0YkC1mn0NrLQ+zegPGeVBiplZRwkEb
P6YRHWN2jjnNw5rvYp23MbRzNHXtmTywBRhhBJrm0XewybH7vVVd4Ej/N3OLmLcm4HKbtg0J8NpR
ECp9aj6WZlecocrtH+3gGJPXeHh59ZFjANev8nNm62iiWt/7g152wT+UQfo7lEKbmykJQfmpiIeu
B04vdb8dWCXRJ4NsfnXPbT6LF5a8/qD+h7vgvf9F4mm4xSU57pj17pf1A/dKofLuYlAaxKnbM7Js
JtVjAYECYM7n+d2tkq7MCN3keE/5xh4KttWCbUNHBLDtS7vPzAf+wJMSXVjV5Fg8xq1nE2IQNlCM
XobGokFFWCFsXApoppRdVWVz04smzEO0wW6kHdzSTVuW97EMSu1/CcgURrQNqc0++cSG4KLbgB0c
1It0hUUkDF0AAUleCnABiKX4Vkfo+ItsJHDHv/eyJ4fmoUNRlWwCLDlKPwF+NfXbzYAot8uQncie
fcOjvWgaeeIuL2mmIEf6oQp4isp8FQwqf8oV6Sn7U8wv8TP/m0uoBGTZ83OeccKWDaPfp07Ysg2O
6wmfeT/j3gHwghSMuNlr8DjtyhFcojbpljTbOjA7o2Nugf3cXoc+xs763KOw6bREv54ZPFylqg41
0U43Odn7h4FfUwiiGgOl6X6luc+v0m2++ccNeFn/eAsE/9T0TlBNaAtbPwVXo4V+1aVNEBVFgcbJ
Qi4G65FRy7P084+EvgckWTeOCzt73tvia5svlCN3Et9wJ/C1TYABzToBwP+NSo4oYMF9LdBPCbgp
miyeF2oxxVD441QWodYuH+k325LgDYtcZ/EtbGeDMjFDWZZi9lMALQIqSrFRTT8dedO3Wkj/0f8/
bxT3cI4k2pKwXtBiiPn/Sm9rSSkHVzh15f/qOBFSM/a0Bvun1RT+wRT3rdEs60Ah6QQBJAh6DX3i
rF8S9vNvrDACwsMqN4uXR/BVTNoS0ydKcrn3GK1gBqqfRjO6eR/36U3UUZl0RXze9Ysp9M1OgGGW
bKD6IbDYcb9xLjL29E2lZNv5KYNBpBlF2Xymi0shckxwHGu5bVtTqyyVvFJ+qBRpqpadwzaTbAYp
xzqqm0FwR4WGmNcIKqsE9QbKECjacTMUwcDMqz2zkV8sDiCsVUTcYPuLOfzGKyGpZlVscghIKtjg
31TALGEIbnmHGx0uTlww5gPtUPVibtGFNgxIeTw6k45G2nW+d1ZZNNcXQK/qLGFvBGLUK8Ub3SHe
ABvLKrXa6+Dd5lKYfdjNEGVjiCUzGEXQz70WNdqNQ4X+Z8DwUQlY8SN+E6KlV6E+Xv70+CtsKaOw
X3/T3IAvMapIT2dORcKKnwErgpE052yPzRcta9Pm/vZ3GyuVYBCWfJbj6rn4CX7Kc2XezNvJJPhM
CKepJaBIFKoX7T1BrzA24u3oxcPjFX/dMKdan3b6mzVN4Tof70O++ZPuwn7UTzApsn/mbARlXFC+
+SUTkaPG9BSmyb3nkXsc9TLysGx0d3XjLOhDi81WVpP1sUj3LZGP13Q4ptFg7V14xbLWcnSDPU6q
amRfkvaIAcNasQtWc1C+pi76aMMhOG/B/JBrGxxCJsYEp56hyRiig7v4YOuFzdlbhRwnvRCiX7wT
z1qLRYVajUCXaFallVGE7RbcxDMfDmgM7iWkzqDXBI2a6K7fnLSoJcIYDWz4YSDWcDacx7lXACRR
MdZaAILzlvZZbghoYD5uw/whAUxm9utRshiudzovfGoPfVDaZ4ocBWHIBwBq/Or/29tG+iqZFOK+
T/DUDcdJ/PBBFN3YsOplWeHqE5PSRm2swGaofKHMED+gmH7hl9FCSK0f+zuMs7GuXiGBsmnmrUU8
si69B7AQc81LRXgDAKK7O8KO8HkT3VrdmfWmV6Q4uDPz9mhOpRFKGBwnkHF7r19JoGprzoQQyq4o
ttUjHVZRdNpTlmnnouW1V8tEtxF/n8+qc2tQxjA98RWcu6reBjuxudtStdk7OswdupJlSf0n0bKL
k4FTugZmo4Lg0rehK6wXs+2XDZLhdk5TI0F5KwdToFRo4XZ6M/sOsBqIaRd+ZyFO1uA9S5aie+a0
YPpfo7G1zUROAiT/ywqKbmJCC4PBImWU6fSpQaDPVtSeaxYk9t/t2H5fGD1YmmYs9LOpGx6492KA
5SYHT/FncTJh9QtHYBeN0D6LDWBZoKhdeQg+xsOsHNWwgzFN1lQHDCkV6aKhH3TY0TrA/RCkW8qy
OvVYIXH8IToKU63cLVWVs3Q+v+vpPyGsrMYkZ75kM4kM1X6cXfMRFB43qg02cku76x4nVnOugQWy
7YOXPbMucyRBQgJifBuXkbx82ptCHvCQIphcEB6BaCqhbK1aoYyOrW0OuCmH6J1ioinccReNlrb+
UYO8KTNAX+I+/2kqJ6wLfdAFfEMzBZiStD0l76WMs2RtNprayI7IBCEB0dvUV1ggrqOY9zOrlJsO
/i7UrW0lnw/nQ7kMCU2yI1TqMPGCG0KYzDwpq4tUNNLIh2qjdlaijPaDbMlf4N606ogE8ucefVAs
xFwCrIthQ6jP6ZRLw0x51H9pg1c3N5FJUnumysw98tD8UnNBQxCJM2bm01jzF0maiBYmH+/D2i6I
unRPO6n8Nfa1Q08a6mCdsqz9MX+HuFP+ifwboedhI7VXG9pYLs4DxrgzAps2xMs7E1BsuTTf4wpq
TFPK6WvWFpuYzCkFCXSzC14IAQ9k5f9ibd69uQu/SvhfVLKntX2pXJo1KNyRIiOaBtBtygKOUqnU
9CBMbsonovhzx3w83mHBTsD4ZIij0BnKI2ABTWe2oBcGbVt7opqLHRS+OSfMoRX+QaaDyZl4MKwA
rm5P2BYBkLyedmznyadXvGjDlQxDL9sfqendvFQFcYWRIBZHxztT3AklbA/vEDa9zcF5A1Nv/S21
lZgalSWtvbhjr8n9WUFcM1uyG/PNSU8QSbR9DFf4ikY1are3ePtsmbs4bQ6u5wt6Mid/L6LuoRmm
tvraN4dPP81m0eKQWTP8Uyom9FWQlkJW1To3jra+2gTOdB7POn4ivK6uQjtz/azwwRcPsY6wrgVB
TIiOdWIbHayY6IbmKirdLAb/tCWePaeQyfHzPgVkuPL/H8uJkcpmQxULnzLBSJmwC4+yQzhnWMmC
sw1+H7pe38+zEz93c5wpd9rm9F380zrexue3EpV2sIXV/c6peB0TmBPkEmHB/BPafDsCSXQ8thKp
OImX41Y2zBAsl9Bc/DL90YSDE4jcmXc0o2UsokhRJh8bViVao3QzO3LhPd4rNnJt1qGyXVVrEcvp
zVm7caz9Na/vBfA/IKLWdqpV4cgauPhAm1yqG0YRMIyrk37f3NtqIMLFgdMXh5O1DazwVlvnJIpp
iu/A5kGUVhV2paWWTS94IdE0IxSoxzKi8YbSJkSnymbNe9wzn2YmFBVFliFIy7TnOKXkvgJuYRvj
3hSEd11EFb+0IedAHn0+SPdNkYkCWEVZTSx5VVfDis4RT0b5CiVJ7DKmJl+SBL5NULgBWS0mu/bV
Y5d0teq48SKb2LyExNxnoFAUZfNKn/rwpHh5BhfXH1VwaUKI/MuPT2Gk2SfwSl/HEVf3WP607H0k
//3xB+MPVeGT99WrtEGtqICNo2XnRhWEBSsjypEEPYuHiRYNIUtiohUgx0wR1ItmAW6cVU6ZVI3w
xxCenVA/HzmGbVkgBL3cwZU5ADJTtB+47qEO6bVKTVQuD/hTvvmW4QiOv7yiw//6c5u81vvLUlJv
BRqCWiUG8RCcSo+wwoHlvo6Z7goqdoIBhITum7y9MNJjocpUPrCSZKrJelOVtJ0e7B/8JGV0MtHJ
LrkDcUpDRXnQ3QJS57fs503GiB3jgJfsJHxAre8k/z6kc38+8t6POcap6bGpDw5aKPfxVEovuy6O
es0oBBVBqqpzqG5bWkVuvkNmIF2jnfdsnBSw/G0cw6UFu/Dbyb/cBZ5xFu+hjsWzoZPmqcDTBSEi
DnIG8U4gF255xlAcFqTHUoEp6uZEmo3oNBAbanzuf3t4MItha5Ved0Cvv303vAMqdG6bGVTUupdc
MKGz7qgpEuhulFO3q0mfMavLBChibQZkV41qShig0KMXdvtZbxcoW4s6tc6F5L54YPzMHiF4Dso6
ExGqkINI7Y72O8WjPSiwDb1fW2RTIY3/lQeu0omBZddwx3cTKmwQp2DOpRjwx6zC7hJxEgWPwLvc
x5jkGcLV4ttpZDZYPENC7j+M1Ay7gBnGYdhEaPDRnnda0JXIeOiL2oQykBGKG39VsETin/oQHPAu
Kh8Sp5cH09PSdtmqm/KKatyFOHoR3JB1YZ/8Km51DKVM9lKGFqDB4l04doEe/ryzSWAz6y0kU2LM
mWLm6Ti5w9aHwvAiuJfHa7wkGhjecqkM2TYKEZ7+lpIVPinTu5WkUMqfGaKKYyll+0HKQLd8H9/L
FBarM0rcAupLKiaRgQ6moOHqtsVVch/HumXSulYwIgV5XBXoRsDY6AMYEmLgA8aQqRSJ8ryjFV9g
qgDMmfDEhSm24zxLhb+WiHHwgQaMUUR0+PGKV2r26xs3BiB6PMwbXXnMXf5E+2n8D0w4diG7jMoc
EgKs+Zri1uUaXfPsdON5FcjbWIOvqtYsULxD8W/+lQAZW8wxl/602WQ6HhzLlvDdHFaHdUE2ZNGR
Hp6DqFcjSLGpMjXkrjan8xWZePIIGCFO2r0E9nOuj6N4zIa961BrgyM6WenpRxvXXWuqZ0jvGqCu
Q3wZgekwQC76xtOKzPDdScSeyXUu5PcHu01a8p/qJJdD+OVoKIJZU0FLIhOHd7MrXCPbzpcUfVem
Fd97fKztl+RvKZgYKMk1mxjLUfAnpZiB6m2iqn7JwnLJZTgEsUD5zllCFMVvw8gVxgcnflc2ivG3
3SMzxrTLYwEFxRQyDv5Up60w2DycshsOrHpf/0Qx1lJMyjq6NxKZ03a0twCqaeRw81xNcPKIF+Lg
f42Ag9RPq561WvZ2BD8TTrZQ3LjnaJHxf6l5O/c+8pEAV80+VgfRTwhE8qtzINlgYy+JQ7i/97Cu
2dfpmWoFQri2T7x8wM8rnjuORGKNvxLVSveuOqbxUO/Xhpw8QsGfK8dX/qNo07X6op46r0bLlQU0
bpQ4QpEKDMQ4DSEEELx6Ula1FTpTaxCy31uU3IsWGG1Y4WEY50SJXo7sUidqy6Yo4jA2vveA8QFC
/k+EhgLtQ+Wrj9ZLXaXsgQguoElB5aflaAxz8WmqNoGy0Qt3RcnSlMFNvUHNUNy6SH7ATtfKV94d
bZLg6IyVfkLr2s50//vXJVy0LVYzvabCeIWQjspy/61Cd9Him1nr87MXLJsPt049Qb5Qn1Qf96TA
agOMLm8BiYToxXOBxsvUbsA6tk3zH9atWXQWYCnamPTwweWvjkKIL6JmQb0qYq1qL5Z4dJ1SU3Ru
eSs3YfNb+r2P6s/XWLWpTZILJNX2Ws7yWJjD9TTIr2cMRZitpUGtQpIU0HUe6kHuQrkWZaoQydTo
zac2VC4ALTgIAGLMyG8GzzROGUCVas90HkzRsVQJLAVzhAc9oPzbksUOVv8xoN+C9YwxCxoWUaFv
iZQuzs5utlgaMQaYeOwe4s4wbZ3FxyH/JR0OrV3EnoBOrjaFUaBGpxeHAWJCG8zN/9P0t11L+yvU
D1cpWJJNJ1iuRi04RnE2hw3b1IAchNmGYdvGbpat3RymbQQeK43sINF5ZG6iudQxYXFsFLKZCThX
KvIyVyfTWsyIrRXGtE91cSEJXZDFEtoNdxwwkDMIkBKmETZAjd0FdUXIvd4Z/ynWdWI04sxynFh5
UvupS+qsQDC1a2yV8ETBLqdEPWdGEilxbVi7TUpT+IhMeH2rvbgsfgD5BbvvyoAtDR/TpsFl/R7Y
GnhyrgYFgiMmVz5ffCuCyu72rfuB77EH1HztWEq0JUmPAmNM1jGE/0riP6RZWWlTJkIFPaKMIhJF
B+GLfIWjbTo6VR7jKLINGCpCvKICdVxaBTnhkfUCsYmsQ+GfYz9ukMFwvf0+Umx1Mkw/ql9exIKu
68jAUrOyJjq2rmbHBTDpdbfzgXaZrROZdIRxvHidC6yvkazapPn4AXhM7fGTLZQ0oe2fzmAKkxdS
JobAUL10y4c3COIPdwHhbBV9TC+UBdksZSYjAf84HOHk+9OklIl3yRERm8LUUWnmP1FRZlC3D/O3
QvLWuXpb5xRgFChL6GgBcGFJmplTsKUfekcLeVwEeZl/iuhO5ejTCSgTCRdYPSJjQ1HEfH18K5sq
3OeZnLsu3JNd2hKLEa7MM5841mPA6bEz2FG5FX7zHoxsGH9ivm0Drj0TlJGibN9zXn8gqIrk5pIM
VzEILEmiZx7fbbRK9u5akthahVmMe1pQX9QhnJpEM3M2RZaYpXG6sQVe/QtPFS8jf2UIrQD3ku83
rhpmE/Fo6sEcBbO/XhEklqUaKTneAxUpbeijex5UuHO+clWSuXKydlXJpx1MNB+w/ALAiREXZC63
5fx3qm0HApSHZtEK+Q/7po+t89+UGiz/9zMiwPlpbvEEVYEKxTMtFGYQfmKfrwGZ7pEFZ5qK0Mw4
ckU++99Uov+YA+Q+jVmD5pFIrr8KUqrKY/r/31uMvrgyj79CbIzIk9eErfZrvdTR/d2tpeL2pVPK
DdHzvk+bWeNA/Le64rLa7m0HlWdWXc0Vgf8AF4EbY5XSq3H2QX1G0O0LhBWLCFHkqmng+3rEzMnM
jICti994Grfps33SpPXhYUd4db2z440JM92gKgEb8Vap2cbuFp51u1I2zS0IgcEJ4UBVsvqmClvR
s+lUmTwkjHcFFq2Pg5IAsBwdDwe3IjK3Ypi2BEYFEZR3xEkwdbG5QFZrSDB1XGLfPgaQ0TGl4A2l
hePmrk7Rw1f8I+fVIH4fiuOI9YD7U1vl2CR5YUfZfFrsZiE05Kb8FpHcMCf7XG22/DBalE3EWnEM
tekdk9hyZRsl7kFEoEPzKywuSmROf37Ziy34rhqCcESBuWcUnpGTO1gCxuML4elX4XGVJ4KwQajO
zxiO8PRJTBMAL5aTaCL0QJrzfDj3trzWkjqOB4KlIBAlLg1Vh0mJgE99E5gDKtcsQL3/qvPuLccH
GT4pSFHmlQuEVks5e3UJ/WdmeKs+2ywdR4/3vMu9yVh3nX4NkYdSDd19wzry7ZcNhgCyqpAS5SlN
r6xWTHTpT0N/t6k+AWSyu87ru0JqL5y8duuRLWYvDcowiftzCpLnqWDf8YN6IEqPnSl+qbctAnam
d6ucfNatacKNTIdh1tV4TIZz/V58OHU2QF0xVNa/ciYatXY/O8WDcSvAly/kpgkcTzB8fW1rf0fl
MGiLcmwjuQI1xXISLSwqHsNGdycdHtOZh4bRscEGqPdtBz6XilNaLs+bOP44rrjCS5hQ7y8EwBRa
jW5tMTlaFY0XPC+qnEu8ylp8U/oj0d/UAr7kHsbxNqgtev+fAhbRxExYJkoScDPJLUhOJQPZpZUY
9Qk9Iq9Fpz+knodry5OWz4dbh/P4Fp97OcZ2g+FV6SfT3Vf8mN5SqhQjud+SzS2CKY5dmGUfjatk
D35vvjN0q0z57sWCs+VY2UbPcOcY6R2fUmTdf9OxxS37y9VoZeNWWnV3Q8yhB/oxgcw8qhTy4c6I
N5vwWBrkGnhGTdMZ9pN1tTlcA8xhCIx4GekJTZ9+xYXdzWVFmb5/Jw+imPXSAIqsqx5A0Jpv08aB
RflsgsfH7hyaoU/tCez3zT14Ip4lpQcGla3qKqt5f9mlc6Ka3EdRvo+aL4s+Pq/5VwRZJ6m8yep8
V7jEdpogKYpow6cbPeD7/UDjexFR4vdW7r73vHQ83qOZMYXDyQfQ79nAL3j8X3oTZDK5Ahh/OSlu
xU8WGlau+2em+4bwKY9aqkVEF9TFukAPywpGW9XwJN6WKz+3Wk8+vJDXsEJuw0nZIHPYYt8LZloI
yL1dQePPayep3rksQp8fTjYSIRb6p2pL8WquNABexaALgcubbegYdcYHPmnWq0ZogyPcXdQa6YM+
Y6wCIJWZOklQNUkdv7XqGtpFVUrrLyhKnX5KB/8ILCRFnVPkCr/uxB/yWdYNeDuVKWT6+pYeQcXs
8eiNkBXyc0aAa14EfCQWFKOOX0FUIXJxZTfCJfIzykMDGRb1I73HuKq3nZ91o6rwY+HNrR8ryxrV
vvP1+bijPmTYWCp1Il8+HZ7+vanKipyf4TmejtPcwM72VOuYksr2kmEXJ7dfwliNVT0dOwAh3+Jf
1/D/OfRvmrVwFc5WnlfJJVoAWTW9Vt7PJTA5Q9xsrFnZP7Rbe0hhou/AQZhkKxVQHH14xMwGC+CW
RILJycaKuCSyYzI7rofpkDbj3lM6RlRIZAwCenc/ZEVpl14yFcJ59maI4BH74YpkUqavHsczGfuV
+yMnK/f2VjwQV9sRqZxYeK5lOrCPY4+ryG5nEic0l8x1jL/HHQ9gbgLQ214Pkr4CLEckY5XyFzEM
baw9vRbVnroem9AIohh1CEdN3dnXFOOnMvxpwFWPxcRDOlZy5h0LBFq+TlW2nqYFBPKthiSMR37z
vWmRpZrW4VHX6bOFe3OUNqNX/bOmtYyvygglLRPV2cH1F5r4xX7h/W5w6qESjI3WpcWqRvOXg+1p
ShESP2Gwoef5fmtzFfryw3xnS727ayarHq2AiYeVJdiCEeVqTqGxC410Pv5x+q24PcdFnKiXtB4d
EYj+sxgLUR4QeeDkWYOs/wH5ivhOfKgV8qb/lGF5bX6UxtYiPv65jEg0m1oACR6gBDlpXNY0JASf
B+a17YD/AN2iZ5ncNMf6rkBV7PtasPkMMPWG3F2swozFYdD+oDYTwvy1J9M49uiMinWkx/Q89MVH
Y6zv37a9cuKZ40xengF0/RslrzHdKkTeB9ay4UA+dSR5rh4D2j/X63iU9aaJg5XZqmCdC5HZDsrB
3x5RhsHeUVpHMu20P4SmGnLa35qnezh0v8UCXpbSDdaS9GX5EeqU79OFMphUaIBKiE6FlJZ3yssq
jzgLloBhvHcVIkv0zM32j7CMmgp/Qo5xb8MiItGFcqqHVBP9R8ABf1Sqocd0LHPd38eQHq3TZJ/G
3mjeHcqNMtGdIzOiXRN62aR3HleZ7PXnP052+ioV6vix+SesPfKcw0WGkCAPvd74QXZNI1hfy8c9
cM5GMZNyCiIKJ02+3abDo4W9RPog+KUYcQPZ869SBt9d/qbtqzQIXDH8Ak8SyFwdMAu9aGdTb8PN
u43qoRLWYNYX9roFKJHZFrhLx6eiqoKGlbfw2s6pcSB9VEqocD3ASyPCS77AoBZSxtuf+NYF7YYy
ZovUkAldigWeUdhHW9u+T+vs9taJXz4y139Jr2WFG1cNWz2o7mzIN5sF+lpXafvyIfEgTAKcRJjQ
QnUMIyNwM+b+cjc5Ui5c9/Mi42IttUiqCsIGJF3wLMo3ID8E/bdxbm5s/pP8Cjhr2CWagEgBiNM8
FRYgdTclShI8m+uA1fKULg+EnNqVA+UFzZujjGEVe9K+9RECKK5pWokFvXQ9FdMYaqfLE7Kw3tdd
JXFZhc9H5aw+qI9qtmubkmpybiol514+DPRZXu7N7TTx8jXNx9/wjFQEy0trUVWySNEqtwVh3i4i
kNn+NUDO73gU95QhY0wUfU5TJ47lBOeL1BMZTyVxfW8DgVo5RSqMt4ZKXJwoW3D678Nl5qNd8iEF
7D9qDENE105xvC+ZGXB9HLL+HUy44Fiq0pzIGAS8j3eVCWghHWaZ+BCcEKwaHCoJe0prOEaQV4n3
8oRrm90zgPYbcMt29bt9yQjt4FEkVZy0kedO4BNIbb4xAOkTXFh+J7HStl3q2R6Q5+Fiyg11tmqO
hl9SIxTDmdAFv46FS5VZyMuGY46gFz/+3rheKgvI8+O3zQXzVV/nnPyCmGMaBbWpocTJAqF34URz
LwQOwQi0cOuw2OLOAkvi3QO85VWOxHxRP8duQruAB7ZsaBvUAmSug75yrDXnQxer/RwN87kHWZJ9
lUwRuKjmYexixIcnoKzjT81bxXt4Rs47lAp3XGBVoAgi3t61ecI4P1F9TAvMGJRRjf00sHhRPM75
mVc+o0izLbtrjLvm4UKlogmWPGwYB3/mkHFPnuu7KK0GZIr+lC0T7SKQLNPMe4jAByWVvD16jilN
YXStj99HZxkpw7rcdqGrflDaPB2qntkPLimLeHnlAwuTXMADh0ETrga0hdOkmfjomg4WiB4yNASW
g5xC7stxdebWf46clHgjlvFjjZ31mGerJVuv3GCIFWdWFLs4dUPc95rL942uXBmRu67vaZ2rkuw0
wDcXhHq3eDisLeuVZNoJMAXpaJM0Kh3hOd8ABlhhR2q3IE0trkUb+6YlpsulCUOjBvR+QlXftnT8
COWOOQeI/ZqVBTi+3HEzMEquO26uv/zvqDrEYwcKdSNjvhRVc5NXz5QIe6DEsdU1KvQUYWzo8uDR
vB8XAlnG4RzEhXKtLe/NYH5eXmiOMEW4gWRDf95M0V/rI+YlJR7YQEMP5oR6ApfOg9+lwm/v6eXm
odMi1o3XlPmCZI7J+Y2+kEENBMh3NxdPRRKbFY9yNmRWpvra2sNRYsMNZ5uCoTKMJv2qVyeS1Fpy
7GV4MeNX6hlC/jCN8MOA6fxt8N+zXSeAlxW7TRCixA4hVd2jubS9+gpRPQ3se9BS4YNn4nulz2/q
3R7o2WC0nrYTZCHXbWcjSq1ZR3NjgqnZdBrhtZu4j8Ep0ghMmayAk8nreqsOUJ1Id/xL2jWDm59M
hoCHzUyyXIja4xWUHYETZavviN4Y8vsZVPy3q2rF2Aotiw4Ow09cALnHPDA1SCrnnTM9q/69nRSo
3KsKoiXjS6n37XT6097veqza27lOOjLxxrkBLiCL1W+Gndqac29UQ/BZOFldcTsWlhxRPWt0ROJB
kk3IFamfemm3DkRsl4FiIX+JdtrGX0xylwNcE65NZrE9mhQLaWFmTSxAPlXsvpKoR9Og+vSpE8CB
VPA/12yrCdMxRcYiNi0khQ8b4KDjMQpaNXANxCrVOW+/bDFIKvOwNMCaCJJbnbgG3Ua5qOdhL7nw
OjeVj4SEXJ8SWL7xa0pIQHVi2w7ObiEp5G0NuuwIif4d//vGlIwXBR3TuAr/oNIOU8+AovkkvUFL
blSoK4SJ5g3y5bNPoItrQaA5R0yEmGSFJpia5BZzhZOygHJRr+0JQjklrTjy9sGuRz4V/nL9pucH
OkVJ1RAt9goilCL5q/vbd7tb3AZTHjjJeGZxCBH2+zdlULKCzXWFcZTI2d245COlJJYL0OohI5fj
5ponlkT4XoYDNXtJIaiMlNNMJMumptFyEgltcC8JrX6zY+D7d4B9dOA1JrR6sb8B3PReRjJX2XIa
Zwp8mc1m/WlSt1mHgO+b+YVlEelwc6Rlh8NQ9LGfwSK/Xq9LFHPxYPUjtwOLuCHJq6aQDzs6f+7u
ViE4r5ysUwsW5MgYbzdHJZoafTczs6dlUNpVTMYBQDJbf08imnnDaIOYVz0zx5robHBBSg9U1nCp
C0Xg61Q362ZHyq70kKZ3rK3ixZnWEwYy0VGPXhGdVFXnqoCrNJLJd0ZsfC//vA+McNLO8wz0wR6E
GeEzOVTkuTiIF27/wRH6aMK13gAPHuLglH/6HXN230ctpxA5FF4XWwxs1Hh8bE7oDdf6KDfTeD0B
6bRXPc2jIANU+hlSEVprDxz60ncTie+9AU6+J89d7VAhg+AOetnQLPKaq6Oka5BtH7SwqmB3MVLE
iBCVm2oX8/7zLZEwMM7MhjNdWw9fup6GQIKQcKi8OeK049KtX1l9vq/nn1M0FbMSFAeXjkpXHlQm
2TJz5Y4w4F+1JJWYsQIM4/fukmCAEqyjzeNOomRdAGbaV3u3bIejHJxeiL1WG7v3wHepC/JeiMxx
bbRQ1E0Rl3ZnxbYKAbpWnBWqdUdhK0Mu71WPhVs8b4GtBApwvpRa3OJSu/rhUjB22lgi9E/PGDJR
znut9ztyItugSn1v9EJU7JxbplcLKTH6V8hY2qG6TZus6vBKKhyQ4cA21rlTNQbrr/q6Bb18lwSJ
44CM7qCeRfy56pXppYJfmjnu0Ssm61gNAHRxfLDGJrEufomjuqVboNc9AJvqJx63jILg3pUdMthm
lDfE2bKt8Z82NWRWtVV86/DDj1/EZ+70881qnIZnfCqEQxYRon/GvR+WHL2C0g9EyceMOWq+KkSb
tYckfHjsD445mpIPo1rNlte35Szyud7wa/iPlrDHhvE/8JfLIVmF7TTm1bipyFlM58zMuPM2KUp2
i0XBliRTFY7ip2xOXto52He9muTmYhZx04Qg4tnh2Rbm6yDQWRUURo1PhGsnQjTpjSF3ysuGSVOq
FaVvjst8JPwppSVnGPEviqculIueAAyG1oBFDxslQVup8+ytqYwTjkeUh2et6XUCEApLqVbsyRdC
ZqjXYIRDIN+zjqwO3nB6Wz3JwG6+ZOj02xHNK8DZeMu/pkDC+5vGMnm565hnF5/oAs4Wb1xJgLkB
FYxBGqP2JVpf937hGhuL5n7y2vEGkXqRA8tugBAwOwVyNgR3V3ljPnk/HnnLZIOno7aABIYZTkDV
6Qohkyy0fSazdOzI1RmnFxyD7Qqi7j5fVE/73V7/9t0+eLq6gNjvyPzbgeqJhDeqFsdp8kJptp0x
P4As1FxsMBahfRwwTeicDHVz+88UmUQvjsl9zdT2x6lsBtAG6UBithIB0bCcZ+8j51fCh0CFn5Wg
rU7NgdQ6u4sZEed9WhPWYBSWYt44vPdT6w0cxNxitfrqyqOGqWusWuJ013DHQjntAyw7i9czxC9y
o60zoRI+zzICq0tntdFKbmSNwguP6ZIy1QZfFprEPKj+sqwbqS6uULNpiNzHp8ARI/CV2CWxqmhe
rt4NeRyLJCwEljTnlLJFWUlHoEaqe0qzN904BYTb2kxS3gdeVQAE/huHMp+ilk6OHgepXuRIdj7T
BcZbfMUV5MBpp1d6t2d85JJuejDFDzYx/Bc3jnVsjuTey6EplDH0Swr7+bi7j80jKQLhTQunLH7L
bsSs84f6vUm2ZkFMGpKdeHdXX509snfyyepLwC8Iz32ukh/UseE4IHBIIqpBulwNwQKGXfgowwpX
133AP+mdpfs01xC6GRBzM1YjMbzR2LDYDAsryv9imbgRtYgvYf6PxpIae7iHWvcRlz3vPg6gz2gr
881zMmJ1FQ8SjRpMycz6j3QGidlL1KJpQYoi7vR8eP5VuFmos5QM1ZQAch09ZH2NcIF0cvqwaAkF
Ew3nduOyqmZyLHCoV54vm9w7JMox7FXwTTVmSN6b+mCb0AuyIWOY9WHLdPso/eNHvbfCWfO8NAAd
vK6u8NCOGIkjt8GLLXdn9uEkyUEnaHBx1uNCGtasFe3Omkl9ejvGZx7D6HbdnPjF+jESoI224kiC
YZ48DC0pZ0JyR5oyoQMT9oLuaQL5wYEy+PADTdp4IoxgEBD7Ig4BVkVS2tXPpR27svTEnU/lLu5C
izkh98abT0iKtVznJEKC4ovJJlUQ5mmOzuFmUVqzF3RoX3d7dhT2OWBqpRbcGqt7fsUZ1sZm5B4g
IFtWEgNhYJrFtGNMKYHaBqLF2O3PwZ1bDYYFtNio/mGHj9M1//iOQdsv7ztkyaL/stJBPdnItBS1
Jqv1ZkqJO7nTsgfFcoTCM/pHx7d8uwhVUHXbh01DacAS7/sbqGOGWtR6nQgr555rpPQ5uhH4Z3Xt
BAaOG17pkImjSQo1Yg9nQA5JpYtxkXVrZ+lEnEJK11Qxd+khlTfEcFHTZymts4DIWvleFlngjvqf
OuZsqZnIhiXODFEIx8aTwFDeLBNJa9PhVnWMRITvj5C8shHx5Vy5G5FmnEhygogqPBonEpSXztlw
vCOVS17RItnyXEx083r3zY0/PzfAlQbynBBVNfpSu+TwCZNFF5E55NkXEUKNihHti/c9huECBd3D
9PaFH3KTgp1dG6mmnjglPD5pb4gLbEzCY4/wwP81MUHXsWdXKlmU8vryGTPzYmwnBsbauYgds7/Y
a9Lo3nloQ5Iyfco5n5zNI/lBXKCxPpj9unJSVFLxB8Rix2rFRg7FlIArYouUXxPqdkUVdqfDjnrK
gQsr4UCsVVoYi+/3f0cLrwDHJEhEJb6wxq5o/eogF7BfWOTRpmH9gOq9Gfjszpn9alecz+lt8ZWW
4vQgZcE6ZOR+h3b1m1xQNLrluA9/mCrjigrXzvC2S7Vzoy3iO8fUHLs/wMQum5WNgy+gRCW0Av62
LK3BLYWYEYnrB2/D/YFTV3SqLx3FVTEF5g/jZ0/4GMPyGS4I5/L+TKDMpOYCCQyJie1QeI2JeBfw
qAuJHSqHWgsZM94BvPEWA9nsX0xt9IKj9bNYdA6jIN4lx6cRZKveG3QjvrD+cQDn6zEn3yOKSjoP
eYQSRrWa8F2LqVum9cN4SsqlaUCc8WQmhOnmatSquQZ0wt94BE4zD5uNcBeMJSv6Cf6jOpxH2izG
VJmWvslNiA2baWCzfDJkRet86Zf/Q68n6sMF+uhyrXJtjtYr/Gq7RKNVuIZHUel1iiQM091hHC4p
+LXkTbPWFPHENbC3yMaL5nHfej521PrzctYHOAeNGOurS2Z0cY82pFPf/CtympbDXw/fn0SlI/Kk
X0L5vkRVD5kUkaqspfIIxiboZ5oTcCIWhubQP6JDrtm7apWeizhOuSKFlzaFkQar8/Jt5I1+umq4
9lOJFMU0jRys6uwt9Wi9AHOnmBUqw9HsBK0rAK0f2rDIEMGj9UM1gBnNmMEjIfkgKbnmkQHczf4N
gl9IgzMY2OYeAqu1ENCC3q6QoGZBDDrf5KlAXPGwbtz0O3GgoNkVzbrUmozM9ltk/N8fLOH0XuRn
Kf4a7vJmPXTZqjvb3t7S82ZLUuCqmmESyZSWZKld1++VyfXfytxPWofQkdm3YMtl6FPU/+g90DNr
bPeUuJga9e5B1haf63+aywlP6ezY0DYEfyqR2Ip7BlaQwvpeD+lLOhfRxmb/B92s2o2ab2XqtcuV
PN6LECK96dBadAVHmgfLvVafc9t6U1wxHuCDKxLE1cAC4GKMebz9tewhOnhTQsqa1ma6wilPBRaz
WYPead8GJzJ+bsri8yXxKQcBHO69nU85/3e4xQqKhtRH4hPEgWIpthkqguO5Ih3IcKakWC+724pk
3TA1It9wDOI14fGVrDgCp9wW0P9VSwK05Tw6hN4I/8RJ/oDjXJareYhXuWnpf1yhLoUNHD8MmwKj
7LQUqrkCdRjVblKYrBY/m39P+3dxLuE6kTMNn4EHb+Ta4HgcoNaFi2FpchdJoLYWodSQLuSFVo2F
FDtso8rfFgW+r97MlOMlW+konvMw/L1PfhC3tsbGdGx7LuJ39RwbAPUb/35G5897lUvPZGKYOmPb
yoKMvTgvU8woISJ8p4w971viydWOv7N142+UIrlYPurCyfsT6mavdiYUZZe8KflM2f7pjWf9eM/M
PA1TkwjC2hw5dv/UfypOR4RCc3b1nJExJamzMTzdGcnaOI46nrokaBPsOempqqdbR20mh+XQmny/
gyhBx5BfOXiittD7ytFnn47XHHeuh6dyqa8wLLBoGGdjPNCXoM1KchXulsC2rrMNvzDYxGrDXbWI
qydTHygGpt8+2oN2GTNzrRiR1VN3SSIs2tqXxugODBEUq22G2yg3ysY5LJfygmNu04mcgQJ9yLGo
Jsd0Ep9EHvc9jjgsmNkKOgYZ86RnfAZOqz5J6d12jpt9SmxB066e0n7Df1lXY/mSFtcXboLyKCBq
B+vQ9YjxurD0uY9SAYlMfSbsMUFUI0yf1L1cddZCedvW0vwKUrnZMCigL9QoGTuRD3GbB0zk4t2W
lX/LM1vsNfAkLHK/d7hT0xe/HKKD2YdzjjaTQ0zVOXTYY66BlGfkKyNcZTEIzjIoNu8MGnilHDXb
Ykp5mHqqQ6OP14ZJNmArXXMrokMGvgWHCEMGZOtxJJMaCPMsmI5O4xbttIDQF8rm41q3SH2Gbkrp
NPWQRsT9Ilp9vTGY3xlZoU2KgXtIH+M1o8QAdmxCREef4cNo7kTyq+zFWWTeAwY2Pxr4gWIwux2i
FFW9Ocdur7kEYz2XHgvxA1BuxqO/yM/UrD4I7LJD9XPoe6F8jBkBj2fzFzdQUgzDcPABKePQOn9l
pQBBT1HuwyhD5VECXtjIaqLpJOOhvOTW6Qab8w5vzFtSrJBT8i0tbXynrXoQYz1eWzXDkCmze+1a
7Ap33Sb6QFQEx34C/kKQ6C/raWgyqOXfH3f7VsQzkavyjnteSfxdz24wUvSZrVkDgRHstiQ16uRd
RWx6utyCPBUyBcEDPcPAEK3YdVN/g06VP7bMnzwfOfEup1zRwzIkv1ZCmI+tHMDoL+REMeCxiTNY
Gq3VpKVxGVOfVgICMWoaafdoX8Nf03RTJ+YB4XvQIFZ25mQFbssDUyNdLUE4VNxMjYC4jTsjTmL+
k1LiVhx4kd5npuagS8umF2fWLESyqIYdNdvLFUxw0Up5UJ6zJJe6wBfHSijMYbpXPDDAZALEtKj8
rd3qcFluCuDiVXIEeKxGFjUtg5QhZDP410RfO2/QkTpJR/RA3bJZO4N8yTgC4LEFYGqQ1Ned/c9k
lEzgL/ktmZFHAzaBBusu9a6abFow9Nhu0vg0QQootqldoRP2In/UjO9qPreHrAe7T2kosA+P6ctc
uEeb2O3Bu42RRNiOSCMAaUzv/VeKsNDF3IEYd0ghqWLkUSdqPPq2oi7m6McBcHQvcpH/FBNnzOEK
wFz3TOGWYa9TAbE1fEKTdyjU7/SxtNpouhPO8E2tcFHKaSl5JpWhojTkDLfBrHkEpWmZrD993Wgr
Y6QWocHGY4Pp4ToYh9NlCpE0BRIfZK6JZh43kZy1DKWyU+xv8FFidNa5b6HdlTqTDwPOB/164qXg
xclccJVtsOZZMH/+Zmz5Tviygrmo02maeFZRB3TtUGhzis+4MUzJgJiA4ZjLcWl8yV+JAxcwZOQU
H75YY/6SGK73zFnZg18o3y49ZDQDpOfgozbgNYW+GhcNw9VobSx/wMvrzd1habg5XQLZPv7YdwX7
OeqY2xVirhNSmU3AYh4/SnBs0EuVEp/SrkvuIylGEvvLiG5Oq1Rrhqkl9AteMxwJYyyBFuV9GsSZ
5dvGNiz3AEfNe+udivVlg/HI6tplZ2PlIvSbQ3vzm9ipJyLfnD7y7iEt+KYBn0KrJXwjV90OF870
raIsxyYVOF8SdPhTMoWjI1a/GnwaMvtpuEbNwe5Fi2It9BKjN4jiKopFjFspszEvIDZ2rmIFs1ve
urvk9UZuVO+oyA4Elmig/PUcixUs4BcrJDuKiBZViEpeFpO4pzkwbl4yVP0eGqnPmkYhOS1AK6X4
lfbnFGcfMGClAYex0uQu7ZFXHQcQI3778qVMsAsH7/XDm5nJqBF59vGcayoVCR81Gne0xpi4oRaZ
5p0AgMjrhlN/7BSfGyU6SEa9VR4RyuImghA6X2fsgvAOKoEy+oGbKyDXS9pVuesC2k9gq7k8P1OZ
S3A3lBlWkUqiYKIEfRfU6GGiys2/OyxnuihXf72Zudd0TM0ldKaok/yQpBVDhbJJz2BkkyFP5qQP
OTzKWPZQHprIQS5CSxXWy5VzXyQ+28G5yYo8D/p+DanpsviVkLQKoCcTCdgQZ26gPGcUhYy/tMmr
POgerG4BYVVcHYkYzvGmBPuA+nWdqBva97dXjdd1l1qjB/8tAOlxlfysXeea5zJhWk+E/bN40HG8
7jW1wzobiBdRWioVwBBa4v1i148/UuHjZJc0Pz6/eaXSWb2ajvjnNX7EiX9uYlrtQbynxTiAaJQA
K+tgEJ8exO7g8TcNSDBfBKJrMhBvtWEG1Dxi1K5hkeiTVdxExgHgKiNT1Xs9Y+KZbktAgFnNKELt
c1UYzKP9tVBwJxjo5NEdI4VpkYMufCBMgE/QFAEe0EsFf2FUtyqQX9t3nlSb7gmIQVdxynmmt4cW
57KXwBVU/AALO+SLdb4Bjp+pZs7Sz/CWCJ82CcDLokKQT81waTES84aYvntdw1n4bSG36LfOKlSY
Yg0tDEZyWD6QvcOFMhxafI0gJtitj4LiaEs/aDIeiRn4J+/9A7yw4hi+DR03CQcIFGuZr7cNkEY5
E2ce0QPhiO7JMoQkx4vHY84Y6yjb/7dSGbS8COd+o0MDQOVlrnA5aIZxNPdO5Yz/t7SMShI1vTgd
NQ+yV74qEQHpX4wu6h+b25YwN2hkZkJAS8m2f5+rxxUyDuvAMM+YCc74SeIZiukXXbC9Fd/rrfR/
k5bENl11JEwhe5wsvXyKI+eEObkGI2HyLpwtEjBWMdhXCHsKQhVFstsyWVFTOxqUuT+aRtPAorzZ
cGt0odwvx1TiJm6+KcwObZ5qboXhwPGfnZLgQt266EySWvYatDPk5hw0qi20VUWk4TJotp6GfFVM
QIRI6+IZt9HGOX5tqzQlvJRn/kRuSWQ1/RSwclaIJCEfi7W4GPPFM0gFuhWK3HKBuQpT8QzRl7Tt
2rdJeZpp8CsM3VZYOOgNBMq8y5sy76zW/fwNFE9ngggK9sAv6zPKWBuXXqzBImUv+2li1nEgpJQL
k4qb/5CofAJ/6iDp3XsvBD6pRUcsHC1EcqiAkqop3PhzUrhe6x2xIy5oUTZk23yI4UPdbHe3VDYG
0X+PuKJDPEARElQvAfEnhVrUYWJpP0u9eAaUEQyTsuSSsiGN2ktWcIBTglxAWMLvv/2nJO52JNSF
KlfK8yR8gnC6jZtTH3BqgKNohQ1vrnmOhtXObconl6cPNaIUpNNzANhyFwH+wE9OhkF8jq4+dbIb
Nqq/x0+PbF9zRnwRo19lYBRHhufNN3JhxaDcKXhMXQhbu0M1nqpEu3R9FyARtPpWGurmTGFZqpES
akmaY838uiWTORfcnAMEUuhoqt4CbwblI9msydlEEdOpAgahXMlwFYsrPAztvoYhzyPUHAacjrJb
J1n05wcRSgBZ9jNn53s6+NEZXlivq+We0HJCWyBtYqqKV8hQlCD7w7MFAMmxOTATXuQW1QR9Yah3
KDGx4lV2npo2+JYcB8HqLRirgw1nil1cnL4C1y4pRL6ghty5ZQbPQ/QBRyS+0P+6xYZ9QpYDytsm
6+IAwwSX99dOH1+rf5ejt+z7vyOEX7KC8+ryPEjnWLc2fpUVCpU8DkrarweRMRtyq3kcGFNBo+20
rKW5VLF+JDyNryIdYbcnmYrk0+l9ONY6W4Invotp1FAa62DxN1BYm08UrNiCSsiwgUAKyi1QTW9D
s3CQdY9xwaSUe49+DLGiYUmHGe4MuDX1hwwOMM7WUdApan6Stzyo/uVs4+jF+URVztqFChxBio0z
Iz2A/wc1nAILzcmLr8+m+dD7Vi+mNPGDHREx4iOFjTs48az6PP4/lMDwOBYT3X6nl3eEYC2knQp6
o7tSr3j1iEpL9Njw8unnmtmYJB16d3SCltorZpHICI6/ZSaT8WaSNSCOQp0DpDP9C2IE8nnZXpYI
vLvn+BRLR+mB8m7lUxO+znvoAeHLYrmjCK9hXekEaQjWFA3tYsNH5Q/vtdhuIw8GAMzauXSUVET2
IizAZLR13EPCXeP8I88N18thr2qycayMBF2vV6AKjR+i53N/kKppADxzHyitiWuF9+9Qbe8UMhKA
AcwOPGpPVo8y1ZVSvVlDd+cQmH+j36kA3Xrgw09G7Bhws4ZGrtbtSpwRPyY2ELL109VZ7ngDYTh5
YfnsSrbRR4NOEgNPXuYb024k7l51/BgYFAuFAJhjBPad3+RAbNsW0BJFpK2QnBxQdFEpdk4hHJdx
y7HYlPVT8ii+qZDRtLCglIr1RxvqVqoxBCNein6NZg9EMLtmCqAhDDv4LwTEcypvVmZ6qD0/f9jK
4IHAy7VvlKLYdptSMsPfOuleasoOeH4oetMwFDZqqTMxBglQ6ts0RqzkOSlkYo1UJ7cZUJJIZ4fP
tALIa2QInCmbmPGFM73s/zDksRTsK40PpkPo3Bo67qFuItM/+XIxRyw1jG7rLIkpdHnd85P8ls0Z
l6xRR2j3WlwfULBbRW/KegVVAiXJpQtpXP2hlKxaPt4PvhsJ39iJK+h2bxtEdM7yVAZUuHydfXmw
dB9W+AVrIbJwPA4N82cQEDQGi1vTQfqApa2NfX1RgHqFItUBB/HHvGb6HqrGoCLihKMQ4WkirfJu
luaLd+uljv2QCAn3jmsAjaxXf5rNB9Ofm2IqT0yAcxJ0XExdIsFhaeae7DB9J/p9mRdydEjlEPmN
GBOAiZhoNFPuzV1hES2xdv3utjWxii64KkwFGn0mSAnSG68fz9zFJkUVjWKzZaB/mgqH1m62E/cD
B0YK35ENDM6CobkM9LKVeY6g3q5n9AuvKGo2E3MHcIDdRGsqcwvVEJHgZe5AhtEkICE1D0C+0vyG
0vqdQw1jDrrHxXbgeDZivXMVEZgf9lWYuDQpXXBXb5JhGpa4JRGhHH480fNE4uLl0/m4+cSKsOuR
pEljW1gM/B5rWl6OihoyP0BngHlRUDDmHG/GpyAgV0A0F+Tyc4hisb5+jH8sIL5HmIzxYBl0TSvU
CTvUQk/aB2QmlXH1JHtQY0QFmH41lnFjrkUwAWZ75F0VRFTI+5bw3kG+mSdtY6VDdPd3zyKplIhw
MTGV295pRpMfr8yD726f4l+f7nzjXbH2H5213lkf7HxAIORtaVPBxUtWTn+CC92l2Ubh4o3f0Yh2
L6peDUf7uInpsre6RF2rYNbxKQ65aGygWSeBkOL3h9PuZRfp58KIEMcCEbP2Se9qbbLwZrVFYiGm
N++cNSa39siJiX6HQonhn0spSzy636Oy/O1ZfCspwoJdsyl0R+9paQsPYicMhZ3cUzjKugto2bSj
iTv9xBxsbgPiY2PgAtdrl7Wd8mye/gD6Spt6REB/zLNxETK6kF1Wl/Ki4E1ubaWnff8zH6sOfthj
6ABUdSa85H50wXfWSQLuX+PtHQ0kL1q58AtGgmnMJ54J7dJPdnePA5lLROklM1ixCM9GhhuGi3iF
sdeaXirbszLM1TLpdLoPQRCJlJh43Tt6zSwCClPO8feW5GZRyyvnYAzFLb42XHG6ug70lW3eI7h9
eUwjrFlSueSnSM66S9lPch+/eExuYJQYnaF7TetNzj2UqaeDuxUFgC8a/lawo7L/ZElmQFYD0IaK
NVN8IXPsKPRSopjJdTDN0KZCFx2LGnnSACRsWZfDmF9oE+CPyAuZnavnzxwBrOhyMFSRBmHMtQJX
FD3Jipfz81gvqPoa10zWOI26dRXtpa9yeIBA90S6YlAHAxH/X4TFHda+0Z/h2fIHOwOkH6YIZgsO
aetcxsf1YjyruNeaA2I5TMiehKkaPR4cAv/SSqEQMd2vXT/O7zcuWsixWp7uav6QwBmmlOnz8q0G
d9wQAtpuuT283zVp05CmBnM4xzuP8iaSUT4Tpzh0InF/fWNFIyMhMCI5J+ZshqoDehk7mMgmy8df
0GE1NFeWfR31JRzxSlInylRZ5yE9f6gJkQo36m9Cbh7ZR4+sRnteVOEpQuT9Lv44T3yYNhA97Jec
9+RWy0HwDPLJtQEAysRbs/CO6GFsZkSZjdJo7+5wwH60CQFHIsTXOY1z69y5uJxg3z/USds0yaz2
6JLSFT40ZpA7t3fD+pZPBTUt4IXTLZzV2y8o5OEGcEXKoCKlDddQ2lzB0Ykz65R0JHiGdWx46Uvr
BcO1uhLH5nG+PLlOOiJ2z3y1B7raVRSBshrofQjSkRk2H0uocYH+1nQeZg8x773JKBc6C5NkVBEB
Tzm5TmUPS9b/BC+Ae6TtxThV3xJhusb5vvDtopycgmfh0y8acpc2HTWP5IPI1oZo4m/uCdqlo9F0
6iQxqu2t4c5edMsK7rnTJ8DZ0YzVWo4gwrw07Tlb+lWHraCtEuaRg16OP41DUI/uC+YMP/nbclrt
GIzvgvRGWpZVTB6r6IhBbfeV+x/K9vB+wymB8Pvb/bQZcBQM3MMhSgPgJhj8M4LKPgJ9HGDmQVXz
EV3yfRhRTQydp4mBVbP4DvbZFy0t4PYH0HDw9O/0QtiSWVtynvrdP/6fJAwvPqXB/5Ft1VTBs0ST
ObXd0VHFxPFznhC38ssyBLj/xBMos+vhKSFuhllS+PqnDxArow4tiy0/b+mwms2Lokvftpa5zdaN
Rx+yoK808V26y4fVqaaZ9Sgc+EU3b1YfQ62jw3TOOrZ6lZTSPandu++V9jFKKW7tPcY4s5lurANt
ME3zEoopbpu1nqFomAcA+VnbXhiXv5Jg6lhWwPhz/nIu/ja1CIsSC2XmmOh8lDdSQjwrXCSQwzhX
Dsfav+go9G+oAOxyxBC/S8tAR9FlmQkHJAa5P0bUZzrz0GAa7i8/6cvN9CC4iFC3ZKmHDXgs0bIl
pFe+jaSjTF0YqaRLFqYLPNxWsLVqWAO+s6je99ZxGEmi/pS8A875mmiEtXZkq/7l1kmNkV74Jbab
4toz5t0Dg524yNwrl6K8VcdXU8tf/kYfX2ymcnAHoeqgprt73D6UVAxhXpstwfJ0CyrI0/PVY8ZU
sQWkIZI35K2DybXNpST8PtrLgq/NsBxHYfwwXoo+0EIW1gxUllq6PJKzf8+KYbuRrOdJtC1mN8Kh
GQzjozRKpBi1gI22blxMT4ymFSFkSRTtq5AIESb0cCbMiUqNBEEaFLzx5TsmQEYVQhCnBX4S+WSX
U5fj1g8BzpAShleAxgyzbLr/aauwrvHWZGN0LoqFkuSgbI9k4IasuCcqw76HN8h45Cbapez9k56D
KkUzHBy/XDLEqO3qKlJkN1g2DxXOkrtGKp77AAEU3RxckqyEvUWBKMUbrIcEJASemUpEaCasd6+F
YFneQ1TUJz/wUuBQBwNzC7+/0wG/KBdYnztYOcem0XrX58+O0jMghuaDrS8BTtlzhVtWebh5OGk5
sDTDVqsIMsxjn0SfxlmVjDCPF5vxBNgQvetJb1yVTebEC1eXUGeRBvJnIDWKp3Ab/yQbuTCS+Q42
vqgBb1GYDz7jRvLfIfbyMPwlfyVIT2Pfw68zfg+CNQZgSV3PGa4TW3jDhSpYrbjfBICbqtBiyfuK
Rlw4xJPXnpNJCYqIttlWo9sMALqno7NYtgBl7WcTX3o3++1XrLIyNdkITdvy2Dx9cEC44AehvJOf
KAjy72dZhCrUqni3cv5KNF1XAa+n3ADhs+0ITelywFDJpVv9LXhSS+a14cHk+FVNcHN/gXq13q5I
5MwwryTDoZr/2Sj2OjxmC3fmnUy/ER1DGvTt7tAs74WUxa0FESwD4QowAiwtdMGxs3HsQRXgG5Cx
fTHs5uZNu/ZL76yT8jiFxp4ckK8NSIthppezRpAn7VNq8ws6BY9jWKuKwwklWJZQXAlyZcobcXKU
ZdGVf8u+5QFHtNFlTUVNVuhk25hy2yYAi/E5pAPb4LJtrlEIYKNrPS2qpjy+lQ9wfsusdDCPdlwU
H6pLGN7cAMUeo3widQ5DyuqdeAlJ3Vq8ZeCE+Sz9xZa/PalSJhhPmkroKZfzIWIaOGRgvZdVRzFm
oDIkefbS1n2YiBaevzqJGzaFl0BuyANXtg9aavk7X/nkBeqTEJ1q7IwKPHsWAsUJQfSwQ021ldB5
wC08apiUuEp2HYbPqU+hyUn221QXhIJ+M+sSg/PrKxnk1P4Bm04wzudMFAg7JuqW/vnMtAQtWLIX
/0Pk3RbTSGAvOBgw6iujAgWeCi2EDRHHZTE62gHFR/gdEGj5wySSe5XIOJs6rOm40kPOlIJw3WVn
SvIb4VIFR4rJapOWeK16PCUV+TeIWPK+X0JWyxEq+7VgvaMH3NbfXqom4tIW9j7w4GpCGeZQ3/+Q
NtnZZCVlHZQBBJfeDpvg5PUIugiwCjLgk6Kl5+rNDsvnb0uwNE8HPxDQga8dTShg5GAnQpCLcYxN
EXcpM49TJWpaEKhQFzXgRYcrKdpLSZCfSp99gcoEXGqmAEK9l3g9tVDlg0QGupAhoa79aIoJzv6i
mAsqXgXd3gU8Qbbrlq5Wj/3QDo2bQArwiCrd8anc/4nAyqhPT0y5RN8bA3y41o0C0dj/TpwTOaYd
LEPsOAHjEuoJ/0vz4n8UmtuSONmGukL7l6gw+3PKGEMMol9KMTTaYrER/QAw6PlgcLVQ20zQ2hb7
X/aH5014ovILMxE/055PX+RDyra9pLbwinh2rY8uH66ZanwnK/ORRfmQ79haaBvo58nEXNOJgk9/
31QGp4TbOfnXPEDcaGSlZZK01b5mXcgQTM3csDXAUSmDNhPRYLfMSMEegOqXY6trGkj+bzcLMyFk
QyjUGb6zlXfk9/kmIflu7W0cbtiS8UVKvchPK9wsFull+TrS/MW0rMsLli2GKbgyVBgMSB+glfL0
/YjLA2xHO234Qhs2w5YyeV634vGPws1cxYKnY6lDsh0rnrUtQO7cYd8QdOZgPQdOworz338vGCgc
Rnl6XvDoxV8YMH9Z08VhZdvmaqO6q4Ewoi+Usa3rvPO2jMtZ9ukdXtEl3Vvx8kTbeeoSdzdXluZj
HfbSwPbTty382BBaEGH5FD4KjbPe4LUlVoIsrqCHnC0kyVSsS7k0Tb7TeAr3MtShcEaejfHw/927
01tdo+ua0TdK8zomQeFAVSa2hVnvKNybExL2Cfja4B6WoxXTOvFUX1WUh63tjmDa1Q5P0jOZ1pvU
Q9Igsxpq+QuWuUJl4/7csqTRKK9y3AJlRMvc6EY1SKjtISkfVAsZc23OtHG4C8wU3oQFBCxzDNyq
8LUV/suANdNaUDw690kE6dDc8KU+83qTgSq4UQQb6/zOm/xaG76jT5uMqaNfZ0mUxVGXnnm3YvY9
wNCgbacI4HtBzInFyJJFI9tUubucn3rauVxuSto8/Gzncr7q0j8lwZhAJr0QPhrLwUBdUByAuypC
a/0ydjgItLn6xKsBXYDWsQ3xLAjK28ZEkFJgNxrussWeMT+41rLZnZ7LA5dwaojIt647KGCxtZos
jmA6VwdyhB6Mj3jUiweV+mxOqboVbXO94GJJ6T/IjRyVgj433BrXisd8ux6P2GSOyNEzPCaRZWjv
KGpZi0nKAe25yFaEwsmLAg0deouUZ05GgZfxjyBDXhAqoa3t6TGuXM2jApMxnB0EbCqgf5Hm52WX
DbQ5m5xupzL0JZUcv/NGMXGcbW6AgFB2O6zk0T/JHc/UcD45TyyyFOXceuJruIYVLNYlZZfFKFuj
0NX7MR92STodmWA4e9IKnD7g/IKnxsL8v4DR1u9cmelMnM8fZ08Qk9RUmLEpE5/I4cIMzjiMG/4t
RYTE9nJFZvuUdR2XGeVEOXVlwQexnsxWTimKKvJsw7HAdjsEA0tdgzPUgQ0LUEodlz2auIeThNpb
+CzcPr/MtHOTrmtz6NLh5KsBk3bMl0Xmr13RVW6sshCDca3RCXpAn4Lvhh8uboseuucrHdnw7Cd5
nZgwUiHHwKouN8SnaJ6z+XtKoXSxxN9wV+2P1bBSqAU7KMlKEQT6xVNr8tJTy5G673otB6JPaJ/a
IpzPMGBnIa8+gth8Gt4ECVmt02MK2nkPprPRqqdJ1umpLRHW5ct04k4F84FJyGj4OY6vVtwg3OFP
vdji6ah6AAKUuz97CXQPJTEIpNfXmhO6M8bHwEn7yhu5eQm+nPHn4KVOLtN0lI/48KBlVpkiEyEl
f6bG/BdvYXWz9mYIAAgR1eWJeOnXYNsBqNtfKYxYFus1TjpndBJBIJT+Sw8Qw7pHWvVCSs4EaUJ/
f7aEZppNhurwVoMr72GGKj+2MjZsxDXzwZNbkMG1mOrCJR0SXTGKFfVdS3pUAaHmYYbtAB/Y3a5Q
JiFXOZeLF4WViZP4BEoZnuEB9UORHpHJAnrTexRRJr4hTfU/oKRSN+CGGgNN2PFJFJmgFYSgwJ8e
LCdULckXZjbC+HV0OeHC0f12iiUyqXKLekDVEWpwws5l6CNrZddF188e4rLLJZES3zfytzBQKz9L
d/CtSAj1LsSusB5Z6QuYq3BV62ms/bIeMGTjk9AL7kn//FpxyEJkSLQhli91s45KUcbwoWsvmvD+
wxc/yJFIBhNgLbCB5NysN1+soAmrxfEVngwQkd13d6BORSv4YhyiFNfMiy9KyLXYWHCOOuEw2n3l
s66u332lVQKTLr+J0ykmW9HyY+ehrJfvyuZplmvY/xfrs9ibys6K01APFFZarW9vZDi/BxTKrAyg
j3Mwa+RUvzzIqKjOprCUwAqVUMUEDX7B1zgSI2Ii8QbniuX5JnXp8sIAfC+K2CW5I7IgLSmPQeSl
+j01a937vfEUbD3Ch4xDHbcjTSLrVsniSdmqxhL6wwJ10bpNE+pEt0ehVfIjn/Flup3hz3UmtKCI
36NCjz+7ZiQK/pTi2e/KJ6e8B+fxKQs+w0bEz4VE1JwaiYa1OEHf3leD6685bf+AjfjmwNCAjvmP
8FAhOdt9HFMSZQGw2I36/fdSnKVNI+B7RGpM5GCUbAGN/1whOatinEN/hIvK/EwiCOS9Yo/mWjGc
lqTdpvOoou7IVRBzCWH2ZWsDMv5Yw4A6TzzJPVulCszIeelUUpWdcpOtEtHw+4lbAcNGpWdx69FC
LuUBi0ZI1B3tNMVNFYS3IEDOwLrg32+cK0U3G2cFv1eyMy3YbDyrcZT42bj/pEHppHSm47xvnlDl
Z3WVK0YsilPxUyMY0QP0myjV+PYqjLe/iJIagh+agE/FQNPGDWOW68/DOCDb7tfKqWB8IHOhgWPQ
bes4sQesHHqWiOVARKOkwQdX1CoARRBPHb0mJndvCYIxdXGsysawZkxbXdux46ORrBwdQM8/YzVz
rw5j9qiSvJnf1jaZLRrEZSIdMA3f0Q4Tck11qYWZOflRV6zgePJ9o1vQupNUmVsfMlfurZeo1WuP
4psr1Jls5FMuP7r1iCdsHt9ZRSn8hHT+KajpiPtFr87kS8CXxhC53rNhHn2X1TM9DEZkePkm3MLO
7KT+L3ZkqnF8SlFcJHqAEdsjPrrdecvtf68WE2EfzLFPEb7KYkLKw2Ul9+7ujcPna1yfmZ6+q3yj
a+hTlxoxS5nYT0E8CTh11nxbzNGI9ZqP9GvGXllpQ4kLwCV4pGSezJAqmQ2cIo9OSZsybRL3+hZY
S+UMoJpoPj3YY3eA/KqpOLr2xUkYuYSQkN8D079Ttj860b0lhUdJgW0R/u4QPF96l1d4O9NcugGC
9aIcFDxiGMlgYPuTz02tmD295xc9RBIH49sk/5hu9R0H50e1Ox3vwzfGrwdi/Y9mCFiERy9+mNgP
oCiJn35jfsqm3MB1elDlT6qK3cDb7vhkQcV0BCFwy6HgJ73Aq6Yfo3xiCoVIrL5PM2gZsiC7Rkur
UM7CeAPn/c/rBlUs+NdeUVG/xyBwpr7oLFsMmLt2XK5TYe1pWRgwQR8gYfEEgqeQWl08grfwlG2e
mQoXuDcyZp7Jp+qGJgzn3mZ9vSbYrEWUxn4VjVru2qZHqoRK8C8VEABKzvqQtV7/0QUidGtFr5J/
kyx1PGLI2aN6LLwDEIVFN5gh/3ej3duHjv4m/4VaW+iL01PSLw707OXRllKRki2EPY3Rb4EFMDwG
gI0/ch1k2+wEjEvpS2c05Uv3b5lwDKiVQYe2xyc4Xj+8fLctTUaPIyuc6LeYeBTpVhtdAZ6gKBdG
qlFq4iEScRaFyBLewDQ+jjeRAopF+Z9DQfAC2OrEvfPNA/O71A5hv7SdQhRGpaNgydGkbKcCvZiK
aBu+AJAKSw1Ja0jB5GevVxzDRFVA4AoesO560wJ7fEK7CAzmA2oCguTR0EKzCO2I/m+QbFCWu7Bq
ifGbDar6J8CwXDQEdXMFe5AlAg+HtNA7ua3vupjI9kmroLd1reTcudLpwLhX6waavM+AX9FL9nDj
WQK7cDZfy6UMuKin23y94Jsq0Xfe+MrR5gGgVG2cysNmin1yD73HronCUVgwYOA8CwzhZl2+c2w6
kvGHR4gt6tvu3NnOv031/N0nxYCI8Jw+2ayYXQS82dGB96db9LcK5vQ4AuqVNh/dSlodL6bC6Cb8
UnInSAbkcplJ/JDKh1U/SbkglJsVRLUXdIeYOld4zmPlpOxqYhK910A8bziUx/okqYf1nZ77JPFZ
ghWcOqi8MV8de9hsMsWEL/4HddQsBKSnFT4L6vnZyQPuapbUQSwNsud0hrPPmMcOcvCoimlG5Rc8
OA4e5uMP6Bdge5jkQcQ/MiJ+PCPHd34zGiZ1qeazgE4F2DKbCO2KUR4RIi4uG3P3upW+IuYhZrKP
tr+4uZUpaKpGAINgLy4RaphkRWTdp+cf7QNoUpSHsmCspXQ0dF8cagVDL9ArUIDBd/2zoOXre2lL
L2MM9M2sjsFBkutUXsNYewgMkya+9fFpERLH9pn9OBpD3wBPURXNiUr8OleBsnBVslLO5Ez1hdFI
/hZKC+dOQhboEBmByJm4Xb81cJOCVDmQWJiMjc44/JNHeFYbnBwv9AuCFW4hu6ac0uqNyYmbS4sv
A0oaQ+mdNzf9T0chJ8/J+FAq1CFVlL3WueeFbUnsLfnrll7hx8lsxY5383Gnt/5+NGUZO+wKxoMq
bGX7N2uK21RTNEmw0B4o/AtbAPd5DOE4zSkYYWLtGNbChsURt7bzLUx0e0mo1plEvXlg/QP6pHFo
5xYnJbWber0zf/Ujl0M7UyQlUnlY2qrOkvE8lnXJYEwrOb82P19EdfZLShuq6Lkb+7CiIfAdTKGK
zaNbOtEa1QOWcyaVV/wDs1iA/4DZ5D1OT5xmWFg0Zvq7QGHMawVlc89VCyLSsx/bQwrN1CikWwjc
LaDwZwmpl1am2qhjLaLHEErvBE60eCV//79zL64X+mosZS4O7ygLHiqvLnjKGQKrhudBxTeUn0m5
qH9GrOuU6jfssZz4jrGz40GAdXAy3NPuICWm+msCzeyk8sb+US97NfEZSQn7Mr5dgbTV8Y2pzRd9
tfhM9dCldAK3OVJVHTazvZk5y8/bSSsfy7vAhJrVj2GI6BWR+FGldcPgNrKR5hWyZpIakByrpe7h
wxiy9BXpx6rHnc0CzQqvP6JZ3NmKKG3z1IJkrCnh78QGaVxzeIAEDEAEpZrjO1TMoEnXREJc2EJQ
b6yBnXJQ5j8p3uS2AfpoQtCGCxG0lIWf2nRnsYdAP90jPnCYplkMh00H7Ygq1FpqKA47iBxZ5HsI
CmKTRVmCzE8G7OR04dbATWLeIlJjV567TYMvPyzeIxWjCuuGGY+/FDcaWk4yV9XhEsGX36lL57cP
YiRrmARxmMUQxs1r5jPlAabd/+aUOXqfQHQJtsmNBzl15dFF/SdJcX5fZ6TYk+JIxebFndkrI50n
X7B3ORZ0bnwASXiPNVWeVR5Eh354j2N6l0Oz6eT/fo1iGEJBhBLg0AQKHsoZ/pX2voHibvadZLbm
irllDtrBT2IdSDqTbvZm692f5c2EX1Rhg6N1GQvA9XkS1Qx8//qngfLyyk1FVvQOWFChm4JTRS1j
6qL6nT3VacMHkwvYm37WbHHJ1rGbz/KN2d6QUXgOlQkSq56BLUeteAgLG9k5kag7kp24H5YfuwM8
2/SP0fdBzbsS+2bw1yx87rCpQXkS2i64HyTlEtSq5QbrqBDlHZAAb+SJBVjNUdn9mRiVUvySiNy+
mBUuPCh3O28357N0X23X1KpRrOkTLmRSyE52QZWUS7VkkFsmnvjOqTIEsNYMZ5fubXSLpH4uYSNC
qAz4Cq4Evdojj2fi1dBxBLd2pdKz/8y9DAWRT1kzDAklvyc6gDl81SuqyhubKAYtJNYKXKRohJus
4AD4/Q+VsnND/7RuJ5oRgAXCRHiL5/fJx5w2uBHPa8XLt0S/E0eAmhmkabk3dF61sAn2Xjglx1l0
600eRx62NRSWLEbQ2dO8Z5h55KkJV+2B5zLXFXzfhifU0+7xF6hkEAuJE2vipCU6uPR8I8nTmDGr
P01Ec1ldj/n5f0596FKSSbSOn2mUvLGq4GKCNatFrBNDBIIDoVeAi3UW6G+CZE6H3QNhVaIYlnZx
WqNJd2SFsEcR9el7H3stP3DIRg0vnZDS3p4VEij9RxU7AdPaRlC63886xSFJF4MRRxc5ZiLOoOCW
SPDl7YjWTKNWVtEVUQswYN4JqZuc0KYpehlVu98WDzLpwokAdJaPco+bQaPSh3sBjA+yoS/2+2kF
IzQTMY6h0L+CFPIv7qk6p7pLsG4CDLaQ9SlgMDCPT+H+8Nvw5UA958hMoPJS6JF4xR3aAC9oAMu8
jW4kz6bpy2fTxSikxrQvrrAmQE1jLcP9YWa8y8DgAywnFBkNZdyDO4AUTSCFSE/Ga4kOAt5M0frF
KiaLS5Z+WPLGrgVlxiO6nYLHx7t6TNJkBTdmL7HJud+yOyFXwQ8/CNmxITk4DttoNwL2SJxjQ9kZ
SHRc5FRmSmT9JgYH+2D7iuVt3nHPqpK038Oi+eu0SOcbbgJwf74yHUMBUveZ/8llRnMygoZPb8hx
fGMMX/KTmNBk1L1eibJV3Xy0Wm1ychajT7lssLjK/g9EQasPArc2JAV/63OBqYLvA/aLz3jQ37mJ
tKbnEr50EGC347BkX+hse4g//hE8+6887W3hHLUYVGcX3lDmHd9qAcswclsEn7rumQaUQWBZFKBl
uAklGCr8fMeJ+/GgiGRuo6m71oMabGasCC7mrKT+3XfSVtnEQzNWgebhyHtI8XdRmoxcGBWMXiQD
slQB4TTzWoAMuOU68QcNKzlBHMJ5qPtEIyscT6r9wlQqstVYCWbWKQWSBXbWp0KDnZXVXTuVaQB1
J3eUGfcFKKNcWHSKqiP962s/Eu8bhs2x++2zHxXDrdc2a7ClBU/MftdsWK396Tnnkj15p+vLQOeO
OfWJ2KhHR7lTzWG9+SEnaFT5Ko5pOcXIHPUGBInNoIWoiCPGcP4DPcmkQVnRQIjKlqe5PndjHHZx
RGsDpHwQBsQn21ktdDqatWtH7SNaKUuFNDSUlqRL0CNJK8RIoGH9J1dEYNUM8S9pASmNzk8g1+Hm
rKOzz8Y4xb6W0nShJvmhmMLLWwOEQ2G0W2qJM1Kogv1AeISVclyWV2qokJuGbXHbl+cJNgLfhIg0
O2/jv8kyH7mvJD8nzq5O0/A+iYbvrQMKjLGjiu7La9/Mw9SikjrAbbzOws/X8BXvXc2Fyjf/Xbpi
DzLmp87q4WSkAECWeLcEQkViWofVPJBJpnGfSFtjIRFUygR3G+laxM8a/H94+nxwBAIarojYPB/h
zPFa2xYugoJX+5uEOaVKxDmVaGMNG0IPTwMW143PEw+Z+jCQFD82iU72IFQwQuRM7L/ik8ch2DfJ
vlvvAi8olcYz84ipE3/gRLDtmcDEN+WWvL+KyQMRJIxWdvn1z9OdyoQPMLeuk8PDUsxkaECQaDeL
xgXg5UkLtgfOpDUbFcLArlNuR1o8P7+mpNXOZJReASFsiq419cAOfUC9L3s8cSKynpClJddKa+5S
q/o9paK7eIgG2dx+Xa6k66vg9KHCUUzwp3rZN/0CGfOJudj4ZVCkexP96xrHIQsYFeIA9gaWip7k
EhwY9DRwqIVCnossrun1RoBMMh9PHmYB66n1UK01nQhQHcQm/71FpzOA80FtvzmHCSjHMsNHBVkB
DLYhyaIwBeX8Et1mljrpzX8bMWWgIcjI/RyjsAVpy6/zyAcctGyPK4Omin4hjCcQqiuFqV252fmm
9qGXoZxjbRsDj6RiHBAW4bKa1+qIfcajvysd5tNuHK6cJCrr2Jhs+lFXdovIByr6ftQidfrvcn2I
cG/IXpB0owQk2JyJVJYXL263e/w5va8jnMJmye4IDO3Ay8klqgNWS+JOr52uJC+GGIMcDin1xmhP
wbCdM4TIRvuXk1yRCXf6+SuKZaoz1ZIFT6rCRWYEikJrp9f4edEFwitAVnNgA/FHwOqx82AjdkNk
pEwYcSxDGIuamXUZKWnoFRf+CVX5dBRlNuvdRE1fPKJ/V6RwOIT2EWjcKPcRNLYd7kpfgI3dPLrE
bkcbGpIJTCedPdg1ubG+hCTEzP/4DhwUJIM4kxirMa/AJj1aG3W9oxxCMeGRW7jRRlNdpRVg0+ls
Mh62CuraBx0ANuKF4T55NE3P4kPO0cfzskPChfOgaqEbR/R/gE+Jwd9xOL2jCIgI+y7QnhDvvSLs
Deb7+UdnUyevBfyHxH3LPUDOKbw6d1q7+MlSodo49S9zYluRPYUmqWYrMGvzVTz3Hc7BDCByYn9x
r5WL4iMarB1cwBiPO8+tzgXbmi5H7XH2Mkwv/lPQgqycbfQAeLFnngXuuOJLc/goTgcYpS5y5i2d
s0cyEIMW1RtiNlytkAOqYpcbgtmbIcpG3vUyYCncW7UNOXGa5ILo369qi39ZfsNd4QcCPiOHAPPX
XGN4lceCPHOo5hSu3iUfF9zgrSOJ4xCmL0oZBAgrxwUSzInHootASN+0NZ5P0U8N4ZDsyPt4/cfZ
cwbSkD3mJghRD/UCVeyRSB4CdXctXn2ttxg6wtFtbo0KBL+EhTyN/G0Lo49UuGOGaBZsNu5fvU1m
4ipiikSZZeFJ5uGp1Op+3gimU0i2asZ02+AUlhe0kb6VVK2k9z5oE5KlIObDMOHRcIIq+FArLit4
wOg/V8dHvbNJhiLQOiSQL85qBwKh32qI/r8jEg1xAIF845HxTKTeT+jA/ZGKQsF8L64Dfxern45G
i46EHcmykQQ+DHo1C1OPn0u3dDbjlhCp6cNSEJM4dSxjLRCWMEarouisH3taL+MGHxyye9DCYvYz
+9zS4NqeeB5oStvROlvx7k6cBTAGrSgPXGPEsploFLScYPLEbQfHwth3j2k0hXTpTth2E13r8os9
gBZ3bqk0SEN2N0EUi6+kBijAsXGJhGMdrxLTwmDHKhrXMb1MnPmNHhOWql9oFQyb9W1KgvorUdMx
ieES4IwQq9nCCahUoZgP6kd+ahsvzYreEODybuxkw4p9kerzp8sXvs2WWZki57Jl6xtzoROC/HXo
k5bG4f3V2lf65JGJp2jS43k6jR7opX5m2X7FSwTfLmAgt353VoNtT+ycWyt11aFFe3O0KwnWokb8
61TXtI23h+5oTqXy43kwt40u03FWrSw/AmoAKvpYXsjHS+H3hU49f+79yXcExPMf6HyfRE0xGdWi
OcWkiPK5O4iD9G51V/nql0VE7FMYIgTbCXKsNk8CvCvATK+7PCbnymMAaRoyKIkLpIajOYub4Jae
4MUIVNtlUifbR58bq5o9Vp/nPoar+5ChkxVW5XUgVALKJo6MUkCLiWHVQGiin4tGSIP5btYjcJqY
w0KRmfWv3rlqmZpeKUv7v4mYKd/1nljPZLjnXqa2A8aa/sfnPmbWmZuNe7iDildUGR6WzRn7lB90
ifVaf3Iq1NSZlRJ/MW7MhNhF4Iwz1Wr0om2z1ojkMhY82GeckMFe6G6zpOw7lcgS0O/j0Ic/v22k
oCIg0emNFdmnE7DS4P0UBDvhLn9v/1Kwo7PchYa6ZlAlmOf1k0TApnKQbJK2rEaUfWXmO3Ogjdbp
hXK69Fu7aEL+OB0b8NjPjQoORgu5v+bdPXCQ1wWsbphTjH+oxv697+Vr+1aCpXhsz4Hjvp8fG+gI
Q8yUEDCgZJ75x+NvZ3a9PePwk6ZxI9xumYMnVff2NhfbqMBLaqq/HdL/SviQQ+REHm9H3ifObbjU
M+5OpCbl31T/2SIvfaUnQOmJTannqHSWS0QF9fkuuLoL7xM0kZoxa+wQFa5OgfC9UiLsujraGq2X
LEvY/nn66Pak+S9mFbpM+YjiIV9g9eni1witfpGrQ4U94DnC7ZkM2lQ8ah2Ut5XVf5DorQfErdN3
hlBWwZPcVT3bYxkN+3qWL67YUj87beBAzZ+rDQarLpJHP7jGRiYmGeVybC8Zl5otkeuzw78rIsMz
wmVnoBPs9LDvx+pUytDq5zyvDXjfzZd2BBPUT7TstG/DgHS8YbOoza4wgJYSDenbIULUOwDGEq/f
AaqKN/eu9f1gA4xohuRyYxAe8jARzrqJkOSz7zmyWqcOAI7XIh6nC9eqsz2wn7MgTze4VBykV5qG
vylmJRy4UOOJCsCmkP2T5CIf4PXFFySeHdnNJOAhQQ/amxFTTDdq9W5AiteHJwQyUHnrXE+mqOxs
fDJ/WKNNMJEfofAPQZPubLU4s6x6d4UwmVfSVJBITx9ETn1nQLUgthu14mWA6DzAnCJslmmV96Yl
tk3DzpsgmzR1zHmy+hy/m7smSaYGNR6KKsFZetlgx5yIgsI2XfpdJajRFGWiZyQYjNTUmvQPgGrt
xgP6gIz3VWcPfovJw76KsQ1CJ0j/K0mkRt+d+ODYFltcce3bs824sK53CXNX6wFaicsgSjkF2jN4
DsX4IgcCkHJXd0CBgQ9Oakv9l070hQ+rXyaRdiyfizH/oJ0ADU2eGffMEb24c74l8IMM0i1AAmgX
IYvsDa826DOz9b8CKt/7cLvsEFbGt2KZkMiT9bGE5Kb66ZBF2nZt119Q9hVQjC2PzNSSWgOfIWPL
lCib7GR4z4EsWuIht8PS8erlAHeAU3i6oL07ahDV1APgsSS7OSOEQcwcMVXm4p044O70z0nrBT5H
Rj+PKrtghINIJf3ZrW4XQ2ODD8xLoz0B4DWaQzrTGPRH8n/oAStt9v3tv6B8dACi2b/u8QIPHsA3
scPgN3hmfHhQmjlMhg4mp4thCyhx1YY8woyE0ijZVwGeiXg1/89FrIngTcALiOiPNP6Jlak2AbaP
0su+guiavq4+bSIo0tW0WD5PpgBZ716bPpMZRytSfLR6Y2HzW4jtApc2a1Rfen5RhSjd44AZCFyz
zxpf4dl/5MPyXZ/Ni0KHUnbN7MAq9w8Yo+TF2PIEnaJb/kR5b7jLM2N8XekjfjEGWXlKLFbn4Dl/
juwhGhjx0a3VrkUoCt11Vef+aRbGYJehNhdvmRzshrzwnBpK87qQJSznYje5wvSLZtbpmnIT76ID
kpkYd2G0eZlsJYkwsSwNm1+9iNp3DGGBQnfl9kx+LDb4sjjalElPPLg1U5RMu7RwdjdISCBF8EHf
4yKxVNYGLTcpOYbcewrUAbSDbKQzGtQjCgErM0uDvYkgUCQuOZQVjrZDYYvdVH5gy3sPWPQvxuP5
fwxoWU1eqIkei8LORBmb398wjaK6C0ux/HjyW2YHBv0kKJyuNRP/rv2BCwDg0WILMz8woKTFvvN8
h39zf4U3rg0xPa+qf7oH9LSFSNV1bhZ0FUjObhP+ndv4iSvPjmEW+McaohUlAi3YSc+S8Far0ML7
pmly7lIlKfOQnpJF2Q3IZOMMR7Bej60I0ANuUvLssfTn22dbK8mCpalzxCwPsmbGtYwbbF4jW2ef
AuPms1GH0D/GgYq6v2dUTOW6a9wH11OL9yX9tEUAechIVdM5QH35/OZSDfI6izyXpwI6IegX6OxS
iXo/MS3YpXPggFbpFC/AuONdWgeYf8YU7tq+jG6xgSwDqKE/DM/MpjVNjrs1eVafIAabf6zuLVd2
R70TXFGmn91Zo4DNB7XMp8Zr86bvK45EeQmNQvvKX4+Ro0gJ9Q8CcpkXdYQ5DwmWyDWToZAuM27K
Yp4PhVW7LZhIw0XSVJtE+AsJAV/2HjtlvY8HPYdwdUiuqZ4Lhjs/eSbr6omi9E4tPV8N74RKKAap
VlcRM4Z9Z0WqNVbp6W41uuwxi3I0lewYzGm1czKO92zBiKx20dWoVfeeo8nLhlJOgwKGtnLUxt6a
I77pY+Ao2JK59OrBt+NnjAtGR8y4dXfh8uWcD59ttye+mZyDnCWXi9o2+wQMG4akFvCMKoTXM01I
eCrfRko5FvArLCKUlu/gVF2RzJux1BxrhyuH+f+Ys4rL5lwy2HW1wtODNUTtGU+z9sxrdYsiUzTr
BJRRiW2srVAJ8meDYxFTbmUiwnC+nNsy9lab3B08tyjc0yiXxch9PmMMu/tQIj0SiSJTCrZzugBb
8o5Ahd7r7Q+5ZRyyF0fyzQE2PGaLfv5QE8zP2hu3ISP1hFJXvPFHI0Gd9k8zaISaN8mG4VVL7gZt
l2CTX2jp+PMp67B/Nd49kvNN3h/ophDLDUyGClFjpjLHvfcvkGnw0fBIqfIllNkjQlhxGiDffUO4
Z9QOrBERQgVTicyeytzZwym+lzWUmJWu+ijoxFcIiskacONlEtgwoHQrFLMmD/2HKcE5wtxiFyC9
B9S0USNvKnEct0XRvLl6/LWfILnZs7RcPekfIox5wmPvLGDrdUt4k2jBZxR20rYT8vah0ubpjWZR
Xq4ZErEhHLGY1M+80Pj/QoPws0MbaxEK7BWu18sgKQOojzyapTNkfEYljMaCJLcoBFRi7kRzc2+7
TrYQNGrHfX+q6gwL2vWZuWTO0tl6YBNgwCL4Jly/XmbekmoYyk6NqPUilZeF1ns7RDiMZ78SG/7q
w26dgPaTOaqqYfSDm4XkUJFM0ZW782Lwv9BNHCKe2wmrvCW/Xfn5z2gl7Ls2agxvPyyndgI7blx/
+6jmvQpzvskTNHOFmtNQ/JfUuV+kxi6EQBPq7ZM1SA+5L0C5o1JdFoW8M9s6fiu1TroV4xibx8hw
0Ue9zg+0fwTj7kHHfBmJ0v2X9i5A6N33fJK96/q34jzByvKZZU4S+CSB1scnzIfR3KM46k5/8gw7
zF+krUfD3IUBnTybQvgP08fS02hdW/TSyfzTo99uJBboYIVrwKDrbi/ls3rvzwUW9UI+BRqQJPF8
tiKBmKFjq4fLyywqGAH7bS4E0z65x5JBaXVhC8O811I7NaIu88JuedvWZ9UqFSNGo6MRmE7I1Qnf
O6KwiQP+uOoBqz6HXaNHJNh2j4SiruMsl8HzxrFDlRluFtsoeHtlhMxXRbLqnk5n5mwl4fxbenvW
kc8zmITEKUU59AVapAGjovnRVAy2+uDEXvw9iKevj32mB852R2i8CosXT9J+AyalI5f6QqMflhlT
5/4dRKPHJF4VvqZMHLLTq7Ecr/aBNRIOdX4A55Ziao/9X9OKr/sK9aiHYWg3KHoB64wKq27v7GqK
1OyXSvmxu0fUZTTaQGJXkxVU4q9Nru47WCPDlwzDITseOJkaRsU8h7yZrOZt6ibab9tgINpNjvFy
9WwEosHQOL/ZKcmjbkNzA9HO7R4/e47UNLp2gR8wWz7wneovMYhFvYDOPTWJkrvOHBbgmH5gL8Wu
nsa7XopaBw3Xcqif/S8Z4oDgDfjgpBu5uo5+bfIP5kVqZEY3rAQGpj8ft9GkQHRr4ampBQwY/p2x
67KA2QJhntfja3HueP0ZnGW2sLx/xHLfMiH1e+JH7T19VDVic6+/cnSTyR3+6lIE02QCjvLZO5Dm
YCqcoeLvjXP2d/oJsg9gmA5tNYzWlZqiXABzjR/hpErNG8EVE+53PmodCNlv6UGdYtiNuDgrLpjc
skNWYl4bj625ny2bKoUvUYVya3OZn1Tzkx4u7JB8MYSRgDx9ciEy8XTL+gqkFA4UsD4yOyF9giyi
f7T4kv/w8aNRCIVXCZAGGNtoJhaoiQIpOw1uP2JheNoyPSF5GKaAEGdgkdULxkdxY0mFXl2p+8pe
y7CuIg8UwKotelXYLTDXYaGRmoRtpZv5es/7bPlhLe4ItvvEKfN+oyEl/5IzKT6tMpfkQy7DR7OJ
7pkuoDhlN712Jya9sQW/S0A1+OxrBydsQBMoQyNSLKqUkwfTG6ipfx/Wh1uDtDJ6zd7C0J7WEeiE
HThDbC1/pX2WMNCMNhfNOvmTA4SzoopHtXKTwpwqVcOuJ3uHxxBmKgzq/bBdfSQ9N0oNqgXcSdl/
nad4J8glgWAHpwpsCqYXZT9RDH2nmUoXFa1v2kjR6DgUM6IxRcZojO8VyhQ1p5Qj5xa/REd4LNAT
bCF0yewIYZKsATh7c27jrjZGO8Aw+fCfVHReIT5Fff3GeRQM7RtJGYBU53RVuaDFPfHnl9SmOto7
zrApfwjzg1Xb45RX/TZ0XOww/GUeN1pClizKoieSM1LjKBL1NERh3Fpyjhj5p3UM+iOrLay01SPP
0iVHBeNo3XcfA3ZcJCgp8E6r+nwzdDDMucWqq/eXsoWwfe0pVor324F2ORlpi6HS2Ovbsub0D4a1
YvbD7RDlXjw/n1ciE3fh14ZgtmJBHpjm72G4yKyVt55lUM2HmRG9HnH0GP2p7PyhW9I/PM/4nqjb
cNqgCwOMNXQKLSNAMPWpk664s+nPsOcmgw8toQzHh4/mM2sPGZjvw/NYeglTpAjSlBFMl3+kC7VL
gKrGb5flYUOBIdT52zBnnJnkh21XIc/iib5q3MpY/R+kk4yzca2guhUfkMoqLUhVzeCnc2ED3kJ1
AGDs5LBVEFpxRN4WNB8sCZ7fBNF445Z3Gr/jyiGSA/3uibAQF8vokPPKXQgSrOrQvAERueJlPK+C
vrz0pPg55xQyuhCEG+62XvGgpgNe3SdrVHZYKdsSiLYuvX9kNtySTwfh4/SWq/QbHyq0S3kDmMI5
H9NLBeftoBlXu2s5uVt77R0G7Fk5CklwvilNYa9FRFu9Q7ncjlBR0IcZy3AowD75cCuj7svRuiDk
0P2Z3kIv+UlUiJmdSFl9NMiirK4wY85EgcR2JijaqJe9Fq2FdruNiWXfm9CLvHIfkyrmlvoLtJWY
Fmq4Lg6YO5HvxSTZ0KqOYPtLX5LQeydVF9m1zJnyeSiMm2EhYPxOGN2YNcC7sKtOslxjyEWI+nGc
hBqJ1FAR96SYjtScclz0zuCNYY2lfLKpNeKbQMrYviNgv5UpWaOJoz7qEv3p8Ly/8Ae/qwPwNSi+
w4K3ITJbi0Vq+zdHWwCTrNCqWqZnpLPHHJ6+3aqH9I56dlFCEkzijLRbJPBbr92etvRQozb7tjZ5
OugpPuzwzgoUxyQLIZJrAnni2IdnIE1eH/qcpcjQJ8epHByTszXKTMpcWxQfvHfgNgKO2V2RM4tI
CWTUcee00xv3JnyKaJu2Bl7hp8ANR51z0AuoGR4aV16timozug2/oXj1ga23hA5XPHnSd5jglbHz
Vm33X6jKbexd+mvr3Ecf7KedK/BjT+PLaZTSasMHMtR6tl643iC6kqvFV47YTOtBOGY/YNlz8/+J
yWJUwwyTiDED0eHrJgtUkyDoYrU4UpTU9Hh23Px1gf5Jc0CLRLhyOA/6WyE++Chyu+6NExXo3P04
nHe+aMSh8AxPJ1GRQj4uzts+HMM1vNwplLZUN8eGdrmi8P8jCWJbpY6/+WWbKayaNuvkyp+ru5oH
oc91Qd2KUG6z6bcMLpLo+pjdLtBrBsfWJYJ3JWEc9EKyCJ5vrHs1pnbC6uW/vYd1KSmhq8H2Dce5
VhDfWYuvSl9w2ytZSwQNeJ67nZ7L9ZJf7Ux2D61fLMietuDg19e62DXI3m1Qlz6STBxgBBAohRd1
I7SdQAyfvjks4Qp/yKCsdkQv0XBFnNyDERQsefOa4PgnQQFrxejf/HDJyaFz0DQc0RaAsd5wT8Sb
evalI3p9Vme6YGkbJjZOsJY7P8a0objmcBNXeuPSUdQ2piJf34ZK6ytfvnDJOpNTyY2NWl+8ahv2
JBvuDaRRqwBJI6ghF3+R4J3abbtmKahXZe09nPM1cN3FtP32GoH4Rku/JHqv80Q9V4DUA2BGYlAX
kUEOYzUQwTyqeVzOpop+yi4rwiLTC7Ox+rqQPkYN1q9ofUFT3j455TJyAk87zYCIoxvI+/+T3k1E
RUyfARCT4Do+QUV2lFKy9ZY7HPt+mRQrkAR26IhHI+y1Cd7a3vJrtU4vl/qIQ2ClfopMBY105oha
09feVNKUvV8Zjr+DUQcy4W9lIo8sr5KmEW+h7xJwsXXlYWeA71tVTwjerjdZMcJmUdt2EwSlfnhU
uoJc1hu8mkmDSSgU34hrnfig0Eci5snSlpRw2KjdGYs0AMViCtsmYrYv+Lg7kJeek2/ij4QmcENg
bRMwyAgDwzrDSW/QzTebtdNLitiERZib3vDd9VTdcFd4Vz7mCP1GjKnbNwho28k2cQWxkqPukm/m
vSrW8MbxBBWt+CRiW5T6awTtfxbiUPGFsM4gw8cKi/Ti4u0RYtghljf9YwgZwlYqBCTHaGfd6sok
WrigK+LfRAbAkw4JMftbJx55kQ0qyubpbqFiWJrVaq0YshuJa+i6SwWbUpj0v7skxTuxc4peLrpb
PukgzrnCabFNtEAD67s5QqllrLyWDTgM2MrcjCd9gn2XfauyEIKMW0pu3hfsNhaTQqPOvU75v3Q1
YP3IprSoL4xy6h8wJfeT+LVARxoJUJQ+NSmaeGG/8SG4QXem8yqC+0cr1E9e6NtRF+XgLZa34mgW
gcEU1CV8WgSWc4iKiuRmkJ2AfydblibeQrk16+JMbMIz727WIyIHztvnzmmn8ce91yIaCigb7UTI
GBOozmFYVf+iqz0/0bX0f3dI3EZGg9oKKIHoM48ff67CT957YEX0QSZszRYktEkgftdnYcB/xy64
cScB25i+CbCfbGGoc8sEQ02VV5B+fkM06mZi2FwxwzyFDmKhV/ClO12H1m/KnP8JpgpByms1NNvW
oiOXswKJgQ3bvIrNHmFneV3tzXzwurtPqY7emrgL54p7Fnm+nSJ1z+jPbAYJG7rz8flCZwkvaSfu
nV6ML/1F8GRMY4m2g/VYty5+Q4MAmA20iW5+lrn92w59oJPqVskzVCNyaX9n+ANwVhtVRTFtJTBD
ckuj7V0VzzeAPSIEVuurM84XQDpZY64hHBbK4sAUoqKV8XtD+0z3Bxkh9N76l5MpN/Wd6uZ3LqdQ
+IEjgH1gFQ8rS7OgUhlg2is9hgjqzOlVCnrsIU8nIsUEEV3jWyzpISS+RXBzyTVOGiZrdOMPTndr
o3iKcF4HRQXFeBzVKfos2tGN4qX7XFcTo4qx8V0Yme4D1MoO7gIef8eKoRVPmbbLeLwFOVkgdng9
K1uSBBT2C7ZHU8HzhH3S4D5kwmfvzhltpUE+zjVtaa6/3O6bdwRYv2BDx74jXrBebir0c/EtM8zX
x5yL1t0pGkiHkNBEtph7DV1WxRIxYykWH5QKrgZBW6PKFKeZb1qNONJkGsucrE7D1BA/jlwBqQV3
Zv9BMYMn2Yf3bMXvNmTqL7gDoSRSnjjsAaPlJvbL+21gXMRq3me1+PjzAv3bMMNNX2+d/tOwfTNL
541nrLBwzvEgQhGHKfrEG0tnFFd5vp1m3w6lbeBRWNqz4nvdvq95idbcccTcxRb2uVhJdUrV+1pA
xG8FjKzv5bBFADez94fsL2izxLfypUdgoJTjz65sLtHNT9CRSb1SYGMGB0Xu4jsHoa8mq+TTHKxK
o77+qmQenYLxxszXhvgAOWofs6V/JUHYGaruPWl3JZlIl7MBEqMNOA1oiROErLtqvDTurDX/2dMi
fMligMtM70bcV8XX6nAELM7Jr4A0X+cgHSpFCi8upwjJwPltaqpJow8sfprGFTejjxzLJjfEVWoT
sgC2m1kCA8NIbpckiVvu+aEjJjzDIFqO6/dhsG+KEEQ3nnj5iXxaupcTOEq74DFTsV/b1s77HthT
+3rfAQpTYHgEotm0N9MM80mPicCmF3hoKyw70xz31J+GtowRgl653mH2KmJdwD6avde/Cf0GrCc8
55Z3yn54qg4SaJfbCoZmGRYbhyfZCbhJ2cbCFkjFJJRfRIt0sNaVlpA+7yHvLUNs51Gn8n+vBHCF
+zccsRm0nBedEaLRo7HMSiFcy7EpC99niEFquMadjAzAxx2QFCju7nxmXhN1lxPHqhn1+z5yH6vz
jRtRq9Lc1sHMkSqhH8qdRvGrmeDh2hzlkLVbdN5HKqRC04UkiqWpIwXMJoyTGIlqXUz7ZVfY6jKe
Wu/Z4lL2/JFdu+TvBDMZM6Ov/G2OMYw1wBh90h9Khy+3tiyHllgxtLRQf7Ut4oGDE0Ie6pY5eY+D
WMJHMWowvaYsCwkhcrXxNZgaHV9kpfbzsJ/YbTYVspMFqE67n+yTJnva4xLnwkrW2ubXX8rQan5X
dskzZATm5eg1QmXgtG2AnfZUD1Gf/eT2DRUi2qY4oJqJ9fLqN2CaXvqnQr7A152rF64D6wZFhhAX
uu3uyrMTb3m2JDzCSGG3Xs37T4fkS6UqGXsDwBnonyG7lwUFHfztMlzWomsjcFfLy9Uf1e0FGS0e
JRVlRppXuqxAuGAZ0uKcEAQJV+OsmEOxfuKHxEAWvH7gLd7d2GbixW0wnw6DfEeUafMm0GiQk3P0
08m03VrW+SVk5y32tokABw0jU7Gqb5I1DzXagFPhn8KEtDAFq7CORuo0I3gGg02v2ZGULqNUag7V
tVSc6B2P2hqFQlJiHYbnnNo3xTu496Xf7duMG6YK+/gODNk6gFyD++CMrHPDn08k4wq+sLj8lUmd
YPuOV/g6EZqCGe/psMuc8hXyLQZdqHlkcf6OvkuRCFn7ke3b8BDeqShhXUSwgLaLSzFzIcp9HSYy
HuqdvkVWyaJkIGnlcQKCa6XIaUvRpsrcSMZqhe4Jmtdnzf2mhI7/X+xgGf2/vl+AZCQJr/cggyvW
GNZ8lRyzWHLoMPjB8M472geeQXGgMQ/NWjV2ArpMC2+CvaNzuE7oCbSLfYH1g3vbzDUub2PinShH
Nz5j4W2XoMXW2EBNSp27Kz1HhQqaZP/k56hh+XwOiccWK3/kpJq+l/J33zOJZE9xKteNMnwsMBYl
EdO3IWobOrv2/Y7tToIBbp8QFt8QQiNA0zBaJkeF8EPjKzUCS1SM2gkkM/LyiOxXiFkUHjgWUzWK
7FsqHh5XUtU1KZjiZM8uclr1RxpmOhikiNU33KMC/O/DKGrpITd6mQjM+UiA3VxVYBB9Qs6jVWEE
YfoV0a6gHSHpk35iVwPvMJcbBRx2VOi2ZNlsxrupPt3O9c1T1k9jlaHQu0p/IDvTHNdGXRdl7cfD
UDHSvygZULMo0l0GjQ1LPLu2GIYrpquHqAPsV+PFFeYC0xAPqEsfe4zy4psfaDVyh1p0DoKXHYpw
vrSVBCRPG/XCS9BYFIyXgIXa4WQyrFcFi+Wa8wwxOsq1I1TmUXo09+K+VxPfNhTAx63eq7XfzHdq
x3cJxh1eDyCda6GhDIdnOOtJJrpFvft3ahipphx7BA/uo8FiUDL2cxgcXDhwkoc8AJBz3M6QTm6C
V74bAO3W57+Hg/5x9Jy+KFBbMKZLwn8wNHYb+OTtKnAwk/ohd4xDC/YharzRfjyUYHRJB7hgWpJI
kafG3DBwSXqpxBdMsoI5wqh11NaFwUUmQxiftuOZMcIP9+filn1a2LllA3zHhz3B5ywQQv8KUQwT
Lerg/lkOt/8WqS402AdW0P41ekiU5a8W0oER8cv53kI0LN8zA+0OYr4eJUunlVBuZlYDEji0UlKy
OgwdG9VTdxUVmBoBV2OET0x+F51sCQXvD336loCKj+Jfel85E+puq+gtpzK4X35WNNu+s4eNfxb4
/sqrclXQ/14H/QnV9ExyDE0sSQxIWXLPbg/H6KYlp+KcLjLbBjMuVwJ9kbfi3DWYPAPpGAx0+cUh
a0FoLxv/2oJBVvI1TOpIdhLj5hW2XzObczUdRSIWRYt7w0cOvs93QoSNTfdnZhUbel/XuWW+1yrd
jtA+NkieJ5uKRVM4rkLShXfGXXSWwE6cWgInSrHMxsbbA9Bw8/X+RJZv0/B4NRyUNeIUr1YObDWe
nKAGqi4R8Xs1oHx1GyFSPa5KU30QfSXwEYwIFgYmgG2+zbr73hJInKi1sPkm8cbPBS08GrDb2kfH
hqgEK2kF7VwGDACrZyCMaZmiINGRaY2zgMG/p/v3u0GXiUKPuqIv/obh8d7GwPOabw5QvTc9cZi8
ifG7YKbOjjJ/XEUJtjdrAuYacRV8GAOAJQM9x3v5jrgLH5LR9dO2TtwJIm2bG0sNxpWLL0jdgx4y
UMcN0qfUotgNdvuhkjnbYykhvnVxduYn9P6lwKHUhBmZwSdLojlqeaJN3R5FlMiVM5jHt9wzOsPB
EfVUibngYkSFquQ/g5xNi69wLBmoo5+YSoBCHIRA9TTQxMba96PheKSPQj/ToEB1UWF32t7nm904
z+av+2aBXcbNgFTaXabOu2wN+EHvS4zFeCQ4Wy5B+xkZQ/IhT/VFbu03ijN+xmZB5Pir5RWwbDFQ
Kxc7MjUNMEwFqzWsBcQfeuys6vfsatmMZGhPOYCSNmzRzfFBrTXpcO2FZ5L2f+3fLZN01qQVU1UM
6c34e92+KHsrR1Hh4fOOkpzngD8ANnvU1RmD2H2qsBsMkP/VsHzieD9eK5zPI+K37PRFoTPV5DGn
5JF6DMmuIgknsTUJpCN7WVUB8jtCVYjFcGfi4aWOHkznjdKS/ARj8lKmGwXtGl5vhWF3aKD46AN4
KW2PvkbCLgH3O5579De0B3ccfwUSz/C4P1ULpzg2hqPYYTne9h0QTnVIkTGhy1gHZ8NbjnZFfwha
ui1PG57jkP0Gzg7RX63WIhxSqIboc8uOEhQcawlBS775HnRCtl67xgBds/jPLGXh44Ct1JRf5Ls6
qLgl87oWIc/32CpWyA8bc/hhp6IbONCdTEKrXzeB8Y9qheQgLgJCVoAdEQNWZkqzfrlsr1WkeuQf
nL3441c9SS+i9YhOeNrmPzIDRjNV+Z4SzPnoC2mmSI/ycY4s5q6AX0YEUR8GytvZwa4PkoQHdJfo
lzk91MXywoOUwwwKzoLPV0xwqlrpnb59Q0TMg8o99uZ44pRZQxz1b4XoiAxjuYVrs4yOD/FXvXUT
bOzRl1ccsiIxSEZ6W6ImzLCXb+MqRGSVTT6ZDn4G8MKdpU0kkT3oWThrRCLSgXnSFTbJWwlYrI5n
kkDQky3gk02qVPgZhSclZvIJUaJt00rV0PV83OwfQVCSN0rHb+H5N4GcoWeZcufoVP9rzHPQ3eIq
sMJxc79wl3am3CLj4OuhxShhFueqoJ/E021IVEyEdOSYbLVpeoUo86GTkG2P64WZPx6gtLfIHXtf
VEHITWvuR9OK7R0DyAlVNy0s2SZPE+ltj0IaqJLJq4zfNDRWQrmCx6w+LjhAX1F/vOJO6/aSUzaA
GW1eZWTfr8nqyXUl4athr9VJIkH5riEhil9yFX/zuyIav0plQeS9c8qDuQh8Bo6TSpmu2YOU2bq1
2tmjJgPOpovOyPOaTwQjSyTm0OlGcGQjy3BZ36SUYBZ51jZGYDa4aLnNSoiyF0UFK24UvJgC5ulm
hrodLMT9v+i8nxilbqbTgYUfl+RT9KTc6Y/JF5eVLh9DNczt7o8BrJyttS5u3aaF4JMY1YKMinn7
NN8mwVpOLNpoqB3L3SND3TFnqWEyMRx4467W9E6RBGjHeaKnFKkzPFp4x0yzAFXqtoczGymx4YOB
SaZgUZ5gDqZokaTrACF+dPhc/lRkBJD0h2ddI1zTypjEGOWmXh0GwCh3eb9LX8zsmoLWJblsd35P
UQZpXSv8k9sLthoyB7V/yChuMZJicqxm8QSVO8PYpJMS2bp5SF+3MDU/h+Y8aFmKladGwMRbFUqu
XVe/LXvjKFOflUQn3d/Ev6a7YeW+nkuotKW2Edt4NJlo7QY8tcNtpzYU0SKyiPKULF1fNBLBMhcu
8QOsksHvtnhs0tDKeUVL1jcnL2mury+ZaaZ0wiHyIEZAdXOZKH4AFBxdILCHxYIzKEXEWf6TZBLN
hzxYY89nVp0W1ByXbfEQVN2XKwO5QAKekrStoX021IBLvoOx40eAHS3Kwa8cM4S9/z0VYU1hivY0
xvLNb3at5QwRNwNQ2NHJoA5xC5o+kA/wDlJki2feYjQNYSr3fISRjM9dI63uuUz9XmEDyy/5o2oo
nMDKXK+wPESB3SSvqd3VbfxttsMhdZ2qokFVDGEmke+YBExcC3qfA3cYWGvFzKLIpTnVoSPqB3kw
F4Vz6zBfM8jgbXaWEs/+gelENozL3eoAEZa61wwUMga60vk2HJY9UKUMwcbtsluuOtx344XMBPMN
iDGSWv/UNEUF6yF72cc5d1O/k5u4s1Zu8SEWmyMXf7058uJ+vYJ2fszd066XwbqsWhpNfrPwzgVk
voZz2pXI3dBKm6f6Kr5Pz5m5rmQKsBJMJCQzE2hbgjRPCVYFHVpCYOIShAqYpixfAjP3/fcxql//
IPUsKAg5zz+19W235KxHmw7mV1IyF8mLpn+8uAD+e1oV8GGcnt3BfBZLqyoly68waxTU3Se5Tq7v
9a2t251t4fcLNAuK9j2oq1C3uvAZvDEdK9TotXne8aZly96hYQHAgQQEUm8t+ul7McaSe7uYiV/+
2PJtvWaumXhBA0TYG9kaNcD2Z/uHYxIpB2y8GsG3re8OA5z/BT7/2nd6GWiOcRdUizG96JX8+HsG
sLkxXinRNWV7tFHAiRGjWh5dH+1evJ5P/tkNloRFHpWE6Iv/eVPZ1UpD5+dVZyQp7Yecg3dWxOiX
L0Pnj5de7jgDCU7ddFcsTVREnxrm0r6P+rclQkVwqSutihJEDhjpehb7SryDQo+A+Oyq7hBkiyE1
zNqJUGkxG+MsFtQkmWdb39Rdj87SgywhbIHkOhyD36fmZDccjILmn3LJHdP1Bfm57bd6Auk+J9pG
4Xxkg2CQKsqMQIdBo7p7UZhS/znfRihysNYiE02O8zcQPT7llZeM8e5VSCFXJ96MQxnkZqEPoRIC
NyQ3pO68mTQuK1PevC632yfvBB0Rtal4/RiUzs87StmNST0kjgHO1CjsCS06HwaNWf3HMdtSVT+Q
0svZxT7vRKeJjbrIZYE2FqjtNkdTUexNQE7KptUvGgFI07nDZYsrUsoZWQivpyRYxGVIKmFNxuKr
ffpawjazsT52/kVbt6JfHiqBE/RYvaW6sTXKGqxffy7UdC+jjUoiXQNMwix+W7Ao6BCiUe9WVjcQ
nZFMNcZnbJSF3HrORF8WfzdWfIrMp47I1FWabIYVUYrEndn+r4wIFS1v/n22YcJp0mHYTi9oI2mA
ICDn+LtyXjhkmFD7bIU8ksMsTIjcY2KHUwWpDz+83IB/hRS+vWhyyuWbluzsac+ep5bwgxBxOn+v
tro5oWIXzbNj+BcMahN39na7Z16dB2eIgt94WRNMksu7VRRAJCkewl2DRakO1QXaikbcyd+UrPB4
CKTghChc7ObdpVsfTVrxHbitmJvQkDC8wf0PHkyMuqxr00tD3Vumhmjq4e44gi7c0DTs7PaUOgqy
Ax2S4XH2YEX2cLLlOFTMl3RpoLs25O4s+XeCgAMEHT6w+ZmGYSn2WvjCG2J0uZkAuCkcd8n7TuyT
nfX6iKWaOWLm4TSLaL7WirKYNkDS6a/KUlfb2N+XLz7aZOxresnCGHSHecrP5QkSmurVSUYhIbuh
4iovw7+rKYLi8UV0trvRGMkqYrWXdx4zkzKpe4WDR/1FLRfiHX2F65LPYkq9ojphIbWgFmGSZ2Cb
rvwgiEqW7ukDDvVgkro6bSnJToYQA5/rsCm5ZptjByiGAsTUrlXHBH5zgFRjt/NRExNHLenFryGF
QXxaIBHL6yGPJRBqONfZ6XeLx9wtQulPPXX7ZLidfd4vhNA18ZMCgnF1QtqvFN4tOIRS/cZPQ6q0
aduno2ritfnpzmPYR7vkbQSvFID0adrx7UQU7NanV8lO7Xgx1lLYOsmhsf+j2Qgt/nfeac2U1Cxg
Br5zpSbRVsfrKGlgLWLHQ0WMeeii+w72l0rHhoBwNJ5VyszROwy2Wy19QltdYt2JFl4GFv+iGmbK
LeMMF+lFp9CCtN1fYx/4FLNCWiD+OSQlY3k9DWXiiOrOrfOxobqHJ75FAAU/F8sbXPNdWdI7xtnT
aDyPE2BKFRgx6hHx+CdjSOr9LyWAWXQbzIGKEPtwJX3/cyDeBnExd+ffnHZ/XsjqS448t8ZhIf4p
1Fzf/DSQqGl+EScbZd6TeA13ojpwybRe1zmQ4G5NgmXVxcTjkvsXNhWohIBA92aCFkDfdA0RWKaD
wualtdwAc9YmEKR+qq7NWHJA8D6iCG857hIreEDqGcRy6gC2J7ZkTw3VOvLixbeyn69FwOl90jon
4WUjLurZp+nllaicxQC2QxxHf6T4H2BpA/eyiCV2uBwTJZEL02h6SXmakg4aXaBiESy6xZW+5yTG
ZYawEFIVI06hcnD7IBnIuvVLIUgOJLCmawuS55RoAp/0UU+1DoNRA0kNKV6hldu456TaBORHotmN
G3vUhfEHWerCMdHwTaCJhcKxXpCiC0iurUfGF2LCpCGiuHTl8pnHzUrSZaLEIuhnR2aey7BLTvj6
wApDoH9XT0gXHtRuLqU5AkFZWFoJ1SE/9aWSdTCY2sKEtV8f8zA1hDxheBy6aeHaRk9/NwuGletX
AdKZtg4OcmDCMQALF1DbIn4TDaPlb0xBrdyY4Y4pEzNfMHBCBIsiEEqK1t7qT1GLms5X3nIvDhm7
3Lw1hB+uCc8105ilNmBh+x/TVGM9LIpr9w8veJwrBmuPWo29wguVSufenWLrjHI37PA51Z6XfEVx
ES7UC38zYbMYG6yFy8wZcjMk8QkRVDmdv3FU2S+d84h+EvONu0qGRkgXhjGTWkeItcqs0tgTCezp
Tz4Cdrc1D/kXsiPuLPjMSbYzu8wkkwQ3iffTSgk0onsDIYsQIG7jIFtZ2i/bhifnKol8pqY4kmSz
+HYhL1Ke2th/r1zOJ+PmM+Wx4K8vGksNFlJl1VHQpFXac7mkiHTGkHe1wlxRcvCI0LWwfdk5de6T
6Zipk9AKZK45vzdK7cmlUHoSUPXTNTef57mcjz+HOdGYXWj3nc3OfoB7Z1tyBBbnjhe+c0KTwD2q
0jTDDm1vrIX6c2/SV4da3vL061gTUbCuRIaSucxE+TMT34VkY9GPBqhXTIGTxgYsKOTTo5uLBTcx
JcGmYDg1dFH1zT5iDuckDBrm5TgmIWkP7hdQj9G3B6iYqI33RMW20qUY5NDHuBVlhzCriHXSpCef
WNkjM5OoE32P9PF6ZIq18QsAieOUxffbsIz+QEy8Bfe9yMyJWdtSiDDBphYZCTBBwbAMD7hvWAcd
hAlE5ZnQvzEYgXjqziFVlugFMVo59pB5SImw20o8jeig3/jtvGYoQa1fei4rniCmNK/hRU5WsSvX
RfRIYLfgEpIJBLukHkV0FG7r+YtxwdYB/TMkVrLA5Z8JveCrDbxmEcMytN5gB/XDBrENsttkItLp
jYR+UZDvekCRZto7FghEBh+BBPqoC/y7d4SZodrwLTkP8E93QehtolWNJ0Hf7+CqbKWuADkCZYLb
bNIgFY7q/5B6HsPuYMA1z3nP+PfrFCgrcBYrViiETqmbMqsJyJ31muQ10cF1/dZ5A6+DLuEFpJzI
dXy6AiOZXazPXqPXxOKxJs0exmBSlmeUkj8/QEpwejbnXmfrsvt8OzQLAISwWL/zFx+x5K+XCEe+
n9P+glHA1YTBpYlnDgzyNDYas8a5UtGGDUZg31Pa5HifwocmwzNmgAFztQBOH44i0nSFoF3qelgV
BOaS4e1DDnO8+AAZqLTfYrThU0OYQE0+rNo6MLGC6ys8Lk/0pvnPVK9sMVJLlrBW8zZ/ATJveGRQ
4eAyccvEjg8gLFo6cylvMY/jd9HKiQurZ44SX8eVjym0T983kRXVt6a5Hmf3/WCvj0GyRXkw/am9
JrJwVVqORZc0Jix0Qi5nFNNlIa3/IMmzQAMKBX5sHFYTyf1EXvK8KrWB5yC3xMNagBRsuvh901Pe
kAPQ/TgEksd1Fe5pOQZHrhQb2ZY03544ldIc1JPgC1JaL9G4Cf9K9mOsD13uDO9O0Z5N/Kv+4nqX
cRX4eVJqI/iJDXXY/JgufBmHNZp4b+cmiwkczANg/c0GD+JJUEIvaK3y21a8OYuftfWJoEweq78F
eKuQXo34DzwmcN7lRlAz7KN6em3XUFvuDvgwSfdTY4LdN+vSN3SBy6DePB7GMtNvp0yQNgH/D19W
hKTgxKwmR4vCM14EdVkyLRN+8t2caKjnWmToH8ML5UxYhwZGcyYUr27knWSGP2d5vMl4HO4y86q2
V1MKVK/rUL5ShZHa0D1qeRIIACtwOZQTIGjhqPD7khKvC2e2chZbLQ+lNtjGwN1sEgGXh6N7v/KO
yflmV2xt56V5BjiJ1qOYzz9QHR5TFV1tdi0jWsfsB1+L5WRBFkNAZgA4Io6gKnbrmB5WhDl0AV22
sWWcuSjeJSKJNemBh+wR6mwQnvSfBBVrwHBbR5V51atsK/NNmKZhacAo+2UPI6lW5vAZ+whFurq1
jog+1CyYil8aAVDLIYlO/pUJuqr7jNJqvwP8sUvqj6GRE6qDgOfW8aeQZHcLmp2vC5RFveB0TU9c
uUfvgsCSFsRxnoCNDUzL8AVd76BoNwF6Y21UnngmI6rvI5y6rwTE7eG1a+MMLojaQOa8RT5K2tiq
jCtCVOfz5tIcVSkCrbrFeukROrJ3xcGdl9SvlTPtHvxSpCZftgjzklbFGLX81eoLxtdPoP/85wu3
bosZlciaZBTJi2Bj/+QqIWzjs6qlXzDZD6upCfySotBNqz2xyZGuZ+axSern9Dt+k2BTdkw7Plz7
RFmXAPzeIZTetg4JThut+eDd+2zlnu5lELB1XJzNQv/1WC5i8/hEtmJKzZLf9xXkB2n1MNVfvE2a
0KmREy388FM/lue0jcD/0UUb/nh/rsedytPSY0Jj8uqR5jyJqlgbm0AFOV1XKKsgtbGk5ScSR3Cy
hA0KysrBvycUHFB7KfL1HqoF2Oz8qZ0oS3kZCCdxEQwhPuxHrksojXDevzUtxzqJn5Z6vG59Ua0W
LjYSjDoP6OQAy4gpUirbPtV1PGPfmpcHbvKAGnihJZaBwu1pHjPeN3BCXtydhwon8H69xPVvSf5+
BdC3HWHjZGSV+vD0mLUzeOk3s+6P+Nyzsqs9UmPSZCW3j5XZLZZJ5MGJ/T7eNDhlcUntp9LzJIHJ
+OlviBkWQJdWSTFgCOWwP+vtJusirLmI7B8P7nVLAEZQW0PYf+VY7P8+AEc8/07ux6i1JsA83GxW
flADGrQy4uxFZa+ZU12wyAPPz5ye0v6m3xpx7FIEsbss5sD3eiBLOmMXPvxUep8KIXqsS5MKAy1N
qSAiwq8Jhvflb9IfTiLkL1W19iV5f9KtWsQe0wtyOX15YbOT93bknxdvnKKPpd5JAwChlHzOt8/k
7RiJIRqlX4CW6Ve5x0k/2FtdPypbcewmyLyrJNPg0TP3Q4EAwv8cClWdB19ONnl5aPYRzcOlVEV5
LA0Gx/IcW2g7ZNoKuN62WNMPsBYzHIe7dKmwRQjzFxMySRNXRb4yIfJsDOdxESPEFs84io8Kmsmu
8FQoq08g+ey+JZJi+0jJy6vz+Hem/a1rbmuqsNauiXgKl9KFRPCnjAcU8ej6qUrTt2dY8c8envLk
Py7v4i5ygVe13PnF19L7axbd4NdgYoJ/dOdszLVQObgWyoNu1obAjgKE0opD8Pb9KtsNM2RwVx8d
wbpz/QV+EAiwkMn4TDfC/vk+3FQOXLK3tpFzRb8toepeQp7XFljEG5n0YGbd7lPXlXPcoOk01WLf
/GAPQeYUbkFAC7UcFZaho60tlI4wHGi838f2EOu0YT2liBo/ZCrf0k5yeUPIWuRygpaX51i20DWM
r1ViTZZZJELM+Cty4vg3/6notRTXEde6PIXD+HxlY+PE6iOJEZunMfIUCjmpT3GLZ4r3F4CublRp
hmJzAXr4eI98wICOnULJ/1bRkurbUpOhhe5c2a80mAo+2O2q0qt6W2hyCYntrvSTIfbGs03xugNe
U9OI32qMH7yyitTuuFrfG2qKYY/oW7fZGRvbwpwv4VeI9MqEeB/zS2Z+Z566N0gruJpylcPwMHuM
mAIPKp8iw8JU3OhSAPC8aXqmVVvy+wjpxTNusHgQLgXbCGOmQPSvcT+Tzf6dvYF0sTLObE/HvcYh
x3OMWwEeMpSa+gEd2pGQdW9Bz1KGXwjQ0iInNbySCAXrboyT6jxro7IwN/gL17IjQTo+BUcS/6mt
Gatllo2TSqQDknHESBOZfEwwif2gXeK915iZZYiHWFpOw/3jXh3sS+J7P4cmEGCmdja5zhZ2OAWm
9HD8Wr0GJXD510ZIeWiNAb/yMHAIdvzaFhwhZ6qf8g5WagSg3OAqBDpop8HJ9IfViwx66uvitJlA
jTkPg1EOE7hTYKFd8qGKrC9G4iyq6MuTFfC1D2orZZVUBT2Ud/hWKB7gWnscp9XdlB1tM0chPPF/
2PBD4XGkSLpAsYl1/gNQmZz1R0I6JxM6wlsnRuISGK2eX51Idz25HQ2p7eOIaZfudPmI/yoCu91C
f+8RKcAXKuX1YQzZ16K6PEo/tu2T1PYGgCs4SKJUIRuxZmnhcqxTMf2fRjugSIG5PPVQKsitLDDr
btLLyYr63KlZmzoEww7eRk6Ans/XGH9pjNjmiTNsxET6NAVs04Je191twpLV4K002YewW1gaWR1k
Gi7WaUCXKjSPELv4XihAFe+c4tYLn5yvAD5DmuhSMRAL4meQA1wO2tZKxIKQorI8dd5JxzcxAjrX
1mCk8om+yAvH9AMDEnJVWn1FGvSB7TqhvOjpnXAS3rMyb90WMfW+TSRuzyusxbHRWMBolSDL7hfG
/7iNfNxNKQ5WeOWztKGxnxVPgYI5kBv/lgF3wcodQX/kL/LqDIu9cqcgKZON1Gxamfmf0A+MyrBj
pYRjwp+jMjYuvA/E8AueJ/PUMK5g4E/TpmU15gx/nMEUngCYHKFBGfvW6kkICwWV7riw8fGxjxyq
sHAsArTWi/GfaaVwBqTXwWo7G8LSeRvaFFAN9nZie0Vzw9Tczm6IXFTCoWsH5xyuNChCTP3+BFxI
6gwhE/6aCEH32kE7AAasoIyhVP0EOTGMOQl+a3HW5jSaN/ytEnre8FaFSux+sZZQspS95zOvu8Zo
BgPHAPepPbjj/PvRGjORY9VWptNusjYM18AamXERSTWUlFhGKEBjJ2YG7fP+cGVZRjxFY3CmhfW/
C0N4ESPBpRyYsGw1WRtPXoifhxzYVrKKwzjatmfvT+fJ7IRlyeDMhyyxfLX5AV7ZOaINDoxMgVj2
pzZdaktYGCPvwzPwleuWMZMEjJSO3lq/YOfX1D+GKePba5svJPcVcIfAAwVRIf61VXmv2gO1hWi6
ouhV1tqSFKFhEbMe9PO+vc3drO8MtNUq8B0ISMOM5QqBLKVVFf2yzKUJJWsv2ShnZ+DEicgmtdYb
Bgxaj5zZDigZNbsIipJpv8tLXVI8gm9K0pHmDf7J7Rdw2xga9gDLxaV4VunhMGaagwQDAvGVqaXJ
s8qIkEc1TEoyGh3UrW6qq8FyAbp7glAPMahWfaH+VqhV/z+FAJaQNpfRb6oKM/w/LGh3Z9Bg/6nh
5ZPaa+uOXN2qc9Ru3wQute/ZvMIi6Q3hiOyvF7ATUQAjADDKdy3ClBDu/s7b50b5TT4Q1n0VcAni
sE9f+MCgG8VGumJhM+EXF9GKvuqVoUkU3h7kphVkeHUxHTVNB2gJrxtwRBZnN8ju555V/7dtsqRr
Z+J3Gm8kry2HKRX+nuwF4efUqMszeRlzyug9JbrTekjpdIeCHj+A/6PgV8QkDpKRGqOlem1CRq3z
ThRGbME2nJ/MJFa0/GXtD9U3VRDx0UE5cQ47OsWumBgV2BWsRNQaDgjEH1AsShzC5NAcVT3xNsrt
7sUrO2snFZ1/MyYfpQRqSca69My8UpRfSey/nR3aMMinH2n//0TjmIC3iJF5skX7grybm4lx47IK
zanxBZ1aWZYyEXjBhgSH+xgsX0G2rK5NLQEnQDEoa+dI0x2IBhpxm25Xiqru39rcEUg8wZ6RHcRx
XbGYjlCf8IK1aQsacI65qK5sz1pMmRlFWSJxrXLly39Awfa14jshAEZL/+iKOLaRAioC/JH0b2Kg
34lP7mvaXMe4yptCq3fQsQpYHrVG1ZuxlEBnhZAyh6tGdOrCILIJeVXvbM26Xb4yKuLwbCFTFT3f
f/Yn9MqFw8LRhLPFuaw55+W3IeyJ+Sf+tbFqt9GLLllSX5CRNO34n6Gh0x080vx66ODWmZu5NIH9
zNz8iySH4EeJGbMKh0pVpRM+/Me2lb2An0AG9TulJ3TRfObjpoDuKJQLZGAO/mRWqtRqSYgw/xw/
RYosTVcHwqPXNjCuLXgtt1uYdZKVoEQVudncIHcMGUjFABEPAovC2xVVJBykE0zZrXQW0aYrVgu1
kDfX+G4KjkEZuKD4rpmXDaY50Pa/wFprbj0ThQVVcpJo/DkGLU1uqc128f29UOToWWEJcp83ySBL
St7wlHDb3cAXM49q+vbODBQ5ibyZIWpoX/b1+9M2h2S0NUst6jZKnUuEBYSG+QwhycxiHWvLwich
1u0ioRxS702WLnGafZwzuCNt8o5Cz0qtc2AExGM4WnagIF5k8204EDGB1TwmTsEtoW3nJ4RIatLQ
SIJj4i60YL8Ev1G4plY9qg57mALV0w6dQWu5UDa7kJSmTFcdLPly7IneS0LyQimDfZ63VB/D0zQl
rj1trEcA0KLWGtO8H5T9rn5Onhmhoo9eyXpZ95IgdEoSnJBIm1IDYj+1ghy+HwBE4u4K+gub77bn
VuQWxqU7Gv782p8uAJkO7SeX+arp73ZmkjWn5A5IsIEJzLkpCeUBQKBia2FxVUiw3uWUnBp8SWzT
yr2Ib//FYT4fM6wcGIdjmZk3/MeyXeDVPbaGiPcs14StEDgqgw4qXqxi1o9oxbTnRJberMrxAflH
S1Sk8bgCy8Dl1YufJ2QBBEAH/qvqus+eTLrChPF0rOwMrZm8br73/rWUMenwM9QTPIjhGUyvVk9x
oBHnIw4i5tcBkjAQ5L8T3KdPt9x8zFo56JrI2mA+5IUkcgoesjNw+ak0xHVk7KvcX/457PN4NfmV
SJuTHrPK0CF/wZEqBj1+j7QCFie2ka9tI6j+0ixRLsv3JMADerzHjVODhaZH+iGbMNsAGMPKBIPV
lg/ME2xBh+fo7AtL6PxpmrthxXsx9EXQREas48td8TN6R7tpX4xFY2QDIfk+jNFI2KwLPJ7r+yHT
tMHJ+wl5RmluvyrVP6LmD17eJUC13O6zVaTbQqqh5DtKD+nnnNz1IGyvu3EfEn5MFa4OVsDpSW7N
gl7F/JfnATUcyvc37MeTcjhKTS9tpXmE7WBHeeZU1e3q2VXTTJn2L6Nw1JF8HHk6r5KygG7HLszt
RPf0jS45XQYQaDoMCf15zf6sc2+HwbXEuZ42KFdtnbj/ROvzX/MZHRGAmayLxEaP6zfk3mxp6WFJ
nyYXzuHayrO87RnzjjOin5EPHgwISuNegzLSpD6QcTonHf51ZK5N8Mu1XVkG2jlu1dm1kwroPM+T
Z3KyzeAvR7AxhkoSVhUDKDIiIFtQJnkub2bXQeVUvbILSGV+wkH5JAiFCjfIZkvljT4d9OeSj3aE
Ts9rosiw/ljbRccfrEwautKKMACXxBYPtMZEcT+saHqjcIgUGiQOge4i7Xtd0zN6dB8gGcNSkXwg
yU/SvZCgh58XVeKd3UdNNGiv/E94aOyDb1/wbJ9dFQ9pnJWlZlSXzaYadp3jbmTFzXQyCo4gbPHw
1UMe5SHSxPUOQ9AlGvTFMz6Bycst53gDtHoJusDUq1VSZdpmyk/hMTx/8z5IF+v6ONJpWx0zAn4R
Qz18Mu24o6eAhlxpIJ92c8g3AQechsLdEewFX+QqAnRx50PHD/xCGOcueY5vAXZC1OvS5Wwee90G
tSGeEBHACIhdZeI5vqUhFRWXGHINbUGG4AampzJinWak84UXo9LQIWCjXEvjMUpYHzN/H6A281bN
nsQKLK4yE6eS2PEfSJaSoGC5RkvPolgETU8OS8IpUvonRnEg0AZp1bVlPPX5fW4KxGM4zoeOjH08
sj1frSoe9NCEkU18BiUUTpwrrzh4TcXrtNvhDWkMI2VHsjLiZPyAgzPqwhWk8WJV1eksjIL9Uyup
VnRc3O5Ic10aZ4UUXq3QsifBSVV1GwyXULKu6ZadwWe7dhOaIfGz8W9Lk9PO8DxrCFDOxcAe1nm4
tkUP+0go46uoeIJKa0Oopwlc4xHKpb+j4j7LKcX/WAW6EWL5y9qQnuWfRBMzzwYhVliWxr/opu2r
FHDFl0fOsaSnXst1kjLYsuReZFxuYqDs8txHy4WaCWsaRAUxGXAOhsLtY/Bo1XPrVdMGl0uFx+k/
khUUoLNizqApSBl4Oxsgz4oiq3oBoFtOTWrwfx+QLC9JdXQ/Lm36adIlYpe1gRYAT432krkUyrif
BUV5HNN6EvxI03a60oAbH1QxMcZwCDp4K7it0fi4S0s7IR+RbPT3Heg28r3RfcEN6cZzLWtSHJpO
o4z86766m9q4MK68EFBj4waVL8xSZ81DWiuA8H3ZsnvzmRDjlHSk5UXDUt2I0ERPQ2BskW4/NcTf
+YwZllFMa+05E23LrVrQ6fnS8bZoKy4+a6C6aKTYKJR3oZH/vRCgcPckoI0QomWBXE2QT5lE0z8n
Iu7r22pllEIV38BvT8p7UyarDglHPCwTKlDw1j/hi8ypUAzp6QmXflO6cADxVuD3AUGiQ0Z19hF/
sQDj+lhfXADKmhsKr/b6jdEP12Pq3i9fSLs19Qobhxrr8FJaLkqziPiiJX+3BiFWp0rzt1Xkdi4s
A2rnG/agmX6uPujirlE7n+8mGVm5zWIy/crAJjEbE0JqER9z5s2WaIWzJ0sLT3g5J8Rx6mH4ATY1
Jha6+6PeqmDarWbXrL0MfmmmXSCwQ+djuMsXz6EtyLMe7SZLWFaU/No2+PIXvA+yYAO4pav0LBBL
vvg+L+UHQrP9lG2YbGgH5zpS7y2jxthyGTcbxtnu1u8p5SJhJjMme2IilVEiDIGqEusN6R64Ecym
HY1SQ+UyBHI0m0k4aylvT6ejfc1it7PlxVgGU84GLyk4lT8qLqYyTJEwFfNCaJ0wbpmzkUVgkBnD
qb3/4cxGTGVxz120sHKc2EHol2GeqXC0UYfrOv7a5hlE1RrDz/Kn9I6zhfNDisEKnGo82uot4Om0
R5yziKOHWe5QCgKt4fsHzl6NV3ZxvY8pvfgmIzTnUYfOklXflCMtQBEu8xtOomXKuy6qlNcpWQlK
6fEoBYY8iIzURg4c5FywNOl6W+qCMkJ9/OjLtJCi/c7FwmyujLY8LP4wxE0Ucr+lHDO84t1ZKpoU
IqpbyeqxuvcmdTuG2tLDDnNjvT1+IhU447U4y5XgyOnHx4+K50LzVvrsJ0hrjHueRePRqhNAWJdn
fXR/BA1EsS4Gk6ZMHxG18jYt7un3efYUZSd6lCKKyh3gFFJUINcwfsATTUlWZMGOCCk5aNCiZ0cq
iSh7ADnT4CoxiBhMS0nNdBffvntpulx2AV05Y8dHFH8nRVeOPADEYbVJkmNlbbHo5fS7PLR0fRmk
UUt0Y2Iwmy2+FMtkvp1V3kNcz3n68gjAXx3DGs1YZCDqfoTmtT4PXj9qV15V3X3lWq/cl9D1OfUk
UU91T028ycan4z3YOG63gcQjYyhE3EEn7qeDFQ/K7bvpNQZhtxTCdcxycgGHjTiLCOmVM+aywn+h
CcdZfxpnk1PVvfFQR42Ekjq76OK60HtO+iL8btda3fvqGyQdD916focNRp1cBR6ct0wNxFCYnAH2
iqetan/CmK+O21kDGrFaQftPOCV6TAB8kDsPHlXZNjo/QnzKP/XKoixzfc40wFyICU2wHxCEvM7l
3KkM+hsKz2D4PDzLldBcU7NMifn74IdmKGfhXbqxQwRTeKPq7azoa5M6XLAFSXhq0dhpiwA6tD8x
Y4H590N4fALIliC5c+iyL4TsnU00m3qr/7l1mYpgk2tKBMChYtYT0DQMfrY54vPX28ADpvEIreTo
ezR3/Bncah7fNpp9hh75OUFsukifaAYWn9RXreSp13wchdhw8vSsWhMKhRTSy8JuMfTqm9sb/wty
0tKjXGaq4rcxDU3t0jq5jX5oEFVcySA0y+QArGD3AGZtVUvKt4WjC+Lp/Q2Z8xgiPLpg67rXDzO5
l6syjLjG1mXAl9myWGQeW115qtnxaltkfHdgcWRsmPqpFO+TGmShRfDOsJP6O+A1TFsKlheVX1Cc
ZE2MmnM8ucmbYQWRPQmB4G3Tf+mkxQmsKUi8dARGyrgW3/BXwD/pAI3979B7VCt1bOHqM5TYQ87W
pi9F9vk1x4rUd6/8Bp9J6Bp6I+LyE9DQ3SoI7xp+A877Kwz6mEiydbCw9zAyQUnNmEhzSPrH0+3T
ylHYCf7kA9S2O1XfnfRTkXfceeNGV4DnP4YtkVLVeemkx8OB3XxxPdm901B0aujiJbm+SMtP3qL0
fLuT1q+iT+4UYSRaN/oeOaN1bHABGl3aQY8OPI5LvzaXu2nNK+caSr/RnB3Zsq7uKIEj6Nkjeb6D
jAz/UmjDo9WCHYMUNPCGA523Bko+9pTZIWYU9TWIQiWru2IgDZIgbbEwGPiEf7LNlIhFekeysEBy
0fuMrr7nUZbeQNnnw2tQ2PVAYz4r0mVJ1SSCx+SBmTbnnPFVwTQrNHzgQEF8d1zZdTwP1bDEABsB
0gT9gxo0mfejwFAvAtnUPPdCRvHqO0OcTBhXkGC2lXutHfLyyqGwBZ4Bgha8PaPkVLE+ZubJwtJ2
t2Y3LWSSNoE9oVtHWBno9MK/1qBKM4dDVBjmO4tF/A+zDNoHX+85cY3wHWArtYcZrvvkxDxgOAfj
DFMP98VfW0mYETJweR+cMPCxcTj/6oLW9WICaJ+4VR+293pUISD8u4L677uJKuR910M+9mJnvs31
IjfY6XLFCBIbKnuGahX74+C+LgTdebXHH42HxU43ATRuTgBiYWbXN1XC3zd/vky0nLRjbKIT+ei+
BCYlKOQQQ0VY7AKvShohrVEwr0mpSJWfdiFS4BpJrUTgsqg0n+Jh9fviewcztQjia9uGj8uap1kA
LZbCjHmhiiQm6vNZBT+XbUS1kZmIW3lfv9e3e6c9zPBA6YtpnwJEDdHT5a9kFSBQghw5NOQD2h/z
EpDG2A5mVAWE4Cu8eMYo4kefrWLjlEFi/7fwUAbfsg6wgcbvcWIJwzA3u6o4EiYZJCOsxe6EVOrG
C+xpnUclABqCyVAmsZQzP7BGfDzMlJfSrVF3XtjX7r+x+ertKv5TsQPsOKMxG6jBpDTXKydCMbKs
m9pF69I67R2Algl7bHJBoDZjHvZVfs6TadMHWJd1+Wj4Tt1f2DNtdR/+H42lcWZnweab9erIfKr8
0GSsZD8KpQAxhTxd6fm3EijjNVXNSE7h9qD4+ZaMOK6CBAqkKHfpppg4IYBW0hijv1YBq+WzMP5S
ROH9e50sJN7HNuzq4UFY+mG1eRNWiCHSqDhnR7BGa9BZ3rxR+SgjH6pn5PnZt3YCynH7Yami7e0v
TaMXKKPefaWYEU5yIEiRVgqerCxNj58B+mXUh93+MaUqHfplzKMyTgAIc1ozjE0gl1ymjzP+mdCe
q8voOliIE1dHUCtXUHdVWapKYSp5YcZaVccZMnp0sH6VXyt6CB83qaw+xJ4x6cXMXtIrqKLrDfKa
P5iafNv+xQl0fdUs9iMksEgrEg2FvPrNilAZ439fi32t337om3/np5Z7ESeDKnhpOJtwzMVkcDoG
/COuPDd90yBTaQ3KcM4kJSIDem3dlT2Z3tG9J+1M2XBS9/6bRg7sMLdwqQ5oce01EYBd1CiOEBET
BT2MKRnKuheUhAy04hCh/xNzDSEmaKR5CgoJ4eUcOdvD6gabS/1xc+QBhY3ge/v+slhK1dntdCXO
zq3wfQ5GVwCSmWbL5d+nm3HG481J4nGD9zIHL1FCdGcLjNYe5VDeMuX74iVmlU1wWJ6n8HVwrxwg
e88XpK50J5ahO0KU7uH+ZxdIK+he8yK96dKzEzz/XmkEm/oFT4QeienrCVaVlGgTbRDglg/jF76G
8D1nrEXoCdteo7+2udpiPn/KJ2rnfdVKT0Vf4pe19qRhgeiCuFERB0pbm07OSzRL/8Akk/jq7g49
S1Lq8kBo2dTrLfLYnVFCNLmuwgOL563s+S4jXy7RWx9B7CvEv2VG5TmHYGIRzh4E0boy1XWr5kDo
o5Se9n9T8+aRpvISgG8T6SiHcB4bHTt+dlX4vAnT9rptDIXUryD2GMs1oOIweX6Ug7DJZ00qxiD4
QsvGWZgnnKT0Ok3/HJ99jr1iZREdgwuAi2h19fgWHQyu+l3Wm8prCih4wrE75TnhCjnKKTuMxa6N
CyYU0Cyi+QjFzZSLShy8sk3MPr9vZgjqzBsyetHD023zmYLNcw/MM/AxMloEp4g4PwAgLNhEGsrX
yB9sXkfCh71zCLZnL4Eb+zMLTJB4c9t7bwKDo1DTyb0x/qTRC+BDzqeBRcvlsD2damy/LAFWzg5N
rquTh8VqbX0WTeCluqtWhyW3G2nDJEBHhpCzmyFDEhZbQkoCk9fqyS6ZY/YdTuw7BqWPjipGoNFe
HT4Mbwy663vd+MI5I05dZxzNp2RplRkMgpi0biLEwyq3op2qzLwCmqzrjW413kuqEGbepUxNbHe9
bSmiGjVkTLSmnpRjtFQFCvZ+x7Gm/pyIeUr6ZLNSYorGnLq6MU9H6gBL6Jk6+ZViUP4zbjnEA5jG
+yzcTykeLfywW7ab2P0D1Ot4EXaw7K9eOLX/x+tCAmBa0G1rKkDhF9qgljA8ZGjNZS8yADgIye4m
PxLKPDQoJHjFewAIrSsY2RK+JHwZAHzFIBA0m+3ktSkw6eGhA6dHGu09AeSyCN6AHQNCZWpGGTTu
2IDxahp5sJEFY9X6aht8bRmnByHQxE+ZPD6nrCY7ImPtQ7RKFpTfB4Qdzqc1XMXkvTGytAvgDkQU
IV2Y+N7fANLMEeQnqoLP5mffzmpjmWWX3NJrFcuF5EVgV/GrgzqjzbTqVh3vaxc5fYLDsJ6tp23y
UNNV5bWpmhNWCIW/fVJ4uoWAiZVCKWu99aWfUclVcT51WmIIifw03KB4o62w9N74YdnAFyBjBrQ1
nXxENmPlqwhp3uatv+aSRKlu6fe/S0H6h4X6WTDxhjUTofqnhT5C/41CaCnkGV5IhyGN2EjsnA3C
8mK3ibSslOgjFofJAELJ+Adaw88l7arOr0kYghBvb9W59TwSWr81Dcf51fdJ5pHP0hjeDnVJcDmQ
p18kq854Mm/Ufjw88LzCdY3olOZiRGAaQyFuSELlta/YFvjDLlPZwhJuO7Zu74pJPuiVCHbg4rtG
QrO5CiAUZpxH6At76tO31GKdhgolir3cz4Vusa30OV0ip9f0v0atUQaqoAWllHsifz4WPH+Qdw1s
ysgab8loQtDcB9ZPmfQ2URkvRasEPBxx/sLnGUzrKLw5FJSsbG3HA8LgFJvyLBtcUN/EMtuHhhiY
gVEwdXqlPiwz8x1uzKDmoUqQdLV3uvDfKyt4KkhWNF1gIMUkZT2aptOcGzJ8Sjai9+evPj1OVJ0j
ALqT3aFJrVnMn06AU8DQGxascZfT2XJaiG+vr/i8q84SMKsR0EmXwHHH6s/FhmK1LfRUfUJl3pC9
GQgTpP/sA7ngZAQLUH3/wWR1GhP61XTAY6g/tRdmQ5IXGdRSycGw36lxN8lxwIvSNq86wFw6rIZE
SEZWSQKZGLwl8QsGwjgNNNc27rIa1FpUg5Y5WznZluagAKo6SPvKlV+pLe2WKAkV9iRMnPbnZYv/
aapzTidI3iMmy09/xCOyl6prbOiy3rVZnhL4VL/7S7/KkVkkyilTKfhTE1u/l7BRYeek64FwhUor
vKxc9XBIywXMqKTifYPJFgz/+CwCCbuZkV9ZBEytMv15uz2Vgl0zuN6s7f7zXkBMNx4GCcY/286e
MUnyyFE1hc3jCipkOR93PrPkX5iVO0IjGbBbvqKpRZd14npB52mc6028lwAam0dy6Gcepdto4Mwt
ZKntMBaPujvOf+MU4z+9/1Xyg/dY4ACGUA31hXogWmM5JY/dwFfMrTyGw4vXgsb286ejmG2iYK0j
APlaeQuu4pve8C5xso5T9j+pbJpZctghVShbg9LNwFKWUoQ+oM3XHY8dj5h662TCnRS7YnUJqpEF
3E8jTrezb0kSmQDrC8e6glUU3GEcZCKwmEu6/CiTBuuydHjQOE6is6TEkrDy/13ZCrBMLA/DF4UM
AjYxOPQRNBvoIBmwg4JVNpNr49tQMMzqBvzc3MgjlYwAoTPmy5vTkNYA66jiM95cr2k422Zh8EYd
5O91ha2tbxz0T7S8oCuSkdcBohT4ZFS0GU2W7zHc8cfshY6eSh2/1NJgIRBPIRiJvp1BkUZgw8DM
5XPXHGLKLFu0iMWTisEQ5xY3yLUICHkXfWiXVrr0VcZUM55LtsvXMRCoSZ+vRo/tkTIRur0QdjpX
X8QW4auj7VXGsIX8M+SmOkFDCAvArl2AqNzWvqh5ttcrfdxfPajWKYfzOroPp6ujpkXpb817G338
laJZh2EItAj3zGSkk3jcdpi4YRK1jdJzx49SRGkPOePPwRo79vq/Kd18RWidXmLOpksTQW/lpAfh
SQlY9f9LU56HVXqWiGx8jNxgFQp9fIloof5jA61xb7D6Cxuj7IDfhq+XJ0q0PcBQwuO1UFZ9AomR
I8pGejGB0fiyMFeX8BfPony2tmfc5H80uXn9aDserD21lUwGyIP0uPhwoBkiDKRPUq/7uqatIHzk
7szz7YvuMKDzJBgzbO7lyAiOCDmVFFONgJc4xutm4FwUCzaEy9XuSRoX+BAvQIkMXZ8YoaLcXD/s
SjwXAr3+PwJj7jxGx2jCF70X2fj8k8ucnWO+ukB8ukveBnzMwqBBa0imPNXmCcQIXT48Q+Iwpduv
nXrYrwV2P2dgQU/yW+eGDRTt4aJ2fhstoT4PtOsBST7trIMhE+ner/e6iZfP73PDKrGL+SFxE+S+
pHihPZAGJTZvfJEXhABdi1z6Udw5H7D4NzRQF1p6DR5QEQsvg4fqjQpjjaO4o/uuDoEIWxzUJtzu
pLALM4yqoR3M4kmHxQCaVbHuSyFZoXtdTD9nRSMiB/pNsGxZGH9ZKgaR4TZueMs4tSM/KAVRu3oX
1QbyO5OhUTz2z7Z5CEFLE+hzfSvSh8Kx/T2OBsV5GF4SUfuH2DT7baeZqAmT33pJzOjFEYz1EMoY
IDQIIh/r48y+Ae/LC75g4PTsgsoEhPyxHgKXGcZyiV7s2ovK087ksHeWts9gWgkzglYFcwZgUN1A
PD4BkPImtR7s/lCEuc+xQQbz6SBEiB6VfmpLzJj/WnROwbhH3MdaxFdKv8OuY+okIbna56oIdlLB
c53USQy+GjcRoHcS3uwD43v9L4FdVujL4If1RSJsvMDsQcaQNGbU0dYMnUCM8tuJU9rJTawNMxBw
XF+Fb91YIdKp1zmMcywDScn1Dl+vTnFKdVxz0sn68G2WohVe95jpFVkSSyya3gB3ncUrFNiRHPQU
f8NMenqP9ezi0hsFUDWwU+MGyCwgEHHtgCmRq8v3m/53Mu0juz/y/hzXjDit+yuntzNfPSAlJ6kr
tfj1LGv6gUgMABA0q1SQEIktlwDNWG5NmDgeeVjIZPQrLs+ZLpqbaytK6Xuh5SYtSAaFt+tdfYMW
VIcgpIlIMSONbQc1rAdrEtSteuJVLnn3yWz2damsMZuT1MBo778C8S3E/J6Vx51aeyyWkZyFIdwQ
hUTviIIX7jb/kZw3R1+YEqJ4SoP71jACzSL6e5yo5FYt47N0eXLWij2wYUz98jofz4FDOcrFBjSa
Gy51xLM67sTW/i2ybl1xkVKtO8CQF7Ra5Z6hOUniOKAnlzee9WgrDoBa640ZB8xNBX+KDgxsUdiv
5UnnqZq7ZTMMiRHLw/xq63wvnAyqjbNEj3jqZZblGHtziEposLruz7ATwjwwbNbEc/NIloBBdFh7
L+vMKJbkVKBOaIHNYwKWGtp1xmMYy/gTTD31pB1TsmA1ZKy+gd/1nObLodxKhcnmzt8Lhirp86uV
Rswrx4C96RjBz0kfs4rZn/UKqrnCvfsrUdvThUrv9/FTk2EfS321kjLyaIlfzNvyH5D8H/3R17lr
OJM3AwpP+n7udauKd6vdm0kpDecJBM1ijd2WAbsEW2bK7gSaqG5S3fVDlfATDfey5cO9Hq4HDKAb
eYvu9hqrDgomu6uVPWwq+eYbCJ21sj1g8veaur0lyalkZwkucDaLzZ1dYvu9kSg0zY8kjDaVVe9b
BQQIJr3SwvGLUvGeNsqRVMA1BA7YQ6RK47aOpnaZxdLpIjHoumzI5BwMA1UGvkAadvumwF1VOikK
V5o5AVjFhWVn0/9tH4cSVaOe0koCnEuBKw4o+R9jZ27QfEsNWbIDXJF1guW8SbmdTfKol5ZJxSP6
KcwtQqaBvBXy2FG2l6c0Xnav4yR/DDGra66kI6geu4dnWJPEXbVrpxTl+PgOc/P5CjKSt/CSR/Oa
IoDoWgHwj8lj3h2tNk2lFoTcWqI0sy2r7JE3ybZXwhARYalzRMzexCS1oagfeibj2TWiunduW74g
WMQruLCfgkFNFFGOlTVyU/Y5ed0uBMkbbK8Du4nwWcfFQGnKz8IsBrMJMV/91tdj3pUVcqO7bVwy
DOs5RPIOQvT5BsnZ5/W4n5BQKh1fpnqzgimoRhcXd5rxw2oqbO+lBK0SuCoa58h84yfZzWcof0sY
rcQRR4rjZFzt61z6L7HEMngK1pjjbnC9pqXKup9bg5ONL5gsos1+cgNhowToqfe48B2RpO5uoT/F
8W6FDM4LBC/ix5cvAen/PnCpmXGFAQaBeNv0iRrugmT024URBtg3U90OtEtv9rqSSz4+MWwi7VUz
Mawh0MbS/pVW7xODQdh2zmzKjHwwEQhuVzuyRPM6XeaywdS/nvgWwNuorZFWrR31JY1pDlaBv3TI
lrx22/Xed+oQ/SDjEr0mOwjCSR/JWF+sxYrptWvedjWuSGxPpoq7laufbvSy6o0HxVBOAqfvfozc
Rdb8rTWNGkVMLH7Pw6e4tQxXM03GuN+6RtnPY3Epp/T17B0QDMXCdeJ2nAXZkB74VkO/WVnjHtFD
xRufL0t6TXNWZiAgi+OH7kqGjZqcFze1DHafX5vTps1I1cfrww14hNKL8Kzi5KCn+ICdHr4QyaQo
x0JD/5fAKP1fQT2tsoCUPMb+ruRLkda2sV5d77o4d5zEx5SKKpuCnEe5qLL+Kte5OCE+VtA4k3OH
reqGpD8XT1ydDOGvXmIjU4N4jk+sReiDl69ydNvJBzKbf77WZDn1MJU49aJrGunWZanZkAxiNZhF
A2gHzU5JfrJ8xGW3t2WxUUwiQPo/UoltJv4ERjPdXnKWimWshSUbNOM4BEzDHsJYt+zV4IaTffeq
NciTEjXP/7kvsUeyLRnu7P9gvyQILgJUslgPezbEkNUMQzTTgF8eqmfz+jvNQHPuhIc1J28ixAHb
/8ip4CP7Ym6zUlpWGhfy2O7R1w1xraSr8+dIMhWPY6NdZxdjgSxg8hV1v7+UHiXmvAcfUTZCMs0v
Xhl8L1SJNwN0o1xdwsCokMC+8KLLuxyULIlFy4pGhai6Foylc+SGLen/NsNOJHAkAI17/RQHFiJY
7Zq2C/JORWKvK+jkuqwYFWqe3RRkQ3XsEQGgi6LsMAH5dedqGlM9yUTdasauez5bfhPIR4WLXQIH
KuCHaijBNBRFEtntXCgv7AlXNglr5dmN2dCzgewpNjDBP+gb8DmLAZ4xUoQbkwhPnG/Cyy17GStn
QwnUyF8zr2BG5b3GJdQnwwvi+DB7vnKvCemC33sa97Vn0sJ/vtNquT0/pLAeYMLS+XL9W8Lvlmx7
1wZ9V3ScJdmR9E/RtzHSTahyOxaODnVRp99soU41VvT64Y7YuHm/iO2kft1xEyVtLULMVKqCORdX
31eWN4jyMfZlDjBLNAsdcB845jMbty2hDlG2O7aokmmBr8hfEwxRhrKQ3qrXz0hL687p0fhuz6B4
PCCvXOgA3oN5qiR3zyRTOsUO3TgwtcmTgomw/Ho0CEp73cQOL+LRkznMTKGTllvxAw9AYz5qf32k
pSlUjb6fgXpFaoimTh6EOdGsxi3r+foOoynR8SYfupQ34iwEDywgutxvNoqDWxhP5ZptkIBBAiRP
RAJinROnJBbkaStSocKVWq2toN19XHOhfrzQUckLd4b3vEycWzDWsevmTkn8kZz4YhXXv4aw/82L
78YOePUC5yut8Cuz9nBo77DX+CW5ksfDLlfriiSSb+LfkimIJj8HYah+GBALqmsu5Qk488noKkSr
uu+BWuknI1iSNslndsS4hyBgt5k3xz/lM74oPrpSsqgF2H7estuL2oipHJd8zF0f+u3wwFK4WC3m
R8HlF6IwGAZmkv3OVlND5eLEIABbDqp72Eo9ntdrh2V27GJFnNy3OoHSfXfjojDrm3waVD0ar0QN
49wOEg9yOhobd4123W4sBztPr1YRGBkrKstX/5cHm60qbtfsDMuEWgkieIKBKxgK58pfY3tHpI8A
PUn5tUgZq8XPkIJ8a2krXofmnGpgrmHk/yNmsfECt3Q92mAm6gHrr09l+dC5UQAQoGlmboc242Ke
wOb1Jn42HKVZB+5HG03ErxlPkG9Wrkde3fj3aIpiH5znX6IX9Yh06IGf2XGlZ8fHt8rk1J67UvjA
VOb6wtyRyiQibyzaMfY7eNngy6lPTYarx7eSkZqdMZAnw6dlypS/Dp0yYlXlQA7MFKKxieTDiuHh
vGpOinQjBBHd54A6agHakT4aliPfG4wOQevlcAR32IE21vcXn8xAzfJgvMBzRmMvQHtrY8s5csOR
UlwTmoZgbYTODRumnxsVbGyvwcb2XDT1BHN6OoBjPFj9XmaC/6zR9CVAwjg4sTxN8gS2HLoOYP5g
ruADWkWMgBHs7XBwzKMk9nZz+1S6R9HEAk4Z1YdDySRAPCBG8DWcb6v5aPHEl6+Z4fA24h46VcHR
1nnFcxCHqNdrGo1iKGqxPO3tCj5qlmmm5EPB67JNIj8AtViD2uOpNLYqkW5+gRJhjYv8eruIokFt
3iR0Upe5lTVjvwvAKcWCe3mTw+38mtKeKr89w92YR9EsfS2zq3ofLDG/d4DvbR1oSDwG+QCoQZbM
oaGcJD1MmxaFOeV2a4A2rQ9P7jIz6/Qaq3KHX2RDssgV4iJ6DnlH5QYqV8HGM8kmEHOO01ldyTOR
Ywfd9iZZAxrj8YFF3qzP9GaUwgOn/llxX+T3zXoCIp8OUwh5FNUdi2nxONQNvpRTI6GVkiulCCVM
01+QAzEN7JDn1qQt+WQGBEncoIc2xqnCjHT3yvuu/lzhyDScMzDi0axV0iGAkvl5tzDB7g8R7i+9
t8NufSD13q18x5K/HGqtiiMXx53SJr7/B9M4rqwkFu+Y5jYecHbknS2x8hF3JtRoc3lu6FSzf0Bw
7bLl76bX1R3Xi7IyKnKEKtgIZWVIUK/okhcHS5PLGlVyjxU56lCRnHZghBKm0i0AhRiS1f63KT+D
G+LYJQCko14HzcIoByXeXlVkbJ7bPZHpazAy68ekxsCMjPEys/VkuE1zqi6Z11qFVqTenAqE0oR6
jSdRQmFkxzMsmQGN8vbUhFdBoicOMT7HtCkLf40porWWvYMa3JG1ZMgNnzmYeG0CB/OtYF1ax3vT
YOu0AJQPMc4CucZk1lltwMg6x8IdrE9cs9qiVg1eG/HvWDK9cSoQceEWQrr4Qr2iCaRIQWpekFM7
Dq0dY78vy6tLdakaQAdXGjUiQN1DLNG0c4xWBSOtgL/qz1T14n58NnBWIuVAq3jWeOFuHo7jY/Jt
WI8dfDtkzj8CLPGwaZdSXGjZ08uZgdNtXZNgvKCU8yIiACq+6Gj3VtTiOhQH5Nkb+7LAl6mHUtBF
Adqwu2sBCKhWFnPtH4KdQEFqfMzjs/P2j22RdmF1E79q/2llt0FF7p5VQHn3QWQS795TVdMmiKkc
jwxTLKD4PKSbROe8leklQYXQgMvp1OUKNmwnsRC7PYRNmqQw0l8kz1gpfMhb03m00Q+6CKK91ktY
zlHdTG+DkwRibI0JL3mOW8G/fmXjn4a/+9c8ACsSuMgvxW8wc+TMQOzdb1lcnW5lNlQgPO1Dtjpq
HcV1BhCUxujocEZuAo6FOJ4yplRX11XsXVbvv2lGhjL97mFI+PedYU50KIHdtsWUB3ULHZXpvLHf
iYHFblfpNvrw292QTC2NxO+8D5c20jBGopMXZArLJJaN+RnLQ04o50HoXFJqnfN7taOLXiQ9UHcP
I7ioUnDBwllXfxf0ZPMf5dwl6O3Mk44JNUnZsLj0/1CBo2vmp4SawMGJhRXJzFxt5mJqP6ieqvhB
DPE1OkNspPkTUrIMp6kAJr+aWdLds/afsEJcUjPtJiy47qf7EQMSzURdVf2ERDKBp+7cofo5LUKF
5WyyWAg7EuXoq+E5zd1Bnj4df3VdGDVPpFthIVfVWDhK9cMmf2Rhx+eY2BXz9+1TlYHbQUsNTQxV
b/9cwMATVIBh0en4T0oZb3aqRlNxsXlvNMojYE91O9gqv60DbnUkbmEkfoI4H1Bbmi2SlySjjeJK
kN9P9ZHpjNM3+xE9Al0916nYbEKEuwYXWOfn9IsK5Ji9Y4SDLx9HEFV3JgGbbBmQ+lwax0b5VhE5
zOzfujl/P1QpCPoq1Bju8IGhCYglJZkPSSs4tKVtBtaY5wKulUsnzKTr7yR9MDwVg3PfwIaUJ6NS
RbzuU7BaRf4mP/Fp+5vXnNiEEdzT9rf6VPfkJrLEjAAsUukaIAUZXwWlXAkdoWf5iIhfzXZvfldv
8YCOG7beFJ4H5eFOf/z2xckRr4EgHtC9kA7m7nOfL9Z3r46/BKeWEl5Q0l4Uc9Tf13hILbUlpowm
JsSoHoQpvWBBKQdOXN+J4JokTHjURG9WbafnY+DQS91Rx2IMgvVXQULVdCqTnXCZpkMuDU0vmNO0
e8gkkHQys4pml4RnNsHWj28xKn6Q600bwgN1/WapZGqunTKSXFuz71/ULOW310hhSl5uEaW8v0Dt
1CYYQVuKFLlfwypJkNM8ead+78yz84TadtqIsFUXoOywqVOSiI89eYztsL9g5O5Mi1oHTlLEzQBk
QgzsTSNIbNp5LrcTP5zaTnbAOEqW0eK5eZtzv6h8GqxrA2hyw1YbOldJT4Gr0VOfdesRm0JfGq9q
lnedUi9LOQ5W6VBLYOqWybfR0Xcq7djoLTSRGV+tAGv1KDp1VVppf6ebetzDwtNKHLSOk8Cy1wlT
hKM/6VeM2Z00lJsyU/NpZvxm0Os2mcIoiUH2ssO2LF4OG1c/m5wZ9shm4ZUxOrcUVWbu12uIlYDS
cWGdGzN1chD+5velXHIg+ONydhBNq4eu33BXtB+J4f/MHAIVXng4FD+I5Av9U21OB8OeBWEokSxX
VWlZq11V3hcvoF3mblfbSzr7/cpNbkNSCEwNqvCihynA2LvgVwaC5Viol62wBl6gQ7UkjOLoAdUk
uE5bMz8yxnZeEFL8kTQ/OWESsQIjqvdJEUzSQNkDZaQ2QvSiLwrKSiNdsPhYYRD/5LyDvSAHRkBy
/1N8+Pb5hissZeWngLElsUr8yE92WAW6WhUbgQBSfxD4lWA6iSqkEnxw22LAzCShf75wmf4NQfyB
V4409ySjJS65oIvnt832DCs+SYamASASO4ZOjzPinPa+Yy8iigjaLA7QXoXJoYCzJLNBBSIlULBO
6m8oUmzuXyZXRmhZjYqRquG4r6/jR6W8CY/D5M4zZ76KU4fD9GnZwrHtlV3V8r/20ObEYQDqGoLS
dnkHb7lkk4PJUgGX34VY/EK1eW+u1R+0YFywjxD99a1LEYRA/FrLAdJ4Sj1JsrONavJU0qoU0ofe
2yaav30QY90xfEn0RYn7NNTNCLALRcY3/iYqpgHeI65wdI5fG0Dtj2RhvLgegV7+H0XipxsujRPU
dnT4WH1RE/0UdQXvPu8PHUDHUYPjxFyF2z0VlYjo52Zcg3wXrucmEl674mjCHjZohhKYWps1gXSq
LQfFympqlLwOeWitzIMFqPz4+NbmbYR/G7iwtDq7vyETe9N+t9Fk0bqk19km2B3RHMNOJsbv0Hca
JuysgNXee/Zbehv312DojzF/igaeHILUWDp3ymDfTZXHvguKsAC1oLA18cPjVTqTNirxb/cMVv/S
2CWbZkxhGLmbKMAcb/pEf/jlr+snqN2pIbPAqdEdiM8GtdU60wg3ax3YqvM0mzG5TA/eXw/pNVS0
gMd30bDlgY0mTBwwE2emRTcFozlQ4U0Jhesobj4fqRh19Tg/A5uElgnPpvKUP1Z0gJEcFyorUyz2
o2k+H9XLUohI9TxK7cHKPo1Ag88uPJQDz4r1xduOE5QscdOJOVY0duceKpc29Wp1QWf/qn88ZYXX
QKv2GNvouoxIZSA77GDA+DC1orsBdWs+MUzt5XQkLi5GHAd4LQ5sz8kVuepqJUS0tIPzUHFxeNso
wNs4NDN5SCwBkhULxVpP4H5O7Y3ZyB13VoivFhEBD99dJpjQw867KijbE7Yp8uw7rwor6UFkljjo
ZVIi3c6nUWpLaN51G1CMyzPQKFH+MHLAMQikfmvWDQbWW9IqVTYNts9fuHJ5zpYCFgevRu4jXP0Z
47vyMtAqIIXVdgRRYqDz1EihpWB/w1rwB9cTo383+qPF4C4fxl2n6rW0gg+ScR5Y2oF30bnT1gZ8
vEwBOm3P1XknmoBLtfm4OVytlCOK3at11nWgJGGU+PzGEFBWwrf+v0KjCzpr6EmLL3fNTtgi+vYD
fKdXR3U6dLLxJMuWc/DODv9JuPkwi4/+oXYUndT6ZYjX34K5sZjHEIpfapuMjuZgicHwv04tAQAY
xSN9+DhzXR/IO//sEn2Trrhm9AaL0sd1bduEaOLe99S/rtjmkPfbVjpAhhacrlFVYXbcDDxPjFNq
c2wkgbUmc2/qksNifvJq7dEGgtVViU2k1C2X8NA0r3Ohsh5iOVIhKH/ckofEzO/IcbX0Du5IlR7A
zh5k9QaYgH8qQ6sqLi12oyF3tfftFFx8HeiRFRfHGvadsqbxJShz0iyvlPmAAFhc/A+PuK0YsMOz
wukDCkTEXD3zVZWTW++6mH1ATHGkbRNtSZ2367Q+oNjh1GLK3lAuZ16LQSl+DXjce8ihW1STindt
Q9+DoL5fEAxy4nvU/S4YCzW3nmmJl1Tj43RUr+jqM6oOiHZwLCgyTV7rTKHu1Qy2gdn0kkMg/Ic9
mqxpvYnTu0EEE06SqpQFcbIPk2uhUk4vl+WnMN9XScMu/19ToWPPoVXHfTiowhWRwkQvx0gGCy2j
QQ234UZvxGLuBUbr0+KkMZHQsjRjlJb0kWrkJV4oOQR1zUHDJnC8dLcSA7dY+ARpGS2tjxgdf/JR
sQCMJiUlFrcwsgMg5DJgXR3apfX6gT7DBezMFXWnxHr1gnFb1I+VwZ2W/PI+hxsvVKwUST9vvJXb
G4bnVBJVK9hwHFAJsHR/e7E0kfBQZpphThmLSJf4mHGY5A1b9CYAJCnTGZRDxqnNkCMKQ2QHnpUW
BVGZ9BNrlVUgTFaFmUh5jDEg2b5PrHltJaBEjC2fTuHC9gcsXqQYg2ev5I+SJS5ZCr4XLs0jScEx
eIpjH/vGOo6IqDPfrh2GAUB1fJ9f+DM0fUHd8s3njPM5P57kQ7CIbZO1or5kdTKA9ueD1/dFpIR/
zV1mJsvTINkPk2dm7SGWEyq6RgZ87b/sgjzo9ztJP85zyONXUBuK5VB7LHOSfsc2doxmPOORoNjs
t0S+RD70RATpKLD9TfoGwJWNSChmJL96iYRnP9c+/fL+3ChOxjkoocWCkeGS3N0dI/bcMMTkhFFx
Ne29KUghWsYj4jOE9nXTYax0Q7K25/lw7/N3P+1QrmRImcxcuFsw8Iv6C5xmx49/yJSgQbLd2/dM
6p9Ykw+gj5ItmYiQ8pIP0frbkErSzynGc+MKUdZJUh3tZnExU0I4hiF0S+vtXzdIhTiqQOkSbGh+
mvjSgsTYYSkjtRFiAFjOZeNcTJNQqQ+OSIaQvnpCPXUaHoG+VKmKEkr1R94U5KjcoPTF0GQ/Io+6
y7DNdm3VIS08AVX6Cof6hozU6A3g2pYOjdD6PZpqRsBv9osa2bLaPZyU5UZ9e6mstmeloX9EqfkJ
GzKu4YVtJVWv6gOhtG5V/7k3cgiuHA1CSjp6zyKl/wX/tFyVd/x/pMPkbKeLtJlvJPL9V1hsQqLj
G6zmD29DXrSwBqj5tYoqwB4F0Zr5yPBVhM3y6UYQuhAk+uD/41YZUI7MrbmqevKmY/Ur34uimZQ1
MbeEOKjsRAltC9PQKO76LbmDbYxbqZaUTyS1RK4LDIfevAyT/n4ixkUBigSJcwXrRjlaqfBFcZcG
UmrtkpoZiQ4JfsigOgemWrYdFxHG7Mdns0C4LXfGa1KWjmvvhWFeusINgtAyczzjZtDKlbt90QHQ
ZNr4qrrrVVEb5v61xyjqj3/b1cAr9fezneKLItPOVm9JIEH6DsRK+diTY1MyKfqiLdYVanXRwFzZ
V0Xi8FQ957y6ENLav8UV4K0WaUvRWsKul88Ocq7mJDexpyY/+6pjCq1YOmjj9dJN2JmLvKJOPriP
r87eSRGpgCIQjZ9tJo89056TpuminJAC2VOwA92cg/NXoLtZteZ/ThRQ6plKPKg35KVL0UruNKIv
zxPFchZm6dUdknP/6Cvcn4/mWbZ4OQKyIoJR1apn7/FxN9+01XOIuuvla7RODbEMryQ+CWkqoYs5
7RdJZ0x626GbgFP7FFXQBu8nFFTepQJSf9PK09ThZv0WQwRllJivGu4MPqRzE4t8deHmNGWit+sn
jUH62Vr/Rvylf1s5TbrCHHzIz/KOQvkexZiUBdT9aaFubKReUiHRAB3ARFkYtz0jWUKV2coP8Afm
dhCq+Lc29CY4HxfVG3ffeEPKFImmU/HBt3KInqRdCcvC0FjhKCSZc88CSGNRRiWNYnFyM7XJdyU/
7G4XeQuN+KhQb/dv2EMMucGidL+3vTDgRP55qpS3s2bgMK1uyu9/4Ro0NpMZjxYlD9pttERFv+/7
UpYSfzn2UK9XRGWP+1RhAGMrX0yqyZYGA7Vb09+Rm4y+9l+x9lAggclc1FJLEN8EpiR14tnqtMoC
WzNyxp3bqQMszt73PzYtBuMhg9LtUmA4k7AWuGL8o0EE+7acLgeztAFcov8PNZqpAEgFwMvPBQY/
PZMUYPYaQ+DigMhtgtG7hcaef/PJ7uZfwx638mrSq9c6KncHp5eXWYA7p8IhtuewP2gbanRDdwEm
XamLV+M6m0BWOJpZLp9Tzp/DbBF9P+qJcRxlgsf+sJt3aF8PHH0vgpXWeLg6TrKULMR5p//iFXuI
WDskedziJi51G/SJwVZFJxY/QxjJqXiQ96XxSUA4vSWw73G8438FK1L8HixHWajGRL0FyiEFAq6k
A7fhD2dFf7sCFRLsMO3SvwFtEhtdoo14NmnXWeCGHVzYddzfSIt2KlAimYwiQo8dI/f/rjaduyPE
Nf6LP+7fh7oOkbMw2gZFhqn2DMnD+UDtWRNDAKVpEStPUN/A+BWWD9N93mvl4gmGgxyBXpQlt7QX
A/5gXLymP1KVzQ8zr2yMr9PjR72WcWnpQJOOwvv+uaj8jgizn0+7TGWfbJIz3zWWHyK/NCu2hVyU
BNea4FnqbrMhEYhMTItVXUxy+W8PBerJttQsjpgoh5A5ESonSdB9nM8OZC2HPkSYr23dTWbAQLg5
5sMc2mHJNziEv3M/C770nxExDbPocg+IXxhC2D9XqY4KhVrGO2cMcxKMKk59L45ZAfxbW8dz7zOS
OePgdowCinPcLMawgytTi6TrpXVjMlb0euFGJFGgdAvOJ6q1bDJJZ8oGfyv2CQFk5fHdYkIWKqp7
QMFYa2dZUHao170vpXtu3ShSRBRiYJ0E9fgTaY2tRHf3Gt5GkfBq6NPqAbbNCPiBeHJEgmR4D1Ol
//qb8O0O5Q4ASu8vOFz4tWBOy3G/mp0oinwbQ3PxWhPpLMCx0/R7yUEFT94VeIYpA79048OJwASH
49VapLqGZPhPMB4270RHGTITPvuoMt/xu6axK109vtPFPtBXhnGnqLo6g6LE0kHJIgtks31Xsmvb
P9UdHYrE0aT+64gQffMowfiGYkSZxOaa31mxrR/kamUzmBdVf4DtVvnZYof+eyffsAlVadpO/ZAd
MBTCrUKGvnkjrSNFkqKsBixodGkkSQqbloTTWtinwcabEsmVeDZutuOPxiO3zM+++2ndwD8LA9J6
LuENRoixy9KdJA3xJH/ziIm+VYJlGsTF0gFAvFeYz3x4GOf9oxNx7c10sENpc1xfVm5jzVA9i4NX
b2yaAq//Ct7l8G5Z2QPNYZ1KShcZdJOij3l4z6AObzPAnRx9V9HBgyJKiw5a/49sc3CPFgfLS/JT
YHSiovsyK3hzWhHmrHU79xQ6VMqCaYXNe/fcsOAGmK56Q/R9AY9pELu1MJIe4IOpZCmCwOPxGx1j
RtUawU5rjQ8bO10xfEuR10t2iONIRwvx9yXcUHcqztb8EXwXoqjqbNQEtQ5GhmSubamXuIaLJGsC
9u+pg1+eyQDxooAsCptwguNV3eXLlZu/QRg8qYh8rXdb8dvs6hm5Juz9GyljnmpDwyhdEZLuFXql
wFWouBMUREmplsCGtqWfEUa9NsSNoWFxuM2HohNXMiQdD1n8AtJqBzz7ConwVSJx4FWSB/jBg8X1
aJWaeOfl+88p3Q8TOXPG3JRfum7GgbVS3p5BpwQizTDOJJaGYx/X6jQgKebCc7ika1kVL+gmg+cz
iShUix1Ipsr7iPaoA5p+YSDBIZSZjgvW8Sm3O/3wp6wdLDmhrUtCM1bE900SPQNxWIE2GKLyofyH
QiVcNRV+PSAZD4oQ3YTuNFDVzUqORBvthBrI1n4vmsrLrZavVHIfQVq7fgjUtN+d5szUxSxioflf
28FjiV1ETt55nkXvcsjUsAQ7Ih4z/msSYV7672qrdjJff7DoeNHLzDSNWzPsbAlshn7FFirtSIjK
z4iF2KAZGV2BOJBvKDFypA8Ye4gEB3W9L6FuzxDDPvYZXpi21ptVZVUCLCNt/jCVs/wgJjUOSEUD
+erQ78zjDW4L5fdJpvd3YSVq7Kub+Ai0t0BBLIwEHeFoCAS3E47K2dicoYyltQzFv6kAYE/Weoow
SPwkOlX/WP5xlI0f27S1cVlIS2AlqmSQkyHnHnQ/M6INNu0UPkz5baeZFkmz4DcvecvEK37umElp
867MnuqicqHNoDWlb5TFbVS3jrLvgEADO/j9NQDo1cslQ1uPgzAro/NyJ9CXnze9QtkcsHbYPIU+
AXOYDT3wwA2Xfc6F1XKgYWDCFNboxDmE5pagEdLX4AoYeGmg9qqj/QFTkhqv0RZKI8lEx71jBha5
xxJ9wO3ms6mOn13Qmj7kiWE/kna+lhv+lQZkAsbJjmx3YVsNT5JIKC9I0J8UcYiUbk4BZ9dC4iZg
jEauzKeLMTqjfol6rB49jFPATt4PQIKAuNXBEAhO+qz+L/dfZVpdbrffMookkxUmhHaxejBGq4l8
pCqeJsqXfyOHoTi8pTBJEHkHOzMB3dRYVLN5LAV9w28W59ZLb+VzQrNk6+THOKjwwty5CGXTh/V6
296KHqXT7QRogDlBPq5SFAwpX5gEiCgkUFvdl7fKEn/+ic6s59fwXzsvLRljx21DLNymbSiCWT3Q
jx7JBMikwfRMWcthsaFFfpmtXJ1fgewOqwbEnx7+gdHJrrtZ7Z8CMLtT0oWLX5q0s5wP8ycW1KCL
A0LoIzZkJ4GORRLh090RMFFWEyMT8G0Z52b92kaCZwpBKHU/Itcdofbq1dUs0/TvNu/+/JMfyqzi
pHUBI/ocnCLUClXCN8PRIMFHadgQcSoDfttHva45DAU1FY5vvgbrlPgEIkju20Oq2yjeO/irGIve
R6Bs7qvNHWqgR8RXUbYe+Gnw9HaSEZhcHKdgzzVSWPsZNSI18gwOALJHg7Al2KXuAyeJQmRfnu5N
oEg8s/Zd/8xL9c/cepuSVwQ8SF7Ws2OFARSB4GwUAqJGBs2GuTlS5vylpytmWvDasxJ1Tjl6gVo/
3faL9JZ/HWQOXT8GJz4FjMRR+G89FuJC3O6TLhxm5oEn6KefsYnNgCbAtl4vZm4q3SqyKzTfDXXL
X6vx5c8wtE20Db8cuB1cuj1eTPwYAvvv17uwNHsoDdPNSDFSSlxB+IuaROO1LGdQgHRsESqMnJLB
U8WmUzt4b4/zQwhUPMyWaqBHgCXzpdQYFii6AXZQsw3zD1sD8jEeViyqOwbOwV5u1pqO9MW+4hat
xPiejArRD0qYvFyndTud/umPGHQslaB4GkY9HFgQQSMc5uWqZqfjt37cbJ600tEjWXytcHKTIYQX
Km5ExEXrR6bO7yvTsltXoSZOQvNgwjWdq2syfgooIFdEIh/tBnCvlJ1sbhzE++Lgc+8sqGekDwtl
2qd25utjD9oCqegdeg8GluNHId3r4blfOfbgycHSU7OCXNvRHsIt0iNE5rNW8v/AP4eqfYSZuaaH
srxlZVSagsh/YweUxvKtEREFAvNUSwK/T5aqBNYToUbeDPEy52Rcc5vfkpKvuszPH74kUrolLTm8
CB5KaipngfDnfB/32dE3xCumenvtykdYfx4+ZrWcUQM6sHujk2ePZhjGD982Pr4gDATtu8cjqIvP
ephq1vLgq/AtpQQQKKzDwjdvQCuwt65H9LwgJx64m5aZcfrVkpDKqnwibwXs5/rDz7bmpOMK/tzZ
mvRebR3oNZiElwIg9T+OzkPmg+2/0GA13eMpwrwavRa44JhnWZIxhl9Vb8NFi0JyQtwYTRGxRPBU
BIgmrEURn6VHCGdqBgu2+wDpy6NZMAA5uVNJlnVeys+F8G9u2cz0jwnV6Gi3KZkAn/cfIBRKngSf
p8X0prfyG/7yXcie1KkkIn8Zy2YBaruTRuVshXNQjDkISZmMN06NwdzGM9yeRDlkaEnKQbEz9pDw
ISbFr1iZRidLOUQHmBW5HafcNZmg4cOCjBWFVB1St3wKaAWBnY5IFuLdmS0DgnbAMW0o3e8GJabU
6kn5tGbVizktnkQkawfsWtcM/BMtifMWskAcC+VTTG70+H0F1OQtuoyPAwI1DPVOmcRiI553Mev0
lBRfXG6wdZdhhhENf25zjQS/iABgc0GD+1ZKbxrJLkSrtdyOn6x+vqbav/Sye3TJWj2YxNfyTk/Q
3mVXskiP4iQnZzbEHLzxuNFwFeyou+nNcQ+fNSDIexiC87On3v8mOvGYALwbMZKS8WkMJ0z7GLxc
S9MD/Qnf9W45wbobILvnx5YEl/H9tEZeQdaxv4p0/wrICnHMB4+/4Tt2QUF58cAbbLubqp3bAYW2
VUjd34A9nX9nFEDtaMPQBmVMLllLy1+dP9kLGPQrmS3f5mWNWBsaPrMAMmmv5nQY/GB7UFgkvz8c
qm1pNMtBu7JmZKCkf+AyjkeHpcpeR9HP0TyJIQr5WsdJJihnTW7UwDAC4CpT0SJ79kMR0+mTSO4G
IUXpYcrA3lizi+wXpcUcmqLgVsGaZKfsanwxIgRcM4afviEORirYU38emHG3A3NaQMDBkTbjEoTg
Xh+3bNhvD/g2qHpqNdKC0igQnPRvCJWI+ZGQK7BLvLofwAQ8z3p5Tbo81570WRzhC47jReVsssHg
l7Erg96NcVrtcuxnSf8lJhen6zE0kQLF2UFLoTjhUsIAYrmQ4PM4NjZz2kpedLOxgyhfl/m/v18w
klrCE2201d5rSxTz7/kIpCVHxdE3CptwFfDJIgKR2pHRrI2a3T3qs/3vXCGWA8iEiJ6AIvMlVeli
jMtkzQdMQlopnjlm7VowDsi0ZO+b8vaRfpc0NSz2p9UzvDAIBAN8bwmzkQW/Slymndxc9ua35nQP
liJLExt/1vmZ15+o9ZCAjBZl5t4G5EOeEROhiMhaqwMd+FJ0ziXnDE3Q2ia22DyoyttTTyj/iyb9
NedjsXahd7UMOezfVjZkPp+Xt0rR6/5bEWMZtBX7e29mNyaxeriLsjAQUNFP+FhxPWx1o5RuyPNz
VRs7BTh/2Iw+vUrDE8YRWoZy38eA8vkKWA+Z1vKbrW7V+4Vaj7lZGxBs+mTXvqS0RnYFvvoZ6qVl
E8MKxJHwbH3bZ9luSmBxBu/dbI84b1xgWEQLy+ex+u8W+vOKPxxz45Lw7biPGNbYct2SlDXuQoV9
RuR5DaRI69NyH9H3Q0Tjo0NTZqoRBnA9aSS8uheKWvb+dTOIXB9HHg7DGEltPStC2DLcYBWsWipH
x5xk5XunhCAroCmZdjjjD7Np0BZYCTRSsmp/dt1VOPX26PPAtEggGQaIgQ7M+thF5R/bLMEVNpoK
4KEQTxP4/PZauoQmTrrNNQtiF6Jx9N46FjuDzECSNzCQLRhtYWxA6a7yvOerKIaFRZFbt0kR6MHP
g4kdEomdl/vufu2ZcDiobXo2hoJwHes8yN9pww85DFe1Jv36n9ykQfhDK96AhMskaoFv4HK+0lJc
ItBfoGsnJA4yxnIQKQ5V1pqvd+joxCZtj1kx78hbX1AEicOEZimVq9gXwpusVb1oQOGtBO4zt4yP
fD81CoUe7jmfHmegKDBhzM3TQcf44yc1eCWbb3NIbAzq8nNjPKSZ8xoRW6x+3BUPqHUBguYCMbKG
AaCApWPYRf+XTRgO40UoqcjrEEJmoQhZotNdTHT7kschI67NWwUaF3HCG1AEH3s1nxTHAaRfKCVt
ZHBeW0wUxKhpis5veHiPU04aKfeQhBwH1mM46TDal0qbiaKb1/2KMjX+Afqeh2nzSzgWRds0LDz7
4rHFf0h6S8MBcawwm6pq0d1TZSWElYEvHQ8nswrX9P1tkG/8fuJcJzbwBFxzGzSFaSAP5jPPXhIE
qc8hoRqB8hi486BCkz7WQnYhLa9cXCG5NmL2++h2xhDqSpC+NnUfWM544EpiNHwF47MYurLWRdey
3immRmMOWe489pUaIWbTa/w9m4RmTIfa+VIQWd2FLd7dqTsITqNaYS2zHekMnNHxVto7t3S+bGKf
iXorCgY0NYJGgktmuakyMMKqio8kBCgAWySjtnqv2illNYTkmEaQvLKXY7v2ge0xj1sZMW9B9aQp
lIino0tU3QybOF/FVuNwg0oshxNi2ye6fvvJxLxXSEKfEwqHc7Wul9ghFUKv3lDJu35vobpTzcO3
sxVrVqD/UvQUhtgkaCDiDAw+g96AVxwlND7ib0KDAdYJNJ3EL1dBfAN/BLAPu+CJCavOQvew8BpZ
JJmxwEXEgsVqp/weKFzMWiBgdDF/exN9Ktu/EjGTZBJCXpGYhqaZCux/OXqx1ORf5rKwVcDquojX
ZQjQ871sucvZjiNvH5eONq7O3flw81deQJ60eO6qCI0agjJfUWB+GU4527NdGHoWcBrVhGSyF5GX
GeSblhEhVPKjWSFru+s0tIk+cZYqrgpVoshHCEJ0xNfFDQQRDCMKhQLeskfJ13cK8rEclyQOPsx8
Xsmmy4LnVTDj+dgJGdTCWy0vNH+Lnf5PZboPpAwr6mye0rT0XcwgaXFNkbDZoZ9AUnU4GcILZyN3
gHvBeY0UCnGGNKrbZVGF/EoF8Twf6QDIcauydtDAWvmVHEFJlAc7zRcQLCQuSYwGEJ/E6hza61MK
iEyiGLl/prgLNtMVlta+CyY7hoUQJ1gq/OARnKAOxyLpuB+JT7KG0Y1Jx9OvqqyP2gX2uILs6en4
6uS+n5JcbpJkW4u5WAb9VmBeShXIAGAwI5gtqlrmBp5dR/BvDNc6H5rF11izG3OvY3kAsX/pLQzh
3mnzynsKaxySj09FmNUf5luIXbP7kioDPUOoadc61HTqPCIbukNxjMzvZOCv8Lq8JOkB+luXt3KU
JKBRC4EvZXBLQUHIKa5DYH86sH9olpPNTyuvZycQPW5vg6LNMFFvwZTGQLGlBXGpqc5L9Rr8NDF6
aQ9vgjFq3ROV06aYj63Ld5IqPnH9hsZmO7A2GqDjBaFctLkG2J5scEL4OJtf2LGXauNclq2zZ9ax
lM75mLdatcNuoOLUKDvXUYB6KtlFLNKI8nMCnO2me2rWSKtCsCVriDrusB4P71nv63C+3HoQ/WYA
Vn3jioxvKDF6Tg1bFnx/kN6trQwk2G4VUs/pqOpa29pRGb1a29hsxhIYCuxoPdyBZ0mboKdyq0zh
u/Q1daoaPZUMNkImh1y30HXFl81TJeb/2bu/olUrriZQZ/mmuSaxgRQtd0iYTdEAJvK4gxAs9I6d
8LJIsf3ROU6I8jh9jQB/avMiXFdAJ5sHKa14WRYSsSrWHsHM0XRIgSbdc5rml1mMPRzMF+Rm766i
7kVhUuA124OUakfDG3ZDed/BJa0Mf/4TiFGk6g1B+4YeyQfsbOFZdMpK+k7vjhsTlJx88NbaNiB7
I4oh60mY11TpwyxN+UwP1pGf6+LDXpbLjz/2XIfG5Vg/jiwqxY+T7Tgg674BVPxVApyc9wvrgsw0
wkZZot2Nnnx6/VShcDBGIRHn92nnkpRO9HOycexsPsX78KZMa6H2SHg93v3CFXWND0+eyOD/FOIZ
B2FnX7oToX+1uMdsG+eDG6HXuHMW51zgB2RYIqfMAr9x3guzYKJFQUtYi/KoD488Ns5nnRWT0x/k
UIlHltFKAbSXsG7+XSoqqYzcG1q5DEdiu2NWYrtD/zftTAjLAE2ZN4PP+RNZ1JiwKOz7jtEy9NFM
ghxOYqcfnVwUWBFTv/KaAajLTGjzBEj9P6EtbkqzJ3d0DPREYhKbL205+zG4LdOJnq846OIkpUgJ
74KDsdffV5qZ+tJvm2HCo713dScLLAFcJmdLOA233GxAlV7DhxkBkaiOim+exvKdiK2MfPHo9nHo
E9YxQDCgSbpnAL3Yz8x5quwUG7g5kA2pmvMozm7IJYG0auMye1hCsI6l891Xlz2OLu7THL0UDrBA
/TuKz5P4FNnylxB2AKQNy1odlni4Vi6W+xfEd33MBbvR9wywkgQkAnvIJ7OGhINNdWXnMpEBLWOf
gVok7K6bQeYeF8QpyoBOTcDluAl9s7WbChfXKgZEnryicopkYRFrjGM36WxCL/xduM7RgEetdpbe
U9jKo8vhHkcX+j7YO01FhOGJXd6+7hHoDOSa6Uo3hhNgrW8I/bje98OH7l3r3wUOMxKR8tVXGUbT
QnDPzG1NP/kWpwzWkkeGazQW26e/tfUIAuNT2Oatmn+I48P313HmOYw2KtKlq6o0XX+5w1wfRprZ
YRYLynZ83E8myq6mEE1hBcUsErssKHRsKBesShcCl0+ZVK54fadOLlg2oST5PX+nK6b/xn+xw3Pa
UXUJVrrvSEI+Ks7p46xvhAQtCyDwn01+wm89YQWlo4h7/NcUi74Q5n+Z5jL+YR25Qb+WFBccMtUs
fFtPs0+3oj27nPcaBc69pOclXS7mg7FjOUptHOzvCSYZj7rNgpaj95kX4+MTe5sn5Gd1u8SvI2j5
dbmBokaBmuF/XBMa4fHFMNj44ArRvA6vmbegCiEsV9qx2qrYsFGxkc8kTtM/SW8cNntKNbVLq4V0
Ou1ICeZI7nxdfSLrOgijr39ITcmhfI5CsLd7FLGSWCtt/uqy+R581hgfDex5F0sXv0rIkG+CKbMI
fv4UhOkKbZjQtAR3werACBbrVgkTp2xItR6Jo3fZSp9PYzgtjVGwasfE9HWA7Ta2j7YGtJEuQTBE
BK2Mekb5cx5N5RbMr7Af4X1ASCYrIrm5KrkVwSvGKHrujH6MVxt2L4k9Eu/bW8YAZzBVHscwPtiC
hfJjj2Y2UbubN8C1n7nWYKQKqC+oL3h+ZLPBCW04RIHs5OPYCuguRdR6w3stwHgn2XrFCAxuBke9
vrWLBk5ADwppbNl3rnold6jqAzI/vw1pEAYb8b2pQ9/PZXfzZqH2fD71vJ/bZuyFDsGRZiqigTkF
0QN3X4fhYy1JcxZ8otgE0S5d17yD7Ft5LHJBVfCUQHG+mPauvglVqBIiTbOaMM7BGPuOnflT8Vjk
HyTWslyeQTAXcKd20Pa8/pKWZwiwxI3k/gAwLbbw5rb0Lz3it1AgRvNq7I2lIJQ/o3r0NELJ6On9
0FojPmpx3lxDaG+G/7aJru9OPsE5dbdBoru8KCVrlAX/UOperbBgzAlPVyNzCq4Lm0judpzErv4Y
txlOkNTWkONzhPiNBbNsQJeQ6RWLBPd0JKLViJm8mWuhqaHB2bF2tTHejbHSxu5e262srbTIIqlA
HhE85w0VA/dGgJ03/1noJWMaeGq+I1PUIzc7ridxYxmAZPhpGRdZLXeW8GcyG5GmGp00kV4sHipr
lHWJWl+ikDLeCfGIg4/+uM7RubEEMM3Wpn7zSWHjGy48es4oIG1O9zvvrJgGCLdw/g86BelQ4bGR
aZCjQTKzU61VE5+QZwXX3zBO4H8feM7gQddJcJv4snrced0YbdARHLspEU2xxiGqc8J4PC53sgrC
D4CkmqTX45LEHZ4cFViYiHZT006UE59JL/8x6M/V6vy3Tr1wUBvvcWStw5t8WU8jRPyvqwVRJ4FA
8ZfO3yNEhiWeR6Wj9Tkz02OCYvDm0FtUj01tqr9kXfEbMZ+/gRuy2M5QInTcMhmb8kk8gRzNqOWZ
jTj0pCZcvSV2um0KYS4Z6olOmULlKxur9wAdBUGZ0165f90Wug+M9MivMJ6HlZPMZ0cQcRTaKP3g
19reT5srt4uYlVUTNO7Lxdd9jipAbQw01yaSNTMful99iOwVcYauGMcoIAFClkyp0R2QuSigE8Wz
tayqh6XeLGX8kQGPYA6XshEn71DkMW+ERCFhcege0m9RkU4o7zxUHP97V5D9/RrchfDRMdqCgjKH
UGBgxSDmK5MN+BY7VfEiG9ookJm/a7DQUZVlvqC7cJUWFqawNiD70lEDl+yNcPy5KU90qtA58VJY
kfX54a1PaeKLh/74LxXTj+6tAI7i5DR5MmXS2QdlkwnvLsEP6/rEcBIwzpywvUTsX+Mh6OfmUI3Z
qjsSshbLIvNgI7I9HVtcJROjohCzwOblz/r0iHwkYwAwAH3tKtgwHpw9vp44qGMLmiG18JHOLr40
OzEp1PHbavkRrZMGsyvtY8PAae1ORzdk9AkKEFl1AmhLJJwGCgkq7AsEowWct8IdHN4A9M0RVCqO
GrrrBFPjuGirwfEo5GGYdW2ypfH5jHqWEEYEDTYgk25+QMX3qUUJAUzY0S+ss4d9MYBYSNGIPsF2
Rkturhf+KvwovK0nsVPx3yKI0q75d3FhijLWs0YZ+Pw/D5z8yPUCVVi9urcOBeJEHwFaI6NYyj9E
yvkTx5zDVyDjBAfDAiCSHJljwYGNYNv5TgYfspwU1LlCzg/2knYg6Vg7HMm/I3AbzbQgpCEfitLy
WSMd+HjZEex8qOV8yK9wmngS0M1e/ez4PR8efxVOcM8g49th0jzLagtpOY0tCLkBpytJqrOruwGZ
rsHTg0TGhs1BicDE02dET0IK7hy7P9dgPk08wdHAgK8VOfQzoV9l86LCZxE3VzsaBSQaicAaGg7N
p+OxTJLWwM0zSSoWFocthtnGyRwgmRhZz3HwMDjA1tYGJ9CgN3aTL0kTh+cRPvZB7GbgJ0godXnV
DA1IE8abcvQASgxRXVtT/qJB/n8ftcKV9pTKMq57LRkGUTLdT6gIerqllDXt40l+SiHI8H18gKfK
hciqC02WaXm/BAXrf3ZH91WIFfLM89IPAf3gsprTmGHXA7F4ki4yMKdHHqtU2smncRv6/jTIU0r4
3Ge9KhUDMcm2Q5QaEsLXSlBzaUR/HGYOqm05Oq7bJHBBjbLfWp3cYfYHApoIfOqqjzVG4Kmm1vGS
U0dm0vGgu37JuMl6GXfOeSy8y5SyddE2NjL2V8YSu4VqlbxEnGfoPEMONEFbSYIQrcW5GTAueMUV
7Zrve5cz8+OjQEU33ADqJ+esAWQ9xv9zp6ZNvTJKaSVvnwNXtiTK6d3ibcjLPeT/ME9ZMyYvpUPJ
OE84l3LQNoNPYe77s5ae1c0QK4thT/JA/jEPNni6RAgGD1tCRJSnfZOgluEOl6tLcikKezzrJ77D
gzPMTMhw8BPnglARXIuwEEw2JTudoHh31h0uF2pwhsH8jJdmZxkPUVxLESssngt4AuCp036tYXaH
fBRU3s+6If525hoH8PIvGEm/I9tPreiH7aWQx0g+lu1uLgNjBwAxDPrklk6DjXMj3RYEg0Vh2kVG
vrSKZtCN9s1Lgo2brgBlmslHPixn4ZQ+b7ym/rrb3M0hivjhDpdFp+V9XTcum9/tj8xCnz3dyKBb
ggixacU+TxBjKTWMZJJ/ILa1lqmtoQ4Vv2F8AJGW3GfLRruRPxUQmXFmoi+89hFs96jZtwYOuDZP
9NqjkZdl6hGFeSLJGxcQiM+GxyZFgvUNCjyQYOSHAN715GYTdJMSiKZgQnU5IAMF279QdBpjT+XU
gjyuRTnQ8uCe9NOSqLwLf9lydFzBDLMuDlse3Vlw9+avMepT+b/RF5TMugwIDODR/QFnxhOKL2NB
JlLhwMzPjTVOe7ae1zzCnBiIpnVPPsCelX+NmxOPsbVWxH7FuZCxnZfIvWEFdxwWVWj7LZm6pqdh
OtHzMYdULPJ5+wiewdPXR4SIkn9S6sV0WN7wJYFMD2RysOz1RlFYDMzK1pi9N99VeRVEWarBqviQ
VjMyUuInLdd/qyLJ5VAHr0OWDqu71URkwicNyN6n2hgeYJsQIl6ymQZACWW2v3jRLfUrShUzgGUM
sol/ROqk28mGw9BgZQlS6PC17F2vHCEdYHxi+UFlBEIepcbHHGn/wqk37GgC/xpfH8ZFz1rF6zjp
oJQ7xv4riUAIhwcjW3foPqmt8bUG2xrWnu0vlh6lc/lmUkhq8g4X1vYv1zDtUjamt+JNpVzUVJBu
zhwWeGPYHoV1mZM4Ii/JQXYO85xUdhmBNfNy88j/fhURUe5aT0otPcJko20vS+NxqkuU5qYIpi/c
kadiYNdXshUbD3jBWaqpNG8Sz4QXTrZG/1xjUb2OcQOjEsQ4P2OQFIj70TzJmd2OWKbFapp97hiK
AhSL7H7k3GeeNpk2Q5m47npThs032kIHJaySybTwmNV5hIvrF+6KhIPMAx3XKP895ntRyBC6kLby
ZIURyUGhLZ3KwXpkXAShPP+YOU3t8Zny6aMIIMSM7zszvmnNQSof8VPicL17FwW410eLPyuCL7G4
LA92uzojGIGHKLq6Lh+qCNRdsbFYLdMgcOrGo+EeFBNsPDaFvGf6lDCtitzuT5HHyIu8dEPhcRvi
ceEDZ8J50DEc7zIjJMy0ncUNRzsPPlCZQs+oRbMbROo5xkQ7GC0CitnArFnx1gBDwVcvW27NPR2d
X0Ps+klNuHIioeaqjIht4ksBd1VHyvE7npnl5T4ZrfRcx2wc3B3aWPaOZdyEv1Pc6d/mHOmrYUPv
9OehHE04ZrzYtmEwKtj5wAp0F+IWXX38yf2OYfI4QGMDjLz8pzDS3kunCFrIeENykkDjkQdJksMJ
59b7N+JKXT1pjPNXkZcGfdAzTQ2oxgoBC/HGI0AS4jV+5nbarZymOi1eHxIuC1CB2L3gNUY5tMw2
dqpsFSAFMLpe2NJwOcOP8BRNS2cxQJrIFajvkE0wy0QGTw++29DYlpNW8dPo+luui1PUDVzcc2eH
YSoig+lD9IwHTy+7rF64qKwS6ay6xPloWblg4UGMnRMYY+JmG2ni3rTRrGx5QkuPVJXjp8KCe8Mb
R2yNZqFaH0jr8r7vmXXgmu6zYcRs34gJaRL70/KfiHnr3Su1L+pE2xfZyBdefhdnya5JEFPqSTLr
n5FJJUsM70wbUp3fLm6gGtoVY+9w7bJt3nW1Ns/bwrJRR+S/3cIaTWCKk6amWYfokfHqU18TPweP
pZCxVI1Ugm16S99NrT5pntkMT7z1rggRMVS1uH4WstVbAgAAVzZI43JM5rmebzJ4YNysePfQfBDP
lBJ8GNXdn1sFc2oMxj7OqjGh5UwDwSlCdfQZJt9MTcW9AIFPTkrMMC5fjs6UOJeml5ZH3Gc06S64
HN4afG/o7gqvp9EXaxLmUo7QAdxCT1EBYtPVtVXAMTImf855rFhNxLL1nRTYKvblRQLSDJmQzJL8
2Ahmqhvqfte/G+pRf7XaK02QKMOV7GmYZQ/GagBs5SVTVPOmJwXvmLyiTgZ0FLqry7z0T2gukFpC
WN9o0810KKzX48JOlvmLyysRNpusHmU58WfKdnABuICRaCj0rFkJBZ8yoHO3gy4WVcU/UsxhlmPx
AdMKsdQBIEpDZQsto7rYkbDQyAoMWu+siJRN2wqzFMPZU1c1FutV7s/dLM0uXg9fKwdxbRYQdi9R
2jP1vO5/qHKbzWMQwO/JoWd07miJnCICMpoq0eB84O1VSP7eFlQkC5Aok7H6hO13F6BKU9ZmCyru
kzeZhwKOohSChjuEqw/PBwIIbSgJOqPI9DhFdBML6Ij2oKDzSFaEjp1qeHbVeIVUV31TXkGwcqbr
Wwbj8eQnw22M0Pw7i6fdyFiqZi2HWkWK/XmnT1igRD9VwtSWI6Pk7UdBtPLr2eChZpDfRCnoZ3iT
uw3UtVYBclZ1rofBRNDCNOCubPiaBjotRWdTp0fyHP3ciflq7XCvzs3cX5rUcnbn2CIs642i0XMa
+Z8IjF9LGznPQwrga/HzG2qsrHbs3g5E9H7WcAYq02YIvwbGXhApWiuioFSTlshGqb0L81uy50OZ
lBHkhLtuXmiLglkCC4V5w8pmLZshRNuUwbLkAVFxT5t8TL3A+e4TF4+dhLLDDGVTszUXUlvvtX3U
kOYCCJ+bnDGg5PSz4M0+t/uUEy0myL04gDdd/ey7jLSGU3E9XRlLEfTsKXbCt85fhjlTGKy5KqJn
ldmZdYQ96F/TKZRUIG4xL5P4E+tZqucWtzVOG86R87p440skS+URvmRHvoTsXQmGlvcFd8xfzfL9
VrOFFXIeBiH9yikiYcn5CAH3bPr6g+KDX0DdyFmZnGJAoshD2+G0VGHPFnfjN5xxdol445OMHqnI
Nhma3CDas9KGjoCd0c+Nd838hAto3d380W1NTR5HBDqYWts3gDDMibKb/tZ0gPlapWGvYohpIXOO
lTTQsFJLX6uuuwCdc+2MFpEuFwJYPnXjz2XyupqKK1+X18TdTEeSTirwtBx03YqfgWHEme6a3gos
SjRxHdxZQ+dbCH6JWAThNtnbCaBU9lSHp75aDQY2Ky78OE7+EfvO1jA0KpNe0rsgGOBrGHD+UXU9
hCESwIFoN5J09oi6x/cohfQxEtsQa4seRDkWhPp5iQGL2+Z8VDKqOT8gn66Ak12ZS3/1oXdIB58C
IegIwKHKXxEwpZ3R9CmQwaEQMb04ffm/5ilN8epYiY4X5qjCWieidLsJIYiDSMs+wKqkPR0YQBu0
j02nBt2hVZGba0xEyzVpJDtA8eevk9UuyyJM3hkRinH9Yc3jWJNnJl/WO/suRG+Cpdp7MgY7VScc
Wj0Fc/hEK0wZXVexdSVh+GpZ1L00NVXyQBRzsCJgRSpdUUza6SrgVPcMZGgOa7rMyRiERD8tuxcY
ZGyeRcCPsJDdHXMLfR/iW35mwgcyFc4Q0Jq2tFXwSw9h1fHmeHHx3uLEZJvdeYrUdlP9+oN6nbG9
x+PeVBYQrG2VX9xGW4kLYxP/6e6GyoI7rQ1a4RM6z/rjU7GxNl42dS5apnUQjvzVnOwLg8hrXoMB
ST154GxAJa6O5xqrEH+47PKDDuxvS36yijUjcLpWnQzSXhSAP0x4HfEMwDlPRJojoA8ADoGQ10Dk
UO+VJlAPw97KjAGcD4Hhfs3fdKXlHEGmakt6725e3icfsFq7Mppcp6fufLFrhQVgBndpD2DSXUOD
GgBtW2eBw56jZaCQzHK1H/4IRQdTcBe8+yxsuHWBgOAIvC2+f7a/LXIs3wf2daaVvEeBg/Ni460D
pyC19L68dig/HcyLZDGSMlB0EGr46CE0B3k+2iAJ++aoh5xMNMhQN5GFXSsKHCbgM7Gsdr6JnzI/
xjld8A8cAAzS7M8NpgGO95kV7pHPMqaAJgU2qAMaVwg8LycHIO6C1Yvz6oPeBJnJFcY+UWDuJ4Yv
YQgyhnyVDeBfTfj9dr8xu3xe3j1EGjiZ2w0qMuwdMJ6xN/W2Uv/dEavEhjYhFy2erPdf1sVipxiY
LIxOE9yXsl/pOJia+C3TGp9ZNYsEwIxB0qajCKBQj7kG9Lb5Y9lviGywvQ1cLtOSdGI8N0zY9OW3
E980hoaM+RIJhlvwhnNfEW7/Jm/fuX9xLTDtYb0DUAe/1F6eJB2YPqw6PfmemxFfNp6sz8IH2EXI
dZSYSOXgw/ZtMXye7yvIwugh6wY7AQ8Bw/w96LBLVMsDpsKvDkZ1fi4JySYLkWWAextXmX+Ay4tV
Fp+PYdMNfEVPq4vGaR+INRl4hP20DB6m6xXWl0Fq9BSx8Kx/J0HtO9UOHbw4rilHCJDbDAZK9aKC
S2GE81YsnxtK9w0Vr8Kcod3vi09/Sz/oXBTZm43dYnRTGOckNA1qDiAJBFBkWTpmjGBAQJ65FX18
9Lad46xKF0zCA/FGcU0bF5gUkChpZldFNNARx4VLko56nz52O8X2ePX+I0HB1H3GV7gFddbr6nrL
8oEMF5YzYupOXylngjoLhlmYJrwl5E91lt8a5fWQsP8jqT++wc+fSKXIzPXDFZewDm5chvpw4Uca
C8baxh/1xkjCVU+2ARXY2nOgTLE6Mm4bQ5l5ig3DDbLe12SVeqluJsI71A19RxkUR7PWLUr6sUzR
OccxKw6YmLwHnnzMDW7fENU8VvYxGiwRnfkblsVbK9RgnztfsYPrpuLXcjyas/yDD50ZxPfDTcNa
MEDyZYLlI1ohrGLW11NLFAPmOMb+Fi3R8hhP+XIxgw3gdJL6RS2JprPC9WJxGBH+tHd5eARjBEEW
KMrhp0zsBb9J3032u3tq5+PsdmuJdQVw6uDEajTllHRXvqRwsLJ9GaBKD0ZInvrU/cqmlh5dvxww
awQ3WUYxzzVbyVhE8RnVSBMoqzgCkYQNNPeYUrNBPKwCA82JuzHCZ5QEMO41nDcHTWdM7BIvVeBO
7CJtxh1EqzWKrwvYi+IlGpGAjjbjiG/GYan8u8HMRByW0ieT8XWhIVzcA/sfsXWS9nP+ed0GDzrl
Yut0v4WC+FhBYtkwHjGaTOnG5aMKlquZvJOL7C7Q50cqujUpkYLuslnUZeqQPCL+QAz6H9nOmshJ
yP4yZ1NxHgvRRqNPpJVinlp6e6madn/wlEQjG7FtfMYhd3QDJ/bGHhNAIyBbiAyYRvXa8RmJuWuQ
VuNz2FgCRcCAMX3avLMkpvtZHHWYSyrHUejNcQx2CMGEygBaLWXDtd4zoWLesZr+wzcJZ1CGuiX0
bKdJyAWj4GnifFS3cIJaeV0mFoqjEiOvrCvofu0hj+JkXMgRfUzP5IP4nTDVbGag+bgnQdBQOA24
ZVHxcjB4tMq3QaNmeeblVsowamsMQlxMNs4NQVsMt84NGMQ7jZwHgMKGQBouz9ftnRS2fjB9pfzA
nYeyy7eKlG8eAFHCplyth8z3F0a+Wmev5SuZfOstHWAFbnYu7i98sGwrYDV3lycHBjEyevalbj5j
Tvt0Y2II7OrgDinjK0dWdGGbyJ+1PE8B7rf0bNueXqhlASYnqa5C96ooxUdOaZx1RRt/FWiz6QMh
wQekU0vpuKgzu4jrgiHeyDjHj7XOBsTyMuJBs3ulXKhvKwhB/k1OqeX5xdvNg5oDnWsknQ/jmt3S
nDnRSZO3/yMUaRK12z/BIN1WHllAlP+E/am+uknXVU2l+YmQ1P3IIW7b5ey81ZgNpZ0Ylsy9F4C9
NQL8gtqoOYlMypvGXCBERnabzUTTatzL29Bd4iLeXFPnhM3pPj09zl5yTzpO02xaxIqWPnIbsjWh
eyz1xv2piALTICVW/uBLpCybYh9K12Cs1ZZrG29HUawfjWCJLG8p+0fqvJhSDAfOFIIClRwZ20qo
KHzzN5lpe4nio4wPp+idzEs/PwY7bSPj3RUL3YFtGm6SdAn+ZgiAUz35HbZE8y+O32vGyCE5dbIq
NssKxuNZ/MUdYiOISRMXYt5Bzdl/+PC5XAx++Z1zIXd9fwiPnEjiLX8FXC4XstUcdWiPj3zSRXp8
mgbzh22tut0DDbOdfaWL77o9ujQIlb+XSENVPqcWrsqSgi9m4e91y2Tj67UEYRP2lf9R+D9qsjyc
eEo40LQYdU/XIEOVcAa+9y5izomMbzMp6ioJulv/CiT31Lo/jCxrpX3yEuarCcGlcFYuQVFB+K/j
YZtq2prdKfRntQONA4QEea7KWGm5GZfs/qgBMiMbFgWAuGHMYWZwYdybsI7Il8QXmsw3LJtjcuaP
EIJYAx6aur7zWXuigOAxaIl6PjLMeolEZ7TZI5hc1aPLZT2bAUq90S9xe/azX8hL+jMuZLngmzal
TdFNkWavOUY4k+wXmPcYNij5VMvQTPkzXk2oLm7hr+0IHnhIipskOKZqyfrLt8XfX4wenPrNfDX1
n9r2rMvg72iXZqcrsdmPQlj1yAys5GET4xpFpq/Q8P7Epa26SFiHsAJuZtqesnDaZF3gvKbLQVPl
OMMbefC3xcQK1O3uQPABJOwIy7CTTS9jdjYxZxP7hGSmbb/Mo2Z097jyvqijO3bZOLtibAWZtfeJ
2I4kaPFQbHG3yhg5Q1nFB+rsAqXrFSg7tOYwR8UzJKbrGeouZ2nv/p2/e0bkLFyKaPgCl3/3osG8
LlORIfY7RVRC3Lf2MyNZ2SH1ehJSajvkZD5jPiepiFuk9kQlNwtpCfVPnTbYaO4wkP2qJ83vyiw0
efMIz/uIqzAt6Si22C7lIiygKA3+3godIFqN4bYUvdlyW6JLyfECetMFgpCz7z9fLZUAHJkgdA3Z
C2MM6P3DT0/FTiS6s2W/I8DAQhUTM/jQUkhmai5g45im1COynaXsWF/lq7CxRnRKVTuequUt/BYE
M7n2E4v2O7hK1YquAlpq83Fbo1ClTPwMRJSkQdoznd9W19M19/QUMJ1eM8mQe1CfLdtSgW0qpaz+
aSW9B22bTLM1pn8A+yjtYqMkmFc2k7CAyo/D6XKB8eNAlScqMn9kis8ycZv8iNYP4tKcUTUvrdnZ
slqrUPL5m++lZpN3v68k1gzog4exNVoT4KUTgk4/kZNzdYan2yaGrEXESxhA1lBuYFvZhd+cjUKD
pZkfRprzuB5inyc3dwrzEPDo+36bLDswLT9XMbmuxgAEC8SWecdEeWaBOvtOjGl2J5j1wfCwpet9
F2aaUqgvqSlz0yTqUHla8/wcFXSntgWmOO/VALtZ92NcG8wdDqne9NH2La/9cEoQGW7DxCUHxM0o
fYcT5ptyRjyV9ApLIS8Jo07VsHR2b/CeH+hGHkxtPtGfpR4gD+pvPh9JdRCvKzQ+pTY66PYFbswV
AkDAB57ZItFJGPjnow49oQI6tYueT0a4jQIzXQaDI8rC+1C4ChAY7H4Wd3qzK3VNe54uwu9IwfMB
PLJgMi3M3qREHJVutcvTLthCM968+nnZTbUFF9tTi+xUuou+Yynyvxmtoy/84ejlEJT/3q/JVtXf
JtQ3SVvL1cAsmGQe0XhOki21EkUE9xFelSYgHWgh3QVzsiAaLsPkO4hCsmDfF9BN7qlWlpg18epr
XGuaVaOWfAsCG78Or54BokjzbPN4sSnWDWO0FMmL9sK4PD+Uk8Ino/oDIVLkEHa3hi7xGiXayBG2
2PD45G5J3QEo6kQuxFmVYA4yL0HyahcQB2XRXRsuZkz3JoDxM35p3LF2zlqDCsn1aDrMvq5X1Ak9
k7LCqH09jYdxfzCW7aLPqR7EXnEBJ1vTxFd43pjdx6ze7ZBnXdnI8Y362QZCodrX5S+7ye7Pl4io
Bp3Z1WIITUmx5nf37+KxZwssbD42nPxCNsGXc7eukD0l9jjEtkPeL09QXpdnpwX2VZRPc+uVNMyi
ziFGHe9Nhpz+4EJ5kbOofm8OFsEUwHWIkV9+UHMu66LIzil1BsW2cSA4F7XnOB6C4kKWP6BDJhbk
zcjCM6kpOuC2+MbydOSLq9uOm0JkTo3rgYatifzrV58qqt6zhIZFdF327/SYlOkhKvZvtZ21o4aL
VIrUtWxabMReLIUP41uBHnHGsbbIpnlVIPzOQOOwa0lE6DfKf7DHeSIwoMkCHv/2fEB3TkgLfBKs
n3Rsnuijlk/XlPQpVqnWzkp+BiwRZZcmUC4nPx4bhgs2duLKALBMRrQWm9ObnzgQ8btNnNlQot9O
b5yhs5Dhl6YuoW1X82jiU5eG9VkVDNQLpje59j9EYsyz46OrfklSAt4qDEGoGg1WN9leQzyk1L9p
5DAhE1kX8AyGAjhJn30FhF2aCmYGsgmRU8wopGoCb8056UV/0dG0RSnoaxAH55VmNnJhrEa8BhuY
YwEyOO2J0V7NdNAmn21YAQ2JBSOy1Gxhd5sifzs5RPZ6EXJuXwNwXM7gTv+4WjEZYuZlRbO1oYOM
VACHnyJlVJMduDNcio93I7C2AbMu9yaKC7Fbl6G+qOL/vJWOcl71odX+3p/yV8MNbYKhjPkUeCz2
v/pad7juYbhI44fmdK3d6ZUTEpDVzRmaJhH+Znm3H4dg1KscOtFvsx4lUJTN8bgEJsy3Soigoxb9
xTdolvo/VlePmXuCtV34K+ZOaeGMEKPF8TiI5ymrtxT02c1IFgVvaXVVg8W7otuO8MkFYdoLQ+//
bl6viWNRWxV1b56HOZgTA+UESaUQWEiM8928zPoz3uqXFo605Jo3xA2G1VUojA5yo7m5sDQJJ6A0
aHycDU3CeAvbRX5tSWC3cv+t3uEOKka8lIPe0YE6Wa/cXJO1hfujmtefxVtRIWH6w+9x9AOPTG9N
JF86K1wetASOeF3qjSIyYYYJWp0FPGlt8/b24apv9Zl8d+9HnamUt1ZFycsgKiJpxDhByF/7otG8
Txd1e7xSkyMzrkN0d1JVKK4MedsTdzVj/4/BPT0DmSu6A3UzNI0Pro4D7MpcADCbeZcuM/eNsXK4
HncYI5IHocgjwPJMRDXKte+m5YELS4GDRa4bKzT208oK3FoT5i9Hm3Fy0wX42K2h+WqM5x9Ru1C9
WFRJ+h0nRloqAjTrtnb5/5llzP1L2dvs2z5AeqPgrdeM7kpO7eZVyOVszWMHHFYAQyDFzjG6KACL
o7jrxicLliCJz6FEmqpkaxM6gZ27zeOWhDTS217KysKBTFuzzSDWnV6gyiGi0VVE8ZaEKqiQvZVk
N2DJ7HHYmEotkQQ0jHtwRinRjYGxrd0lqRlX/Yy3hcqqTfLZXf66wSsra+sgktGGijHh4sQpGBNQ
wFw/hoeQe/yjQpQhFdTq67XIJS5Ye3wFEpNLJwqlxL3AeZUJDnhf+zZD4w8acsF1CFlN9DJSUzLn
keFWroGDDf7mSae6IQeEoxHMPkAYxz5KgNZHaOodO03FtHdhTgDoswLTYjhNw94ALi73Ze4i8prP
bdk1oWdDPy33FIWcKw+f6cK+RQTRGPsErRwYg1YxqMtIerS9SEuo16rtwbThaIa/WV1U4LVSJN2X
LJul7S2Z3Lgg7EhgB+u6FxQWvAIqsZciyAfhy3YNafOxfayw14PaTtlHVRt3CqiGgLRCXPdYx7ZV
K9sBae1dVeOYxh/hwI4tw8FqHoJvQvM03kd6nO5GatM6jFWZDcLw0BGc6Dg7LZ2Yz6RgOhsagwMh
EQKTSr+l09UEK+fhcIHPCcLTUjvD126rLcvQt9tVYZFZ3Xvsl/2JtY4va+e4UG9Q5PRrDI5K3ddI
oum0K4inaN8qoKbcMI6BLziZNey/3T095HSOxYwpojDLXed0FRKSkv8vEHNLEAdYwTofZujXsKsn
ivu9GoGkU9DD8t0Nm25AtSxoN/HRDzaDfeznDu/0judGesqqIgy+y79HR66Of87v68knApa9be+0
QC3EgjQzzS2cUK2o6LVt4noqdQfD/6mjfE7lRTOz1arUXiJWuowBs8VeR+KA04GFHO+WQUC/w34k
VKS17yFgF9dWKWj8UfBPi/ajlcnPdMCnAwXwGKhHiYL1W12gml+yWJ/UpYidDvOpK5hidxHdx4B2
u9Fs0siaenOHtCajMv150mg++yVsKmH0rWl1nb/TD4FTBLkx1b64pGkAntep3IbHOBOPCED1I+W+
n8EhDV2cbNbStGZ/C43+PdXm61pOZRO2EPOa2Vhfvw8y1Dz1hTJqXgZLX4VBwkjsI+EwDpIdx0ay
QhU7dx4UHC2keRWFebyTx55YFxyO+vyGS2cjquCEg7lpdKxtTuATxi081oxuLGEebrDWF89iz7zx
jOGebNrsiSBl4EFvCurFSeDi3sH6XhppsQU5T2P/VrVSItYgJCfws9O1OVPU0fQ17UnpAUG0m6R/
IYE2NR8pnELQGGwwW0UNZzO3lQ78D+vNF1FGeQOkuVcvYyYZCsRRo3/04WlzD7hroYLOYGV1ij6N
OZG3GKPLs/TI80H7CTvh7OYrZu7EowuM6uuM2Z22k7ehCunaxe6udMw5f6ZEL9DNnkPmfc++SX9F
5NPiFwHe2in/DO6+EinzBJSH79+JsNOpAyxSGBYXKd343/Ir+LvmCtVMmAUzeL3orNrrjz+yzQ6d
KjPBl2Jcl/4hszdVSlFjfh4x+VIZ5yHPI08jq2EloqyqvezOt4MMXxyhxQDUa/rqpzf9qMaUMJXJ
sOAn3wqToC7AWbdKjo0cH3Zw9X6b6fzhr4Ebh+xQ9iINMySiwLQIWvZBcQ9CRZSZ8IuWl0dxq0f6
EpZto63Zo942doN0ntVcGQ4H48KfYr8hWUi68Qm+mk48hai+EP05FBiMiwv2aub2EsvAm41SOFvf
aU1WK5MrIsJ3Ft3bq1jhdZm4vbzpJ8OOo6B4EG+4A/W0pdHperko7prD/7B/XghUJQ2p+8yfMlKw
PlVpOlh8ZwIROnl0LI416SzPOJQ5tOFrGnRnkMqGFQqnVjzJKEaz/qeX3IY5swDXtFh1FgPaRAwf
7en0tWIulqe0m+AzxqEmSpQH1U6oPc4xuf9WO0xO4X50roxks3BEMthnO4fLhjOTYhh9eTr0EXdl
kAjELZKylXLsTjsU7Nz63xQ9b2OmdgyOwna+vBSlOMCxu2VDRYlWHHMUEbGCmCSq2SOkYKy5uSQE
iekJ2gWKLTmUJ6A6Ywzfipz4d47gNlJrGa2eDWp2TilMiurBwNzL6PcML8KHeriF6v2bVKJj2q9W
T4V1lBtql/RSAGuKW61T715/6vY4jZDP599B101X5pkKSet1C7TPEg5QQEWe+ejTvnKDIm44buOt
PmSISLuqNdsuMbAcbEGcC7+3eNGCGyhxqgzbNeQxZm0x/B0RuDvwPpGonMcAByjBuRfuP+zd5oS0
3rQ16nnbfqPspTizJVNpBD6IaV6GLo6KollB0qkhjZA4bKzLgbxDiT7UZ/UYoQnVMv8MHjlBnIYq
VChmy42PqV4HKdYzhtXzvELAebIlSX+Usqgnclpk9E7KgZng4BVJuETd0OIZ8XNZHLsw/6Qdo9ot
2EoJGjpbNVOR9woIYtVu4+TcdYL9d287aZHwCp0Cg2yUr4oDkTVA7GzojFWL8PNyvjgy3RpjV7mO
F/j+6cnG9NgV6IlEhxIBHJ99JYbP1ju8fhog/cD/2ND/0JvcF1dKKPkoyXBBIIXXR2g2ybX/YYQX
A1LxcBCp7KFbvtOPFOY3jDUcMn1E8cEYJXw6dOgy62bnBNRid34FS2J5Sf82XNztWaQlkdlOitdx
UbijoGpZ5WjP88qvLpiSx+lOq3U8go+5L8NkhwywCCEvUHCvG7Qj9fYMFhOLx2MwM8ICnIdWK29t
qGXMxQzrXRepQyfdJausxSHQfJShx0stAf1BiQJlVPbUNqQxVpk8rw9jTTXpzvFt792i2O1Phvqe
m+qCEMKl8OKdLA7zS8cUTcuj4BhBICrBeARqLy4vW2lgKte95utVSvgESn3Wj8Ou+UZZ9PYHi5rH
WuLrquztfv3BzwE6HMg/H5B1ry2iSKKbQD9coxWVZZbL6lBgG/Zh3U4mL1R/AIhlI3Q3StoOSkkR
CbZxLhHblejzpWHmk3iCjbsXKQMGiWG95CNj8tSdR8I99R1zjEq/FTeOQJ5jGl1fL0UflL14tnG3
SDNCEczxu+S7ziNa2DaUsRe0iDRYLkC7niQ8vZVsorPorB6yH6z+BRwT8Wn+6hEf6PMZZFtP/VZC
lng9jcH1RXpVwfZj7roSOy2CRq4ZvtxfonsmnGz48kc2wQx6HsV943uVQCat8HNYYu9bFjv3CaJw
MO+6FjDVJ+Qv0I1YQj0dG6LWLKAj0jMxojxCjwKBvxO+Msy3fHOer2RZ+DNg/LxApWIGm1xnAQy5
H+k2zXMZHI/Al0oawhrsnn5z4N7pWgABcNMqCJeIvJEX6KqrgtQVMRWBSuGTZjwAXg2JoSfuDr1K
mhc8bLZEEL0fGkm0ItV6Pe9FvSaSM/gQCBGDXPliwtbtlhxUmi2BGVTOegAiCVL6XzGVOomnrj9l
4oOFLDKAV1tS4ASM2Ql0MkreVGKxWobuq78RhtjHKyRxDXWNFSVQvneAvQkwLVwT0e42HLN4JjOr
sGyVJwONFrzUF2/hULDdd1S85qbDFD89Z8H+57KL/51t0AYwtIjbTbY4iPYnDTPvZiiiIK6929GT
Fkk3mDI8dIUgF4HIv83fTNl8nHUsCoI4/KtVJVyGvEyjVMNe5KlQgg6bBN+nw5sGYcXm0L55qJie
iinbNqwC1uJtELqRYg83Qz2YN39orPw2hrKCQmlg5oEhxCQhx3W02dFVrUMzhYW0bRGGGpGq1BOW
CRRudEf+UxS15ZJ2bwdz1TjHwSybcNMcKY3siebgiRflrV57aNFfDH/rC3KNgl4kG+8oXlAuu8Gh
HwK5F2n/iT4CC1a/Db3t/kKOd9xIqg8rWHMCM3DW7EUcC8WncmuTftndvs0WjRG/yz5Q8mgB0AUT
pKqN57srm9SA21GrtxrvIjCIEPpWQfQq0lWkm0z3wnrrXH+OuAHysLRT2AfqeIAHz8zCUu8n1ukg
qBYX0+hskc8bENz1CzZs/aeCxwE6kfh4pLRq4fK5NNsx6rIoZ0Djmzm+w36A7BQSNldjKJV3Czmi
IBeVVYOR7Uh3GbvY7NZmslqvTUhr/twEIKI3W2KizHIGguzRMCVDzAgrw2Z0glXJvYjhnvk92hG6
wrMu16qCrcCmTklc052guJFI+ZMvBRuAuQII8M+b69+stKqbPh+bViyx/E+nabxzpyLFrU7ptnNE
9qRbioPP1R4hyLayTF8iWXjKZ+tidqMj9CH4pE8f75BE1YViXeQcRULhLRkU8t3y8gdhQXmk4sLA
+3D3ERi4CiT4Kp/mqs3PtMqnwfszZASspAqhDvh6vnUow0mGzpTgC25xyJNeFwZCBcqywuhbyus6
nLq7X03nEIKfUnWhOi7wtVEK3MNopgVosel9qhr6ugnw+LgL5prcYTaWqtwywoLA7pt5Lr7UBLI2
q5IhcNeLMNkX9r3f647QjFGvO7L7kZJLOoVVpqVApf6gx9uZOYDoYyFynadX2SFJbX9hKRfgf9hx
dOXftfHKq1g2RuhqRZwFc0VCUegeqVtgDJilBHve0X4TxeVz57LewLXbyglmFg/EQTW+LPY5baVp
GeTnFNlNtZiq7fx5rjBCfMCtXP8X2Oc72K9m/san0Vl2eyd5ABBEDwDStb06cflFAWexGD2utSZt
kjqyZKiVXpmKO4Q5m63pH9DCi3qvTzS22WLtXH38v/3E7E46vM/tLPa2meJ9IK8xPBBztGXXhkfk
SVQeo+j+uQ0Z0zKo4IweT5/mxEQySQBjzKDwc5OYkCNT0JLODJMlQY9JIc1BgcI7R1flVU9rVd9h
EJSSFv/A2DKanorkpIiF8JuaF2QLZBjS5Fpe/MLzV+jTGBkdGcQKQejZHhSMxQe5wLgWh+sEW4tn
p4x6yzdbUIjdqvi00PlCWuUuhr7FOeAENiYF/ATOWXtRsDypaWqh+TMa03pOI64ZjyNK6ncXTWdr
cg08dXsFquPC7oFm8bR3Ja9cy75PZErQagIcSDOtFw6s0Q1yUNQNOfe/AtafqYamsXbgLNvDc0FX
bm8mUfZS+ynIzCySlrn8LUtz48NSrQPmjopQE+geP/QVNCjjQ5hlr5GvHZXmgrilcZMZtYZT0zrd
F+2AMGJDD77puwDkKotq+z7MZ8UGYDXOaotPvZrwMwnoNMkwbn2tnNKrl652xnQAkO0+6V2DCv6O
lZT9MfnOLD/MVTS4rSp57rKxjrcnZAnPPpxlHN+d5Ook5t0FnJtldO4W0EAATFzRX4yfo8aRvmgG
j6uFb6jbKGZxL+Prln1kr3bm5hkUtOZNyrpJIKgxXZOkQUBgbsXMDXsfc4mxEEe1/CSqLIh5FZyM
WWm33jk8Mpup4E+7vs8jNeFAWGRZ0NFUy2aTyGPM65SeRw09SGIuBLaTh+IR6+OZ1w7OdaojBPra
tCubf8kbIgs1etegw6ij6m+moSvSlWxf/FwP7uV8VifjSDXXQnFhYO+aka44BNLrfjuZKUCdrkv3
OI4t/PQEz419zSdyTD02jxS5VO19w3cNZtoq7U3oNQraj2tnvy0Tt20XHOJHvuoHNy0I63iNBWs+
bBgDK39NGW0tCm8vo1LEfbUXX8UI+cm2ZjMEz/Du8ahkBmaitl4Nk5G+NqMiZbPPW1uptBcvIRjF
gVRH8azGQbBgDPESWfdkt39S/ZcfUWAw85OcoMff8fHNmST2e43d0h6/vwcU3xzI0Xlr72dAPxpu
RufRRFU+AV0i3EgR1ixhNIQjfCX5xHvmYrZpYrACDA8+I9sO4bZE15Sjwtd41txGDyRUJrpHDqp2
S2kkqAHDa8NiASMbFJHM2N8W2sEGXu/LYkWSaSZj5W05ROFAiNpE8HgmvhIPfNwgDB/L50fsX/Vt
iJBLOJLRk/ALyyVlWJVddd2ZUD++9jZZyspiwcFWWJQR8Hdiguv1RFnD8ffd0J9osGhfu5YxGYN+
sNXrf/kt8kxm2sI4LDj79p7H8MUy0i5Pxl+1HbwxDiPR9XNbQAzZuHcua3zBpqGWYWypEpZZ5PL5
QMTgbEPCSVimN28FW5VKYyuHrav9eho3+yzWxKwxkMi+STpsZ+p/kAVdW6+lBfaDyWPe0Wmjgou3
fzERD/Toh+F63rW/IKloCBROPqKdjRPKu4p3QuredYq+9sitJjTQx63IWH3IbapZTN9O1ui851Tl
+LPKc/ssTc8yf+lAMBgA2L+adGtgd4eAFFX5yOh8P3Vs6VJDyj03K1UnoHKaSn6l/6ZHz8/R4Gkb
C/aIzSstKWSCgqsFzqEcB8eRS9N5Q4zaIPmBvzk81IoaiISTtk6XwUapg6gFFo6bZXnnQ5YcIVIP
oJrMYrPnHbWe5qjcr2a/9PU8BFHFeLa0GrmB67/pwVv6EHyImqtO2FAVebiYNkoaVAnn0uElPoEC
Rbtxl+VuCpO/y6pgE/KUxnvvq/UoUt6DLCtT4+NWJZ/m8YViaOO0/Y+A+bS7ummux4xPZblucgn2
tpIpFWq5i1bpVGWHd4W35mPWZ8bK8pqCqmCR0FeZGzb+vtnQYACUmyCO36boadKpWCpIt8yrHr0Y
Ri8wTTVpOiGTJiT8jmQ6RFXaP3ZER07pD8lG438Yw7fG19OI3lIFOr8zR3NIOWqopLAg0LmBydqJ
nGq/2xJJnDUoiXss7CTOdACBdEf/q64O+LeWB2SWtSqCJImvbfrr7eUVcmISMUv0Xk6Xmo7YQlX1
kb8+eCsl8teSfBQHkadCwfaU/U98Rb0dBPw6gclGE0dcrvPA1l/7B6V7w8S+CW0xeK9mP3NtLkUN
+LL4WV6/WVzxiG7fM/FNLbQ3bf40II66vezk2CDegSSzq7l0j4IW4sOmpa1fb/ZJ2R4NM2nCx8Lq
nTms9tPS4cfZe+PxuuMHwA2q+x6ncTqHeraUwFPwXf2IEkG8Bc3oc7eAwGUrR5bjBomzxNU0XrtM
Gaf9HVb1EEZmNQCjMThtrPgtQIsHZBMkjVC/GAEhzpoctnm46SsXGgg21Vx5OHYpncEosoWdJZ7i
3kcDu3M6nUqtl8OnhmRi1uswuR3oysDR5Bg1cAKHgLcYuyHP0T0XRMWPrXngrCOIywxdX8dPDEiX
psCK3orD8sdgKJ9gm3f4U4v1U58xd57VvPu5mwV8bIM/DiVQNECtjzVXwpZ3qZMEzu5koZT1CHKx
4UgfBmvGelbtaOYp9ZZlKz2BtRddwoG2CPP7yqofw5Lc5AuUSgQYXy48K9eT+OiY5Oc0HCmOh+TX
hcE4h9r6D1QXhtto9VgXcRE0idUlarloJwIu5RgTdIGdb6jbp3Hhix70Vmxg+YXIkLd95XWqF05N
vczV1xGLReaSVsBH2XLbusPjcUIbFtPxgLEhntxX5betBR57sJSrd83aViBMku0U3DfWYonp1sBu
ct01TKkFG8KAe3ZdyRjVuw0C3bGJByIxXi1MyMieojARKtaW+dcI59p2dZG24jKc69jePmuXbolD
0ehjyAMVryQHaBF8GMit5RGovFSE/NDTJCnC6e3H2JvmJCNTWYI5kIJ+dkIpto/Lse9PJ+LxNial
hkDNncy0legd4qsGVkB+OLUjc6QzYTi9niHP+z/LhanSIDRMxuR5mTAi5woT28mhzmJQ9oyZySRd
SqjIS8e/Fq1CqEYXL9K4Czny+JQJdJl8kltY6HdxDzPL7mTpANwqOa34bQxXOYWqF2GbePLHSV6B
G7Y=
`protect end_protected
