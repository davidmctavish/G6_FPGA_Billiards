`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PGDTTzaJkZyq/Sx6vP8SWiPHxPSvWbMVjmG1+Q+wp2bqoQkf1EP5khzOtWbnSGP5xdMzxulPNEU8
KdGm2w8f7A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E15qksIbH39DJNFmgugZpdiapYKk83QOlmyew32sk3TqZk9JLqKaUierYaSIavwacgtHdsjPHKXv
/J8/pW5NIzZJFUIplGVdc++mr6szt/e3PhJ2w1n9zGKBPzwyBPgi6DOuvv9doiNez+oXAXroE6Pb
0sE6klWWAQLlS9V6BZc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OpoBjOa3Hsioae1ijGqLzQFaDoio5fe5RPWuiNLQeQH9oJI8wiWkmduQYHtKwHxiP7sd8vlm7z7i
O9mm3J8LYFom8Ql1GCqVpb/CMnyoyIlNiotSYfLcgGOmDiZT/9fFAf59cyrJhk09aVeFnxNMvD0k
zKR5GRn+u2hMNV+M58zby3j8ms+ZgMNNCp+G6jWRrGD0zpEklBAKXtNmbaoyz0nBRB2VICYUFdmq
a+sEUymrHfzeyErOo0F8PtJrYDPJoBNt/prCB6cUpvFqhYgHvE928kJMiQnUBM9+sV9cZKavOhsu
pdFTo/7i4WxeH1nf8Nn7MRiXHIMJPRe5nMbUpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BImwwUhQgG8ZtIHPWHApl14MnHbyskgXeHF5DdyvSRkvuwqLfOwIodJ645QrhFbLnN/A9oFjKWwR
k5Ue1rmxq5+6DgkUmX5mWYPKHQ8qV2icmN0b8FN82yqyfMp8Nuw/lDJzAYGFxrD1YiezK33JBN9K
kKEkDpoIcF77GUlKhTw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eU//7gXqNPSzomcEyiVaVIbeicWqyTBbsuhCTn+1ScW6dkJT4INx3r56UgbqrsJhlfTYB/8cJck/
JY0boNqVM3XMIbA0XYAP2n20vd6O1xRbHgNTR7xdYcXnMMebASBbEENMBJu/PITAJPYuqFuGM5c7
vtFijEcUNg+50MnoCYyqzNwLVjD2maNHBQpy9x8if3gdDUA5jMSCQv0/0R6XdIw1cyTiPdwPyWer
+lFZNEHR40au8Uztd91wzAm3dkQnJEl64jhgzQ4noJaSUWMm86775TOmbq6iuehBnH90SFsc+N0d
sOjgxNCNIjxVzb+HneNZ1GP3mqP/bfAai8fAHw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21712)
`protect data_block
hzp9sYOYlFgtHvkOXMVIg+JO4acpW7KELlblknJsKe/xHKdI2zXRDw9m6QBQRKqfkncDAHaM1JTp
Vu+NhsIH942sLcy6ZtKxQlpMxQ5Ai1fWAy9HVJghhpgoPG4IuHhOCy5mJrf0k3k9rk6+mjg01iO5
8Kz7i3BtxlZQLkXi19cpSRW7bMqEfgwxpwfS+kQzhTdTk8Myl8DTn/zIXM1V09Ap7Aqm0mSddC8x
zHFojSRKpKyzLXkNLXtNqeZgYhE63x5VoyeqAf8UBZ8jmVL56Mi35Y2BrxG9McMu1KUMaRhPKyOc
ptQtSr65dXZggN7/yBNDmuRXmWmrxe2j6eOMtRKcqOKC93Fbw/qHyREg/nQZ/uyZVLWZbwDBmmmB
Azao4OasJpW/pma9566avdirtFWTbdfUYzVQ23Yb9G7VJOzffxiEBhWcle/K+PYwyCwsiUGSAEwt
qHSLg2TMYF6wfgdR0X5Um7ncwgjzVD9YR08DyH+aCqZjaW5hsF7HtLi6CONy4Sr+Pi7EIMJN/sHo
9XCja8CqVxKh7CXJS53u0UNdmDWyai0QLOHSo+j3SyX7D713WHoRPL52c30WtfgUi/R7vNH9Za0o
EwX7niKlmmW3JlB2WXtXN9bTBeQBHPYg0pF2+ztbzKSA8jNxH5eCRtePbOpFxmaOxb8Tv8q2VLLy
BcHHAiWpSkN3REaXTIUkPmymdxWejavESmKJtslEghVU5B9O4ObQb3bMSAcDsKfY179Yb8eAloDB
6eBpmh8EiTzh/7JYy37g//1g05BXYBG7H9AB2FPCQy0uIBloXwXsHTy64YE4sx9KE92b6+Itx7za
uNuIx5mLk45vv72VTuEIaplp+HyaBLp+nga8nhHjpoTo0NXnuRqxxL0C5U5e29Y5miNWrJb7Pjof
CRA6p2LC0zTA3jxFtf6y4Ce6+ZkbSuwMQRGhIjPmRCC4aTmuC8aquBp0oVdLEiYNiqDh8JNWXCeN
auJc2Yzb7WzSrjzjREb84nLdTHpA7Ud16c+iCuyxtcOd1DDa6wmoun2KVy9J1JCvK2UWFpax9Akw
zPX2x5MJMa9GlzeWKUjTBbjuCWcV6HpSVXEO7gBDAeNarDUBSpVWlz2qcnBNGcM7pPEiXQwE3FRy
FWFJltvyl3K8r/fHaqelwyikOKnjO0vTRe3iLmhT1LVTz9ceK4BGL1NoIjksVRmEiwh5df9mkEkj
tAadYiDmQOWAxHiM6siLU+uf61q9QAxsxKOQaf7+oUb+aH2k9dEDSOqn3bkvWVc3HBBnFxmp9HL7
Ptebc+55d0FLgPXrkhiVxr45o7kdAi1NkO4kWk/MGBlbzzBnUi0zoU8SXeu9e4Q/DbRyRz1f3di+
QPWHWtLyAatF8q4yAkuTh+IKSjeoCMedhcvnHVWFFwgL4L9vLNAHlwVfk8bDhDADtdIi/dtNYkzP
mck/V75DRoOWK9R1DmItMjynTLWT2f9j52wfjCEZGVuawzsKwv/C81wheN9wn0z39SHctMrQ1t0g
fuDjoGtdz/9zRfNskRwb9nfSE7ZV/vUyiY7r3+k/hLFc/d1ciRHlBuAAss2vP52jF/Q8D3KLYs7m
kJ3CH5ymFYOCfiEPAVCWWKi/Yy7Kc97EfTLz/dPMDDQ/IauPJpOyw0jNlarLWPumf8ArYKdHpbm9
36/Dzu7CTjbZ0Y1gqrAmLed9NV3FyIx85vZJhsKqNXs+Uj5j/X6oF0O3pvTGjmw9NQUy3O1PBeK7
PMPrXmQtnpKxJh6U9+y9NS0/sPMmwweFwWmMt/5M1RWfK09AhzJXjXbq7ZnDiEbDjkIgy0HArt9u
K4788021HZB5Scnw9VE5OpJA5dJlxNz/ve9GMIFyX/RGWgdBvHp/4Uz7MnwJd6/JDaxw22XvElwm
eBbVwwgE91j9GqknV9lJuiTX0sHj06KOBM3gspRgPK32g/EeOEaoUeVRAFbZDuuM8/209Kgikc3Y
pMGr7GfpqlWSwUl57/QJ4cQeStvofEYtZwqtOYJmVKTDEBAoQ7hni8VN/8Hda5RlJzHR5kaZz1kL
vetnGU5vMbcoEA+PbOeJSSmII5V8n5m4QzlibaIBmnk9Qk7S1WV6rtvRAi5I/nLwjhDEldKYwNLY
L0WQG1hSntIbTixGdLY9Xhg1eUEs7O9vUgtPewZluv4GCqKMXbFpA3uZZy1rrBpwmjcEBdk0/AAi
LXwKZeCoBQMBtb2ZVqM6Rbyu/t913HoMobHfPbGQSyh6B/nTV9kHP3z1x+F77RmmeC+OfvC0BV1U
XbgKvJfdvczJw+MgEyrbFvIGoAPhGJA3imhx+famOGm9wcsaRPyIxHsifxU3BgSIkU7XRvY5TNfY
WJQ7xPk+VBzt1Jn6IWwhdhJ6X2rmCtq9306pYdPMHLP0sUO9uJlyVT9yQkoOhjCpfYMfFRj5sNHh
EM/VeVzV5zBDXdrEFFQ9TPQI1W8QEc266Nk7SdxrOiXVR18x18mTZRAvqa9bQm69pP1uYzlyHyO8
fBOCrNOBXkZf2efqIbJLSiAaR5diUUsKYxQ646ETm4xrkfJNRCuUe9fwGRY4nSjZBZpsq0DyKDln
up/r+NMPFyu3tojqceZa3Spq+SzeXbWB3GARVCfqw6WowXdDpl2xzk+b+aT5HE1jM6sxHbw/cNHZ
h7Pf5V0AOV5G2dsRC0SRBjRwg1S7Odig/3SVqy3B2FDsfO5XVZT+45VsNbF7oTIuqyFCfwTcjKxs
8uzNJnvx0I9GTL0jyslW1t4oYQqTfPcFh2qZDliaBe9hUbQWDp2l+OR5WQCs7u0LiiHT9GrCvWWa
X+eXNKTkXqnJh2ph3hpO4C2guh5I7/7nuxeEjIvnG8chy0CBogAyXmCpTp+ny/60wMy+cUb1fMzd
Igc+KVhHhOc5JMUdpNZNKV3nqgW/WE7PH/w76eWo5PyGFKsV72FAjVxQlfXU6lYxPp0jXfah8yzD
f0DE36IYCXE4oJBd5kf/DT4nRw4qOPA9YvGx50tEnnbOSreLPVKylCp8r5M7aV+wHz85uW7gOyzd
iN13c9AYkYPYyQheFeT1a9rB+Xmlfn1kOIvfvF0C1fe8WRqT/kgR8AJTfYx8EBaLxGLdsHT5xP/v
WKP8nN50nnM53n9G+0cgGM+RCSJgT/Cba+ivJfkjS8YATqY1E4sGKpj81Lt0SnXl8TQc4Hs6uTDT
m/xDxtzod/rnjTH1ttgVwoY/BGD1+KqzshGeTmXIPizPYGRVzAigtqvHjWWmoGjMFllEnzEJw92p
FQDV3z+xxt33PRYgtb/j8niz9ropkPREfEiws/cI6mWoFuw8sXLYLnmRNbnXlL3f7KyBL6WMI8gs
a1gZmPT4NY45zOs3xf5fZg91cRKTbxo5roZerNCo4P/A1VVvrjxb1GdqkzUbo0HQ8T1FhJ6SJqYF
W1qXZcIpkWqSA9zQ1dX+EJOojOuFYdabFqK/g1pgWnUIVgQVZRjcf22rfwKOEZaEtj1vg7auy/Y2
g3xdaS6smPQS/QZsb8YGb+elP25FLTaXMOeO7u2AIhE4zigSjGzMmDi3wfmaZf+SbDVrMilQjHTL
J6bGZRdMvVOM4w2WyMkV0I6KLgcg4tazcsit+VmcDi3yjxsa5+9Afxqn7iWEYwu4MYLfutfHUHZL
6ONj4kq8mEamTeyQmdeonEYYG+Uef988hEEGf5l/YZ9nGsbjNtB8fL3ErgBiWLADg8YBUg5c+nIM
PucDVAKszqJM5RvA36YcgL8uwid2E/+v9Ttu/jDYE/RSpX0twqOCavIuEQC+HfVnGjb1QB8DknDR
84Uhandp3KEo3rlr472VIraPA719n8cua1VqNfYRFKHowjhnRL3EMMuaYpFixy5W/nSlESQHJFm7
euTLmTAoKu2N+QbFJ2x0sSZjt+1K4/b93EagYIwt0StbejPV+hnZRAuiKhu1UXTQXHCfgNNaSVH3
qISaxgdeYPmToD4AAC1k5dVd/FhmCqNN8INaFmJWL4VG10ANFdCQA8Ss0Ag/5fGl5xN1KlXWqlKk
Lxbv0gcimqOfQDUn0zuXyqOlEHyNQvmsSlgHdAZiUyxRhzoJ1PCWjV/rFU3oXwEwz52dr68mYwnB
inj4vCVgeyMG4HCqyRqrp9qdAGJegjraItGG7bpno7MSHH5tKXx+Iy/WRjgNRaLeIUzfzx9flAoB
4poAE0yHauF9tEdt8TJ7Rsl3pWMfGxzzo9zR9NLXtOp7yu8KS9TTkvYxrGSO0P3sc5y8TBMww0ZS
UwCY6pmKBNi1eDZaGmy8fvBqgEFIb6CcReVk2yGfTNxZC52wwr/R11mIEzRlMW8DGavsrv+6vIhj
FZFCCVfw6P70REBpOru4FBzsV3w3B6ElSJYMDUEYlaPBeNYSUoGKQL3SERkPVLKHN719hgsgi+JI
gD5W8ffBrUMIjbzRKpsiDB3Z+YryVUZ375XTOIEY6j7I8afgoc6spAxBbd13n+XGE7Y+GlC3Z7Xx
7tQ3Sxl7C4h9H4en3TF131NDS9NuYCao8FZvC27fGlNawOJpIZTBiuXeG4QbnIz5lr6d9YVJVsvl
LJ/ROuWjIfbvgKHu1LH4dnLQ5wd02iBS8fMCm/Auw5zLC8svBiCa36GhrdBzObfLd5DG73gblTk+
D+VIMb5HQHimMxFerchWlMsKsBmWy0TZYl4cjUGspoq/Sm41yKumL/BYU3ynAzJspaIwl6NFqoZX
01SC73Yt/C3szpEEaaATSSjqSGJn+FEWKNDp7SS4cOEMo9dh0vG+mmFwRqYzJdm5AlubTX/1w2lF
rOd1HrX3rLhMFgEp6cwCext8LGINdKfUb+wZqbwOzfLFwdBx/AGy0+ZArZlb1Bd3it6swn7SVrNv
uWNWEXExmBKsrcXxm8Hqxg1PtVOJM2mNVomUNlq+p33M4hmi54VoT+ZPakHR6oM3TbcdMKm50kv+
Ug2U+YZ3xXr/kGekKaO1HbkiJES9IxmW9uLZrG3TMDhKDxrpJzinE4XjWba2bzqosE2y6yDyr8Aj
8ZDyAUywvVjyhMuyMYsUo/6brsv1EXUAGXy1AHPt+qRvVloI29/QB4VDVHaMxw+zN5GO4BMNCKAc
JquTBKH0GFhObXB3L6PCHQIraBkMiJ4MbBzDsJTvBZLKLTpLPmUomjnF+XAuG6ywQpfJw4VzxoY0
71HCwhP74eqRorKL58zOWGkSGgUqYw2tJ2khLrUjezXie41Z3wOWmqTKkx2r8iAj4eQsbsVVhZeH
IsyGasJBPgQKTLZBhg5xQWZGkWMcx7OjMHWX2regj9ieHMLfsQHkISTUM6fvIgxVeZ0QldAx5MtK
PNxUdAP4W+JGFuoD2ElomCHl8NMio32XMoEYJdRdLcxyO+PoBPEAFS76IdICfdczKIBnG95YIWcm
gmWZvLM7n1D0G2qDtzu8ILaADC+oKBg20c3BXMyZqFTvcuQacbWhKkFjxlzCZ/OqYelSxnACXzKi
K9j61ROBb+3QjPuSrGZSqhzKWRLJWf2RYuFP6YY5PviKznBB7pWJetLAMP76ydqC+QrZEwVOWzU+
24d2hY3xeFOFGFdue5zcH1FXwKTWYyQ8jsuV7mXnXOq3ASA50q94wgxytfU0gullLyHNTBfxmb1n
RNcBjA7Glms/S2UYBF0tWFBakKmbffAxr8HU0IehQom4YMA3T+HgA/Oe/DSNj09GW/6E2PoPZWNI
yrTVAgqQaaR6HbuYX2mgpRcFzuFZGUVYvmip32wt5O2eZxW4IWxVeHL5lTWl0rb47BTB0Sn8geFS
05gpSF9EGxa4AtrKM6r+V3SamNrlYvOrvCIAswMism3NNtkfnY6w7wC/m/fjrJ38542jm0BXW+pq
BZb0yXFJa+MqbXoWQpGivCSs6k5RNm1NkZrzS9O81+ePXKHXVmdLswLTP7zZVhvnwC+MeaZOJZEI
s21gCrVAZcMcL+vZwBQeC82QjBtYtIKgY3pfbw/TlX4uMErw0/3gdR6KRldlae5+doZECE4Pb7LQ
u17JxiZF+cVXSzSvxe4dHzDBdy5ySZkKH/xwR2DtVBnrmECy5zAEJX1c9MzA7z1H2UeF4sDezZDK
ZauCWVDpo/R0APdWW8C9uL6kTX11aZYbpraIFDYFRPeWKs+ddERkWkQWzJRXjGMcB8ylA9O3osp6
QOZlA0FR/5IaZ2vngEI1/Q1ZaxbtBWidB5/DL/73ta9TzDgl5eHgeMUi6mTrFkSBpWHuY7Y02SsV
62y0kQNItP8JIUK+v/RoAVGa1KHy2MV5JUEHMASvT1e+V/TFSRXTKvmu8fW352l2LPfcSo5VO3Ey
CmzuROUpzl+BxU3MUTG1Jtb4bkrsXozgkrigVFtr6acUmVPmCnf9hVckEcv1QRnMD6shep2ndLcj
LWtofZwROS4Li/sX9TjS4cZg2k6EuIeuinTIKBpNzQm/q5zW/yA4KfTtQEH+RGYjYZtTakgWWxPQ
NWdgwVXOvUDe91GuLmkoVDX70eK/Jx5JqtmjydSteZSrOtUUrXygDLhLCSuLjM+beAUMmmu1cGmJ
GRI/Mi9kCs0rTx4RMLNmfuzRGibxKzfj0FUIlBAGBLdIlrirprWdnttU6UBhBscCrRVwhse2kKl1
wfh+N4VBdhx0R1oGj44jGo9xXpWlw6eyxmJl3QzSjDMFDngmvG+ZkX7Cq2CJW9QIJ2qwpSvAdJYC
MFmOpaM8f4uJLUkbDpwSWrSMCBmaOkbEVpF8/QCdtMRbxJvg2S1nyYGpTQNHLLa4osvRZZ2+bc5r
rwf1EsR86C+a82YHY0ImI3OwIa+547KKTU0T1g0DKncB3rgRPhEM6D+ITtgDNwFOeDL9qWe/R19r
f69lBviBlbqJKqYwfwgb3ohBRZFSpEvZCc7yi7GLdNvbMuwEHXgr5r/4rxONrR8eer3Rdeu/Zri+
VLMXzaHoYPyKWBw6YEC/ie+zbmO8fNv57SiCBi1f1pjmkOw64Wh0VRc5dY30wzdLSH9GRtXrYdHs
Xr5mysiuY5ApLfjc0z4HYbvXZPAihXGYSJ8FcwZI0+4ffroE5LhpDCrsZfahLBP4UKxJbYZSE3BI
/P+DqO1wb5YIGzZRhqqVeBSLhCI3Vom6ZCUSAhmOjAGN+2qz6tiZFpGG7TtBfB6wVZzNnDejhq7e
RqyIw2mXZb8DxIDc+RyAVTkpZPSbb87MMFQaFIsdtGtXk2fUOsoJkpuNk1CkL2PSeKo0VJcZGu1S
VR+ABoynKEvtxiUgCQKFn72We3EYXOu4IeS2uLzfT4Lwq/nqrozHmgel3Xetf9l5V5gPcFg6/pcY
ZYRMRCKeXFWUCsV9M9sYdGfuMOuRWQ1L7+FoEP4C6zTyWVa5YtfHTLAfwyJmiL/5wp2Argj+dTQG
RMG+lnN6eQC0sv5GcBXBNjfIKPZOZ88e2bqFm/q+44denrmRt87zz38DM5lUkqjhszV/MrsPurOc
/6WNMk0MUcgD8vp0L1oZkXPoXU9MqTfJwLl5ZqC/VVqxBbuHCEtld8mI/SxmRfYxfS/UVlRxiVwI
R+I8Ccu7PshZuhlpA2P/4XM/ao9dre12y7qN1xZ5EGxfz5dNZLVSksjqbh9Kr04ihBw7ciM6DDkM
1NdCqTRgM8hrIR2P1vMHdgXJZ31+kCivia5Jp7xclMMloIuzm3xmNmbRAU2bqErPeyH3AlXqR2lx
uYq/Qho7iMS0P5qlFwvcp7xFVMwmPsMO6/UJ5OMqPx3+3qHrlN0oOJq/PTEStsP6TNMIB1rRs5gH
DHzSa4FIgnWYRO127lxxKJfinyrLOHFj2DFwIMYp3amK+NvgmF3JTHkmjIADcCWkJk1cMg23Ni3P
wAre84aZ9mAGUSa4Ba8tTofKD9NrSO62MecoLpITf/d43NAiDt486Rx8LurI5m4raXZQiOSyqYmP
sAKxgRJ+l88WYVqqlNTaCxDKy8rxwK4KFfl9f4cAAUbr28Pip7GAJheMI+wRzFY+4QhL2Ye1fCCI
znfB5DCDhwGV59SvwU9G4k4oHwd5Ik2k1kaT5FGUV5ElC7SLV+Fjtwy0aGG5BP4pBSB5eJP3z4LN
e4kCZ84zNVgdb0p+oMVqrXWAdKy3ie+hP29YeoYsaApcZHl2U+9/qM89lMhnGqVQq5hBh2nBIOKd
5Wfu7W0BYtuPvi4dFjTmwcSSZcFqwGPTR5Fa59op5AiUP5x0+Zn72jcNAoH0UBfJyRJXx+qEIfgl
N44ROJca6zTAKjoFQP50vltUnhZSK2XoaTZz0N4uAMlfIGlW9hxMAfYt1ov+J57nza4YTIBWMfGY
n670pJUFGQAUhPqcPQXhfRkqazDQDvw6ouwQj5Hr7LOrwdEeuqSGGxgfPLWMmPlkOnszRHa/gy7C
ano4tE/ksBQF4LQnzddnW9MBXpz++EVI2K3R0IpMt2yRQ+yG/lngOe0EaWsdfS3KtZ8aPuJCmKbg
TpQrNg/6JB5bxIkye/GQIyqXou/C61eqRKcJTSY0js9I7P715WGfAugHzjpaD35eRbK4csMlCLKA
2TKEsZTCqZrGjQvwfypLPweLhcrroXLKBsMxYN0plew2Dq6W/L/tkqUFas6GmglJwnYE8xloFwjY
iW9XYWQHzG/lfIpAWWGmuz0OqVe7eiyYg1rZfUKins1uY6VuB2Juc+XXO0SX3Kt1tGGGRncRVq0k
+2pOtVlpSVJ8EEKie1CZDEdKHK8tasmKe4SjRmrFoPskdErREpsBnQ73m84z2b9Vfd6avAHGgGd5
LZjvoKJpbwbIf5aMTX8dSdHhd2QipUEXM9giEulmDn/AXUfxNidOXGBnZDfJKiVVxOaKG9kRC5BU
b0+12fgDQfteN8Rxocw0bJ2ZdSSVEIg3cHkbsfVnTyRb/QpMFglco+RfKVOsxrb3bKy9uVKMhrQT
XUJT15PvduiIT24Pc2N2wkGoUebqRMp3day3Wp5/83w2iUiEAGmXJ47OOgZKIuIyuM3g8Ucufe+l
/Dq+D8VlhG7P8uGKaqNnisrS+cxfz3x6BNeH9UY51c3VgkKQ076DKYIKFnDTiM6JdBYVvvQ6iZgc
8OEQXD3paRaFBU4TaOoQEk1axpidAVW4HhZr+KCo6d/FkziPMJStQN8/o4Hu7kMpDqtnjXhegyKC
/Fs2HAlnBFiow8HO3sF1VasF91lTseKteEX3xW2d0PWEqHuV9a4rUD6vPFB0dyVU6VdROD9qJx8K
GdXG0qZ5v5+/qpBT79wcawesVx/1Dhbkh4TO+krtC6fyCSSPJ2lLEJwfPFRqt+3K2KtMj+Cmg47W
xYHN1Cc7/5DfWj702e9MLfNNQAPYbydymTCx5Q27yierGFuxbDPNXoGefPduay205Jcj/Ed8FdKf
hzxu1SnzBQw0uPAoNSAYWtRwZz+Ys6YBkcW4ns5gd5tC1GEatz42onLxEVQRSn2OH7+WhTeZCNhz
P/hqxWp1riM2ZPWE9rVFZiti3010nvSque/UIQzCxxkwb6XlFqOm1E3QfxONijFwqNfrHY5y9muh
YRVxzYJBGHu27qCbbsODi+OqNQ2R2TLAx7SIChK9e2J5wYphn/KcRNfDhELxYaEoAtZVTVnPBrA3
9qGvmbua4bjexzrMs4nXSpDMI8wIWOQYmKFtEGx8Vjv4Jc0gvl+QWFBM1fB9LLbYiRm8cZ7vpRXc
XgLwBwJ6hN6oPG8aQeZ+oaySEwk+SF8uZ+MkA/4NuJh/QjqRR4wH9SKYaat0X0MTI1liSLeutJZR
PRhhhmzaVu7gpr72V5U1K7xLj0ou0whx7Vx3NjXod8M4LEblJIMdgjtiNaXkvft03hsSzm7f2umq
irW8MqedL8cOxexQKptk2skTKItURu2uMpQ7h2tOxkntgyBczupAUFixSLRCBs5KLkCCPQKAuBEF
KQ8F9Y4P5T7yZdKga4id+tbHooUr6k232d/VZ/x7Wh79rJYslACMkxLNG2eu5uQVmU81BI+oHQMk
tIC2JRJniD+k1Lv0P6DJzFUbDOa29QXKywQmJ4DFmz1PA/lB26fZ0QZnSAKc0jSzM+dwpB8C865p
bKOxbzWuj/1SXRAELLvMl/+gAQ7vjz0Te+tPck4Pw5V7p7L8On0fgQ3GY9b2Bh2J4LnoZ62qjppl
vmysjV1QDBl7FZ68b2ihnMHdYUYz26yElSs/JTzmYqlGVHlx0VZTm98sk/LtYLsY+RmzjBYS4ORW
IurIXsO4uBQSs1pE1Gs4PNyOcsdVzhGM4Mnmby0ZgZx60SW5zs6JTb/heG/2dep4NiegwC8xFY3C
uESaE7oix0LVGLzJCtek/RGRZTuLuxPXb8JdthZBmZjyFQ/UBEvkwXffVIRl37BTGL1C53xajZOR
l4PAWx5zHJJ1O/lFogBOouRbGtR9ZqCEAtCJCEDNDDoA1eqMt6DFCn6O5VU1NqMJ+5wULVl4SYCE
wHDFFzGvEIjD6JRD8k0Q3YwVpP7vJYRlRvSQDiaeXX5Uytt4cu6rP6ajBhBHi0lVqaFkdwhwF6Qy
Pc1ahd4AteN2LRw1RNz81Ppz7K4FW33XoquvzIoTXQTYinuiOBBa+uBtCAxpQFP2hHGC1SYVEDM6
5i84jIReiZAgI11pnCIOghWFyH8IKy4Cwr/HNqRM7rn4p82+Es/p1CVIsEWVN1/ljZDFQ6IIdcNO
OE6XNrUW4fUWCJiXT1/vn3r96PZ2+Ox3eAsB5imll5bJnPGmnoC89GuswdCtnjSCZk8Gd20QXCQc
/S8hUb7nGFYSgEoVm/PCB+6w4q7oxwoJdkknN31YVS4If47FYiwSrdAfjoo4JPrwLmTWONM1Uwhj
Jr2dC1DwTbta2zcOJhlB7DW1fmYDCjmtu2f1AqanHoYkuABowaqmrh6Ro4MlhxzVyuWwJzfueBuv
LWTli2yjz4Ws2c99Xtzf8zbc8CloOYw9DiaaM8n9GmEwgjO4c/aPz77MtZpFqR6ZTRucyrgyP9Sw
ljtoeWraLj6jW2yn6R8+nTzMjLkqQ16JhREuY9a8uDqX0yeAsToevkYMtAhDbS/BJs9mhFk46f83
lPEFaQQysMw778te72wgh9zJ0aH0a4P1CSMLGKq6OpymdshvdLo+Qn4bNtNwj6kYz9C3autIcnzQ
dFqiQu4bPp704vzMgJx37LRNnSzR1olBj9QjoL5KQn6vdf9W6bHtMp4K21eEfWMvXRPoZFPv3hw3
9fw1fIqLfCuDIcfzMs+1z/6yo3Ks4IlsVLq2FShM028ALXEl/3U9QK3K3lUDlZiSp1mLbuX1C8wb
qb8/hpH90woMB0OZzyDgLcb/537wHtHSlqu+P3L2RppNCJV8wW+HP0EQSNF8l99kM1NMbSPHDxWL
Mz5PXANgJbeOJvKWyyRrBCVyr0KSlLkOs4cf13fXMrW/hjArwwDFoqQPHDCm262YGazNimGG+K5o
KxM1xlbVuKk6HLSAO1GRksFHgIvMRrk/RutqCpk51DN8/29D958F6kvBRzRipp+kkO54D3BVH8C9
4TuiDVXOTI/s4WFZSyXXYykofNkBtovy4PAHgOMBP35dboX4Y/whV0Dt3TTwYr72k9uAyT/P9hv5
DVChnrunsk+HQFVd+4B4JIFOsryoza/beJUZwFI5Ybp91qz/V22Il+QUZRRenM/PWbmBNbMx1TUr
owwU299GE/VedqFbzFWso17jNz01QlPdF0UoWRBiq2mszfO8XkOyiPoi+pKTBp+gKPmUMkEG5L97
xhiwSzoinVCLXVsN9QZeTloldhdgoc0cEwtU6OUvWU5N/I4MyXpU9IKLTePGDxAmv9u7YFD0Bb2N
MJElPKNi3WIEzRq2xCNMrFpcLdhisNlDBGZWf5WMTH/XUJQywNVz9Nvzje1XtTOHtvQM1tqiTR0O
GLHy5zc93g8TlS2ayGeZFSTKnZSmXxnundauSn6ocuy+dJQQs9iHHmvZVDLVcvHZhgvQlJ9cuVW7
n7J7N8Az0Jhnz2xvAHRNMzpF+MvC4CwqR9H3eNyyNBPACEV8v2LIm3kNcse4QNha2h7NRPpZUcqE
RtiC4UNjLIpyKzdaUPuFOUgytKl+Dw4MYUYwXprzygIpmE9ZzfDtINUyJqxGY0eO9mgW8Y3KDS5T
sL549tfrD9IrhNoMwy3IHkKe5vPoq6S2UUk4mnW0gcHwAA07poXhOP/fMUGpeK12Vd7FokDTCgLG
wFGYWk2tXvNeZ2xArLuH+kKG1WZDTY89/j45DhXSNUQI3suPK6OwQQE3fYalfB+if80HITSIGeTx
Wkh7VCu8gLFXYoZcfSbWfYLog/ExwIRWl+/Q31SyeK/PqCrssYQ9BRkO350JoGM4JV+/emSsN7Zi
5OludeYJDisqwuCX/KzX4DKXT0iVwBbwT0S18eATHO0dns6L0oskAVpyEQbwxEzRjU5sCTpA7vyq
mytjGT6pulleSr9h2vi7fsBHXe0HKBg4w1EsTgju0lIJrkqTKl4tFXj51C+vUXdgfbyX+uQXdur+
JkjbocU6VAJppr3SmrJ7qnjsbgAyrncq4PEuSgSufCCGxCibyL/yekSjHiOMBSKWUJS9CFgCpOxH
d1K0KCntgh1l7H6yoBUHV3V6demq1BrnxBxagGsrrapy+JkF3GuuUnIwMLR3c4laN5cM4hL2mO1u
oxdq6+Kjudn4HAbpWkw/gRfdg4RBIE1RXmDBFzoV6u3n+yk80hjQ5INsj+etmMxL0fjK1dAp8y77
2KSNCGp7gLoH1oi+LS2csyzlYTs11uk4Uq4+t7px7JTaMAhNU9umz+8d8nho7g5exwZ8B+Dijkqr
VHHI8zmXg7ix39re85kOQYzPYKoJZAVPSK+kDrSbe3p92mRxz3TpD7xA4SjZG59jRNTftwv7H5+X
wlL2uIEjE/T8pldJ4W3nVNrMRdr3RYz2bDhnUO0cGSeFCQcAgSf7xGsjLkYox0ns8dD5JGUVVi58
JGwzazB0YFUtBey/Ph+lxBjJliyBOFagYJTh8qAjlfwE+Z5Ntrk5pZ0jaWuNUz4EZrSjJuR5xRPM
X+Ia442LQz8YdboCmK9m6BGCIGxHk3DCgHw75EwsrxAHlDZ1M8FewWeQlw9uzesmAAW7XVCzN0A1
0KONjDFEEhmxgLTMYtnINtaXe63lLU1DIdICD/H7xLBLOz9M683ST0VPEt9Hq6VQjLIIoBsqZMgE
5/p5PomeonCt9JtQd0UJbizEt6lL4XC3azUKrWDdC7CHj9xpwFezWPHFjZJ0QDKiAOBrbJPQKDVL
sQeC9pbIQQvL5T+vFsgYO5/geCHH6FOLLmBqhO80gcq/bb8A008LUEOdK6Mc2fIlvU5rUC+TsvBu
I4ApJtuU8iZb70uBBH1zy+t43xZclLapY76gn0oxrYW/zGBNcdoz5RK+usd1tqNyxnEbkCUfI48T
c+XXuEVPb+tEiO+dwrQ2hDYCAm2oMMe/l8aMtTZslutEGVwFWHtwAdIZ5SX1pTI1QNimSxjGaa8i
pJt/crYyX5x1HIYARyC3Tiv2gzmPXaAXlRpLfiQeYMYRI46t23nMFJNhN86THoe4vmAXxZkpnUo2
FkonzZK+g+9Wdj7GN095tPaxf+RdNIFxSA/PcQfwdRJavZ6D8ASU/Gnvexw0p9lHQAHbHF5RrdEq
NRsEUazKXSW343Hoo0A52Q7hMFneMY1qBvslWKatEjTwDiAZlQmOHZBzzqHcThadKN075/GMZCjb
19b6B9i5T1+iG410IX6fShMFT8aM4tiaYT8OtsJyrNRMzrtN1SjVDCH3wqza7Q4eR5kVVtI2VByY
qHNXwQkK6UI61PEMNMgia1omYLxaZH/dTVE9RE9PYP/by0SHw+qEtO23Lffl3u50e9NVUZwwEb4P
91e8wnx9eJEejqN6ERwj3VbZ5eyo3F94y5YSoUYIqG5JhAg1161G8xU2OiswkLHSBAuVKokt1JNK
xaPn/EqmCf8CooNjkevkypftEK/sRK6+ZvNB64+8bMSfje8awe/HwM4A5P0KO0E/ewsScXsSchJU
Mya4MytuB8m0hreXuqlCbtXqtgmNpz9MicAC6477A4QGWrNz1Vw+4fRGAsNAxEgxxFWRsS2fwopg
1cCue7jNwYGLTXaOIuXQVEFzvm/jLEK+7vZY+QKIhz1vonCDF0RSIbRiWhYrvwYkLKpelo3P/IGp
xTS0wtlCuUjcuZEJwdpb/XK1NfiWRciEYEPT2HysI6rn5rk9iKiGNjmzPBGAgR4kkg7jJ+kASkHv
KT7DSAft5KLieBoYr95ywMZg2Q8WJa0T2llo0426SZea29Ga7BhqAfcc1JatmC40RKjTumZze4uk
zAIDOxEgdGfyCocCpV71+sm6kDbemRRcAfyuXaRdEuus3O/XqmMXDn3xvrjc0zbRm2v4AI/hiI0n
PeyR0T4YnF3gHuDKcwyv+UjBacJxiC8Kqm/M4lQi+DXdWH6N5RLmSRGBSFceoFPm1dfSvGq8cV2y
Q1GbFpHKmTnS4T/6NPZQCMOY1C4fPM/IQGPljy3D1DsONRDOFTzWCKVQ//pUSANcMy9sadbrVlqx
xIm36IF7xeQDv26NcBUbScgYkC6Ymi21MmZYpVFg8FOorRZLUefBGHGsbdWxa2wyc1Pft3vWJ/Kz
HVICe8HTwrXgCIv2zHAFFFhdlO33tIAZYmzen1bo7h/bC3TdsQDFMpBMtDWgMTckBmEgaGlvDfEL
OvUBRevkfVdC/AHr7YrPWrBlGWEKkDVZTZ/Os9UevJrIH7Tozck59EQJQwQWX7AHOgouQl4fIjys
s0/mMdx1lzS2pswohf+lFqCkh9fwxKdP6H6sEeFZx59XYnbbwx5A96OWzAiR5y+S+zK9fx11fNMr
XzKSTNfx6ZCjrBKych9/AMEonvIVu91tdQxvwC/TBMKrYjgHjQMLHPJ915ywt0dQqCLpDtHhQe1f
vpWy9iaVbNXISYAe4nmFdsK/9ajq1x0G8lkN/VnEtw3Yo+2IfF99eHoEzFj1Axp8Y/1+pZleKOac
TzvsutpTvOjVlW88wzXuKyY/+T4ll9sj61kMKkS4KxQBubAuikjftNwnyXDGK/9wyXgU74KoGTkF
OWu4V8lz+CEaUOjHHs4Sfc/XCcKrXJJDfd4nQsjx7u8DfCEZkKQr/S95OJEaoz+9gtOXacIpONyg
Scvv9AQd6IRtNmIHNJO8DudY85wB0ZUl5OKaeoT/yLI3F/l2tEr2PLP0zL1Uc65NQ6AGO7Aj/uxv
lf/8QSMtaNyvl8AvJncPMBS8qaz7g8ULCqlP9/SSwdSZ1MslI9WKZ1SddstMIhV9k4HOe3VSiN3r
vR4XrcXBYmEmrQg0UpIUN0NNE77Yb9LYVoMztKxQULbslB/FLNCAHm/Y1sqLqtegL701vjEqQr1l
Og7YxhMDdnvlngjIXNeO9mmA4KYo1zNmwUbJPN52Gno1yW0ZqKii9Dj9Z132FlH7Upb0zeMjq7aR
BKl9SNEhvep2CHAvG92HPszGLo6ude+bAJMOq8wsuXfay6awWWZiTibcqdVoRXdAlxwEBfkq6abT
tcR73vBi29/QDPapR1JochVg4CkgKR6uHEHgGvKqsui7PTrfMAgFlNUaY9qiWbq2TcmFS82pFtaf
r8jI9OriVu/tP5OGLQD8Cc+O139k66p9zw04VtqlINpAyF2pLs7YYoML9hxwAkD6qjBc3il/DNOd
yNZrCfGAg6ic/8td8uw/Cc8Fql+7AvL5EIwnGUX0TQeByY77k09eW9M7oaOiVGUyDkaAMM/PnPT4
gqx/feGM8lPhQ43bZiQt2y6yjVowGqMqqGlu5l8r0zYhqdnCQmnCxiBsIHgIVMFdZDq29P1L8qzN
EcW2D+mkszIHIUunk0a67gE+zitSS0HO2udcFr38nO91bglCg2ooYYdcz8dVJa5x1EiwS6j975GL
lFKqOLzsmTwTHIVsY73TQeh/HygBrsfBuE+bh8uE72bw24abtG198i5A1QxV3RrvkrlW5S3MdtV+
M712MnXkBXcc/m/SC9WvxAPgeqUgQUK4qT+p23MzrSaWNkBp2LFVsOV6pOuxdOvcB08QzYjY/ucC
j/I4R6ASZospnkRSoY+jdzKzMhVDQWBlacIcDMVv8yQaNEytEG8IwNdC5bvPqD6Cjz2vrEI6kAQV
VRFFfcjwS8dxcHMry4rG/OOhAzL3drMT+BqOFegzmVWnEuu7KyfpB5HvGj7ROIM+RX178NVk7uw/
n8gb5zXL04GyZgylZL2nhDfkGAmdDxoR9UWGSu8iI6KHka2QiY12WyVofddWQ7h9uJgP7Inmah/o
V/UnkX8FlqK3Z76bGJ/QnnAlrZ87G55JhXtE4rrzkyiOACVoHgGABCD0xUtpxMe3K7znwDMKVZqW
djLfIYwd6a9rngh4g2q14mimaz7yIqMOMJJkIFFwfmvy5Zx/BXF0YS3WQkvVxqMYyjQfcipcZ8R5
ayKO8oaT2mu6JBFep00cPMyjUIGaicisZf3BDboKWX06UDbrzkIA+0DDJ8sr9fNWvFe3ZevQv0J/
OPigvf/kaV8B/Ts1pM9GViPS5jTRbtFLAgMxuRy+uRdrtIQcnMhHogXL5IfqfVq5duVAXDWgAkiW
ghDlbnmWDwujbgko24soYBPElJKUsHk2dN6vBDWyjS471m+91CXT3E+BBvXBCh0AiYcoP41AHJiA
O2QSFYUaEPSmngLVe8xYtzIeHQbDfSJ8YIJO3n2g/vK94/AeU7XIWRRF6RX8vMkB3CfB/8yQ3t4m
7I1MIQ2P7Dk19M0NNBujKpm9CcmajXUfqX+62EoX3C6SQE76cFvr/jzpnWUES7phl/QxW1ACMee7
1aailjvRPoEAsfkAjgSQ7d3u7jigPb+cve8cEICoGMKZaCJ3PJ1DH2eP+us3vNPf/PhMSU7Z705Q
O3fgouIbDjO7OeMrM4BEzjc0zczJVZQzAF7xeQkqB4ctVIqi3e5ULpHBXyWwQB/qA8UQKgiKxfn9
5kI6/LsH9n51mvBw2xNfS0dATjjmaQNKH9ZB4MxvbNCv5ZmdwXRqSch/9KUvWW7MGZaoPDLhOQLy
m5fedgfHsii78dyNFZwKvYA9UXBOaPQvwurbPKEaF6rrCc6ME1gyWrIjlO41NEIfQ7CR9ojWc1ry
O3zwZbVzEbGMy72rdDU0Oi/JK51nwxroxraDXfUkWfCuWGLiU0Dn33z1+kdCiB9IR9XUaBf/7eXf
xqq41BikPy1BIgwQvxYAteA+A2eBqQvu0YoClW77WkKvQ/RtHluHrPJ7b847ctju7IL8KoNlDhrD
Y9/Adr9QLJEZXgxYLEcSKVh1e6vEgym+G96MuLJAZDsnolPgeobRqvaWriafFXYAU8vPi91gmlrO
eoiK3z/rI+Nz6n2XbjSgBuYxbe4yTidyoDMVaCAb44b4dVJ4bSeUw2UEdCEJVwPfnXnu5FebUL/X
8w2IvpTtVYqhEbQdGGMirRHGvJlwGuTeyfOOWVjVVTJSfg3VdbGMGMO0oCaYdAHxayldJskTbKLm
mLxLqt4oStno6CXUVgeHi4moC0yxlZYVh6FmcObJCIE1UACbc2VAwmguFQxeBhSxeYv2veK0Znzw
J5KPzvK2SqT8Qa4eqg02fEMZioI7xkyufXooZn2B4oAwvm8ZppDbeZ+V1n539jgY0062QEsBDI9M
JlmjghmJot3g8Uj/wL/dKUXfUBMEgOIIfoPtxqM08BDJCzTrupSNXeZHJRUAS2WkI4S1F4rtznvk
2SjpiWExKbhmxNoHWoQFecLjAltM87knCOEFdc/Bzhwn++2BtZyO/UAZcjl2jm+4YyzVcGuDVp74
/y0DfBrrRjZHu45m+fi09w2LeS6mS7wCu1E52gdy5i4jF0R62S3dg+CwJAL5hwwr+CzpoiUhOlU+
DbvYzc/a0fRtdqYDKUmgq6K2Vl5xFUbdEOekzFxa2OiEGSkpVhQb0PQshrzXXFT17sv8b1ZEqi/3
cVtlxJflYflKngy4RNAuTLfv/lWi9DX6nU+M4X/RT8ogNybXPiUyic63IQ5FGavByPO7aEiFCRH4
BefymatS9rIe5sGTprBe8yPLHt5IOO8TSQ+fts3+sRWfe8vcsxPbJZsN663DWNIJjRiOSL/HedAA
/tBl2DCez2j9BxXa30lKIgmc+k0OXYmQZWyNIpvd5PPj/hJfG31nkSC1J9eTPN4H2yVasheTRqoG
MQX9DQbJfuOpYHsdbOIigs4KNWyNbM4yGy9EL0yuHkg/bnOzkF2JBe/9MWhxgwnzcEMsRMN0PPbA
88lTSlmr3GCcsP7uZmG7EsCY8gGJMZ9+a1lbAqjvkIDvUroZi9HlruZRUhuFov7cxozzD/W0xWNw
q+7ZJB8HMUBbohAwhJ0IM5o9z/llcnFpjHIBZIwcYoE30HxSEb8S49xipYV5W3s/RQYAuz+Gk1nx
GsjnhdeuHYD0N3+geE7pz5hWRD1Eujgbf4bsgsc7+bq3PfqjYpzyrgzGxhTXGInW5GK1YG5pS34g
djUCthtEICt87bKmC+TRNcbeCOANQAdqjMLvurNKy++mIrK9P2kdGE83hHZLscRtiaPy3Jkm0Xid
lfq1Q2FomDzDiybc75YVwOasWLZg2GvgNst6Rzwc7fW280LS0abxPM+daX20EyPOzwiCTb+efU8o
65+J8Zb9BPKhJlblFUWzMaFvW351arTeu4P/qC6yVLgmwWfjqMMRSdjoS9UZyZ29tXzRe7ZaPc2n
WmdICxy96idRojcsgjfhqljBeP+/TYMq3R15L4cl3nJKBKQlmn78jXK6WXsOmjNNu0KX1sYa798W
m0iTT140bi6Ep+uqPvPPXaSyh9KATxs4H0dOWCR8UeKIj/lHbCFYEPPB21q7ooQH1AMLlEvdn21h
nRpyM9gYnV5Ej4iD0CNCuxHJKrOIsULqWhNNG2y6p+RDrpEfun27+xqYOnQcha6oli0p9cZPgeDM
LdGiGnqjh9BYVfUkvToXVHu4Yn2HjuKBzncgHeBId2nJRM0CSWpBY+SRTb0Zhl7VJ0EpqXZFC3z/
PEif7vOm/8a4/VfMtWjNoG7hQxtjHXB3qYuBwC+7BwZ5S2e06bvxiqmHm//3BVD1QC8JCoVK41wv
LNQD0Tv1zCsgV/o70h/TZSF9wtbTeQqA8FmoA/KFaIk26Pe9lmtQPzKBhE4CGbk5Pz8qVRSJ95iy
IbhdrdfplyqqHXcXgS0WQzMUK/A3oib+ubZBQAk1xjcBGdCVNvtvz8G39Dw7EjiuTI1XS9cHCLgv
JVZhRQttx70HnWC5Ge2nREIV06wwh4aqBSfWD4v01ZBjLE7V2WHgz8ZEIfNJQnAmmG0L0iSYZ/ji
QdkwEpfmOPmPhpKJjGypH+rcxYk2CjMfjvte660p1a1RyH9eo+I29vy+oU3IkCHN3SBLN/uYNg2H
rT+fh3oPWRVEAsUIYLNafqg8kM77SjpouSe3Y+6LBOxC4s5NEHukfSWxPMOyqbTooP5x3IrwzRva
iPwtKS3ORx8tmucLRYazfa/uRe+0XsrisA3/Bl1Q8rEoADuB3GhxVAqVOzebX/DmCyiD8r1i5XXc
zhLesix6Lao/CcePqPVgtS/6iB1kNeWthgn6fEL4BVpqsXippe2iN34iWiCinpIzzR71WOn8kZRX
RlLw0Oac/sFpg03CaTOXg80Mwh72ANfCTSGiibO996J3i1gpe/VFMsS0/eSbhj7ZQXYTiyqEYBsv
MrbogJqBky2+esSHDFUJzrEQYLWuSkamX4pHaMFjDG2s7t1nwq07ecCvvk1HJASn5jj03Rf444Ba
UH7OoDHvGm9G+bC6MNPuZgZjLyGoqwWrtu6FnVeNPBsDdPjS+cIjKxKl8yFzSF2TjdjDobQUNITH
DlDzXV8sp78r5+kFPSbI2YZQCjrRGgGRujvVMVWGZA55+gBiAZDO33wBBVg0HH7EzCUNBun01z4L
Uw0fE4/iFaF7fjpCzsyRpEyaV3TGkT5r/YLsh1ev6n3ryfMZaaI25k4K6uFKWq2YMsox/vWn68Zu
rfdas2hO5MTKhRWczvKAQCR/MrXBRVzyIz1HWrLWOTT+cz1pBREn3Lmft1JVZdo410YaGiLOnXO1
y91Rq5CxmJNBfaCMpvLgRx6XHw5zSh40FukC6TypAQsag3cM5WQiy2WmxW682Zx90EUuyUeukqzF
t4TJlxNgWNVBXwkueddgH8srQiuufk7pKSAbiLDsDH7ltLRB0FUXlVcdaglCmTaD7ehtOKjMNN7a
tlNKpBickMrQCVUJxTUc/nM85uJFKyl7+9jghKkTfIDJyqpX71e1ur8GW5rdx294zUfejz54Zseo
uxpBTPfchZ5sFEgs63sc3WpqZt0wfdctL/oayx4Om99iRyyqY2Sjxec93CeCFaPyPTcDBK4A7lSa
grq2ZIaBaTvDMC20IuwzE8Y16Pi0hsRfTKVESogVHkderSyUuUYgMVb3UAdq2Z1fwolNWKmnNlKn
YAYAajsM+qDzgdoilrs/s6pe/ikZF5Knj8Z/Cuyyv9kMvZB4uvIgf9nCl3q8JO6mQL9sZejtPndk
7cKhlrDRSIiPyMRSbwl7AWWXTPOsiA0vtmcpOHQq4vkWZL4FL23wBEcIiK8B8pe2P6G4+3bSP1hF
0K7Vnp2GO2/qZgtavPgKd9T4Y9kj593RYFfKQOtP7cxdF+2kg3bnWuDT1pmYtRBNHmMdAVr+wvw9
r+DLPsHWAEB1DO2+9lTJiYRPYv977yUA2x/d5MbUDCggih1COD/MABf13eBP1PTxF+JxgJLtSsj0
EoK6cjKdxpIPf7FwFJj7MtG3bX8+i5mh7F70ljMUHBzxEimSWX5xgswWbondHBKat+5BJQ22xu6B
zlNE6rLT55j3XtWXj90SEQYUhSRbcetq3sngMX2dwAWtMJ/hrCovhsTOoApHRUKhawnJ0P8e9Vxy
RcRlcYGEpG0Y0u6M3VmUosiqk9OOszl9Eglx+KPoKwbtWCdW7LYPM1kiWDpUkAwqJkxD+P+m3KSA
KWVW6hHf5iuQgHW9CPVz/S+nhencvM0Ica2cc2WlTCYI1/vmeQfSmJ3zJF85hBMZV+dlX/kWEjhd
iBDOJvswSz6pMTdTJoHHsvHUqjgLzGiRXn8O+0NLWJdnRyE+Es6wv6WelMNXa8dD2bgLa7YNe27R
9Dz8MZjehNlMCY7aAaZap8CCgwsK8IO7Z2gl7u/G1VE7Cv/21JKE99mFwZETuxomMdY1Kb+h7qdh
PDkPFNlBInqOPRYhmRqBejvhOnNHuAfr1hn6+1yHM9Jf1BuRvoKT45dbX1dZIA3vFY17cksI8SVv
I+SnhTApRCY03RhBpHO6z5lGpvP5mgZd3EggCVpx1g72xmnbMNT4VaCe4ZH8gr+yrdSx20Qm+Jku
9YvQk2yJvcRCSMUXkwd67qSE/duYaPdD0Du8duj4pFYOtJWTyGEt4EA2+2+Sf/yz3k/T9S1CSt2u
uWU7uVY5opOA4u4dGj3gEFm89ZwKZCXmgSIj0P5RfnlgxyXZ/8SXeo8xeCijno2utmIERsmMNHjl
9etWf0oBi0xeawhkX++oWjymBxthC4Ov35Ad3ryHMA99kmFP1yMVOraVhQrKHTh08Bq0vl6YO43y
XH5TXDXRKzrTk8nX6zAGU5Mh8NsNOyYzhyTkDN/BoV6BCBZ2Smjyi4rJvIEfq8jx5QHuzYnzovb/
QAE6TGn80GPIIyUyMLpuDPslQr9Qox3OtrR9Ji3kZNJzjJq/uKH+HUoON//fz2dIPVIQSLt2dY4t
uNy/a6pM7c2ada9oujn7XtrlCd8BKyw4HkS9Kj+fIMgzaURg+0B4tEp8SB19Hgu0iHMwuuO84i6H
51nDt5kuDQt8yGcLE8CbfE35xRsMP+nFt/nO+TY3YbneBOQlz6BVv+OcfUsH1IkvQiH60tOEFAwB
0xtGkHzYtu4XoAwyn49iR+BAlyGWFvnpGEBTogOgHBAHs1Uzlct4Uxzt6ZCr3mfPYTS3cFCOIyzi
FHpwBV/i6SvGIMiqkulInPwMKv2B4YUZdlfAXbtJfxdubVpS+/l2X6IKvqRTKjBafC569fFIe5ji
2TFrCWqvyF36OTNv1cH8XPeZF7IAdVAbCUYKUnVQEp7IraZfojz/O8OIbQZFOhhDE0WkorNdpIZ7
NT4CZblELK8kG8M2drr5y9/feauHKRW42gNgXXsJdpm9lGqqCciQxwzAHHeyXryPk46J3OBMdWrR
AKgJmdywC5aOwIRHqOmZHqOWblbis1AHiOVXVlD+pdLLFYcGvQmwLpVc/NbjLViC+GfStddAsFYy
1xdZgEkaZsqs+6339QrYmFdvwrxUYaTowOKsQypWwsXk/4LvpwJxxpdBdvER416jbQmkOZNGr2kF
7kh8SI0ZWw6rNxksXCCwVmyFQ3ZNOwlxQieD9idImc25dGSPucOKD/hR2vANMO1TBFBzw6PRiz1Q
NwIiRAaMb2igJLJkX14xkh0jUuvgaT6lFoKGr2ReJeOSY+kH/MabyJlEEtvNa24WMTOZ95XlOx9J
YgaKcTbMoa6VTZrawaIJD24R26vkdPVP4DcrSi7z3nMp2tqyO0ckHlyg131u2RyG+9YhMsYETFqv
CeVBM5Yp6fEMtRPBmHf3L8U1LYYA07BeQ3y1OVRd0Z4sudXAlr9qiUucF0S1yEQxkGToQS0MKGmw
ysvOaDH2xfWeFD/ioYIaQKWQWFag4zdLk3N559vgOGYv6jGNwFyKn1s+K8LQRmRsaJKixlJuNbKl
BwnLolwFBFkglI3IiOcMAv85m/vRtH6hemfCkGwcGi0AoPzUEJJ3DMWb3hu6D0pdRHtBcWULZ6C/
8KhIJ/42UVxx64W5UWDXe1R9uIJkDlyDBUZojFZDYHIJuvXiMZ/6YfOF/j2dEFSua77wtbQApbdF
tXMqO1DshmtvgJIh5clsHflyCpYmKakth8DLew8wpVwjlJpNDczxutbyp8OwJdZej5MWxsibYMCp
H/STbOXxuQBFXXaofFrMN+mVnYa1V2PKtOu28sH71lfUJ7LPJj+U1Ck7g+mKeZVb/pPcgb2dqdu3
0R9vXSvFrPAwWAeW7l5grOsQ2Qjz3+NL1XLhfHhaz19ZXcnfZrd8sn3PwImuGU+PW37Fpdt2qRRN
UwvQkiLYGStgPDRsSlc87EzOpUmjbYLIjkNw2dI0IJg+bFCvfsc4jEOImi3UI2TDgJvediC9Ox6t
sBmNgwVpRxA8/6RCzKxR8cpA8C5Oxdax1TpaGMd20gzg+mqhYzww4t4DMf6S7N/8nWXgQBCV0mny
SWELq1GLbcj7YGrNkHvIGzI5TJqsM01IrjEHXaTNw9E9eWT9YH8x8CgJPQVyS8xLHEb3iX1Ut+DS
4VV8FaYy7RUBSXFfgeL05j40ShgA/d0yRF1BEJhvM3J1ASzjbq+SpcGm+QDtVGQ9tU/zrdBqKTk3
DAUIqUkTRlofiRUT+DDgHmbPsXyIxHOG3ri1JpH6bvQRqkTd18twxglLmUaoqTsBCfePJPpbE8Z0
4m/RexLEsvBcZSzR+ImBLvl5ZyoCR6kZMKJZsVTMaDngW/b2WmXc5zz078LsXUPs+GxO3kI4je0H
dJuVyieNJBrgcRRHVz26qQV/n+qvc/Tl8AIHaWfftDkqxhuhjVnPi0yp0Kg5nHFQdiIaigFwZW4O
RNCQt4bsBiGp9MDKReI8bzHgt8ju0eMzDWK5qUusZ8kV9fwgBYC57ZqYEtVCA+rWgs7plCd+6kWO
iYyzAkRcvLbLUDpqmfZufRRP1ZRqkowV1BdGohbGhn7eEOM8Jf0s47QgEOZYpATvE2J62qASPLvS
lP5SRnpLrf8wpkzpJg53k/HZeuCUHej6yq7eh9j56x762+rXov7f0o4dRIx7zQGba+rpmvLIUS1N
R7pnX+AG0Sg3T93kI5bAfhym7vWi9PmS7te4AMG9tytlaNdqMypOkUQ5yWdubPYqaWNRH2qt9lXm
ZEaR8jY9iG8PioIZ7KSs3XMxVZOfY5ahA9seJ3iBjdbjnrW4LO2+3Rsf53+p/1SNDoTsWMNrh5nm
KUr8qFyl/iIey6klf24tYebXqznRzjFMVXaGw/LeqZSMWligzKZu/z4VxePQiqqJB7btP++pSFba
pklWjEdxoRqfx1whGyuqoFQBmd3Ve7mywF2gEnQ4W+ce7EtMXYR236tlOGU25f42EHNTe3We2oOb
yJmKHhid3j6BFna3Tqt1PijFQt0lWB0mvndHvPwwJOHy9FvKCjtU+cmnNYTIvRUx4xQdw6PhX/Ur
EKcLondl6M7H3G8dJUK6UpiQaxj9oG3asHq+vKGER1gzRZ8x6VjneejnrxnjkFNpulTtRDEqg3H4
DHqn7nezW/otpO27WYu6fh7QZZRImuw7gtekaZ16hmJrdvdBCqsz1sz11fIhEfHod5UqFQPCnF/R
xX+Y/1Ns1nkxaRiio28gDFzGbTN+7p0cZS4gFbGdyJu6HSSSNINm0aBBtZ+AtzTntTrON/Gk2b9N
fDqWpOIILdj+gEjh4Gm82ZMdaqlWNs7cgaB3qm8ygggKIbM5eCAXty1zrqKZlUJZTIYiQULJasVS
l+5xrtrDxVQ0AEFQOjV36w0K44Ne5yVxwK6uXpS5T2dLJEagM6iKONJXEznAi/d0zp57INe8IEok
GKUAEEZ7kmX0qOlciWFua/rU5v+vYzcZ8Xlz5fw3MAJ+1rViohBzFBpw9wqM0uFxLm307cwR58aN
+V3h4noq9id4x7RAwB7R8b8+9L8QyRQswl9jbZBhc9+kI7d+mbC45cnJNpTVlhqDvyWO2I8uPjYH
6qxq5qO+bQrGhRvFQEbsVRpGgxAeBXMPIX4WvghVygdT9Ton9pfzuFLngf5tavgmuQNWumH7HXlv
IWYjfM7phwfCHz+KnI0eIKRpIi1EXDtVICkl4INyDjJfJA72+fJ1lb6yIk0WDHvx7dx40rMtkoAK
pXbDn4K17fOQYluEIzUH3AO1NmqHRy/1ZHtz1ABHpC4G+KL3C3JqIW51x53kMtLdRKsw/KbvZ+7r
7A3lKiC6NJjvMvLmHyg5XFqzVItCEF3OgKiAn9BN8o54KC5chF/3aVP6xKK74pgYVUsJ/F9Xs0Yj
YxaE151fI4frOg5b3MtQHzWJDwWZlLwH+mVayjmgRkATw2QFu0PHPDPluQoK32rA2CC53m8K89Jb
v6fEsYnssgal0LE47aqIo3ph/JxEj2ampDDNJqxKR0tq4RdwsWPwdOi8pYBGJQcX2KqxaEs67Gnj
0k9QGWXE8y7+X30pJ2CoI/HKfuZ8clewip9yN22+sGGUh3VMw9JhMvFyeKuETf81JHdWI/CzCaVc
HZgFJOuG49N6IZD4cL60zlFciDOC1vHFHUz4VLVnxaLR04HveZxOk4dtEOilT0z6a9miA2lBzeLd
eXBkumMpF0Fi+PgaoIS+f59WzIqX0g2B3bVyOMKHAtDgPUoqbcERTuW0VIJmCwBynH0hz6U3IHL6
IB/dTCg16d0PU24ZcbSZpgRcrV8wIOd2pdYJBvOc4gq5lPRMqP8x/wXgtUYdPUaKfbJGaclDgnGW
+Kgga1KoZsKl0yM5kRmzCwED3QWIxHQodTCXvBHeh75H/ytppNz8dU8avdhUyC/R1QQitgA6HK2c
Q8b0B6Z015cYUzUSWbuoQOtdl/5Z63RjyTHryJvNEpZqW0WkaqygXXnnnlOiLMf0D1JFt9yQWH+u
aFkEqGw/klTjcUzYc65D/6ZoL8EzotE1oaXvKY7pYVerWggOLQkLa1LZjB09yv2V56JoCsCNzCVu
Xqi9x02pbDL9WbDWATFFsY/9tTLgdX0I6osZpg5imnGicjIrBMuIgOEVr50wMeZ1ejlNyEbGoKbb
CYhGTQ4SAhpy2zSL3KQmFxXYVM/jbdAh34k7oC69QGiGcqWTnGevc3h4M7OcV0f1obMGiOoTk+BQ
qtFdClNXX3a48xJoSZVHyrfqjyq3w45YJNjOffKmVtzqQRX4ggRqURwgdX93fAq6zv47jjrarVP9
5Nfc8KC0HeowP2F9ggJbZ1l+Rm/RB00T8yRpPYEnBcWMyCQizM0caHuFxJ1Cu7cVuiFVQP2x0Cbm
vH+EZvjjSeXlapXqOMLSV4G5KJSzBp45F3ZERRrN/XKZ9fPg2a9s1jPPQlWMqTDVU64hmGbRszjt
hoiferFZ4C/bflCxXe6dDYD7ca+Nn8bVkKOxIsgOhuKrwztr9K2q/CcV5YG0OVewRGeXWaR4h+Go
E/qox68LAUNhJx3MXw5k/dUzZYzjLmo2ZFHqt0XvO8ZlV4mloOu/O1BVWvwfLVYUO93Ph/o8wVmr
ta+FiAgd6H2ES1EuGf7RkRar/FfOdeMgIAtwHcKUhLJpctYDZBmWr1pzRYC6/EYHqfC1svtdjWx6
571J8PnhiGi3am1aTNkNEMUPQSZixBkUgdsYsh3wGq1JuU2cRBXbfm/Jx2YotRrgfCgBRLE14RJt
m5gqi7e+0TE0yx9Q7LmaTh45qIQf06hllej0dB/Ztebn9p0v3ZpLZuYE+qOPhgmVvmULUKnzhqYe
fdPWm53LQrsbVebZ57O+2xQ9IV24+9d/3yzG8eIgEZCNCXrssgvZQ523dPIMJBa+hY9rUjI4z7wY
s2S4Xf5IkeCgjcWFH4NOZPo+sIvT+OdpgCte8NfBKO2gFpcpPw38yXI9KZeq44ZRR2AKXdt5HmXw
7yHE4c8oPhth7DuAwDiVocdZAyqXJSHi/eFSA6HbKSIErIbWH2kGHwBlXmuQrc6SHVA+cxeIMIO1
YTdcyy/HeMIad+Mjtt3oRRBZpapr14PiDVEf6lV1T/6jJw+C+C6XTw1T6+b8fPiZ0uOmVR0fXVbl
ONsUK6gxJFRK2b8GfRf+Iow9cbiPTw67rFCz+iHPglHj4CgN3OHMeqoKGJFIfiMXfL33/DiTUiWN
tVPSqzxSbuB6Mxc8na1omTAWnA9tHCr8Ea3XAf2vVpXIs9sc0etrrNIqiP9BApV591+UBGZhK4Kf
ePPpACRsaRx0BQ+YKGlByulnTOdlrOTK+TvdvV8tr16vmMz6qYjnAhsRcRbc5jKmnvllFjCVnomT
p+5pcXEsTiKTLRO2j1NLvkUszdJza9SvaR63ziE8wCBo+Ak/kQDK0YEPdVYAsxpcQXs3Pn9gy17B
Yni4IxhGezXvnArPkI421jEK1bkA702QU6IevUH38be4jB5npb5N00lXPJdhfDy88FpJl7fVfgAq
nBY95qW8CZFq9sOkswveqv3VGAhbVyRk49oEKTtrZXTNOOC5cvS3u2IkyuOcjgbyyhmxt3qXU8Yd
LYO90PE2Sk9dl78LeUISg/I6/i8jSu4iATcAA2VybCmQA4H3sW5Xw8ChXlKGKcvFSjMSAJyTwMEp
OLxojaPRGdRj5YHIJYmQckCST+go+A6elAxvHaGF/d6x16sRHv9/JszS1JWLifRpy2q/ZCR/JOFk
neSbq0q7UalGqj6cYvNnyu4lkpb5qsmFS5ma44Ks1fRnCFI8KGSm1r81EGM1Hzli/Yx4zzR29/R2
HlqCO56TnPLgDv0eq70DTBP6S1WcnuMc3wixaDq1+rhfXyPonUQb+mxtNiQTgoVfJUc26KpGCame
zAEtWRwdfzOewvtJKD08cZRIMOwotjBc1y3tCD6SPfwEqwZc/bMpvvBvSiHgx+ioMnlPvKTr7sFK
R5hQVGzgowbQPDkMiadumpWNc2BgbzseG44qta1Pf5YUuBVMhroLyQU6aS0EFnJIMMiBuAl5u2uF
WeWo/tcZQeGWvu2GygYwwx/5ryKFdCnQbSdZN9+0jPu7AMJNPjgtWFcuCZ3OzD+3W998AWtm8G6t
35+Wv8nxaPthqOd1KPWHWYzTDDZbqvWYngegGBUYeJD2COzGIovC8MmenbAPTV6nvFItU8wlUY+C
RsLEJ71nnAwqryFvr1KJaIQrV05axc+3fCJSFSUkxVBn5gN3eFWIaETHJcVfR5+8byg+PY/w+5Xg
yql7FbE+uMaqrfiIUmh4eebPnhGux8uo+MQLnAd/v+TgJDq4qgSUTC0iMSeiy5my9ZLc3JPjfcKU
RTK0VsBySfO4K79JvVSNV8UejviipQ3I5ThZRwUmvI0jIEAGUHZf988UFnrV0PD6UHkh3p5BEgLO
6Ne8am5QHQcgNoeL7x710Gj3/cFfq0ESZ+JYyOGt/rclhMoNhnDgEqdfhzKogpb3eD3ueuDUum7m
8Naa5YgkVF/0bVbNh5VO11VSVdiEP03Jje3WNJwXsjUYuJY8xFoVwk0r9rtIuh5z2js4IQgGVVxe
52CbCCllK4GQqBtJxNqC1goc57qs+W6aD4DTc+DwKDVB9glsV20+mowTpQV0NRKOQgVs9k6ylep2
WFq0E7dQjDofmBk19CpdTYc/2wxqMPWim8nfj5s6pKQKC2ZYjZvun8CqkmzNZVUM5VCnf2p88sFA
ksTcFyK0B8e/qAU6YiCjbHA2I5kqNIMxY7Rds3zaPxdBRupSD2onhaBAye98yDiwhstrAlx/Cg7Z
vkTuJVlBDU4Y6AwQQ/G2aEJ3vndl/riVvl924ffc/FKfTJ77kDvZJWOTRg0e0UkoLFRBni7WLZXE
oxRK0+msGc1pdGPWQYCb29XTAWZIv2B9HzgbXpXw6yrCDz1zbxTJZd1HbijGOd+dRaX2/QiIun6w
zJUXxWu54EB4cUKZtDeMsy7ZXheot5odX29D04dzW5bZ0Mr6xtyElQcXWil6OKxG2gq0oxdbBOLN
7QtKJCzPMbFgW9HSAoSXcwpHdKEXjrPhZLwf3mSh7yVqdREbnPPeZ2EvlNzesPbDFpm4XCNdnUej
n4lQ7t946vxvNjg01LsAAQJI/IMAQ/y8UmU9dGyhTtwq93AnHHsYWvbABJM6SecZ6M90EbUIHbE5
7bVs+VZS2s8wj6cjahtueRprxzg9QgXjPVy+ZXR91mVpZzKo043WMxOqR2fhopSiV1dZXA==
`protect end_protected
