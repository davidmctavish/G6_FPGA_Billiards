`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mc8LZWpn2E6sYR1YLaosWODd4R8lfDfkxbW9iPFEBqsWtP35J01TYRRqs9J1uWvy1Vt1um2T6jv1
JlkkiibrVA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GorlH84xkq+O2R0IJ3Iu2dLtvY9UAj6VcmD3wwrWgIw+hy5d993212Du2wzDWnag5AJSAwXyV45R
HkhJlaeXaZ+7FsBEOsyd0v9rE/OShKdnGxkilxzixfWFGGDfZzHbIwN5CU0HKfzKre7LurmuU3SE
4DOsIgiohYc+iSq293k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4gX/j4N9zCWXNWpuoylh8njGJ/Cs4ViHuj1BVGvvVUH5rYEJvzij5HcOrUr4xpiPcyxJp2pgicr
vda2Xvjfaowp9GBbsp2bqx4+SdLarrcYRzu7qjsgVpe14wuStjhXgPMOpruayV2Xrme8lByPPjat
GVyxWn+8mCEhc7YLCRx1Nrk2fjLNwbTFlr1igdZeJvWD1vXoa6nzWR7EeDEoJ7xGbehAGCLtAhd1
QKp8MJuF3ffb7zEjWCZ7cwwNqWiOHXBeB21wN3BwPW2eNbu/OkVO9EbShzuGhObJEWtTFowNJmB6
v1gvxnr67sQf+yhFjajVtcFCHvqOGbc+RZyiNA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o7wAyMhTsNjR0WJRPC5+P6xs2vNrYznNJYpi2H4BScorqSfwZJtBZvAokSr/uZsHOeA+Wd6UnBsl
FBv+O6Xq7TahQy0vww8ocF3o2UhC8hCWTKnLe2cwGDVIcpdtcKsqjUCBgl9+Vd/BlHt0R6YZ+1am
rAdQtkxzxR6Gn9YpuVo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XYMDtQPJ049Dv5lrLdkZb/m0PaAswX7I3ZFBAEeGPiDhSJbxBkyMiZTJzcBZN4n7U8eFzRsLD8fM
3EUR4aWwHkgj2d0Kb9xwBnXfg1kxMIBGjCSxiOMV7piI0UoAWgwtb6nWjrc1wNyka3mDGZ4md0bk
2J5jPBLqYaXZtt4iuYT5wfkVRzR36ixy/lE4ZdicZKLCkXYBgX8XvkGnQjIfTnuDBQAtl3EMwcmO
Is3ihOmNll7yYu/rXXJguLnPdfMt0veR/nj7zCTb2DUB8We2sNxDvNF5qp4c3tReEX8JZSpTYro8
haypJLC3AjECJETXooFSIWkfZ9eDD6qJZ6Z2tQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7664)
`protect data_block
UBoQg69vIEtO3a2DQpJR7MQlI1AwoXfpV/QwlsE+LAelpAk8PJRHgaNrlJdvWBq/H45GbB9e1hQV
cBkl9++p9lFI0jzk7WDTcyQLSpFOrgyAA19vFB+VcQgEbZKpOmiVXExu97aQOm1o+l+UKj1TkSQ0
hsksbqnBRVcm1WlRUd4QLN8bELGnfjmwG6P4xNK66nj+2WYFBvE+3qf5VQS7BPiS2jQV6380Jhpj
pwYF6ByINXVm6krm2OlHLh7gHOBMIw4BvdRcTNXhoC0RnCV/nnKNPMqwPPXoTrlMiUfxJCbdRfUT
NeBTZiG1xdI4temrDjUcv8noaDdnnJLyjwdV7giraUINghiAO/YVaOoU8YTtkktGbaP3dKf2uasH
YzKPzFk/8p9LtC9k+mxqmjnd2Wan219ByOcnUmzVO9/KJRKIdoFOzJqWh4fW2q2ZzZ0dF4eO7YPL
zKdfCPdUy2RECaZq4as3a2l5mD3UiWlB1hH8xCqRsrEcoF288AQO5SeBC/ssl3yeB+Uo7Ef7p+6o
wShXNrMDMtcWOSKhM7BDiKEJfVJY4OBycBfzk0m2bSxEtS4ARQiXSr/ASOze19Ne4PSiDVUXvmQD
eXa6z1BWwtfRCnXlS/HAAbd+Lx2va98xeftz0ccGR3MKm2A7Lj9lKn/9IVsDRKiPbvFEmRiRquva
zT/O/+WjeB51VFQUKNrbHjsE/Hd0vlPPAjowymBTwvH/FLpBDrKmc71deqt1orcAwGjSNBWlFXMu
lb3Qd7vyF5DxFEch8cXsw9Jwx2DPssU1CpyAEbmiTszqUdbyQC/CRxTWH7ZG7lwsrKgx/hNmPp7u
x5sjOQ0AgkfkefCIa0HTV/m3FH1QPSdq0Fn5A+WT1MYVWB3JKoGgKxhggqD1H+Q5Bw3hn5LIZ5df
idXGs656fpZXrkHWgbblUhQUv6sOgZ3stUdaPKQKNnn0afASdAM2h6pugSjFouY6VFM15+pso7h6
dH5EIm+ItRg36+EuxS8BDGXymwcjoCxsUCtALmWxpFpazRkwxTST75nRPNC9d2LwUYDuSJlgScoj
y4ibVmc0lac1ImOzuI9X5q1WtkquRtV6b73E050fXE45E4jQkG4eDvR2aNBWKxJhMOMqq/lTBDt3
oAeqsXSdLDDtdQmdDHYsSyH0vwGuLBTa9JM/xfEfGrwooPt8dAIjfVqzRrUdcyb4LylBjpRPponU
76m83Ze/eq5eWLH4xepuBWUACJT22wlIFc9IjlkXO5Nj0kNCTKIX7E77Dpgm5DhcWt7st3twUvXu
/xnaS9FZ0IrhfKx1ikUuAOTaTAvVYwqR4C7smaWplVupriG6ZDbOsxjIqKrWXlaH8aPF41CR+PCr
n0Ese+8GedM08RWeFswlXxUDVImDmXBNJQzqi2prD2qjqOUeRtn55gJdcXkAt5wjDYaolSv43LVB
ZbJFDHWSnRabKzxwlypsVO5NEOeFMCdpRaRk44RUbWsW6BPV5bhs9ZHTPp5ftxUW2U/Le9YwXZQt
DwQAbHzLaViXpnI9CyJSEvQLYCdGZ/yaORJ0qsk1vFDsilKX5T716qLnjkBW7EgQP8Y/XY3ACRQE
nrdool45ik5Mt2Sbck20dh0eizQ4CoYWlHmZ5cuhyZJIzQmknuTJZmYMME0PeMHAuup8LH7w3QeI
lQQLco1n6VyQ/98k6eT6oxzJJsbzMOVAogFaZvzv6Rm6oEdA9Wm+xh/rMKCXtfjrIQT58XP5nN2O
SOVeCMTBfBxoZFo/NMXMEZtU6qqjrwfKNsR0e/PQ/j5Edy+O+KFzNJZEsN9nc/c4t1XbMT65axE9
cjpOFeA3x+mH16VR6GMx78okqCATHSpXD/o2rqnlAKJMmrFXns17A2XErjb4+ZaHp4zJId/lxhUF
vfoVw0Uw0uutyaVIWkwUgjCMqbZyFymof360/q7o2uvvoPP+qXvvt/DHkS+UuH1VRYInKW/+ceJl
5n3NqzWNK67oEf+KSuPd2UuQtmH/HJy2oNagFH8yUQ1nU0xwliQ31eXRKd657OwN1nnPojLjTdWh
VxcpZ1bs/Ke/8X0w+Dsc5ogg6h+6poRv5Bdg0LrYYavKQUn085H9Mdayj5eaa0sXApalJKcYBA53
IpHM3KGsrGRslb4nLB7QeDv8ejCnWmggh8RRep4SFFWm10r1dhyBFuLoDqAcoK1a5MJSYv8uHpMr
HijJu0nlXza0Lb6P3qdRfHcy5hiwAH9Lkm7RYuKLRynHLiSDKT3D3+dsc4XUtfLAdmI+BG0y55Jx
AGbGOBldR8yJDvRGyBcVDn5kuulomAoiS2TQgijyXmrH1OVYnbqYxZ/P0jUs65DpfDG5O5/jDX9Q
mQpQ7M3ssXYVrGUWuDUc9MkqQ5IyfGB7ADZ0sWw6fv8hep8Mnzy6S6uAbsHY1L5uYXSigVblEbir
FucqFrnVd1TKN5msb2yF5XMcqL8VsKLPZXzEOR+TZmLV87N8q8wNI+mDTaYTiZ7+QFweMRIg48bR
62BeyB/lrW3n7jB/xr4SEk6KxJ/CseaOWyqup+Lf3zS7aQYGQm1ftSXkXJl0KLE70kLmrE1lJjS8
Kea1/TfDv5S6eaapVGubcafqJ3btPev4fBGb5wTZ+us/+vMlN3bXJt8+A/AqiB+x1ISilPaxwSpF
zTUGFY9xzcISku0N9OgjUV05r7M25yyN1M5lmvvjeX2wUl5xI57El76u+Z7xFpgqD0qdCzvxM3ry
HXmt3ApCAnf5kQRGRHCF7huX9xIimTnRBS3PYTtk60ExfwdyW86XEgwUKoAAPJ/9aiiRu3h85irR
tsIEZ+5GSdnu3QK9/OyDNiiqc9IaoofJOLpQ8nuOplEbq5iLw+iEwrzZ1wU0U3obrsLeb0OV1/gy
IttgwzsHTh4pOqv1VsDvPIGrFQ/xM6uHfEwovzY6HwJrsjJSzPzr5J3VViOLC6zviF2gEz48XVm3
WWSQlyM0cuNdp7VW1Zl5CzmkZGaRw5QeCQpxKvytEF7nkFM3ysbQRg0y9wt/ZmxXncupEKE0AT11
WZow1X0fdlQI9diftEYixI4oBAanxPouwX47yyTCiZVTgdZ09qeu0k/E4juw20GvgaN0UmEMZ3Tv
pOHArs7IiZF5s+COXIf9NjWQCn1CA02gPq97bQgXL7y+R1aectBMro8R6ZmA/PujSs/ms4w11PGG
xDUg3/vGEP54OpqNO+i8yBJpDRNA1xFYoqLh/85hwlHLYNbo3pnod/d2fTedOJ166h38FL/afAez
KIS4Q1exh8VR37GyQRzVZaBdCd8qMmh3CnKI39P73LFLe/gn5p/QgVNUEQWMcpu3ey2cuWswQ/og
L0LdWs/wVsv+e/bwPMnEq/8leQ4iez7m1aLqWESElCukBgs2bXaRtaWeoobLKSxJx3McBYVgp+sN
+9RXGEqiC8Tm3Ax9AlYcnY9N9tWxZD+MNqb6HkHlH6Td1NheBIeTRrn6N7aLBN8fKXn/0TNvr4Zs
S/J+e5eAUfEvIYbcUs5hkkrzLR+FXE4M9nm2u8fV3Hpzs0HMCaasOYPwG5yOfi33UI+DR6VECcYr
s94aQKzInRi5MlN03GOIz4cirZP2hGqRLsIqDxkWGhUccZacO98buwCvLU584TRfOYjguBQROUgt
cK27efjgXDjIx5XpGl8dOB/iIuDmSahrG7sTghzJ37OIIfu96yIBBUOHXYmicC5tZ23tjwpN0Inm
G8wwiYr7bZIjE5eGrnydimX+UdBMEkNbVFM4bbzX5vy4QMFmCM4XSTOHLslOiotrM5qoGGq6ytnK
ICJwx1gMi6UFyHQpW4DP6sDEiGQqJmsYTepnP1ELxj9e4bif3ShEKgrlkRkZzcRoau2xVguCwQQv
MLMZDy8L5H1ZOMz+JoBOapcBjygfUICEy5a8wi9OBU26Q9SovBFQnR0CFr7NQeveZtbwfVNXqJXj
WC4ZShMZsqxzdV6KlOakR+mue9nq3K5GUrfFptMm2VwP2h8R2aqd765aVTxLiSyltUObMke39C5j
QomiYKcjbRqugMx/U5dw1rVIGCUHaiNrufIql9oLuheOcAhFeEAV3w3dpizl5PyEYBuyb5esrlT3
PPYcd8fQ9lCDcNAq+kvOUZdHZOB/ST38I54wBNdSt4L2mEa14CjiYFfPJfWMMmTUsgefhWxQpPRY
i53VtIkIVpnWexO8vBldZlOw0SuLGp8hPxRfe9vOZAmkBM4oPdsnjlSh7vxXGV1Tm1pU1NJABw3a
2Ig8LLCgybTlRwbyjAwHFnzgQpUdFB1127kSTiz/OsGJSHGQLYXjun/qfBIGxAX/H0HJSigfImUO
yTQExfc/GCK5bZ+l38tRR9dbpfivIyRSU8onNLaB4quozer1u7PAp505SKW8ahCrujMWiRPy4aP7
rjYNgjzTNsgaDRuMrYBHP6SpBwrc3V02n42ZEmOp/H5c0C7Z4nb/eXd9DlUiHVpFOu+aRvNMCbq2
0FGq/BTM5bWWtxOhaO/asbFFXm9EstgLMi3Lt+0BfeTujMsotiTlJFqsSVbr+A7kUofc1bIYqWLj
jEmntLTPwqrOILGpPmCNm8O5l63l07N33sFFrXXL2/3KtscE1GXhxicoq2Xrh3Hgmb+5X57CHE3B
uTNjRcCkRqt+8jeHJs82zf1+SiTe7pvyIc8/FO37V6rc60PTYRFp/uXAGsPwHpyuMDrYiLrYu1/d
88F8nvnvprfN19w4KrH8aV9i+IyzAP49mApzIVKXbrKkJ0/fi4QEHcoKTJVQT5iGEReDTAYFcSlE
M4J3cAM8wOKz5dQsvNQFiFyKPGtdEHsNBuPiy8aSslmBAlPpN1N1n/y4e8L+neEJyeC1eSxxFby9
25hnJyGCDUFx2jln7FiNiMg2Y7S1uN3min3AutzCdI0v220Lrlgq8WO0OBemV22j1sM8DXHQoxdm
0FVKC43ijsA6bJG4iev+S3/njHSDa6I2GAfVAFHUCnkaFc71mT9YQkAF0dGrmcmJ7ejX/hxb5BO+
fXxsIly7tL3qbqcp+ikskTr+mIjTZ4R9lSBVR5lRtDu1TeQLQ2pwX081OveA7axNtyWDOiWlv12F
dgmdCOpMd0SZaM7se35vUHXXS1RUpIKNb3WGoKF/kALiJsNvK8nvLWoBEl+ZkVV2fmImwpFG5j8U
aKGKbiVNUSELOUAAy6W/00/fHauqyw4vbBQddP/4EhBoQhtnYl3zZ6v8AikiMeCKe4rcWd3wJv28
5EMO6Lqyr6YA5lO09oUuapV2Zc3jEju+iMYRRt+e1iLkMQLG7mJoIV6tzfQOwpMrXcB69DLFsn4h
QSefLejkiUw2tjzFZRwngj31sVVlHBZS59KrOqR6NMfR0hxGMyncUjNj+bu1PFS41B1tAoh+adA+
w536yfW+QeyybmRyGWOjl8Q6eFp0cHjCIiV0i4MNsn4ngHGNLBop1eA3FZn3IwAkV45PjacTGOLO
tZl9uEcHPq2u2FqsBtohQAXL2dTZaHBFteuCb554YEEYdb+H1+nEZMM2Jf0d9SUKG8EmFEmnJqli
9wdWzhPcfZlBfUpdbQCdEZYUasm1YI+S2gBiVOW1uHvhVMdxeM7Zmzk4HdRfkhwOI3x60Ir0USnC
ujm8mzvWL8XoEkqCb8pPuNWJcy04N2yPw21sAnz2da+iiCGVfXV1TrF5axGiS8jrEarShp8imF4b
FBpLm9/dmdLDnZc6rhnb1fQrvA5YSRHr5fGxJpG2SM4RhpI1KeaumrTNykf9kpNKcgzF3Zdu3NwS
PNMqeZdYSbKBavfBFUISqfcI9Gev3elUW/BIrz0XbiKovopoYyygB3qsI0DygZUMJApXC0fhsgFy
oW3xZiZyEwvriBo7xLMGqNmt4pJVKSyWzWwZqrQfuR9QzbMQg5yqkDMOPwF1K/oz2v5/jOs4jqKv
TTMc+TDs7MFUCFu7KCwqS35al1r2rSNKyHS6obiyDesbDF+PcrrPZ1NWU7U+kPZmWmMmGDL6vOHP
46bG5qhDTe7D89k8vi7PRcrKLWpwO/wxgyqsY3C5aCXnfo6tIAQ1vu7TWfemM/IGebnRH2fK1ahj
bxnGS9Ck9yuIjpNmy5Qr2m2EpLSprF+x+o3/blf4m3a0zuRelXW62J68tkUNWd+pgghJbyi3ttFS
cAj80QjkVOCzvhiGKFqdoaFjrcE+8yOJ8yHb1DMuNfXCOg+Ur/YhddEEPcdv7cpbjytg76NMg3we
KORzm/8XpeN0jTewFQsu73iuktbxkD4wiFVSUOgj7GAdA2jZ41i49IYycCVBrwnJgfNi3ZkAfsoY
2TBqr/j9Y5qdK1Lm7QDOR8NAFKmVvlgHGJsKnYdUTvrkHfP1ub0vsQ9vk+DxqTLRBn466U1avB/0
JJC/QMLc5cs87bImdy9A4ZyQYBqlGWvlUS1STYcNBoKb/o0ZqAnxQiLIg6qOeZjrtWlWKn6G7mJg
G8/LZnAlkt1EaMXEet/ikYov7KMrz9BwGGV+p2MDLSfx6ViS4FmLC05m3otc8kqTFpVefTLaCsOS
5Nst37Kd3wRixC4TKSTY209GPKsH7ubLaUWxV6jWW/7k+5R1lwppiUNZbgCFFYT4lKqR79XA3JYL
mYVnrAnxUMXjgAZjqcTFrHrmQI3yZ1/GccaL2QOpK8xn4cFrRMn1CiNDIDh76S8YgEXFgZKrdy6L
5hjbCYbHKoTQlnoRwgln27MMglC48iAMC3YONoyORRDcXI7+frvQvUETwmY/Iz+rL4Co95Ip6PEt
cmOL+XeFdvHBu7bLTEnhGXZ9rmdRN9SWWvoi0S+b1wXiB/L382L6QJRp+01/Xl90y7Ng8m+bJa9A
TbmVFuxk3Xf1ZUK5kwF30IDfWCFKNpkb47/mMqXSgNZT3lwXlmN7ZN8UdsEJ/lgBv3CbU8iA/j2U
EapPnX5KNDCnpluONr5AAORPIbjRgaxp9EqH4fvWUcHCq2wJQ7Tvkv6LdBEkOYMSUQQ+y3pQL36i
9Hcaqm6Yud4Mx7nn1q9cQV0VE7y1HFVTjjiIMjEergtrjNXVWsb7dTvzf+ytBi2Rq6CV2QqNJ7JT
IwNSzaO5hopEwVos/HOQIh6cPmRfAdxSfztf9TQEpHYIR1yV4qey97o8EtQ5OAD7iBpUvJhs3Rye
N/kahL6Kimew1rFhWfSPc3m/Ja4A8kFrB40uRT+XftDFo+YicJK7u/ZgG0dtfSSIbuuHUcZ4mFvm
SNjwyK1pUsEHb3U000mr8M+mCdG36mnR5TP1WZePEktmRYMzWCadXnR9TOVynf3nfbGtBBeQf//R
+QrOU7BqiwOATob4Cmer5bo7a7ZTA93UtfRT5eJ4PFYwQ0Z8+zoWmuxTbrhbKapYszRFyRriobmW
aC+PUkHit9S1t8cD/Dmqbi80xJnVPqZbQGC5Gmw+yLO8lavpMQ33FQF1S9VJWUbmSUQnUHGLVxkM
ZS6hURdLTssr8Olbta88e8AugoeWpTk3hfqlBzYKzip6/59as3Mpz4ldGIPsvtuxM7af4ZpWn+pQ
yB8GLPyDCvDqgfJ2J90Hx8NflsF7cUIIDTdMNAgK1XeID1uENhBl9GeheZzGooGdU8s0Jy9GmjDY
G9oM/aXwBzixm98Nns0mP4qz/UDVwBgN+Ccg1bTUpMGXeCoDS2BCxap+g3Cyv5uiBn5BnRDw8Ebx
kFe3ZbBIJa7kdz+grDLHHmthAetpGwTQ0JA2G4G+eiEYvty+4z5zNq+8H4qxCvWAHVpq742SZdgs
loZ3+CW3Lx5jiEXHEZKk21xabjb/jQA9wwQwKLm0yyTUmytzBTzDxZ2DpYgD66tuh9G1R4aPIZWs
oyiIyNKD0JggGyCR+qBpn91Kawebg24hKQJWlBkuRIukmJK8de/NXkHavsp7vimph8xStABBqEPC
YsvHMIzaBIxUGpum6gNAm/4MANqvGGn306qFyqN19UdITLPxV+AGyucKspXGghhss2WjMfFoavzF
LE9Ffu9ZSAiaKRz3WERIt2fFqodWa1nKmnP2axsSCCdWnFMiRkVYKdIHOTQqLm3JkRVh8SQQUNIE
R7plaVbvaCje5rVEXvCY8xRdqVyB1Sekd98mKEWCiJqqxr0WdAwx16oGkCV4MLgucPqfu9hUP535
Gn9lM6OwO9jgYm9Iw4G4ybm5bY24t2TGlYSqqgY7+6asYxeg5IK0osz3cO3J/LwYBC6K574knQgg
NqmsEtJgVVeHJtpamMlkzJDV5kdU8Qy3cnzOGZP4rzAAXC94wwyNU8aN/g0AQ3nXz0KfWiuqNh92
zZM4XnUHPem97sTweu0oFVtjOn1E6dCH3x17fY+0MJ1XPSEittzRDzOY2PGPOQk1SC2bPkjYvxWR
egx2nwc5ihDay0zyhF1R3rm7RGJRssRrl/fsLU9vXM3WmHmwYc4kBSQqBu2+eGeDLz9dS9ct3ueR
CUGkcNGrMzjnhuR/ds3BUdHh724MYZjywRLjFZ3wl9Jo2zeNGevHAlVPJWDdrBEiECjIKiJM+PjR
x9cDv0P6A/ZdOeejQsduo/8JnSAKlaeqvWl6izCQTC89UUL3RIvXNvBLUmrCpuvtY7SMw0HFaLMX
9ukBS26K6U0Iv3/4NOx6d2xjc3iDuJ9EoqtJoHagFWH73YfDs3rUXgwWZTgToa+YKOFYh1NQz6I+
VzKJsRcuZ7AlrqFEsXhrS+grEYfFlwxJK8vwIjRDUwpKiXP+yZ3Hl5+1M0urNafEIZD8ods9m2XN
M6o2+0yVRiJN73C3WJ9cTHNU+tNSezneO57gHbwZCpI+EYjghMaioYcG1llPJU6XKBepGIoGV1B/
qXjDRVn3N9lEYlzQQ1a0aBR4jmXg0Mofg8pCOv0qjYJCMWDRCADvPbCesA7pUSeZnd/27v4KfIz3
EFSnDNHDi6sFwpPfGXESataFWEOkNz9I9buGHdszeUaP1Y+sCuZmL0OySph4YnygtsrReZfvFLyF
QSGsy0/nZ67T6pvmBLuaawGISMPtYg31zy3lUkza9F6sCefqxMfP0AM2pitDVzgEQoQK39PFFV8f
BoQKe32n6tU9EDK30Y884XjEmPhBJICNLoRsMA3pxjzn9AIK/5T7NkkcPmV/BbtZp0C4qpqGoTVb
TebZiesNihRawgBNZoFyWYkng2B7mUfQDpCUxywVFWheMuoLM3tdWCni8qzYzSFXK36o42NYLJIF
cIh5VdJf0k2s25Sw8e/rFRwWQDU7+lbvPVMLjTIVSP/cM3Pu+L1AIRd4N9lU1bHFrChSrdtXYbER
KyNB7uJxEJLUBnY3obCulT14LMNkX+A1oCqRffhQh1MVvS+bThfVb+VDAx1nzmaqcX8nZr059uz6
xz5B2jC7cwSIY6fwmAAo3Dm6K1TDUvG2naPT1/gN8ECfZRrNLGIQuvkiRs6ia12HDedjBUay8RKN
fJBrEh7E3W9BGaFYJc1A6daSjvQbnt+DypioQ/znjr9NrmUJ/3h5cyK7288/pVFkN8LFn/5TWyNj
1jRjaQ5e66CfQFNvhDsXPSRoKbehGTCv19TCnmZCK6T4GqU6IYg7xnz5TtwrfxTu2zGAdO8wEO74
zE4hFofjZsd/mBNpHcjY+0OYnFXd5MoBDl60O/rWnVKAQMPKn2qEpD64nWq9dB4/h/yazJNwg9g/
Ipw7yq5OaPtYfh3HgEXOOSvwAVLqV/4etcwqlZXm+e4qf6awwsGvdJ/J+YExqnkQ1jcJUhXuzFEE
XMsyIgrOQ2RnKbZJoRRBTQ3jqnINAKpgOzsMuc7Bpr/9GP+neNiNs1TxpcXUbCjSNQMFaqi4E9Hh
IFl1KQzVlC7BNM9p7c6JyfpcAR/hybfDo3zMzvZpw8iiuZ/mvOEH0OkZ9dT3iB2LUdBP6uPayAxG
u9q1ibJ/vQFMUKG2xopbhcYTe7FvfmlFHR+lyunOdORgzqFmKNWl/n3ajXUHdN5pRxOyTitdKWuU
LfShigd2o+9L4pPR+tb1rINCEKuRITtEkJQJf47vutmWKLjjJdTJ0gqw7fOGSJyy6HHs5yWZfO0v
ejz8h4lGA3m9ekT4QhEpliziIPqShwx/Q6Tazua3Z2AlcuEDbSE5hlmoHqB4ATkkpAzFYdS9R1Gn
1ulYf2HTc8f6AyBU96KKuJvDbcks0m+CiO7EaeNoRcz1BZyedpTanvEj4I3tnU4CMoYAWDrxaPV6
a8ENJGgLn6Xj2205oN8oaRLFIykYz5Kzx5Q=
`protect end_protected
