`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AwWbkafRpmUgr8V92aHEZ2sY97/tHJvETsM1hSGphQtxrQq/xYaEsMaIXwwIvNrsNqxAJaVsvRvn
JMezsz7KyA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hq7YGrjuSDXZDCwYl5lV4kV1UuWYLCUEpnqnkQMEJAIC682Z5TUa0P809XfzdZeZw1MaF4Vc1NTx
E6ECjowP8EjtZeAbczyq7rEitVSULP+P4HXfxdy1uBiRfy387pIjihUCPJo8F1EK6Pr18BnW4UFA
z5m5S+Zjb35YdVVlvZ0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J8z0ebrW8RdhwtS+c3+yPkwDpT9bxR90BFVWq4BuC7ZCtTRNs5gJ78QUtPbGYYc6lMHulIHX3Olk
Uk5QYrVS2ruhe0vDjJ8oAWj3jtIdRhE7qk5zNEwYcs7UqxZLtwhp+iVK5tkcsM8T/h2S6icKkUoU
4WL+LwFYG5AwBUW5aSkMRcejAOXf9e1BB0YZ7XaNi+Q06conYt4i5JKg++dFLNYJQfL9vQaFF8t4
JibkWrzEEOrlLoSR0jtqLvCaF8fNssW3ksYb/K3sqRCy6Q1uiBl2mFiZdbbfvufHl2+s9ozqn8KB
HzW8coY1ZgOdltmzg2pWNj6NHJFP9eRfVW9tTQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
djyuBIY5lgB9Uah20g7An2w3eBIDkloASAR/7QYa3ADm6slTzhRhNLKiMQbhYssniSYzEU0NpSS3
u7TRZQgLVqTBRl9WE019cm7QmiwOrZYXaKpoNl/O1nkiwyUY39dlYBPhtQx9t+neH5MAeuBRFnxg
kwXgCqZsJJw7WPq8dVM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GYo3RT7lBroRGVFGSAVwtqGNouH5bPbzrA3cFwK81BiaEmyyuWtTT2RJ2W+EAy3bVWR+pGUnEvSX
+fSQUpVwxaNVk4MhOz6vAEt0Xy9vBe54e7bOYB0bV5BnrKNIN3K10ipZSOSaImlVVQfNj8BQx0BO
ttkRmfedmZpVm+hWOLhtlW4L3bUeW86pm5MhoVtyWf3NOgGk1SO5bAkF761GXDhL0IrsoHAbT6DF
dQz0U22yj1f8bDS5bG2Sy3oxiHmYIZT3QNUvwx7rjUhlmZZIxF6mtpWUP83x9N6i9qf0uiloQ7z9
+7Y6KZ9G20JjYodcnBkWdgbus7Wp+iW57er5JA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4112)
`protect data_block
6gGn+h571+YsuilMHPBJbr73+Q6FWgUD5B1TM3cuivdUulxEdMqnG9Wpy/PpETE7slHiQIMRtv+0
/mgRZcxzg3xSxjPCIhEWQqzaM/IRFODjEVABeip5KK6cd4q8pbxlS+i85z6lA/zQonBc6sSif1dd
d4PNW5Jasn6A9kzHYbufQC6Q9lM2+DAAWTY8pB42ThtMzPEz4weaIomzy98EECmbQsI0rimWvFQH
YK74RGZcfPKcR/WZH4L4COC1AbP64+GtsJxH7/3K78+udbHK/gUaazya0pN956+h5dQfJeGGZNRB
k5h3y6L0YnQhdm4Qi8gKwnh8k6mUG+KUqNv1ilSa/hgPN/VRHKe47a39534rQ6Mkx1zkInPPdmcs
PtUF/IpWp4FGn8Qp2Eq8qScRFsFHRUaIXag1TMik8IDWCHKBaazWTZYpSDZgX4mPutgd4askcx5Q
ky4rvN9GGQfrlIGTREWBm1RxhuLxvOvbqhNQFhufsoPTFTXPfJv7cNYWnZZan+FB2dk4ryHKznGO
gvzue3XqNTQTSw+B/XfZC1owxcGXMqvh4FLv/uZ8gXv+N4RRyAoY5aYPlDmzRimkYWwrFM8c621n
fuJ6Byyrdbjuz6acIz5G1WpsNmFF1ITxG2AsfV+74qDcWt9g04flZ4tuikInk9xfUH9CS9Gj9oee
6AMwbYg7rkNsQ4xMIcV6jf4Fmov9BZyKwrDYaWQ6R4t31ETDzHSG0AceXwViNSzjRu6AeorzFm5c
0Di0S6jmiYn7RzqT+SntD+RriLTJl75AfnqcARgZPRbyjwuU1274AJKcAZmSHTVfduJ8lau5woFp
2Q0v3+A42MGwc1iXjkAqTg2c6/un0pUEyfGdIpXNv0Hu3kS3/rZt9AHtOYVii2rFAuB1GXagQ53I
/1Wp1H7QJ7bQqJRmGaSGyA1gg8NdFwg9CvGqWwTtE3rp+yDNv6bu5Ekwc0kDecx/WTC6ACOKRNZH
pkOU0pr9mfDns0HqSKbpmSOs2ny4nPWUwEt1euTXEPS618pitaa/t26S9l1RLGV+D3EZr4g+odzu
fWgl5Lo9J7ZXpldxyt7CteqDbjREsaPgqRWCpbHLBrgCi65UgzuiaFVDHEwBSLPmerdolHGaS9I8
2azHYYkXW9pph/XmgMUPQ//pOK3gm4gpjnWm/RaJDNcB0pHw5WZVa+aI52BM3xHYzEAL2b3ElhIn
LJS9gqU29t/Y2FXrdwxoG4X1MVMdTnYBQyZ5SXzZmTQWQmG01YUcCyTTpsIQyP3HW+ekuKHIj5/v
Nr3mpruey98UTyUz67dCDG5BqmPqTybXHdzPUlU7XMhDQOcltrz5D7p7lq0N1Z1Pw/hPA/vmsKVM
FFAxyQ1UhYNh5DI3gT794SK62uFgeJVWUfNzRUSexgVSQACps023pe8J7cHLBuhOlwn9MQ2CDtSx
u7xX5dPzayOzYx0dVxnfoAtHuobe/52EylxFLPYg4kW6I8okcXwhYSbfzkZU1ypKHzeX1ARjW19G
YUWIqXEaovGiHOf9YCHmUg0iuA/mOcZhwQaJz/iNEkukX75nXiSMbclC3zQQcrLVmbTioJrDpPXO
3/Wu7uwY3LMtx/WEq2RlcrPts3J0gpDB20OmyPnprG00byZLfyWw66wOaTq+T1vVq1SPgzrGpwnX
dXI+62ovEYBf3slre/2BbUtHeqUUCx+AcWYxkisuMgsDuyju0MoRWLYeTY/CHkiEAtWl6cVLpqOP
la+gK1iQCTZqcrta3wAAGssrjWTcHU7VzLpsbMCcO8U2y1yQEWF532f7OOuqa0hIJwbY/CAI8eq5
L5Kbkt2xxN5eH5ciSg7FxRFUzfJW6vRSrOCDI6JZ7D06L9zkrCNCy3Sg1Hqn9EyDnPOGXWonKx9j
2nSrp19CpkrIhp3ql154p41iVcePbh1dxxxdha1te2jjUhygfriqm85DKkfb8pQnkkQwosWoKJwE
roQss+J6LymbGgkDYyGj3a2l1UHKg7tWUkRzmq5lDuw9yqJdhR7tEc8yrH1ox6zLFIP+YmoEcQQZ
yal2gdkh5h5avU++pozGddPX6lQQXGD2ocN531alzDsAspxB1ZAXPjJzN/rUf0RMEEhmaeJO84V7
9PhHKTIPBy1Yr4w77XFaBSyly6Qcf8IBGDJawyy02Zy9ZvZoxqyR09OIuWENklyLHsSdEJzVFe0p
1HUPgBa4NeBG5pPt0Jc+M+eedCqei09/MReoLiNWJ31JbS940cWfFD3FI6OPfhM+umxHajOlm+oZ
LJyOv/6AtCH4zXxO6+oalNFF33Si3Ew+j4NOYxtVxu+jUY8sE1ylryjyvHzaBUaw63RZ9d73eVEs
qrM2tAIAS9XG6n4gwCvG9IMkDCs55X70omqoIAnZ4AdfovtSoU0Un5UaANAcycqujrnF/MWtmGgr
NpGJFh0XhHGT4fmHEnNWoLxwqfcK+2d6Xof58FQTnzlXok5o5l/UtpQG5WFWcMF56GiwbidAVeif
K/twAggsD1bkuza/lW74DFMmP0ffZ/2Z1Mm+OTtmJLcHESTVuumqnwaGJzJa79Bylhi/H2VCHhXe
evEpQPOOjHmkOJedTkvTEBztvOf/i7BH5KUSwfon3hgzVfPAJMDc0pbqUmPbhEbbYvzF6DeWY6Hc
K8usDf/e/rqbMbwwt7xlv/hszdMJ9DRcxng5ar4Yel184qmX5W9QXQ3MeDmARbJGKDWzzHkX3EDV
Z83he9RU0HKbwjlTrsJf1LWoPXcPPyUADnnTsQv85C7pyJ/XFtIVUqPbSpsNRsfVRyV2EngJuvsE
KuxsNcz5Hr0PawIzgtxmPuBrjpF7ZwQSidUlqdnRTWhobiR+Rel48yFkfgQX4ovIjkI3NB2+HaKv
sNYsC04wiRujHE1hiZptpzrdNjeKApWfgoh8JMU6HornWdYTWeJ+ABBz9PI01dXLaVWf5lW3InL0
LUIUPmV2MrBdsRq0OQoUfH5xRqCSbDikzsfE4CAhteDHQjusLs7X31E8Nu2QBdFwcK85I3+qry0o
uO+m2JrW11CzFGWCKgcXE50oYKsRgOoOTS+ndC7ZLMuJ0aYA2mjEo7MrP3FAqLyMbodrOLyqAzFy
mcvo4o7TzHqA742vb3hJT+jQKBcqNEYOL1OmW8m4q29SlRPcPKDSjY0nDymFRhZAc6lL71+7HVAm
O2GoZ2GmO7FI+bqa2HEZAvqaOMkXI/ywjYSAMRiRJ8rFnMHSdiD/23FPQJ0xeatSLfSMWU9ktrx/
JddGAay1QW9I9gCl/9gfR53siy0tLVU84IybK7PU0ByfL7mz/x6myWSJRCmrFqlBNrYAQS8BftNd
zIJn04TZZsPGusyn6WwwjsydqxVqAQchRiPlJN0Y1Oi7J+gmGZ4vfl4ZT+jnnWHHwOUJPTVkaJly
omC1uL7c+WjYGMqQQq2aShcje6Rg9+Vv+jurN2kPv9kvtXl2Le3vuzQhH+tIM/xJAiPa7ZZPnNdV
IzVImMHPBaiXFJHwFwIwHB6T/4pD4iF6C41xryBJa2aJwO7ZkS9joK/Vq8XtbcY4hCFQxRXYCH+K
fjAAi05t9wsTnTqtNMYzElKkwNczcInCDMpIioF3llSEzcof/AKQJH2bcBRJXFYdF6+CVebelYRs
6kJIDeRdSyWFQcaQU8lpho/KYk8kQ+UwGXFLC8GLLF3VVC+6XFoluv362dkIvslbdOkkY8nTuLom
fHlDgsTZk78sQaHyOb4C91+Fo396YYL25k2JV8SiC/bVdb5BFYQvnEf6uPb9E0Rd8G2evA2O9UVH
UPjSCPokP9jAuRVLgd6O6lZKBcyAIoM1Bjn59AywXxo4jIhk11ENccEu9XpugUcOH78g3WgtvvBS
Mv1z/4FmDAgWBzW4nxiwgS0QHM9pttdjeya9fCUcT9p9AkqNyXv3HuxmKVmLKd1KihK1xFxOuoiF
OXfd1mYK7b+AT7wDp77pAM585ZlIdY97O+YgFxBz/vs88xD/wWKp/lqdCOWk0a9eeigXUtWVsY7q
oIyqeJHuCxSUrznjX0KWGjl5QjaQkjK5i3xcGHcGKXm38hkwEFkOAEmhbCGbEQzwHGfD1WIYh0hE
W7ai96GcAvr0BUU72XCum1U1J32L/ch7BfGVGEtYXuPbGlY31MXx4yxK75e6NR4HnHB4InZaYrEn
TzIGYIP7QDQnDoZ0TjUsQpskUzVUHDuGW3bj0adV/0QYEbGd+HIOGsB6NnkjQ2ZiRpPbLZi9VsQc
8IUFLTApzlZovXY2GrGUKQdXtqRbNPWCTSi8hfcFAmAb1qIq4C2k4iZy0ntkjcELUVK/3C6KiXgt
/t/dziZkmIfiYGHXGUsCxhK6K/E2k3CLE7WFHN8R1yj7+s9H5EdBbKeuNhaM1nrmxo5a8Mc5xmCi
Sfu3vySMTfP1zKHbXjAv/5fjGJk/olR7KAZvYOkF5rHiLHWDTZBR58oRYsqHAeNkQQJrsH1LpsA6
paSvrNAbHIQOTvsQcm/z14QDpolPPNOuNm2YLnEA0lId2KMsV9H66fATCzA2fITFAYSU+/CczsyY
87F6l+quK9VqwSJSHFgEkVGz3nR4H7D+j29AZBvq4IgAGrkvY1KR1QoP/wNPhpZYIWxn/ojemlqh
C6S3K+HI1M+G+tXJ1iG0G2rDtPq6CW3Gz57q0X6lu+7GFpGL+DAsmiLCFng2+O6ki6WOD7KbpOy5
vRqNE3QJIAmLrsiQ28Mppdf5Aos/ydrvZnvfUoojKQcsO1pCIJSxQREz40pEWoFr518D6lUwj3rw
oQjzdiE8Ksi5mtVLAR6eXmlUn3gS4BSO6WhelegI0U/Yx6Dfjxfyso2COr8vKfLrzj082OHyzBZL
FcH1rsU7hzbpIXpbeQ9XZ62ZA38spjibk8uGyKqMrE5N3Y0VDYjNZMHHx9KWXZ2gtWN+81UnULfO
WO2WXfDCUFa4W2NMwPSkup/WuYfeRYyG2lb8iKWHir+PRuLM3+0dle2s5FX6k2uPbDCy9e7zlMnH
DLeeS2crb6h7ATxr0yf+FWno2/H+1tAau5hfaETKoC1VR3geuE0KuNtO6DzIaGL/HB37++KYh5AL
332L1qCOMil8Xihru4PWZ67fvI3b96G1VWALYtLdOno/olJpIBY/gdZws4/RDJUi0CAUcAk+KTgd
t1oUJk+mprcZ7ecQXKOs5DWjiE4caZHQgpswgHszz+eHs0P4jcjt1YsfMUUOAEkKTg/dmfle5H1R
/PvWH5+a+QFep+6Dr1+a7pJyuNI+bkWNmZk+p0Kvoai0AbTHmRc79HFwvMLumB8zgf04ZNEXPNG9
Xmw4Rtfc2x8uL4yONhYgxWV+aN9yMZu6R4pfFLi2Tf+RoCj+zqugu2zCcc5lghBWN+Uu3OO8x6KT
caNc+Lh5IyhYdy+lIVwJahcJcLM/8GFvK/3nraIn423NNKrQrsQIDXw77AtXjhbgpYkcbg4kZmLq
qJF4xrapXmY=
`protect end_protected
