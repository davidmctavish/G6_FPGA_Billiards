`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ijw7mPXRT1pNoLg2oZU/N1EGzVifLbU9Cdn5uq+lr5L4PRcM4ABxEl30L70XZTF9k00TvnkF/u2d
Zt7NqyvlCw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EnBPR1CJ+sKXHJQOWPpfUePtXRmoggIjQ+IqYHROTJFHS4eUt1oER1RJukmaXVw7jLTuRUPrPLhu
GY8TCXkJ3zcT1Fa9G8LSDdU30Dz5CZVYWTf4ovjsihy77YiML1+pjuOPzvLe6MRIa9zPGvKkO7Tk
/cwFVpYlJSoUy1a2eT4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VHlBH82gZ4PaxcOQ9hdpymWj9HfxT4Ke1K+CiiLK0AS8i81nLkkkoqf6+VHeFR9ggzaheL1du81L
kxAvyL1QZoBooaZ2sOpjGOzgB0aNxVkhUbsiTEYUSDMQWWdjCiC2BSSogcGDhBvqMsI0b8eTfrTr
xwgD8mjq/8y5PJ3i/T7nECkXZ+dmRABy+LW6uxW8MXb1POFZNweuT5k7xL3BCk7/spD2KYxz0efX
62Tg5vrThJ8xrNvYplPhEDELRoV6rTxP1MO/+cjNkz+0a3gmKrlbLHqPu6WX2Z0ciGsSDC0Cywsk
RAO/mh1O9NrO7KUs8Vihu6t3ayCJBpx91dVw6Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1BIwRXmQ1SbYxYIxh3JZQie89DbZ9Eu43SQR1cngSAFAumtiqByMxsH3sJrChTtiTEFFxTo3Y35I
LGJOJgpl2BW8QU7hpA8uzVbC90t6tnuF1cf9w4Zx3JuVfbew5nMjY+rvdYadfQjUIfRwngxNVRXZ
xv9IEghiZbHmaps9PV0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lNJNjzPBDfPgGc+GwkA+4WmP+sjpdMoDH/HyI9njK/3GSo75c4vODsrKwhlQ91OyQEhqIWv0Kjac
l4KoBqFdFLRDorgTOJS6MMeyiQAuIPZBvNzYPax03sTAKMdvo+2Mmk79TYs/KzU7RoKgsHVRLJsX
4S2Coup21syqJfaLjEwhEWw9tSfIGg54DmONp60H0c55UxrRnERgVrEuOxEQDs4rJNo1aoeegOAQ
NAAK42TE/37PY/zybZevXypTcxKUcWPx8OtjIuPCDgam4FFEp2f916bBxj0AF070/6enmwZleDao
MRuZCcDhbvojq3Mq2lOmP6KbKYahIKTZ+9iRyw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12384)
`protect data_block
9R/da79AQvgUhcscWvOrmx4uUKYbtCFEOXBRTI1Zaz2BALWARzFPGzGwFwrxUYZ1njn/PFCb0BL+
HcXW51nXAIRlJaR3knFGjvooko3oANYuAyy6DTNn7AtCsTLN8BR6+8p+YA0yf69YZPIb53cLJvud
y6Fu1L5zhWWLGrAFolO0LbnM2XqPGpHZaSJwcBcDiK6cXg6xzkDe2doAje12lOMyPfdoZkLUHHTn
fuYKAPqamQXLKGAGhHilgryoe2QVR0HLmtnRVot/+MKzYSrd0fIUOZ4MyevedOz8ONU8WK9guaZH
P6EHHSYA2wLWgA8xm1eDtRLWckpMuABkrVVA46JflR35C/E8sr0qplmKg8dcpm0pniwL3T7Q/5SH
ePBhZCS9SfKeTRp6hOz7DjOBeOv9gwqFdGSlrvpsyhVYw9N4VwCo7kccHwJJomfYXIQoHEXXBGmo
6PGehGjw+vFKQNvvk8aR9xrWn5OFK4a9QpKvj82YuhzzF1rrFV5C472MCA2VRXqANQfJ4l+ME9Gg
dwwMOpBHKkJJ+Ix9a2ZPGe2Twsx64Bth0m8XwDWzhWjKdQL67046Rgw5zGvcbihtPF1SrgMxTIGf
fN4rdrHOQGGvWsuPPKpZAZPmeckflppxy6tRnHi/bp4YqAfafzUzVoFM8gs/afVOt7UYXkdXa0J1
xcyf3iPsHKM90NSue7ThJViTzHmYOQlTTnh/aP9fB0FtqqfVbgafKCYJiq2+mdXezWzDrdYA/O2U
5oGItQ5yq2Zg0HkvNeK6b9jDbghlfFlIMimVeJgx0TOpw1ZOuFVwHsp/t0Pb4fSyFQiBCbutseBk
DiAdWSkNWq0XVNQp+GUtaJDKIBMfFr2wQrd+WTrsLlmFRgqXdc8F06EKjwaO9po4xX2LqMZm89Xb
YHGWHthSebWz2/ea2+8CNaP5c5CUwQmbmboi+KFEEtncsMAnYf8SMm4MmLDdUisQXnLFt/F+IGZI
Lo3aIZF7cJZy/nzbkH+VeJdKwDx5UTCzJWsu1et5sGFdlQFWH5P3aItd0XgD0yt3FDV8srPc8QvT
jYMkPCnaOkt/7HXUld2j8JmBkI4z4soQQFlp6SwbpjY7nbVik0VXbjXkmPWip5qzxdNrDmTWocYQ
3fKShcbNR4kBqAmfGN2cb0AVTv28cyqIcNwfWKAB4iybXme/95ZznTyVi/f/SayLDgGS6CFyln5H
OnUb2s4PBumrmC0w17wPryb2yj60+Nij4soVc9AZQNv5m8BotF4BKud2GZ7Z0YqCBY0QHDhYENL9
6XgHw4hH6ab13PEWCtZf0KI1T9j1um+i+XFDgJMTYDyWNDUaQFpg6XKD7QqHZ1Q6V0z/TSTP8t/m
JAR0YMU3/8UIe4CESpsYf7TeaB2veTFpJMAbd5bMjkOo4l3d1OuNwG8ouiSRME6G5hp4WmTXvFUH
zV9fLuxwXhybhN9RqVBuRhu4zVPHKBc8MiEYFix7s5CrKiwV+prjQrZTQvn+mzz+vmcb+QEpnp88
954/gK/G4SpZjp4LVhQZwGOONmo+caLF0HZXg1BkEuSbHoRP4xD6UDc1fN4Ox4FWd3EHs91SNRNn
7PyK2jpu+ZQLeIMAYpw1f3Mnw09IF7mjT3pElewQEZmQGxAx4UornUt650w/iUoQqY+RB5vTTnGX
eDgxlVEG1MydEo4kvfr8301AUdngm+Vpgy5dmRvzWl7VucvrKKVH+fosl+4kgXYJg2wRpVqVv0Su
V/r7nzTF+TDDT/sID6WQGEz1BP6RaIhki1OkP/UZgg0yIVogC0vTWK8XLV/Bq13GlAenSUbfIA0V
3EzpOjei+un7ki4qVmo1mKtP+Fykchw0o3ON/wkQxPAdtVOrQ/4SMyJ73/a0eRur0MBNODUGpaT5
OtzlMWNxUloNRnyTnPCBkpnDA8ydkAEEoIF49ey2978tu41KGJKYJ78nWQteIWGTR5NGbXi9Y8/e
aylMGrUfxNwOLVIzygaImfVkmUF11IbSXGOSzcZY9ZISUQJA+xi3hiouYMEGxJjn/FT+mBKY9YtQ
icq5pkk8kQzyhzNj4mKFIIO9RF9SdmoYlwdU5DHW8yKBEMiiKmA+dlc0/tsbr6fX+xHvyGHfx9TJ
0B7kvNRgdMM4iUcu5TqmKB+NBZqgb+FR/Xs93unVX1Lsz+gk149ic+JK38xs2XmmyZ1We3khMZHB
yl68Tuj7wt+vhI4Jxmfxm5lEF/OzPAo1GFx3pI6IJTVtT/Onom0ZlrNDJuVC/qt90M/0qBVdv9Nt
oMdUYLHhrY4e/tgMMRJ5IDHeYl6vmS9FNoRePWCyun/ZnPHDSfN+TVc9l8YRNP4+cFBsBdkjKovm
iPblhZ2x0duKBfPwZD2arXuFgbg1g3el/cB8H2xlEZw050EtV6oNXx7NB0a4ekYqO7652VevGGmK
Uc3Yrg7/2OPGqiKnautDEFl+m3V6cc8M0zOXFsDURp6r0araGsDuFJ043/4PkfEVpikFwC0xu4yr
XK0FkE781JTDyciZBANwTGj9Dwi+MXGfRyKg9uxRozFcRwWnNsh8fVYBtdzrUU/gCN1ce0PVFCOG
Qn1suXf99vFMg91Obl1YYlPMx0edlbqjRIBR9HELmmCHONe9A7zOl4FjHEzaen0Z7c6wgwmzuoA0
aNbOoM+KXJDCjETk09CCUzv2EKm1SilkoV1luhPX0Yh8gwzHRklisMtyQNFyzGdeqrd+nXuqDhBg
EEyQMTxgg4wOycLbiCh+7lzk1qz8CycZ7QbhujfXWlsXpXx+2an1ULyrABqMcwResWAAfmiVQoOu
RtzLcUbpHb/QiexQaXHMzqMk77mL917VUviDFZ2ci6DRf7qirqCsJtdFdGeNDKS5KwLjOjEQmlt9
uxK7BN/Pv7Fqq3r36ryoo/X/hnScDKgDHFD0Nhu0tpjLMh6zB4opjCdvW6MmBVYHQa4DQss0f+Bd
TscOqDMqpoXjNbXqaYJ95mlQLQAZaWGoiEHOzotF7oaTEY/h/OmTckpzhTM/sD+mr03ABAOB5VhR
RMGQwT9m0jd2iwOCTubbA+dxdYRYO61CXH/fli5tfYX7xLGkePUkrzVHUuWjnF2xW51OcU8Tx/4Y
PPFlHIMjw954azqoonlu0WRj7jXdadV0QcSfjjrHuwlg6HMwNTc+LnVhIPWhPDev+tjjQS1q5Uqo
azfQmJgK8B8TklIskvdRDrC1bChiagl04+a5Npgp+O60nWZ43VPCZv+ULjCu6xlcBXlQbdW/HB8a
asRTU+RISBUK3iRVCF5FAjFiWhehRYtrzt73yGEz+Dyh5DnN2YdpwtsKaIINItF4DCAe1qHfvW43
WPaQcFe5/DEXt1Dy/Ak25hyjPt98QTRbVelETu6J99GM3F/ebaUfTamrUV8QnwiCXwuFb1rHJNS2
BzQ52mfD3RD6FjjR73Z6EWuhoGHxnByP8ks8G3yTjrzd9+UQZ58wphV71IxgmeQJcKUJkOtm9kA2
pSkFclpOoUSEJ4okR8PN+Yit1vujl3DXS5yX7rsl+AjRLkjeScW+3n0O/zqlQw6UHrUqXtif1tOU
DfKKPEl64suGQfG2b9NDNWsxJpN+P32rTdmNoqmueLuLvTpZCwJdy5DqyAuGpv500b0kzTZdzq4+
iBAsdMFTPqaK6RNXl72OPD9XmI3tErywpVv7Pq4sQ9DOyG4SHAxDBgMaE3If6dRjeynJSZFE9gRW
O+zROo6IEYjGF68+r3KOaPhty8FS1W3GNU4ImHaOh1uJoIFBtV1W0STBLkYgJd60Ip04XOlW8U7a
XID+ELLF59+uXCiA1jtlSmvlb7HwoWaqhL8lBz+waKDwBihMZ9+5PIVzO33vvN2LIAv89yK/1yuj
1NvwBLk0SFqJ/vaRhTeieGKPHc23GxOw6Xxt7XTzRENuPbke+YaRiSL7vUPX0QD6FkCLz40TcHU5
VJJu/UX7C19D/Wv58R34aleWvftKnKFkHi1VwXE3/T6n1nflD1KclLyiB0NrLwxzOLCXZPopkw8d
bYRMm4AuSrq1qYo96sUvqZR5dCCaZ9mZ++3iIyVA4PrWjXEoApTUnePBixK4va6dpBC5CZlA9lVj
kadZVEqfnotc42kp3tgLATW0FhuFaurA5OuzlUgG+aF/PLmMTs1WPAJ2xky78SfIfC7/JZsF5F2z
5eiQf7hkAKG16NgR2AwOQ0INh6OfMPc8d7rU6ZsUd+DiGbqy2JQW1DotSWJj98e3KJeV9Dftov/d
mqj5T5hyiBnZpvvVKyvXiTGRgoJCXU35UwqMR/zxJM/YAYmjHSxG1cCOy+Mp10KrvQkRdSbxRJML
0nIXiNh9PKhALJH8iPJ5cstLJbI2pkGC23lbovu8y/kg8tXUYonORpBWBsEs1fsApVT5aZ+QSx7F
8TTEf7Ra1TbCeB3qunIugzmn9UikKOWwW5YCf2m+XWaFNaTo5I/S5TMqiVjKH/HE7w/+HZrU5Ydf
01WcfP9f59b92JoRGtSFhtTSHujbnmvA+qaR71hPQBgzIPmb6Fc3N3sNbSJoRm70qOCxu8pHMj5p
ULnvvj2K/5xZ9b+TkUe4Hv2g1tKOMEPZkytj8WYWLIJ64BCUIGzoyPWYvjBczLz2Cx93CRo5LFhD
JRZcmZI25GtNdnPVq+tp5HPdxjJj2ZdZEihFZ5irImAPEwkBZBSxXDIBQV7fIN4LQ++LFq3Ti1Wj
9z0cAdKjaKa2Ujhtruj2vcZx0uH7eOuU2qOzfRx9p6agD9x+/sPNEP90ix3D3qKRx7F0v3KN7WUd
tafrsoSLsccBT5dN3sMs4Ff+jhcSBy6MhE+kGxIn8LW9/VHTBXTbVBGdUabzXrOAcqUNDPTE1V8s
0u67YKK4KBbSaGckR3Vwa2BJcqiyG7s04b/EIYZe2npyujLUfpY3GAWmeZqRaNufKgGJZZnk0aKH
kFsetKP6+DzUm5Gl9H6w/vOY8FF8cji61oKzdmZEdmULX9GfB1cLaw5g9kUX6hYdUZ1TjDXs2Xq6
jI6/f8K9zPOhW/fHDEbgmynudM4QMvJPUVyCHRL8VGgQ6dEpFtIBZrU6JeBGJq6QDNiqdjbbJsoN
uXihWAsZ8m7ICMLIzLmrKK3fuWZL7ZL7juOg1748kuMqdizZn6+qi4LMDvCfsviq3duzOFTjW/lw
sv5SmYcqRmNu/ZFRCIjfPqFvfA15zzeDWzaYm6qiCjlgpacAC3sOoYPedToEsaQninNxN4ZNaAGi
p6z3KWhgN5IKrQ+XaDaEaPvB7bLMyLiuMJFfDFIrvux56xEibW+vZXp7BYBozDvg8OsITp3z7EAy
J1iGOoG8qBF/sIDqQZ7tnYPyH30cuNuV5snvXUj6KFKz/eCol/6w60Q/K1Bus2aVHCGbLLTBqpM4
ArOrMFMypgaAgEKG+OGXDTppqd39NK+ByZCwl9WI81sJFepDDtZ7RqlvdsFXNV0jrkiCLefOqFX0
pvl++nd6aTupRLu6GHuOxHjouMfg0VGDlPN+DU9z6svqPLlXPUQKYwXwMX8cIBmNRg+6TSE8nKGa
lx5eIuNxHC+ajzjJerxKifDrkPf8Nf3PGUP0h2ZNSq3bUn4mGxh3KKpRybk8rSoHO16GZLmp7DOY
iMxUihBXff157D+KGub3Z8ZRPBqSPu0OvshP736P8iZtK6HK+PrrcVeW3R91dC+xgXkfx5jIDVrt
qTsaEv07DLkKrO5VFgP0GBTAcyVgq2ZYAeLwhuVVdBP4YnVHTOh+C3HXn0hQw1VuPM9wDy9pJn+Z
PA+Mtwp+MLGfZjT4DADeFyVjWsK+HplfeXbdsc5oxS37Ny593g5IqOtkDD1AZjmkL1JivDwRieS5
ctW9jR9zT/Rdr7d9q356tZuIoZClJsWnUYaZT57i6CQfaNs1lJyJ6PYD/xq7IM/4IFry+9URu4Xl
j+f6ouKkXA6nHokqiIDI9aso3AF+1j3+fZfZQfE8WJWVSbchYqSdvSSliCHANmCBmmqxolI5aHjL
q5snmSv2aEQSSIOfLLbNwFBoLRFcI3oBR61ekIB2cwx0ztFLBQ1fy/hwFtYz8L0pGGXQl9//LeIQ
2y7jWT0q+dcGmRlyZ3F7QrC/h60uFXWQzH1GH39DTQjTfTh2fkLzkJXdPqT21d8ath+HM1Qk0+2A
hb3fH1QM4sU7/x8O/MvRhY3g5XlYnu5vd9uYU9aVs0ivojxK0zwrQNG5qm69xaLEY7KkOc3FJPYY
YvJIEw8t7+lA4Z2QFx748syqVzSlkyB+/cwFMeliMIXMEBSKIh8y+0xgoqsDdIgWufd76EUcktgt
HsZ1YD3CnaYUGMAv3TFmdhRXaB3vm3MxL82OPX7SHfJkMVGW9JcG+l2TUEGV9156KYGTe0cj5wwm
cWXJ33P+2CNLzA+NFSumwRC/y1V/zZpW5n1LGIJBgGMIJSCzob9Fj1z31jCWsKYCtT/l2ZbqRSVg
xJPvAZgayQbF2aAlMkhzpGmeI/OvlQyCPB9b+TSrJ7BFKjjokwzkX+WHpX54BcB77W/H1VU+cSDv
xUFLeZFGpGbrif7r3X93MK3Pv8TgKny35LOG2jJYJIjD9Fk2jua38mo/w1uJHxHhxQDFVKAG7gMc
07hv6nJS6cx5Nda5s1bd17DIoLl7rhDfMCLfN6B0cf4iUcTRecZpVCWOu8IOHd7xrKdM69bcKifZ
QioM5Hx1eXr1yUsTLtWgdoQbLVsteK8iz3/TIt0IJfWxVcNxan1YwhUF/iFzOCZwRV84FAJEgpaq
lMQNPnBMV8Wuy7xjurcvX4mGIvMyOSR+X6FeP0jouLnSGPR1yiOc5068HS/tuMXVEFOtYsMnNW+l
EHHnHfxGtHWvHH7MMYFmkr8xSyM61LPgdbWNowVXH3bY0TIxxUCp8ekEF4Y9AG3QsDK5HsKfLVV+
js51gqlV9glMSPRs8P7zioiTolbxj4tAx4eOyOp6svoPy9uJQDFQusSjOacGkwC8U+8X9Itbg9Do
U9rFSwuKyImhrUT91CzQaRSZ9MFeIhwB7ZQIZ1Jss5IzCRWZz1mSZd8qdb8s79UXKAx1+c6PJYRS
USIga00egjEsJVxbQptU61qAkO32pBaxqDtsOhKEAmWI7rdcmEBnbwBgk28PL8RW3QQTXPHjD6CX
/6nijiGS0sk467yGnvBgwCPdHHa8R0bU/GqDpvymdYwBX7wLuaNjLTDVNL8/JYUs99VbJlKA3IMP
3Ras2yA+GXHPzV9XUO9qoBUQ10g9IY0IQy+T1BzYXS7HhDf9sJrTS2ZU3RxV+SYKI23pvyjpg5bt
34KS+EgyCLdxo58112LuRswy+QT53e0VVZBmw8PD+XMOt8J+SFrogzu4R8ZyyG92zupwTn1ddHte
Ns7ezI1hRHiYT5RnXvQcwKphT79sfRZmidAn6zXUjrwp5+90NfC3jcvfq+ReRIuW2+ixJNA1NQe/
1DnpnVYup+tWxp1X4IDKLmIO9V5SSIfyB3ydzzg82AFOwQJItXVVGnwEAgOi5ojBDuWSP0EV2gw2
4+CLslaDEXXy8ZXwPTbCgMGTMKmovgVVbdbC5ubX7Qb4aTwWcDO1BHJSNKQwqBrmhjgOCvsC6jzG
J+fQZAuj53CtSDOfrX0VpHICeDdH6278t+bP9xhYGw7gYzhb61kz2m6P0M352WkRxQM9nNddANMG
s5DumRmBIr2QAj7BoFUBPV/QK0UmbDNd5TvRJHeiwG1bKi/rdSNnxrrT8RFsZj/IxajeBz9FxT1w
5IRqjR5HRYnGOmXzNdPy1569QGWKzWSBxRC4BRPQC9esGH8CZdfRMVxkV55PCDfuDZT0UEmPHwjY
AHhyrMxBHPaENM0eTYDmbfy41ACxl8ZFYM12Jgs6iZOn8Ronue2CKnhUBPmsw8AuFx6ezewFRiud
Ef2jKr0ZjbdEEvlkMa3YOP1aJiY0SYxtU830H0bIq2cpevUmb3fUqXGR5zgsqG/wX+xpz2UNffVD
liBbM1+keSUlsR9v82VIArDTDOAvPpCyUsG39L9Wvy24lToiQSxCfUJrfd4IQ4PtW+WgREEEoQfV
4PMgCfk/CTUp3vfGoKvAgIr4O2ynSWl5nqucz1ZCH+VcSbIjEib25/DDMQnuQuwcAhr3gyfH0vlK
xUb/NZbYPz2djAGITHbeKFHyZ5BMGMWVUby+TzRk6E/B8aRmujOJ0wTpxwuEIrEgJtCv0OlVgjvl
Ue6895OPg7gGJnnxFOE5Lxd1/2EOYXizqqoteg16d983JOIBoiIJxLsO2a4gVoAv9rf35xf6kpP2
qyhWy4zsaDq7YXGwWwcy23Hh/2aj9KOBep9TTlKAaqz5bH9oyuodG5OQ6NmT586A7HFmTk/NLHiy
unDF0l6HlZkfuFQG99+gQxOigmUSyTOxBeydim8Xhrbz4fC1ifcD+1gc070yfDZg6CvI/q+9Ben5
pl3LHsVAUr2jaB6v8CatZQ3Lbw1jOzlIJlL4HKfmYKaofD8cShjbO6HIHqJKOPREZ192MmPDG/Hr
FlNcOkQaoNg+Qb1vLi8aASFbbiGUp2Q1lQ/GMbi9nBDO/H5yeieYPhdo5SKFuuxBCL3HO1vgzw05
mb7QGIEBbQ4zNP/nrAZIZLnzqY5Na6TVXtLz9hCnI471FF7NIRhQkqgJjrMjY9s2PtSXJxRDO9Ka
p/YzrJsry1cJaVpC1wPGj1UPtrAcK0jY35ibgG16A9mw0O+U8nW0XjOBtt/qZugcAvBp9O/wWkUN
Z23y23VBWQmg930aXQ6D9kx4sR6SFdcrHhF6iDztNywZp6TSsiBdXjkqicWDFqJ9OI1Gy4IsUe4A
aENVFCUPBmwCAJmJ61gJl0U0O0LOw7QMsyJHlXppRpqc9NCN5W67FGmrKXIHIcOdsbCMiYXVCyIo
4iElkoYroexuweeYHZqXcGo3Ptu6+eaMf7/bCyJUeEi2ubnYOUl6DL9iCGuFm4m//9qjb1DIj2P0
ciCresygCyCaq3wxMIpozfBf1/D4ez5CcDPGNWtns31r5c2ZepRgIyY41ZJs9+9RgcuL6jrdWYN3
e9VuJxM1OsAE34gEjhxLWfCM5qyy6s53pp/eWBMpMzf9E9qryFAqY+9f+ie2r63y2e6Vc0P9Ynng
uPzP+FwlMNLSkjcChm15IdP6F3ONN5Pk2d8yytn5YgXs4A8f1YPoAeBtDb9W7ZIPj34mSrrOY0Pd
k9qBtp3dRJtum/8dUiS30fAHRzR+3syufJnECBHoU79mj+1bjdglCEJP16Trjg4754Nm5uRzOrfR
KpWDyNUKpTq1Wktn9UbF1bLLpaMx++QFp87qAPVowSeuKb5q9gkdrQHcjl9k4ysFXP9sp29yH1R9
72Ry/wqxq7pnaQNxkQCjwqOH9vH95yeqA/VQZMdSxWhN4aIDvsX1/w6UzQaUW5T38yjNvTMcknQQ
hpCCHhEGVgAhIIYeojWxqTSyiqOQQrH7YHUvpkJ9/FAh63H8mXNgT6ivdfiahEjxbHZ8CYHcEnnl
Kerp910jgQxbijX1wZdWPE5LS3EWzRcZuoPg9LPrTw8x6bU9mu225fq1EcykLj9FQOshMOIJBF4B
RyTPvgEVCmFsgKU3ZuG/o6qXDrXJGdHYcSguZMSM/5QuKvuUgvenGXI10MxF8vpwrWBSWX7MgKse
Sx+bUN4DlEeMk2RC9VXwHE5MbbwjsMr6O4gz9M9iVwoCdwkKe7CFPIrvS05HPCeKtN4KWpnpzihW
Tq+6f4gAiwst78ToCYl7wY3l1DMx6DfHf7vgp+kIrsWmAaZGKJGeq+J9P6H9MdYcxT/8THnjs0DP
U7D7oGSaBiSCWfmn18KJouOKPuru4A0+Bxcjs3caLdwAexlsRyQb8S9MI4aF08CFLg4rF7GpPdfx
HxiH1R8oG8iKZ8Pkq0hfV58Xl9JnoB+ZBTrSx6q4n+LTN2gCYK+WuTZZSKI8WCJSn962WSz77AkQ
ZdOMtJxLhS6+FU9XhOLoE/P9/kWISHzi3xTaD49y4tjXNDb/afEBNW/u2jYzPsJDHWKv+vc4+0AH
K141LIqECettkULN0cVKQ/Bs8aWm/hsUGp67u8EkdzbWm0Am2yWlc8d16VxVqn+dE3zK/TvWUOBl
yrD6IKmHmx5o5gxmv3tyHy51kS8SBWd3KytMJz6T2zhNAosGfHBfuAc/gwgMAuXh9pb+Mkn5HOHt
sDn3ESuBJinr9///Twt9jo0YtPlTLhlNbrrBdBoov0gMXMawmusQz6byazSKfaBHt+0A5EhH1+Hb
CTKztnr+tKcmgOJCGCBnfEXU3zQMvlrJvj5posIOYuOUIjvLJXdDHBdiyt6iE9dfFb8njdKoO5R/
e1N5VOPivyInkDHHQyR7rSPfssnn+TtxLRTdNTp7DM6I11bW8YaI4K8JdYBN1NWqY8lzMYW63cr3
Wkl3MPoeUQrTHS0K54td6HUHxXMU1Vay3/ylNxzZxGcivGfhLRHYgqaEhNKM5SQaBvoJ103ztC6O
SaZYS5Bxl6w5evjBul+kjqcI0Df3/94vvau9+EnBm91LSTwzOr62ls13t4GBB9bF2W0DvK5cTFcq
KwtwH+FtObAdZc1Y4+rus7fUkHSFSSIzC7Qy7qTkcmFz3VqoIK06bN/VJr1sxsT8FmaB/bet9cjK
jRkzJ7fVcYpCZZy6c3ELwfk7C75NPJJbbfv4Nx0V7zzqpZ6yEGchAL/uBZao6yY89o9Zif3qAhpb
tkz11oSFrseG2aCdFyGIuyILqIyRcnitqtAAHSubV34Qj5luDxKQfEHUUKQggV76sVoYo6Kx70Wn
LTUEGJ36NB8JTZXts1j9jTlny1AeB+xkhNUbEfKLRXtKXdOU6dvRbvgqFhfa94RfSDxU6bqRCkLs
vEcpsZ35/1h2IAawsnXYHIy96lpKfo1pc39/9RwjmocjMaCVx1oyLzMFgWq2PbWeTO+oMKrCbbyV
4xy/B3eY5grxK97U6XQgBO7S3i2kc4wQxBpqiTo+fR1ICqIWxXcrWowhpunAXn7TIahDYYd9ZB8a
4DW+t1jU6wgd6hNYS36X5M98DSuCL6utn7iXUJrsz6ddQS9YyD+d2QZ9MVu/dX4DSJ1fY8vNa4Qq
T1Go9BiwU6c4G++JzBC2FyehaO4xcog/mwe0P/FkM3pKd1LgRMrveJSlA8NIRQZiH3ryYparfLwd
RBssSoQFSvrVmPMe715nPJyDjMuuAf1azQ4mJcjB7lSluLeDFqIEboAT1LC7jVJC9jwIva2UXxxk
cVRJKpTooDu4MFfNbcmRDBytgRaxVBGsnyF68KlnYNpxaXUE9oMVh9bKwbaLeeJIeCiA78QBYuPf
28gqo0vtIrK2le1iu9kR3R6uwoCFt9qc0iuVmYYM0Tf/OQtOCoydVLXcLE/Ds2knLfEGChM6Eyxt
i0nGMQr8TVvYLLVTuoLYoJ26cUwLBu5MTUAuPIikAnatOFc0/BcyqQwKXq6ov5hSTq1nOkLl4CXs
4Ue1LySdQzYviL73UT1K1ByeNAvX5JgV0QmdQEdQkSSVBwVz17Lw6BNsRLkzz8uAj2m4vA/FW5W2
foVU/MHN73J7hJ5aMi9xVUfrXHfr/YUoxjUCgfFG/WQ8qhUmypE81TTJDD/UERAxpIuvrknxw2/r
LdwesF28NMy/CAvhSgYtu21QcjvzJTlcGvuITcSdMjTktVDu6Bzwfg5IUmH5lU4T/nWmC34WtlyE
/fi8dJhZA7CaRy6rYjFCOl4AooWtWKeyGIlPJw2uPxB0eVJRZNZDXQIozzkRlC9CdeMKThPH5O1r
myQ+5uEm4cCGfqASM1nBKW/semTxgjj6UPG+6Edv+gWRlapTpnVTjkrxwMGL/EBO38keq9q0W51O
LN2mCrviu4CQGDbMrF/sIue+S5/tAcu5hB1WD4+unWxei/sB7b6NzjI1UB3xjyvGDnnSBqvndnd2
XJIv43GBm1sAJPfPQvkcuVcMjMmoQ6BgrJpaApfw2ToG1V6rhTOxcq60rxCIhR1SdzzLsO1CoIJO
oUC8zSl9hnfXKkgaNQ+NCNSyoWvuLCJjXdJNX6bHg12aGpAsGLLK3bRuZrrAwGzpR8ok5KRQ0+ic
wgnwDOG8vvVXrPkAqoGQokoPtLdTwdtlBMaGalE4GiijzxarWT4i8nf1G6pg7CNhE2jL7g9bYH0U
xtxO3Chkpae3YQCOocXt9dqOrTgGpNcbLPniQfAljcOf5y4IpcrNDB6036EX3IQBBVJrVK+JKvtb
uWNvdN3ThenJDPNkmW2EcJDoipXi8LzAL2bpO25OlTk9hbicz4I4yKv5KxufWqgUBQTEEsw4ngqW
3+yOlqRBeOyjNKJcL55p6BQd/jV4+nb4OGO9bfMhq5c73ELmK9C2fyG/BHrhKJP3FRyv4mrOEdER
4aIC7/PprD41BlS2NMqa9FAFYmQIlAE5/fqmIaVnW5wPAX24AsR19Mlec3FZlQpnM6yvGHzcYf8E
kW93wxKbJlS9Mf+eQ8pkOwzWh4EQNSE0tJnkNvSZThVIKKGdh5/2hrypJXmK+n1/u3ixljPt4Tqp
MTI78vHWXyn1tIln5THBjrM8DTenlbeBhQBx19acatDgko1YA2BtEFWU3r7mG2ZJe5BvVQz/QTJ5
FMOaTpRfk22ZTBWkImGW/4UtnXGLs1gdrSCDc3kXs48zbM3PfywLb2Elpbt3ubqEdHW9EoBAsF5P
1Rq31wAm2He673Z47X1nlO6d5dnahe8Jhyj+vpNYnzYpAoz/7+HLFFq7hGbZAs0YbL4EiG0BMCpC
0crSiTsjpBL+hJi2PEwQRWAiMa7y+U7GzFATm7w1+L5ariwXjh2I9Z/mJKBkdRNs9U4jiztZO5/a
4hWSozTQZZvuRuWVlm6u4QxoGpqsx/wtwf0SIkEumnTo/+q07b5PrvtmKsnLjE4Ei8/YlDhOKHbS
qS3rRGrXpauaoNl14NUMBFu72VCI5cv9fQhpJCy19rUzZgsxFxZppOhmLQpybCE5alty6deDJO4Z
F1tzKxnbpXWaMmBWNByJEbpaSIlRc2onUxaq5BpLijh15shnPxX8iFEE3xXMTV6Unr2xRc8lFmTx
R5GipDUPVtCDHE50tRJ7pCd6EIJQgA+PIOshnYfWtiVhDjDwEGIEm368Jpydr67/CdE1rm8R8Tdj
0UQdmXkYuO/Vx5gsECXafhCVL47QWR7GLVJJ9G3rYacVis5EwejALGQ2+y1YQ9lofAH5bFwCmh7G
iJksWnNJPq8napHQL2OS+Gttf6Kx0CV7Vf/juDIENimUmQD9FieIqjU38mH0xlFwJkmlMq2vavEi
DDKDP9finZnz/ogOljnfMUQHmsuxEpd0IJfBeqMbNa/SLEVZ6fiT/T/fAlHiLh85wsG0xVDpyuQg
MxHkdmQkoe/z6QMqTGt7ZuhbYaK9n7BWRgQSZnWzGYN24vjrbem+Ioj1uh876Fxo2EJVsTvSN3t3
Eazr05bfF9EYayeMwEgbuk4BXYJ1voiAfCXxCuQUqD9ox2rfg08ZA4WxvTv6Z0fnQjE2yJbDYkHC
JgRR+WgB5C5EShAwWzbwwhZwVnt8D/oQKKJltXf+oopvvxVX1tFjB0rXUTmhX1DClU0KGRT9fClJ
PSG7z6v5IRVK8gCo7WDxxNh9RPp03TnD2Ny3SrREMg0cgWQYBfonoyCF/4uAfNLumd29ow4x9PRQ
j9+X5m+zZnAAXDjYTdoMgbCcQQgMmzvcfEM0MJPFQQKltsbyaDfCpH3y9KZJQzirU0ybnP4j4yIX
QNQlYnKfp0PCHQI+kHnjr0lRgFsEe2EezeFuTXEUSUb5WWlQ4ZiuipBK9HOIYTKEdC3X+8oU2Mb1
xFJzBvurLxhbdV0ygPcZNJbdM7Q3Io6LyT3D7cJrSsvbnHpeRt6H0cs70Ca88BLRddagab3IyiGs
D4Ctjq/WUeqPSml8798UFQ1I9gwYIE59qhvOKAeB2Y8qZAn+E011z2N4dPEflHs92uqN0FeGQTn6
B6IZe/r8PekTlNG68uwfWOOQWfXn2HPBeLv3yBA0xiEcTFsd+RD5hff/zhbIM3HVVr8f7kw4XetH
fzOeUc6VHirDTtc5LISewaj491uNw0Jb1CqASFNP8MIipgY4BCgqwGzT4d2pyovQ4nkZxcrvB4WD
zoeGzQLv1kXm39peZUM+/UT//z9efYPzLhmmvOSsDS6exDAOs9Yq/e6r3/OBIpVZHWkI/N4cOBHt
sDD7McsNRzye5usqH3YSMwB8ev1Pa4EJLchNJlG8RC6t+XqRM6wa6CsMUFOePUCHdWo8BDqtQkhr
DkhbW1qztzjHOq5cAHa/jJ/bo+XKwk2W9Ipg1Q6NRSxdhpqTbD8Ayrvhh91T34dCm7v7XXoJxKcA
Bv3nKSYPrnpGDocNnbvBuJM2zqGtGg7FnDkBVN8PXb41pFwPjD3BjNi/bfmkDW6k24gAsuPPxQtF
Y+sxg5HeHd63UYjJUdzDNWmHVfc8WxoSG4BNJmyCOM8uRVESg5XZWYwEyk73HFXcoPtlkTbs03VP
oIgDQnvkAsOoluEHo1+uXSCS20kwiPI0RhBGVrRuwI17OXugCse8yqQDxJ7HpVKYN6LoIRI1FFFF
VDPzKRTeVcY5JKSlVqqlNNrhph80cTUAE8fsQioyy3g1eBry3OGkKxiPD6gNStkrVyUy43uhqR7s
xGem9Es5jbU4GRq3XJrWtRxfLC9FZh90hDfCdUbcWnsRM7i9wa1JT0gXbDj/KAeRWanzDCSKiCFf
i4t3CIXyY8bBU4l02UlShZUNHK+7ZdsV/4VLrt1QGWwXsv19pEmhEnhivhF6ge0lPbkxvcWyNndt
uujvdIlMJwGaLWLiZT+92xSfrO7bYZsc/7u4QMqEHXVOLla/msJ2CafzYvaCYZabFmzsEFWk7WxF
qR7rxGM9P1qBP61M2vEVZflJUHLY65wm+ja96WhGmhfHt83gvkxC7JG3df+DykUyNjLeRgpj5Ukj
evB+CGmaUag7YF4ujDxw8FFzmDZAQzdPIgAcrJQ3DVHCsqP/H9t0h6+XPlfP/79iiUkJz2ywDvwB
GJXC3ZjF0KG6Qp+Xjp63YbHNN6Ocfl8r2kE6jIk4KcYANuzSeA6k61Bc4z8xUi9TX3GMrQsXK+uN
Q/jO4bC1fMw9adXk0slcFlVDUZNv+hTL92ThWKt6kiEu8qqKgFqb8uR6E7It+pt/gzRNCZ+OIvco
QxOXl6qnMJMnqvNtuDxWCitJli92H+7S2yv6gCcg8ClRUoSBPxgjewGZAdQaSNp4V9ggO2iHtcei
j/TUqrFafaPMU4kD1pctn2TTHfjXY/F0dbKdRv9/7tmq6eQp6HkvNDjkhVxiZtz0Aaum/rP5p62y
NhsCXNtusGrd+u9WeFA0LOa+im9WNrHNp8XzfXLo5h7TaNkvQ2aVaw8fecs2WRwsdJijr9sYyVNI
LfDqBI2P7jAAmxJoiJRxUvuJjCOw1DP07xac0nxhOs4we3Fx80C0XBoqhcRGC0uAl/lYvwl1L7oq
R5WHzXSThZXncgdHZdUP91u9kFAn+ki/zurtoyGt6vGWgUpjxfZHXTVys4+yn8oQkxxlszgISnTp
Uw6AqEh5er2m4fPtkSxPirpVQvXk6E2x0hbLAfuAWJIsIE2JECSIOD47XKi69AOtxS1nAoLWzlX8
2IbI3jHJitjcnHiVK66H7QjD1YhEjZKYB1l+4Sj3VP0cj/2JKqg3884sNKsFUNf6yCFf3KhKTbj1
ajy3nI4DHkIvc5V7kEUJU4E5nodbwWCdc4iOcufAycD4//6fsDdqcpgfF0OiNTd5WDbzIYVv85dK
ZGnbe3rZ3yAezzqlzAfkeMS0dN6xJBrOPhj8i4FQUbKv47HzBdeLVU7uAox2wogMaAqktim0zaFe
IOkSPZNYykQOdeRnN5tYZJ3/fh224D4Cf+dZsuajvT0TfvtHYHEWHhfS8GTLgkrp7u6Jbut0felp
pNwY7U/Eh16o5pAUJpHPzniJS15wLxEL3KVYVDGkNmjBTWwIOJ1RSqTqYsGs24xHn5dUBZmZSWgL
ef2G0bVhRwQ+baNCIEw9qfwTujS5kASi+4moYxx7GWttOuif7a8LF1UzM61cDo33McOzVtMpyRAM
Ukg6QUUogG29HQ7cJ40PR0+Oz685iZfThOVx+gXAWmRwtSeHCaSkhaZqOZs6SvWLAorEnfxCW5Vi
JqJcKKusRCVenI0kaBQ5RI0HezsQAZc/spEGvGj735TDLTfV5TSS00i1BjiuO0Y/jOLSZyN+VhKp
a3T5g49TLDotDt0ISlZxs2sSkvw2/lZYIvoGIysnOb5rYQvrcpQZB8xXu81ot954IbHkl+A+Tf+U
/KeRCGC/lMeDY6eW/TkT7GWmYxmfARsGQDiAVtDuim3k0tRDjQwKLS+lx21yOwFBWFnfM2dXLLaz
he5p8FUfqMAPvlz6cRLRSH+THeKDnDUdFLyWWhfXXZ6TxaNA7jTOhpHbXHJtmy2Wnlevpqww9Ck7
yXBHx7DNqggCRkVfWhb7
`protect end_protected
