`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qk1+dk0SxlsYMbLxtSYFB89S4dR03Ktohh+MjH1KuybVuXd24qVvaSWoyMBJzVgtpguT95MODZU9
6nOHOr9zqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PnwqaCvh6J9ZOxv1i+Yq0LxPfr+MsJdN4M9WBJSL5iBHbWP2MentI+Jptwlu6j7aLkK8G4e/BX+E
CcHwwBsj+xenNZJeuMF2Hc26iLnV3Xue4OQbkK/4EpMHhfWUU38ZvF2nPMTm3ngHovvwKy7A+x0I
B4C9lUstEGalPOec0do=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IGGr4GqcU26NQ3nFhrPtd5Wyr34234FvpfTUJhNz0nGCGkWWE32GQpecgPam8aJoNIa2BM6Hxxdm
eHXroBrEWrmAY46uXeB0qf/TThGCY3F+X+J+AnSJyAJKHLtXX8g8ZbgtR1Qqslj7+UuyDWzo7Nl3
DcGux4hbFy3/L6eV+nV4tJx/DBTZMPhaCJi8BDucBHDXwucbYkKD0EsL4OQiIveSrcHvzCTd2Pa5
sDblAtqny1lKpLYBAxdCC6Vl85kY0DKb+wlFaB9QpJOYsO3LAcOjCRCZ0nTnco3eGlXDz9wCFEaw
lpBopv7pDWTQqyXDMcE0WwVqjRxZmroCGET3qA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QHkyCruxyUUegutNzoXAKakYWf/MWpybUE9qun9H/L2EImY34qXAsCkcfnlctVpCvCACoYmmtQZa
9X8Mk8OjCThrSbpbZZO//dXGn1Tf9JGM1mRWZAXBXL9wv04fbV0IwZcmCitVFHarbmb6PYgT7AXE
oL1MVQXNG4/1n/bQDBU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bZm0RseSCPF3k7a5RjuQnFnLj3Uo+8WftwLpzLCUR1Nf6zYcSdDQVBo7y2T6an2KvUSMlozfLv8m
Oj2X9fLMJfIDAHGqZAIoYhTkR5YXdlZ0htX77C7glIPrpcHK3mkLgBRmmZ9Nj9ZbG2BXwngbojsq
MvgHrcVwBBmxtDnZ8JhJUQtcCzXcMJrV+ECfeCnVkeqwsGOlShebwpVHFu5Xr+6cwh0hHP3V0htm
iGK+B2aldCGrKFI176DiiQoQaF4UM6a7ZPVZdVzdkbcRW82EVw7MM+qBdR4GzXLWyXCwkA6Y9TkX
zcUAnJML8a0LITtExNxSrqeFQiSxZ7fYCSNVkw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16240)
`protect data_block
+5u8id8dlSH8wH6ElzewSdPCNLn9CRVIpA54IOPr89CZSxFHlspv/O8nc2K/v8oPg+MosfKC8KfZ
WGCwemK/G8eQjS5jKSEZJnP3BRx28N0RJN/v6asyS26LrdcfdcgWpGSzdk64gfx2++pgVK8cMOSs
ZeGxPUedlSTVvdk0lvRZYHPOiWyIFlufeor3lYTV5NI8+jediXMLXABE0yT/FMlG3hpLEJaOo6Mk
lP9zluUOV/HqGXePibLgzX5ooxP4m3YAPWq7xl4tqx4UBIjDiSUQU3bgTcvVls/8G6yDgf8sBVSH
ZaUabw5dw75xCnddrQMqyXqDbJRL62hBiPNPqktxEWb666lij7+dUPENQv3GD4RT6nmL6XNracKc
9RJ/bSyhwT1pXzSX5rxZyFHkWRrd9cV1POMWE4ZdNzOK5HyDg0fCQd7rswYGkNRvsB0zTOrfFimY
uDn7ZtkCCJy+349n86OPBlFim7xkEJ7H0UwJolsKGxhYAaykXu7N8HW53yKr4XAP8B8RgLy7ab7C
2m67e5JSvGJCy6NeMUrHV+MmMlM5L4G9Xfddo+EEwMzcfn/ML7/yjOymNoyRJuUwuHHhdeV1hgyI
sdoFmorh85jp+aJme2viiHl9l3LhXV8QGsdlewAN0xn6/Cd2lDK8S6muLg/yxezSEm1lak3EL2lj
TGi324K3P5rph5eOR2SRmm7sHuLh9u/II0HyBagwvyaIx12YF03pwejjkp/R3IhN+ffQTrpjWWT/
A0pUH4URudB4ageBmzuHU4HXvolAFlpmAIRWT0RqSyjUcX4EjaOaX/LG7D0oCT92MWMJtx1vm20a
CI1pkD6wjcOhrU1xe5yngnn/FTXzSRCFcn7pRzEb+fTdHmQ9VEsGdnuH3octOvvLGVF52Io021ps
0F9IThyJITu09c45/Pn8ilgwKyUA1MHwMjFr2W+AZ6iNyjyXINqHV84zWV8GXB+U/tbl9q/JNx9a
t9T/c3WdG2/njKN8HRtZM6Jgk5ogk9EsE+rx+t0WRAw1YIO1BlxQeFZHy4L3u1aXzWBCeGDJmhxM
tlLjjFVtu5Ie25RxwC1HjDc4chC+fXpuFpN4U0/wkkt97gewjRAbQZ8LmcOE9+7QDGILL0/35ACg
txt3CnKnsfTYmNEJc3CWuwNcd0cfy9qdOdKhpHhtxQaZOJSL2c2HQaR45ZWIYMlR3cWCPmxpTvbk
lgfCLZuon+yX1fUNQfp3n0wDnoY5gb2ePqrhg7EG5BiKFyv87thNYDukAjHL3x82BiRVnNhv3ova
hN0ki5dNIOlf71xAfg7zZCbegpOPssoR+1Idq/xZ8M5J+HZwYJlhuoWlVpWjwkgLfKt647EcZlsp
iOFDyekHhjJEx8wdMKy9WugKsmS/o5EEeNpY+vE0LjM8kGujuO4GFQXB0yrWAjmbF2miz2MKXx60
tYxbiyABIlwpcppfBZJ1ZcxrRn6TF2ehnYecBR73gpN1ABXVZsukYsATct5a3VGIxHoQM28l1mto
Vgcr+EYu8Yp0Vsn0+oxHUyiUVUs3d1zSABsRZKl6O5OjTi7jTXUicHvy7f+YBbeA3tBDmxwqHCOG
BikpjVtTz1LbDomuzMNO3+annYeOSSLabebCgpDi8hx9njJF5WIJAqLLCYlYQfn+eaKy26stpc9K
YFS1bcuvwgjadTzMT/lWvxgceC9OLg2gyc5+dS/VSZ/Ei/uJN3NsPycSr9yR+OQkzq0Kzs8+zEmt
u90+Z/9+z5Zc77wm8gQXjbJNXqFAOh7pyFIKYhGZ9NH2YJZF0DAcRpx7Sadxq2GwSEdGOrx2ZUA6
A8fvlUuxmVN8QpFnrH6X0UItrGjeaPqJ12UGl7yQO2ImuCjaCx8SpjHoVRVFxWg+eXRKClxLnlbQ
Xjy8OrxjTh9nxTlVQZwJfGT8hpig+GOwlML/rlxdXoEfiuHyhMS0WxDVPJi0Uw9xJk+QHWcDJXQE
pMDj3xBUriBl3wTFJC0fbUlsi6sVy29MaMN2Q0TaE14AUIUwn2qKZ86K+Sv+WdnSOEIDNVCwb+mc
VLDe/2weIT3VyXeXIWJSTWnI/dx16s+saCS56bgYUIg+kk19mzhTMPe+/Q6qyQ91jcHJ1RJ2RNgO
0IrsSMiK3m6EYxAz49QXXzDkZdl9C+2VzXirXYiD3yylhyElolX5whG9geg3mgrxv2SxPmQqeDVi
d1S3FkOl+Gp2mVXpu/QGECagmfvwrxrb7OCqr6XDJbTmVfxBurh7gD3FbnVRkd63VJQUBMveUQsQ
P0yEjGUID6cWqqkm61sRDOP8eq3ECxK2fTioq4FWRYvrkVTOmA0qxgGmRrRWDsH558yO3v6axW3A
YfQ85xrz9A/AxtF4mLN39BBK58OYgUS725pYWIKOsoUJItIlk50cWBhCQQB6nWQ72s+SXICYB4It
Ux0eEfeDoPHfEpRQp5K0PjvLWS1zA/H7AJ456z2jdARIitLx4S7puoA0FLandBV+wEZrCxmFlH4X
yqVEBe9YVbBQ6vKT8PbBmcDihFDJPJnGBfslHSP0J6BBOrZnsREEJzgqgXxYbzJFVDzQRopNbUK6
/KeuBzTqIezJr3iZ+vAY7EPYqN2oFi7RxPrSv+VUtfYaly/CcX/74tYEfkFK9Knf10dTa7kZN9Og
51hucmjrFVOqHYIfkzgp8nhbvnwOh8Y9LvqmDcM8/H2etc84MjWTVMsbpVndjzstGqh/qx/feKN2
4/0VnTeskb/AgrJBOH8Y4bmn9xJnwucMxxJmVAfMJiv85WGxdrrboMqPxLSmLYakh7G3DpcnAMeP
dXCPYF0I456zpKuqFAekJsDfkwLyBCQFamq4nxT+dfoq7BAuOicqDTN3gCV4r9jPqKAsi+8d7odf
QM2VbVELMwKD67eV5H0BpTsq7zM64bMxQSWaLojctNElpARg9cFu2ncLu7dG74YxuG1fXO58vHie
TXaz7yuFq0Hl7qO4QCsfvVSjeN3JZVlB4kFGtuvCrksjzrnEgla4p/gSNacVFbr5kOtd6IQd/M09
NwC6dXN3dbIi2tlABpsQfuhbtkswzlGTLdKxah2ISJBNI4maIH4yJ819pZ2fVIRf2aHyPChxIrMm
sYacR3Chmv27i1qKfK40OvtWR6IMttNOW4sFg3AzbgWPvMATsDW8laPI0yEY1AH2EFuYaRJr4cW/
kAZj2yw/Kkw3l49vgTzWfqWR2xyvP4rculbkqNIJfhO4ZEnDlJs5IhtFoslU3MxodWi+YZTz1ot2
ZRap2XfHxEq7kkhMZA73xBwRmo1ZzxHaN31t69/5yAVBJJhwJxF5aLM3IRq6tsQ32bxgrB3aKIGH
D4HmasxE2rfbxMxH1ptSlpqW7dCj69VpHiUuDnY63r5wNyIWmoaf/8OzBdFYyCVX6ZT1pD6bNjX+
GIWEblrZ9ZnhijWJZlA2kkIMfXmfh0w4mo6ddgUxK7X7R8Zfktr/Xj7FYHqRta0eZICLfB3M0okS
NAy9f2NMoK0tJLw0n8zIBa7qYb8Znu9asN8K2QUFsTK3b/Oq3aKe8k0XzXRcDE4RoB77SdnVl8J6
BJ+WJcKOX/pHKSHGsvgri7nlfCRNY293ShRa3K/bJG9iwLGNjqIvqxkXAwok7xzw+2fbpLxoycX/
gbnxxg1PQrP9SRZ2j+a5COzA/7DWrpjKCrX1/y6IFmD/H/NBCUHFFGp/8D80PlfJrXCHXyPMoYBO
w/ZEO9jA7FR7F5U86O2zeeuq5EkTFsZIoMjTdtQV1EN7wpigtAqx8yueqcAlGyAB5uIFMBOgzegu
AqzBKmNdmdZ+TGMo1JS6sDv69BTWsmCRvj675n57nOSKPxi8TKCfSjXEpvMxQEnGHya+AVJbTc2j
5qRKerfsZqevBtSS5rAiqzkZbUEW2LBBy/SXGiAsvL9/tDdxUUnZpF1TtPVkx6P3GYAZ/Rev2yc2
HziJBsn258wghgO3bRiuffUQT/sczJ3VEzXVzk22taIV4fyD06KTLiyBz/Ef5xfVhFV9ctBfM6m3
9l8/htoVY3B/GpJtccXS/NI+SthXgU7Vhfpb/cTbyjAf8EOLZr+nFpjAv5eJAfYr+hDrfmmoybAb
2g6EJvVpB63MJOh5SSSXGa4fM5T8WDl1Epo8Vkc9HZU/pFlmTYj9cG7rhewFAbRLLjBMFu24jTws
H/Mj8xvZy1MaISG4Z0AN8zZ/hieuqq+iDlWGrJhuSNcbW+TNElaT+MyijlHZLl8L1RsilmuidoO6
GpYr8jQGCfw/+vx79ERX2/6RG0gbKtzdWgduUXGF+ImQRYIEPmZZh7LwVOBb5Zp15tpt//zQl9BY
SIE30iqzL63lTOuWM/BK1VSfdR33c1KFE5mdvvSuMc0ez3cIp73nDktOiNRPhsLjPN6NWTWLgI3B
Ojl9Kt56sywdGscQl4OilvBi0BTvjMLf19jNaw4my9Rc768U9Hu2nLj6/7eW0h6Qc8MwlBiIprv1
Ois8lirjho/+unyK1s2g2wOZlYUu4GWHpUM7xjK0yV5EQtPbKO42PbwSqTVlY/7GzSnypq0lYGCW
wbGDwq3GQX83yseqD21btYEkI3OWKWEABES1eAiqte4enXj0o2IR64rjVtmWHS+8BKGbRH9vYKYm
qq+LYCUHyx8R3pqwmYflLeZTVyjVUJpyA4DgIrYmSbbUZrtE14jawPMDRyyg1hwBcwAm5Tx94TE8
tzpYCaRnB96hfDvocDYgQvBcuzfyc+0xlGf83xO4ch9Ah0+2qjPZYFof6MyMpTKnzqjVxmqpQsx5
V/pCedxR53RUfJRvRkMxzTb4lMWaPy6F7GD5ICPMDx43mo5XFds0LF4sQ362oa5b0U5BCpPyNKtl
6PL2e7DBnuDHj+TSpkyoDIL6JQ36tDre5xSXF33ms4a9ZYiWMAC+PYs5V548VJ0NVRWP4/jCZFN0
616kqRs+NnLDM+GUjN7uBfmt7y7+GiF8u8hhypLGluFp5p9SvLgCBFU3IsxNuTnzE4OSTTwijcVD
JMW8c+WkL49SRJbW5X11DPfnPSUS7vZkRj4sIMG3p4g8u0TNSu7qc9qn9nremUvgZxJHj+D5LqAF
bxONx3Y+M1hV0XC6WlRhXSF/jzlmTcNZosQWQQGUDChy6II+fHs5fuCKUFh1XjcVjVl6jMc9rpmP
zcHIqb2O+B7PgDaFVcv0d3uNosgXAvz6kw6URpaUlmp/W3v9dW4Z8y/keDyuPkHqWqseNOrnx1u0
a8Mv7DK+vrpL7/OIIyqp4VcjGGy6j24hOAXoyCNOcDdHP+vY68GPYh0fR8P1JvQCnoeBzXod4K+w
GLwcHKY8GrwRxlKeK06vxA3j5GNs9LE1IC6wpDm6/8NjFMEce+FhDOADgGjHjSVpLm9vhctr1BbJ
658YK05WrxE41qxPbQ6RYGuCAjWw981MgKb3cxVsvjVJjqi1i+DiqATBmLsXDrQpyYIe1MTXrUS0
2QuDGCHFHGDFYBrJEcD6bEysKc5DwjsTv4Ei3/LPOB/CPmfMKjrK49pt1YuJ7FHzym4YCa4nPfTq
6ojZUCrzUumIvwf/v/AwVuTf6HGn5AnoKoC222bm71D9WVvUCVhNszvacq/9xvdL4hTLMsWlVoMn
vstOUG8SZisy3sZOQfDPvAQLwy5aCyGqRQEHYWhScaQW73NjFEBHcXaFM6D9ZJjI3esWdOGGYUQP
gEsDRriDWN+KpFb6OPf0vZ87zo+wAYj18bj1DCCt3L2MWxSaAtHPUxyDPSzWQB5dW05g3KgaHjHi
6x0P3ZQAv3uwX8cSVJYsVVVrj1o6EE0pEjb9YD3LByZT7p5v16x+G6UygD/gX5O5x431JAnaASre
TdhKMxN3W/mG4X78+PRWIsd1bIsk6/Bsq7QAKM4niYXFhreHYYmYS7guqA4768wbdzN2NtXL/2JE
0Ww0j073s6eJ/qit7KiKjBlro55SrUSoSXEGy8dvTSGdYlZlJbFY+Vg56Q8ds91C0AMW23pmLpGo
aMyR2uJ8o8bPG+fH9qL4pSSZI0dFl+rHyh75wVtMusZrwrCO0tHI8sZE0PdWiRCUXoHg7VP/EBzf
fUjdCURryhwii1Vu2IKGt6V2Z/VYZFcSDI61/dkujZmq6DuU6XPflmDNTvuGud8WRG+9DVvwF8Sk
C4ff3jEmTJE80K4VZBWVcsIyrz3sZWYDHbY9WsFqN6f3q0nOgai8E3dLXTncrmgoXO/2b5M2bmzk
fFIDbV8NBc8ruEVTNwmeFNQr08NWhNKkvCJI5SuapKMHi7L6NSOvgattEXLHah9FWmAjcXUL3K4E
u6CrxN0GaN9bAcBL8uQM4FjqLx1kGwzEYWBG8euwoc8DDOeBAuiTBEn0cDRGpQLYRVFbcaVReHCt
LqjQsjojLUGhVpNwhFQ+1Lljly96QlxLliRBHCKBCs2lXArT1vH7k4WsBKMDA78Vg2LkHF98Sbzy
HEaXpJZOQgVIOccQjSzlnA79fgopg1lNAVQkrH6uTK7yT9iW49MV6NcmkVXHkgf1Hh2PytJopti3
n5L2QMa0fxHObE5VwEVF82+6XWFB6Ubi2cyPvySeN6GKgiRQlqnxWIsfxufQ/5ZRPsW2lbNtxmJM
WvjHd/RWAoDDb/Muxp8MblXCytBQLloYq8I6OlGyLZWtc4BSOCKJaeEKZ5VLzcEb5wHLgl5831ab
8jikOIPbbU1KiuHN02aDQC73JT+GNH4dODzmBkux7sNx3wzAkDX+o+6xb1TqNTAZjEQCkRbFM29e
L4JMjHscZBIvBceMkdMeOCWswqZIGtrOHAF/vz7xRCNwOl0yZW+rhiUc1uTnTayeF1vtufJBE4c2
Q/DD1pUkOnRU2lyq8BRO7skeKIVIkk5RMA8K6qKrMVTeXZE+gCqKj/XezgVzmYYzr+azY3guFXXw
kZL6eN0W5IUBPfsAu4DPJL4m32CWjVpg/pjkNksIQ0Vs6yQUUNHl1WOSPCY1IVnPWP1SiIEi4Y0E
ypQ2VRaWWf8oRknB4cGB3v3EtppD0MPSIePvb2X0WK73eNkbVAT306Ia/fc5bqPxDbcG0G3s0Y2r
NJwKMGHAj0As4B7LISTaKiBps42RnIZ6oL9pGGWWu/DUPkAp8lE5osBlbNLgW1NS5zL2ybJfxPL5
EL4xr3y+2BCl2zb4H44RF7dSUxUaIz4kbo+i1qZ5mnRIp4yb7GluZbnMp005RgJ+CrbcmjTGP39J
GlyCpW7U4igjWNgLajvb6nrP5Qt+QyTuCvY4KXH6LP6Msmx2vMWpP9kisqjeYkKMjiU/PHPVOxJA
vx36QSuA1cLsMZhK6ELX1/jmtsmhQHBrMhPJ+ArCLFO9lfSZSvfz96rwrrcj72VzIl0XH9VBVQl6
NhuIPam/qU4NH8pEN9KkXhjjuTg8gB3vr/ClKfxW+GJJKzWjugDZwqG5c3ewx+g4xVcYt8megcGi
mwA/+lhnFO3b9FcCp58FOd+xpqcS2OywVjbQYwhjim6HIya7sesF8pKThcY+8vMiWZsz04smQ+jh
MvxrfYAm2cMlMo6u+NcrG7whnUl8VMgaoJJXwzTvPsqZMUieIfNFXUSNBzOcwjxA52mtLtUI9IBb
9SmmiXfMGFCcx0tF478d9H6dNGEuh6+N98e+KHBn1+JqfRpYr19Bm4PAvG9zf+CeCz6xbCqXX8RK
qVdedCop04a+EtK0lyd4iM7JU5goOt+31FncjxYC560V070EP9IgU18/4P/aDtmpBOJcT1kz2FxO
17m4XbP1o0533g2wH+sgZ18IQjT7N0iBwVXlaARHwSe5RhA34L4yRv3FlDwXE23xJljjezNnqBeR
LDkCa6RwDe0VlkY40GhGkfRxbioHIb0WjpX2XlarCV8LFKR3dAx1emcetiz753n5ywZ+TRTVG270
lkWNBlPcOrqZKwIx4Jy2JqnB3U9L3XqfTkXiRy+N655uNHgHOeLJm0UWZeMpV8EYR1ZLFH0Vhpc0
mCnhV2SP0UqIaknMg65kou1M7B8oA4Px5b3ePNy6CzHTSJLAwYjfj+1IIDP1fqrbVBRD+vd4xMZQ
xQHs5eePUoCC8ogWQOySLcN9G42nOYv1qPX+FYp7TB2Wv6l/gXonGxgG3SuKqbwM7k71y+4RLs+6
sfxrLVduHx38zhuaowU+aIiv7Obq/Wpd2pm+58EuJ5aVLg2FCZv1h9sKd3MtKeispjZ5e3eV+RC2
Sc8hEBcPhMZECwQq+zp/JFugFzKrPTcXPANYbrifsto9OlR8IggrFfw8CdLDIDhsCX/mvKijrJti
DGDNqDYhfJikOvJZ1FaV+rjv5N1+lty6HOUkmUAVcyqFWAs7oSVxSA/SEu1MfxEfjxhoJ5JYqBBD
iGNIkvOdMxnfE/HAjDD+KrKtNfT+UknomxTlRBCKCVNf+4oXWlnuRjBcvmgs5091wjSZTldMvQhO
3qiVqUpRW9/YAgbhijgu6999cZcSJPoZQ+MPQrekKdWkvt7WhFuBR+hoWfGTo5y3UlSuOsKBV1am
sk7PF5zqewh/I0/9MYEAvax0Y3Hwbh5ePBMQUxqj4YCxFW09+ZuSSlwMrJIu+S+qAWeJoa2SQ5rT
pYuA0+7Qi7bWcGHTmEEQeB3gYpmW1TDnJpcsxQHXc7UcVPFqPWjQ85tFII1G0LhxwlEttH+xpt5O
d52XYNPw8IpI4hOIJ0KFe8y4UgyWUFt9SCBlAHEfv77TyH0bX0+ozbaWtqwhDaVjzzqXzSnpWdip
DuIAMWzfodMXv5TaILv8aRq8I8k6BsWK5pTDlXKZxRkDx5W85R8vd1v+hdoVH28qamLRp3klKs4o
zrLA0GWj3AL2am5vIHGPfBGfd7to2rJB8sN+G2byJVmRVRDtxO5nThXGsH5LyZYZWMzyGzpPTxVx
8QMRaBfwvGtGscCgl5+go2yhTMlBkpBrH4qT/V0aOhm/I+yj4FY07AB7o899BywkdkmCtsYhH5Ql
B/ZANCx0v5sprbujMq0sX2m2JbqxTUHT32kuhH9MfHI3WBa4ZGuoyU9KnKAJ8gAboFEw85zdYrqK
is2j7WPlWn/FRI0JwcSqj/9MjL4UdHigwNh6iV2Bg22fA8JQyJ+R2QBkpUzLFH7gvB4tftnukZZ4
Rz3kmRqoZja99ym+AJIlgL3ba3nLzY/S5vzby86axBZWtbEmSg31fmTFNODTNgval2FxuPqsDDKC
cblTbcVMMGXQfc6zeEV4CjmBMgFE88lvyz/QSHloVcYnnY18cTWHMWNw/ZvCfKtOaIXNRkyGnbKM
oL+HnuEAhb53hqVQblofcG7V5oUtcMtRhPdOxt7xHKyZ+sRTsoC6JZsA7KDm8ZSpZAzEuk45m3y/
VY1KAjUScro3FNiXtrfVFAt4LcwZbwg0Q6bfpiayRKvRAlXYbdRGdejuSJ2i8CVVt9wWj8BDF2mC
quQistLpSlRsRunqo/z9mkrWZdHpn1X66yLoeUnNLEBvj/7zPN7r5fSEUyB5+0XBrGFMVL9CJ/BI
CiaBg6kJYFJkZqOp74ycr03DKnDrtfDXedrwSe9rYc9jwFyej40zvDG+7YQM6SuuomBMsMyuQy0G
o7ie2pgUnqqlcPFGLDRqFSd8S1o1h2S/dTx7a0cPFBUZscOU5biEXEFUPcGqs2nDCH4Wkcy7M1rR
m68cf/6d7OFDXYTOWscGmDO68k4KUs3jKUKGAMA8xG4za4k/8DGLJ1NR4KB9WhlM24Ii0KTEWzIL
ZoA16Tm8uUzw0/8b1sfwgkYfaIkuRC6WSFhN477eD95PPiWPRSHg/ekOTAwafYJTEKFnEplfWd6X
I0U4vQD4Ldrm7WV94n7Ck4i/KWJkoNN7s+t3yrF6YochbRb3bnYwdjebnwYrsJx5Zscbrx9UYU3g
CB1slqNxC+8ZL1rBFxzUFJTlv5Ksbeagqbu3DlGBbJiTyLYXrsahfzTfuF1zxiROn4DALxkR12Km
PDKiEr+9lEEMXYV+tfuC/V0kaBqhh5DKn8N5ex2U4WrCXJm+JN3tU4/rpQmG4okNuInbEDsio8QG
jYyp9cceuYVB+Ua+ccmCITDPitzZ8EhsPE1pOAxDPqW4rnqYXoKxa2KT458MeHzOjzclXV6v+STB
pLcjI5EE3MzS/eZ/STTqSTXAoicwp+wcPZccKFQWtqbHdU25Y0RwnP66L02xtfVvPrNHYOOUPA+l
KGzAJ/7qZ2F/yV/wAcOM/GyOvnHGPtu3VCD6nra8o6MGgbGMvMGKU4PD8a4g63Xhm3KOPHwRS7vb
XrLbFM7xpBi7eUigRNvBWQ4VsDHlnE/mWDYJjouru8qQO6Q2/HpzOkEYfTiM+qGozWtJj1Rsn9Ry
D8M3lgas+GIMGiKiv2iOAdkqXy2ey+XQ5Bjj9TWOd/w41YJkeeac5JmyJJC8PDi+3d2SivxcSsBb
nF9Jcv5fZLeuSSbrhOCMchhE9XwYOI3FN+g6wdt6CPMech4stz1EXj/h167nCwdW6VGl5uxEhb9L
0hNnhAiCGwI92RVP54OI3nAWDTbLXp/b37Bx0n18ASQpBgX75wB9ZPQ7Xoml5kM5QsMYyYLnSIqg
SdEPYwX9N2cjL1gq4GjbRHnHw5ugHgkGrrWDC8dGCDhCViwwxYi8K6oDhR/ohdQ/1xSluqw6+oSA
L0wtzDF7zjZy/044v0EmtyFj/cd2y6m+U1l4wDtLz9L/uAI3ccCg9goZ0BZqUdSX2Rn8kuumWj+p
+SuM22S0ZsZq+qFALQiXhLssjFOb8BmULNXdqVeqnm4fkx867L50rVniUBjoAzDztRczRoaVw6BX
uWwhpzGvWy4NwUaEQfSX5pVF92+1NNwrG9F8Fp9lU/0n2E80a6uiECmMNelUh3/k2NW9QSp8dvPs
d+oMFZwcg0e+zuY7Mprz4a/WYGyXovRXBhdG08vKkvTd6sfEyjJ7/z7Sj/SyTy17E+qvsmCvhub2
K56zWwcPhFGVFHppxRFYuEf6Npq1xWUId9Ta+mO7WNrdB1DMrd7X27iBc1nTK17R9TfiMP96BQHo
hBDgw5dBgDzuo3BP++CQ5xFSJlQ4LWpSe9gQ3wzt+BqiL/r0l0m8Pp2Ionokqzcj095DPoLr2Ugx
7gsGzyUjEFp7DzEWHd+JlPWwqwFjSwfLVkObIFKCcBxkZo27WiS6FY0pD0BcGS9M66kTbb2E/po+
s03vMB89Bx/arEh4+Y9yTZgIMFZEWHsxYNybsZl39CtiDRLV5qZzpD6Jm9I3wRlULjwNgK2n17JN
7tfocvVcJ+e8KdEnfoSJc5UUmhgCtDqXn0XsmlCqkA8w16d8sElMDgC3ZqAFUnC2T5ylnxmMOS1P
+WUVG9WQ0Hg8VnyhjrEAQxEXf6RH1T037lXKcW+rnK3T6RSMiHJXbiaUmuX9S9dUQXQw66eSRbJw
tldYQ7Qj0f/Qu2v8KOrnjNvMMa5HPnWuoptiH1pI0yBcnA5Aa+Fd9L4TKOgyUKflpMLMbPhDokw5
h1+ZKd605OQye+iiX4bRdCI42uzhQlLXSsxuj3S/7mM7ogSpx+GArn5UskcQk2EtgqnkxH1mwglW
qJMg1JZZbt081YFQOtXzrdUlqVNkUPgvh+RtHD2b8rVQSYeWrRoyK5g20u8R3h8aynn5A4soiMyT
jvUHM1aGFTozRFXyQqS89gB4iL5Idxizc1pTWYUFsan2gpnNp/CeNUGwZQrxpOo2TRcoFFyX5Khn
I7ZB3SgKCrEdSmEPO84B1wsdc5n6wFrbBNnsfP7sb2yRGSlZQfjoaWTWOw67Ni4ohNuQki/IBeZi
ABaZ1ZnFs5abZCxui8IVAVW2DX2P4elr0CoW4rAPaFvin2rVHX9wHrwAjLDwpOE/BYWfvxeAqCXe
6L8Tbj+z79pSMzld2YpJKXMGrMHFA6kqroDoWbsjer4Vn2fn0kgD18saAvtjqXr1wrU42kRntb/z
1//bEFJoZbq2akkdZLcVLfr44NF6eoZXUOT1wykjCWkk+zuXB6YIySX6IvTGAZYAk/i3cuIF9CoS
+Akte2DdZ1uduUArH/yWjaTIWer5CNlqqo3tw0THSuxj2VQ7YPLkZzI+fC6Xee6h4z5cYw8G897F
vBPrcNuNsjtbw8ITIjvxsotwuruHnQhGLGUpfdAMjdup+k78L/MugFkvL0S02bAsC1sIUegTu1mE
AZkhi838p3X720XnAz7yc3MNzfcF3z2RrVa02NriYHKVkw320RfL7AG+OuWt49hdFg80qxpePFc+
T2goOgSeUfBgL/1qdkv3TJgWi4KQw9HPT+PD0/GE2PT5Nt1qdQNSySG0SYVQepN/LbSH/lpyOu4z
NgkRJLMEgd9rF1d6N/AZ4T5GtEpPoHGF8bEvsmqdZA4qa4SCSgN43TPWI4acnRVME9Sx0Fhm2LP8
eEKUiuLYFer/ZBL/ufcSDS70h0+0wTihQzVj/K0prF1KehGawCyzKkdMsAzi2nndgZnQIvSg2oVA
rM9rsYzG4AoAp9rEdddO5riIGPPcYJiZGADngat/q+GukxBdqygHy3DfXILBwtq3AtZOY/wZTx20
o/u9IKCgFuQqn6S8CTfwmnl4D7dcnJ9juoYuGKa2iMQ4kn8076IceJ4gmsHa1Ft6uz/XPIg0hqh2
KfR3juM1qhKNWrBRd4qMaXB2OSmR9fCYN7sTSo9vu6fC9DEpHKqgIROuP6yD+G75qeM0R8ukDjgj
LT85l5shKRh2ydxyRzo0trlfjPVMIuKPnhOtDAbR5oseRgS10oKWp9/RdS5bwxdx41R4f8R/fuJW
p9mIZnIzA8uIB8rf9NTVASAAuMq6amtoyk+h4pAlgTaI5eJqQfzZBCOtEeEivMFsBQrP5PL08q87
C/7mF5W3wSKjK1Y3hhRdGqnz6sLG2wt3ZSl07MezUCBunE5iOwYvjSjahaonlRL1cn6jJjpj91Z0
i3cuwsXhN8BzyM51Rv5BCt1DudlLMOzd/TcGIRSxYpUdbJSc2j491ChQfXfI72pmZPoHqTiMVOMb
DtadcKjBTY7TstPJBzv7NEebFvmOhl5uZ6x4VF8fV88KBDLQy3h3U8/6essaY9ZUI3dtxPbPuwer
5TT+StZjKK1xOV0tWijz2LsMFkPBi8B15nkV+vhieER2crXAkyHXwosWHg1WXRX32+hd6CWUmC85
RC0VZvkjEDYlG3cEqNWoiR+2BxuBAI4PN18+e1ns4WhI1JMImKlco3aVPE4qZh6FkWaE8ohOn0+r
+aEZ/NJW9uuCBLZQ099oZjARTYllVGDOpbRl5XfH61JD77zwua12/jiQAQ5EgXp+sKgPZRBTs+y2
AJxDu1bi57OHcPid1peaR3UXezMirI/+yrGJYuBk/YQIrZx0nnML8XhmY0tgHnhwRxKLaVb2Ne9U
M/yhDnU4nzKtQl+lzHsOhTLvD6ih5bNniN7PKpuIG+LhAuBfb8UvPHFnAwi/ry1uF1+UeIAblVPJ
bKEJdhPmo+oCG663UIsIDJDASD+CaF3AdFzp338b1Tf2lRMp/6bSM4w8vtIuJeMImjXtku6Rr5JD
pyuE1juiSQuF+PG7sQ4sSkL25KXqwKY86tnbj2Veio1nWslmgDJj84skUczuI6z9K3VkwbVKsv3W
odn90IqT5Td3w3V8Z/YF7TF3AkZMXWaFLp2daWccQ/wb9txFDRknjWnnUBm1JvGPt4QOQMc9/7py
4/O3FXDafETMgE8Y/iJ1VD2sHW2rEgBAB+Dlr8+rNwp3Z2Ayl46mo6HZk9RX+GR2gnqNCSSwK4hv
sogZdpvvrAqbOaDwx5WR2L1sRVfy/W2QISYFrfVJWBgz+f53tNPjhppu2i4WNjLO58Sp5A+hch1S
y/LrRzgOYWt+lIapNZ3qK868b3MMsRLmPEA9ZeO72LbA1H68GegEEfjqwKPKJW6otjy/znFbRK2m
83e5AqgriIbSwok/tu8Nm+MvyEkAxnqMROfOzW5FaV6KIMTC7tPY4j/dFB4ls8QuJSgruGA2fqAk
yDkK3xmehtO6qIlRwgfGhpstmnUHIlcVm1QrwvSw0ciWWuf4joSX3k1GtujletoO5+qVEi0onoms
MZfHaE/ElaXzj3cQcE3UnS/1ARtTLZpyJWQvWXbszA/xSJrT7XTmORiC+NKFnJJo0VVYOCF1q0jG
UatMSztqTmYegExov/fe4YvSO7k80aH3/nMuJoMo3KX/OuEij09erIB5eZch+WVvbaaaTa8JFah/
uELMsGi0UUK2goqs+epifEJlR1f5qz6Wo4RYC9ln22Fi2FzuaJ5EgZ2TI/hiU/m8/2MIhpRfrlSG
WRiWvJ959+sYzVN9Z3ZElaPGRx+/IboUbmDozy3MnL17HAuJ6kXPHDbZHjSm55arh8+GoC9/Jfhr
vRqprvht/mJiCjAmrjUN9jy6kA2vbDS1fgmFNsr72MTN0mo4UraDpJGI/qD64V59mIWKhbu8Yo6O
I2oJ0c1akbEpS8rrWRpEFwLROPttYcU0HLNj61cuNQejDlVAM9+KgU5SJDmABzYU4DN75Syzuwg1
w3yC8tr8xXWEAueurAdOsAeb//YpDAAesl7IkEc+ZIWcZS3tW9EPqiXVmegKeR7pReaiapnuWV6M
UEYiMb0aTpazMCcPh9DKJLiDPSPswzv+ADE0zIB6o13S/ScNq94fCJRk5Wd5fctPjugN4ZWRprVc
JSuN0XTxsMwKV8ftfZ6R2JXmClUa1msUulofuPghwnt8nKho1EIvDH8OAgBLXnra0Ni9y+LhUw39
boguvg0Tlvs3NseqGJ46NqoiWXcn1reQoK2PJBfOdhOmnHSe0ULt7t85PPv6REjUszjSUdrAt6Ey
/s+kYwd70UJ3BOzYVocUS+XgVXPY2WU0G8Rif9NcPiYVqR5ue6ghkQXdVSwKERQxYQozYIOk5qLC
x2WM3ij+hU4VG/ACawdtN+HhZyqWix0arhAgZHPXyCkOQAy5211VEUXgBBqTxOQYkq5ZrCf6Znuj
JQAvhiaEFsEGYpmRLbZ5d1BKEOCdrrhEo7r+ka9FfUh+HskeJMUl8F5jEbpoTGRZbUPmoL2+9qp+
DXADF4owdLPRJi1GDgt++T9KO4PS99PYFgDWiy6hZexZVu2Xa5jx9zC2pzYvXx0VLzRPBxovpQ0+
BNwooOiMjunvE8q6YG49hJhbourGtN4L6I1lhO/C3ql6oCHUmgYQ0zxe/AtrDYGdH8P2QdYTv+YH
xlMS9zG0vhg4OGILcPptbTirN0AwrEV3ebhqrxAh8nW5eI30Aom5H9zNUVMpWcpMJOCHUIzku2OA
+t2qVGsoiZM4WW9vZ/XNtzJ0LtMqdUNxwg4pRHqlD04AolXn1uyjhYXtPohTvPVpcSbQbHYA/+Nr
SjF2NNECFi4MdauC1P8EpWWtioYAIUaQza0najG8KDO1Q0xnUYj61+dTcPfALYIdxMGrHbCv0Jr4
nEx20MPqsN+2zZ2nMXwZyaKBSt7StRCzRXsG4nbE79z3jmEhkJiVIu83eJsNN+/EwLCyhSW+ih+r
scD0txngHR5cZbU+st73z6ZbRM9Je5vQ50HAT6kTaMHDM9CsHMZo3yuL4DPAIC3xDORp9brZ55/Q
2YvSVnuGP5ZpCuDdNw9t2LYw3Bdd9X+sAq93HNXu987j7BNW7wxmnwp8bjFdQmQPLDD01qjwb0w2
IEzY5T35E7FFxFeRPmWCmhMES9lcxmN5ytnaMTaTvZV/Uv4wyO1LvBcUErnz7EsbCAz7PgvVivuB
9f7gzOuTUcsrFBW7cRrrXnVdEegwkWZDD8Qik6TmhYRuQ7ZPA1kInVO9erZlbSdSHQkuHs0ZVE9F
D2XomG0kOwbSraXNfgSXShiEbS1X2nR7SUtgffMg+BnZ147eHC2eGDiqu013+kF8w+0lZHR5R39g
MLsLYgcHewU4pA/PBtYXjs2ussZa+jmgbYRQI1OBMbHWo6LPxZFUvUI67bNOwj+M6ORw8qM/7LSv
uc6jZQCfQT+ucTFUXcmLG1Uqg9+royjWqQGUR30VBssEVVzzlayitlINNKumF0tj6wSbMhqbD62w
y4jG4z7DAZLepq5M3+U+Tu1n+vnTf8rU/F0zrQYoABF8O7PKXIes+l5P0ppqowMbhyFpd9nKPexU
fJrjzAczvTrVwXMJ3J+CQHNBW/nXK/SP+iVodAJ83yqNLhPWVmLVg03xqfChUC5C0KD3DjZzqYIr
h80+O22U3sdDZfajQNWffd+QdTQLMu8v8X/sB8LCrNnZYTVghv7eYd9wDjNNPSNQJh1x8x+L2m59
huesYExK081r3Ymtatpx5U7k2W97wS7g8rBVRn4VPyhfyKHs04zqAA+PCOoOcn1ibqS1BwgaXo2A
gsgEC+ohep0bockSJ1tuOjAj9Qv6ktweax5xVNqAkIqvPonFrN4fro1c66JfWh66SOi3QPrhMcry
MZtb22G0kH9AdHbKdn/BgEXhfoxGWAdqROA38CqASwJ1d37to76cWk6lOz36wsJhTC0Izz50TiYl
1FPfN5wKZ+mCvtZISxWCGpnH2De7uFz+z5aBGXUzznv7fHvr/wN63PHtE+Il3qDI+WZGIPrsEJhS
GZA4uuKd9Nup4g8lvHlYhHglAg+HHof1pVXyhXT8Hc4j5V4rYxGjnpdmxczcxXZqPS8kkuPgR9Ou
EwREjTtEhfH5xuQfLjoL6Bw7SMm/ZkFizUGE/fwyuSlWQwfeaHQwEsEneNHAjKKFH/Oc34P+WoFN
3w/RUPijEAT0MqLVxLY1vNjrdLg2tbzqdkX5I6M4q+i0BkJJNgVx83n8QQH52zczFKdZZNd5CSIK
boMqQEyWN4vkvgZORjudgBT0Wx5axu8jiYu0tf8ZTBY41lrg5gzQlvCsaNTXqPgvxOhy8VsoNu1V
u9sqpCxrKuigqBf//JJ3PHJJlHi2NvAF/cod3PtnGmhKjVj+Z6S/lHqFD59gAo8ssOAcnMG9zvvs
+4vFuaYb5YqU4JqfT2M83XuZvxNuoRaa3125RHX2Lc+2OusFw3oc1B77mmCvrximDqjsOQ0kf2SP
xi6gVX0ox+SV09kWtYg8UC3lwv51B2cdJtghd+fo/WAsjFdr+C3KcrEx0u7Y3/Es1lMa+BKMIQWT
LCALLSsw9+IzwJuNTbMU4wV8qV3JDzPYHtToenpMjg5po3LUwxQKl6DQqngNw4MwKb+BwYEVNmUH
cMqHU/8zeG8nRdut+EWEXDrWyY9an1Yn0fMMgO0oQ/qEUo3qvBARu+L4kBBEThWw0/7HZjeIY11q
YFxCHzqZ4JI+ARbOK9Str9Zg0r67S74OcFSEpQWEgxDSFhsKvsL5muPG35yVM8Ix59DioONIxKqM
v3HnjlNjgeNJyqJRalVJCx0B4Ggdh8ySUPQuCr44v5yoTR77EOCWOJ/3ibEo0qS9VjzVjm8t6ovL
IwQd0Ao4wzaIY1qewfm8szfz9cFl7RuhrZepcddfDNM9F+ceZoUMWarEaBakrWs/A+TcALq1i4rI
6M0kHOKr9OuLwd4mpAE8IErB4M7hYPrxpG9FtXNtdUuahbBHEmmXmWa6u7bIh0i14Uh4J3SasrtL
Oe8AVPQnRe6i2WEc7eXZHlOBVEw5zW3wLMciS6sbCCtL0CuVptvuSWUp2qwxFrJ9VsxNA7ROOGli
0/4CTtJfcnI/G95+UGodjccOJiZ0/9rq/egisJ6RySwFbaht1jUtTqJkMWMDayr/RVXU8p3FD8FL
WRobM85GMwEEEy8iEMOskGOnIdeEANKMHLt9nRTKA+Mm625Cf8AKqvPH6ISn/TR7GWRFzBPdUNJA
8TCDkKFA6L+z+Yq9FSubM/8/p6QiNsqDDHgyu+rf9Gkc9acz/zj6+xjtAqvcfyYT0ksmhL2I5JB9
W/3a535zAvBbM+lWNM0T4c5JGsjZLTPcSbWOfGSpfIiVVLVcV2/V6X4D7gLAnpZ93RkoBDtExjrs
71mHYbaH48kfrMXDoQVC7xybcHavvQHD0nOazklq5UJ/mXfpxpI+iyhnMr0GpOz2+z3zE5adO9CW
8gIMd3p3hBCpQi7CMmWPTOtafAvgY99i5EGJLEMo3aTTsHkvEQzRRPVoWkgn2qJQ2yuAOUUbk/hk
oQ2iYwiqs21vuCIp0wrHCYMpippjao1jUWQFtksNPi78yy+srhf29MPa8N0UjQkq9WFJMrPaaM1w
cRTsf8gDEyXZJAfTCeOAkCGYvQxPXCRhw+NLNE2jP2CU2cSPFdSVbSmkzXpbdzzbvxJsdBa4D17M
zFNdQqCFlIWNkXi6K01zvUmi2169BmGi69IMaqP77ZgCdp1oVsloxnoXdR5Ac5Ju0oe+2ESFgFSL
s76YSOp60f1u1hNQbKQyanycQ5Xnp7DyxNWSF16WWVwthuvclxU5MPkS9MqLSzRV1r921xhpAU6H
LjLidoGY3pF/Dsphg8gqwwr+vqIovDxZ9KvFXag/1WOq+hal2zNqXltQLI84/kmCI5KV3/Vqy7mw
uA3VUE5xkxOi8VOkPEf3BZcl8kQGkWynqElX2z40e8OsG09l9o3Ih2kAA83DOQgROc1tvzkqQbqm
exooLZd0tplqDhObr9BBEilFNevN8dwOS2wvlj0lkXslqMb9PiraI1nkGs8XDbpi8h2hQNUqhE1A
KQIYsex7aGKGBWpdlcZiG2s56cxRrh6v1nKF1EckQWCU8BRxSFDgrma7XrqYopUCMFf3N+79kWt2
Z92cNcGU1a44qU1Dp1oHziXBRcMx8VataRaXxixtPfennw1s8qNMNDDY6Hk33mLXgGMzBC/Y19+K
dJjavwGwKuTHAuPWKOTPfe3xqOTdg5LReJV0VWVrELDAZe8awQanDcAM2rbHUV8QLMm5EcgklgE1
IvqsA3ktC/iJlxWXAdvHWPYpGJZR3M/yuwyS5RJv8plNmEyREX/r5HSV0hRXrf6t8xRMlP/96CyT
RvjKR+6gfJByIg2DG1d81JlS9FoZ8DY76WwpIEJGpnQdKgeBPFfy3LkESnP13LcWBp/NumxgC9cp
8mwFyVVOrE9GI6bHoltxqOP0sC3OrlrFtXr5f8Jj2BxtDaFZ+MLCTOtNFBQlG6yfq1IAuQ9/kCdv
kNGVzr17JIbNxKxFPc/6WzPk47s9yLpFepXX3/eVt3N2UWSJv8h0gqEdYTM3mUkwdHOYHTBvH8jw
9jzMl9qr5azvpNRABCEnSM+vO2EDGMPyNbw8PNFTjUPqsZWcjBRLw0K+qIlAYeKiJv6UE76j9NTM
+F27iztO/5vrEjR8UXrZuQnj34vSOBIU87i4qJyo2TqUneGhhTHvoGixCSk1SpF0jbUsiQ4UhKjo
EOLMHfc0w6d0A7hAnnyJpcBrPEZq1vzXG8SRQ8rCa+pwKp8K7Ovbv7AkbHxq3pvsDjlgV8G2rfto
2ZIql9l9aS2yZ7YH65ZM6B3rwOf8Q4D6pnLLt+5g+oura+60Y++5VT2miyogLuR/WCgIx+XxPeYi
shzg52+ifWw/J44Z6hhFUYWh/tFuo+rbibga9i/TLzkHgHyKE7Sxom/9c+oMIP5DlLayCwIU3mXI
L/hv+X/+dp4iyQ03Q4ioqb6VsfHMvZN1OXWdloW+6J9cMLBnxEm36J7XsbGjvyE96wB1/xPtNbUc
FuZRHULZeLJ6e1i+joiN94ydHmk4fYIN7jh9DeSUw5nQKHki3+UBS7KZouUVvv9YNZRcj617yVZx
Fh24Oo7nEwBjKi6lu1HFaZgRX1bQQNkqypODU/autQ3up+auw6jHsuVnkCksgaScxkektBraIjGJ
54iIHQwYEFs5YL8qdFjzzRgqzOi58neySSd28vth2uihuHKhK0ibV2ahQNIi+1uCK3IzHg3ZEVH1
3VrqWrFQEcE47rztEpe5svQVhlZDlkcTZIpNAOhy3toY4ZOFKHB2MgPxJ9hW7qw9odDAtrc32ASK
dKBjkM5AsFNGpRmbEe1tZmrgcZlITnUE6oiJDWflOCVccd6cnMuCDbL8Q2HdIEbq+VHixDQ7NM9I
LmqZIdX6dMkKecsQwB+mM0N5BDs0oXc1zJD6sffCWLbF7xgyz4t98ZOjfwYWGKho9+Kl88CuWjr8
hpd4uwbcf5HHA0VqGjqfY6Hgz/mUYmNtIb0McE5os6+K7UYjqbxrV2WkLo4PsD5BMHjN85KqGXOG
eVZtwi29nil5QcWeLc0+9rBkYh+YIyNusEpYbjRE0CpvBrIeNElnJBFZuKml3bLq4nPXWsLaeIVe
m2U7H5vju1o/dUCEtZxKhtOWamBR6QzlOhN5gyTGOiyKF4czyHfU/9Veuap/TKaV4/KvkXB8DnZe
bRowuyd5BmAkX/1W7hkbiQK66nGHl5PZRjS0b7jhvERLr2b8jk/r1pbVgbgB97m2A1Gu2ten5qUh
y7QWGGBKWlL5mV5oeL1x5RHFNAErYx43hFJVRIyM7G6oId1sKHb1ksTKwLq4EgQn44IeY2/QgYO8
l6dwcjuk3FSLitWz1Q//uLjpw+a97MOzJEdIY1cQXymQMZXR9CUZdihiKD/gLoqJM3Uyen3n5725
bWaY8FjopYzXixcRBmcXxKhjxntHLyb9h8fc8/+zF9i+I9T3q8PgYYWatV7DhYT4AwgSCvLEJjkc
JBKFdpm7d+oiXS0Jlzj7tof8rz+izsdoNcwHQR0xN9RTfxAG785VFFx9GTZxLD3yDzml6j9MYJRX
KISI7fpPOmb3Zkv2VBg//Aw7/tnNhvgOq7lGMgQozl2HudgZlezwuzxN6sXh1YkH2VQZn1Ki3R3s
ztH/Jl341/EO23snXRM3ula0Vi+4Xr23MKfC30aKS2F1850r2pPsk+EnJfnMx86eOdiVjwTuuhg0
W8YbkdkVbM69TtFAJf+48UuNO10YJzRhkw6a7P9Ig8bsAV9o+inp1qqLAFrE5DjyRha64iJiQGX9
etcYsBRgmzmv++PZITaBh8eBINMsEKQaX7Z/bdOc1FBWOIo/nBzFWZiLr7rnvWONtUgn0U7q0r+W
stHY3zvmWOdNDplbnccOUyPRXiDfrb6bZ/uNFhopnKyJ6xL2AiDpNrrrLjJDzaKBTpQMUBUtg4l+
i3bXsTP4kePbwaWKCeqKLucpCpcj0hOyaxPu+R+PaeMawvtrRm1eABXai44IZImvqQArAY+sg7h/
HZahFxFvFfzmxPcB9zZLnM73pibBII8IfLfWY4Vk0wsxBmIf+ElwCt1Z7MEtJQXBXlZoWuDI/TId
y5VRAvWp5auvkeWX1lpwssjhTgoZRfcS4EXRrd6mcTUbH4r6trv18adOvOvg6wmftHDYEEvF2sqh
4nDPTCHgUy/Qat9JwYQYfvFXBZEOamVZKBwDwkZNymPyu8Z7V7P6oQVG7nVzCdc+A4rPyEGFa6EC
cOHnGRbqVh18FWSZCkKi4NostKLl5fmWLnbRfmw5LlyLefgiVMXSlWedibb2lBL/kScOXp3nyTCx
9dqxAohhSMTvQpntAEcwqeFuB405AGnxBRv5c5aDfkof7YR2cxbViwJUhiLMFpkpt1P1NVZKz6k6
yNrcqBCuk81FcxS0ghu76o8vauXAur0ItsaHHbT+iJr6NLLm1KgoNrRQWVZ70FWFCagWXHZQBp6Y
f9fu36EzNYd6RvkA8hN3Dr2+CBI87TAJwWZE8gvOaP1LZpua23n6kYJDsEkWP1E222ZrJA==
`protect end_protected
