`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GplHQla0/m/CwlfewCN1SdUpaj4cuYlZ7bKQE8x/mBHO5hfpzxYcmKgaqazxtLZECKug2knLjhMs
ObxNVk1cAQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OeRsX/GllKXguMkeKw5EX0QVQ1GCXeGgs1qHv0V5DaCN7bl5QyYmMgELN88U4OFCYTBZY0r1Dm1V
hCU+zmiqH0rtgyr473TUBJEAPJI/mkNhEUiDthjCwJNSX7J6mcgCH7fwoozTX6am6Q+Qw1AyQYRA
/BdkmSjLYHFhCHNOtEU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nqoVmwPqq6CMSmIhdUJBD81jiU0Hzx0e4tXRYZc+/F2K8w3s8m4Uu8jSgfOKTIKRn6rFRK2qUkX7
f18wMF5ipruP0f3qhYDfJRluM5lKPZCw7Od/pRYx6qErmYqyXbmIpW7Q2LNb7ovaGP2Jgo304/fD
E41r8pCOQLqlYeKmNQYOSNccq0Xq6Xue1PY2pn+ziFFdKn++gCdVHnXsHFXEpXI1sUrhRIPwNTIZ
ZKApPTLgVE6vEJEXozTO89ieQ1VsTUsF1taLUGuPhY6SxUxTcScBHwPZt4JzzmSVA62pdSdvAUKF
o3LA5gSlDKFxTX7uvpnfpzVoG4FtJN5vfrw7Uw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
El82/FQ/3BPaOD8uZnQXKqCbJI6uVL8XP9kNtBxJi330wKNZ7PnX9kFKSpIwlVMuBTpKI74IZWMg
3c06pWKE7mY2HHCDahU5habfiEc2Zvrw9K5+EiQS+T+cJsf/bGf0o/8hkatZgeK4GXGXPR48moDJ
5xrTJmkKpFqmx1uCNyM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iVM7GAi7BM+FFWo9wXjdrLm/uaRGfmVjKCnpM5+SgvQkvcAIKvraBC2k9IEsd4NAb22Fhma3QqRf
OTCyN1hxhaj9/n6vvT7cq2Ppqwf31cV5+xllumebu7oQ0g0gRxL1DnmyzTbT3dhAsBrPtw8U8x7t
vO6chTc4HH2HBVRQmd55GUTdG/I7mNx95lFxNHgX3DKB8qkMaMsyDbZ+jcr/jjTv4eE5a76ArZRJ
3aeobOfnQdAacawwdVx+FA94sqT/Zj45ieeODR7TfF6zktmHvVN3KKU5Ukt0yS5KhLNiXLOcH/2Z
6j1HPw8w/tqm7ceVS/dl6hbfwRfrlfWPRvan0g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14400)
`protect data_block
e5HkF8V5ACC6etq6M+WDp3IzydQAmYBJjppbDXMo5W2o8z19FxOmN8EjUnVpS9+BHaz4BWcCmz7w
iKIApJvTcPrdhT3UxXWlxM652o93i88geRcjhx1Xs17sz27yexWmTFNoFOJ2F/28XOVag15u8Fm3
Ylsye3ItKmq5jokaOE6RrYZnqyeez3MfVXyvp+JvaxydpS4dY9ikn0BI/+Ttxsoonikpf0xvWDnb
wkpLbkETbFM+ZcX688UnaDFgJnWzywmrCQJYokm+RvNq9MK1X+1vrLesNZN7fJsgmNbGuafvlIDY
D/mrTbxZBSHSAg9ycmAWGqCRs4Gx4nQ4T4SiQa0dVTcvY4WKohhICiz3MZrRoZGwFbUZjdv6Xge6
Nz5YztN5ag3FNO5FjNOzCoxR0FQ8sQw8AP9GgXgC4cT0m825NrKsnrXd7hEwac9P2Mszf+DAIySA
/AbshfwdyUPU8iwz1F52wjFi9hPMfAhR06XIF03e2cDlstgtundI1X9js7yS12hL/isCVFkUFHZZ
zL+ug5yk3Z1aTlvXDpl/V+ongL3fDnPYAf/0Nq+tdwnhahBCG68+k54aUriwvgn6Bdn7X5cp21dt
uNKMukofnrjc6USEPVPo0LnDZDUP9jVvAxL0GUAbAOop47VSl3ZlrXObi75I5vkIwfjNbmROoEfM
QyyW3Ck6kCC4BWNCXJHkYei/iCPNYD6nVfamEdbqvaV3/v+66vIRaGxdLfhGgoEp39RipZNiZ6xl
5O+4PwkCZ0LOC4mCqQ/ftJRxaJJXa2a6nRtdwiq5nyDLolMWvTBuxXS052BE6lLDwYNKlFH32jRN
P/DLP3H4EV3M9OCiXCIB/0YvnaPgq5xt+ITXWWoi7Rt7R20NsDyaexoKfnS45n5QLHZha9duatmO
XcBpxEpcqr9DoesXRRPai2NxTltYbcpRnr846QQwF+l9lt9gLG2fWBrFPNGhWiOZvh/CEYzG2w0T
lwJaab7hW6d1ZwfmMhz+8hKdUfUHBj15/MmKo7Fo65JNXwfdROP0AFB6390ZF6igsaP+uK63t4p0
K0tfm5te4tNOWE34dlInNrvo9/lOfQtTOiSsHKF7xIhBLHza6OR/mZFDBYg7v3Fg9ZSft2+yyi+s
AjKNiBflt9g3h1h11VnZsk4j10sctivkHNjO3DndWEXG0bHFjBkzxb7EByP4+noa4NdafViqC0Pi
T3kMwstuQwcvqLMm/xvMvCK2pyJgLSPavVRWGnu4auWGpTQpCM4BLdLsDmU+SVfk5NZg8E2U6oin
elrKNqPyNxML4a9BLW3evnz3zuFNw971AxsYef4BQbxdstwG+RWJCs06rO/vfSaWrHIcyzDr2dbf
07hyVopHbOMLgu2DLUx1DfQ+nE1SlQ7UYk/qP0o7s1Oph50+ca7RlK9PhCfvOB0WjEoQAge0AQNs
tdM6aovabE0TtHzZgGTQ+SXRb/o/bWdbJYaV74Vi+xfGGI82zITKzmIsXaBAy77YgVj8B1Ev81Ue
poceQZ2X1NabvsO8MRzKPn5ggMydyl99ZR3H4LPcE8sduB4MeJhSTqiAVkpn3e8OEg7QdMu37JJL
2z4ECE95aqWCCAhV6HGlBsAMxRB9sqUcKz3cR/PaV3nV8HE65LNSjimlw5QtOklmBMT6BkiDX53J
Lp5p0HeJzQBUADZNh9+iACA71LAgnDsoEFLcketxy1m5QAqZmf3WqMtnplI+wdgMRpg9KL0QEjvX
L2ULmJ32XMKE93FcUWDf85mNSyMIQEIPWq/lY725Qad2kV9U3VVXqr933q1O0iQOFy+PaK7DRB3r
HnuxqHwOPrNcHY8N+PfiBp+ucGY9CTBmWF6wiOWEECw5iBpWEC2ABoLxIB793C38AXhUhWb/cBrk
cYoN1+iRMFqfXNn4s60gJ6Cyw03jhpoocSy4uW1v/r4Z1xxYYppzlpfAEl/lDzVkEmb5WvL+9VFa
sb3iuc+LZMwnaToaqob0ZWMwl5D4Ypb2VHuOcYEfG4A8AwVzqCcF3GZgds8DDtn1atdzv90UVz75
rTUY7uUFdMY+zAz8VJiqigYZ3gwMn1Jj6CDfbGHq8oQHf5NGVUx9j9EqApATYxDZLKkUo0hFP7Yf
LlsJ/xLYsm1nzbgX5VMDoAVnbwP+f4zRv2CeNLyvD7ffaiiYyCeSWDPY5zEIbvS+gRxZ6tcvMRWW
JmCvIA4ZEVWl+gmP9nvrzNS4osFmMlsiKIuZjRULcsMB+NGwIQfbM64HSQ0UD8wliLnGU5FBmiDI
O/Kc/v9zLvaRA5AX8Umo0SmJBnmFJm0ThqPwBDo88HcCwvnV/XlvqeiZiQQUnb6WoDxUrZcMewEZ
ty2p4RhZjfuXsSB4+k8GSq1oBykoWcUXtOkRX8TZDuklP+q3DIle1Ckgf8/tFj6DohABk88z5txB
d0zHqkcvYNjZ/YnfNGTADe7uq9B3HwD/GOQ5f2k/MU/lIKeMi5GxsoXdKKh7DUfiyv6qRrHUc9Rs
EwToUKAmJYvqib3XdoWgVxVhSiz75kVgFEziR6Hy7oEQNI1KSek5wSgGmRQoEj4ddLF2XcUfCjcK
3hiqt/BYttldO+EXtuFufSqhEjOMngOuNVF4jYxAnbMYn66IK2xfNtQEjJP4XucdpIhf/GGYoIro
0ov5FnGceRD4/+dT/DNuCRZQhWFlvMdrg16dXdJkFpJwJ+oZ2MnNNOAWfk/LqyTwcTBOuWcOEAp0
JvR4VQHx8U/P53H+qqtP6NagiFAD+TiMKn0gF4jTu2CSVtYH8wP0BDehv4J74mIeigVgjt7hqjaF
BJaowxZeQvbeAYBG27/7lo9dUTduNN9PZmXcszR0rDFbKBNZA03jwChtmruor7UYzKY4G11YLM73
hSxyQlhK6NPbDMN3ioG1NKlx/Uex7YN9Kwi+3YXf9afqanjcsqiqqsmfRnZB+8jo6VxSXZKlgXQK
9U278UjZfmmR0dwFnJswa0pJpQUk5QaBEYwQl/zGL1hIBB3UpWCFtbVWXoBu0hOHB2y0/giOF4sR
RhFEsUVisd7YWPpFNmbfcJgyP/drrQbURg4zS2ntvlu8iNOBa/d6wut2aOZT9/e8yLo4f780XY70
u77WbfLsbURFHM2+DLlmD0MmH34LG27rZgwEM9FzfZx1kZbrTnqISK+arYwQFbHI5WnCxwhVnkND
HPzK3GQDczZvAw4C5xKUFatqxANyISXM9l3slKXksob4hzxW+N+IMkyYpQfF3IJ/lRY1HIDZCmEL
837ZOcUGBzZMacdChz39od8qc/53/VNZkXCKrHSkrrvXEKWdoqmPCbWcT5TG4/qjH/5koN3oHM/+
keM5Dsx6T7EH2UFoLBmq5JmTJqLfMqmAbYRPgMwBSO2wuOqdVfhEXILk9UvY6nlHGn8odI7ySTVa
jV1hpmO1ipKFrpdLATlHpBsQjLY5ki9lEFZhAfNRLFdcwJrIuJv9dO5JeozqM9gkoOL0hAR90Nas
fwc1nH637Z0Q/5S24vc9I4Y1ugS49rQLy4VYEL2CoL8TNtFPrqz6npbGvLKe1oKNWrgeBzuPznGz
QeknBxG9tn1qkghv8j43irxiX5bTdV7S6t/Np+oNZrAdvAzptpVtoGJqkSfvbt8iXnnMbaiYk2eW
nGpiXA6Mo8nNAkrSa/MdGXVEaZQSFsKVCxsRVknxCvX8dDuLe5dOVt27B7fc3Xb/dOV5Ev4fcENl
4pWkHPlY5UWKT5XWf6kF7ikYGHdkTXsYn++ZCGVJgnTO7LNLaVrqGDwHqyohtY7osEIYHDzOBn5/
zXL9g/5k71wNvIEyzCrT7AIXkko7i5ErwtoToefg513EFbSIUBEvi/raQa5K32DCx929CtPWE6DC
AnjrH2PpAGdZAdCkyBPc+GvLCIxcuEAHZJBuR+o1ybMNE/t4nAWKH1MscTbPVaE2wPnaiRfzDj8P
VGpFK0kaJ4i870DLM0WVaqdct+gMG8JE7Ba553PNeBG7l/o1jTkDafEoz9grSsbR362g79RR/QB0
oN9FcM2a+9ASp4IHzXwF0etkqw8/rHa2/eywzhe7XDEOrglNXD40yh9lCAbRNUvrV5YChGLZjSWY
wuvkVzWgfqQYLJa/7vhNZeZ++tbTHjionXqU8lqlXgZpM65Wio+Bynhfc4L2i8m59QvAjhn6sdOM
3NwQFIq9t1CUQvEEzhD929SR//63pu2NqMWx1cAuBzWGb7uBnJ9iLGjr2esE+iK4anTVmclU/IgE
QZAYMgXKkwqavyfaQwLEZKO7Jyg7Ul0z+aI50h3BeBJnDllnyBPud3NBaRs1NGQuMd/F2zXpDQoE
/eJSgddyig/c8ZSwezIDTlMO9QDjLrgirjf/4gXOzLt5I+SjtIHSMlBJqhI0r9BDDB6RXjwGjNff
+q7ENEPLBrTynvxBem4epzTux5b1lmV0JKQkvcWsGwyLeM4FL6YsX5/eT3fedtA3kbeJkthUnMnE
0BCS0jgr+HVybHyb0d08yr9al4xzYejoSAxv0Y7I7TDUHZyXZoEM6rmbqVp0Z+DHaSZjwUu6MPLq
GmYVIey7GUMHwA9EiJexFwTvGMaTnMYEBfeY5m8VDcPxB3D65La5cJIZFvVexVStutpxnnMrpYKf
vZ7s6Koh7JRjFr6Ll7PDb9AzNiA+OuRKW1l0uY5ZNRkel7ih0Di9YeG+b2IvRPYAN38bbG2u3iX2
zgHvTnsGRf3a+rbK9MVbQAJ3ZKa9+dGhn1AFphEjgUBpU0cb7vr+vqmRWl9S9gydae2ntq4tiGAk
T8wtAQfQBTcRD2iR6vDF2+2/AUVKbMAfYJoap/3PJZuEHfF4v/P47gpZi6BoxuXszytDFiK+4yY2
Z2eIi145jNnFcgvRglEYCmO/bpWjeucaAVmPAHTdI9+ZbLvPzzI70HVaoh7YK+U5IChyh5sYdBWw
C45CtrL7+flu/u0KJpSMpuEvhN/Ti8/E3vbJ+moN42ZmpNGHW2E8/nFJ1p1n+L7lVTXmuVPlm2dr
RN4JJIWWGTZT2t1Ld3opXINe1tLm//DxC5nlffU2M7dokvjr/3ELZ83QFGXFUIA/+v+vwu9RpHFh
tcbKP/uFtvuNgG0cK22zami7PfcY6jyCoQOfW5OTM7EPZoUjoyef4CpoLrqwKvgW5xqmHmyGL5mD
t0oIRZuAOOc2ucMZecLXZ2xflHHWkb/5KIaoqIHIbzAw8lsbnFRvW2fmdpH/QoQgZEchmQ1kZ+lk
BoLVTMO8SnROlAvJS22kvBubpHwT4OQTw1qyzWgFD6ZhgHN3c1OJHiUA7TpksP+HRTInmwcaQ2yG
AZ941btaoN/UY1NwXCoAGCqDnn7YeH4TZbjiYyPu0cX5Cyqw/S5kSdleSAGMG1O5FoAQJIv+YDMP
T93UhcNLrB85/C+aC9mNQVvCRp5ThMEfeoHuAkV7CUNo4MMmOrzMIl8prvVS4BVGQY/GlxcjJL4t
nYvz/CIb5fCyh9wpjgS7CeYMQ+x/mdYfxgM0QZ2DPGtYwZDP3TwbWM/p8cYwdBULdJFg4UA4YYjz
NOzmx1+2dm9QJhvk0s57khd7mjbei9s3wCGX0Xh7nHEQ0fbWOGrhYVsndIIsXIKmp4Q5H8ffAblm
ECgqBIqypFFt/0ggXUapqWZc6ct3xaIeumNbOg0VtPbMf3oXvPpnsx2eZeoAjkWxCK0vAziwDdpw
3ihu8ETiTXKkrw94nJbE0qkI+/1Mz1Piv8vj2xixqQh1KmAxzjdOorR8O906jeSFaVvMkn1AKgMH
DVfLwdHKBcXZv5tLfHPeEs2rHs1gMenQRPmleOIr6SOuZE8lBOaOQ4fmQSsnwQYGN99BquIfmeDc
Sn1ATQ4YdDxJSjpQXtnb1FjHwvVDNEj0QPkH+/s2J3wtymB4bIkgVmIAKk7abEAH002ymMRDqixw
FahlwaNzxBUDaYoQCXlI7+nnqHTDRi8sfkqbB2/Imp3/8ikT///c6mV6f54j3JmUAwQxlfcxSKfK
gbwfbpk+6FXgxt82pEWBTfc9p/1scKpV6lCeweHlZsGXizryd4ONqSkAJdyHmXIy+YZvQmH+Do+N
DJzRhEbze77CWBqY0QADcKIBDDM2vxuS6pk5SpHhOybphP0Dp07AvPxrn+i/lZUPMuAOFvkxtWoE
g3SOhDDnNGqa3mqi+U29+IjAy0jMgA3/kh1Jj4LrdTX+Umtc34PGptXNMyibUOVDYdxhThAsFUhw
v6u9yvMULfBcOxm2parjCqY9OaFR1MOK3kJaLm7w2dFd5KkRjj91mTwcrMcPEn76OymjDMVNzXd/
6ViPSlgkn119xucleWETFMPy73URvv8b0tTfh3AtKHeJ/Coxr+D/cUyy9pwETgNwIYNRJsxk5zj3
RpsQr9gOEHIcxKh3Zj1YTHgi0tSyrfICuC+ngZuv3/6UHHPyZlHcAkapNvSh9JvheAcqgbnQ/81w
55HupMmIelnI8y1Xu5KSBcIVLYRAYmqZZxam8yklA/Rmc9qDTtMftQEOCMhnkN8Xeasvq7efEsAW
YNCIPmkfCRVx+D08yQ7YfUmfkiFtf5vGGTR+3aiOKfVbjOYgXg7QUNhHDZFwqwA+Mw4hA0uoRNZU
YOz7sy4wNXjeir2lLvxfk3hhmzc4G7OQJgYo1JkEhqfVmuZZ1usZOUHe3r4QvF2/HdSVXEIXQ2JG
O6RkapRgmbvn6runrtsLYZrZT/rr0kRFQz/tkrkOHduAzSjGFRcxL44YjfFCdEuiuMfqPGGQhH2d
T5BseumVrunud/HIHbSZZ0pt04ER1GqhyDH1gWnfkVrr1onfkMbS9FZsg+pO+5wJ9cEaOuCS/1HE
+vIpcvR/+vewTtijDHk7ErHhQGjHyCFtpAm0SPw7looi7fRvWN1p30OHgHkkkiJdjj5d5Etsqcsl
+L2KCiTKdafZXkjFLAHqSEqGHttIQj3CaivBfXjySyRRKGJd7hjNvcFbL/JboQdI00rFfn71gKxn
doLgSp82Z3njJ0wwoj0Us4mDmrMy538CYxtEdI1b9heTBh1vQOTiDkPJuS3G1lNkXO8L+LF7vXQM
xiFwVhRkyPEF4VSkce2ThJz47XLrbN6vdn8DE3TfGpEIpoWI/rGqKI1njhkn/m51FARRxk/DEMB0
ZwgJ9L89hxhSsojol2orfBH+eThR7vmjq5VB7LGIbAJ474aXK73X2f5fMbXpdTHO4u5T1WcmUpq0
fuY7+k0p/F+CjeeBV+uWdAMly2Xl8kBTEN8iyGYovTsuu3D575ibsATvEyPrcDxLWEInbVduReQT
zry4jk2JOGrWDBmuESU2CV7znh20tD0xZhjc+7DPBrd/FV0DeO4hkl7LrmL4jXIgOBaJCYI5m0SK
ELIdZJcbGCo686wfUkF6bM7P+RKUJIqbfLbAKq/JghWjLxa9EWONETF+9icGPvsOdEYe4phE49nv
gj7j3g4Fse2lqqJBmhAECSWtNjK9r85ER61JbrnatOCiKI1Pr3tONjjGoA3PdiL39fnKWAwCoEdf
kDaWDwNItcTiknSZGwOhLjaiWDP8yil17XpahDatt/UqdGiji5UG43dr3S4cCRqbWBcQVEbSb23g
d4aL69Wmd8J3QMtX5TdTE/c7h0pgOvfdtZDEDDLyGVXMaVQetAeJy4Z325idzzgr+3z6drQJYsZ2
zWO6D+9SRtMjv6GW5M+tgB/yn4d5trJ7nCF9emizg3y5NYQN7uYij6grZi5h8AUYgXUtaC+0HxEB
AGd2anN7uPkZQRiPQxoVZh29IuiAllggdpEFSo3gFOsggMSlDQeMat3cvxmh4uUxABkY99uPjLbg
2avZOS64w4yP46cXlz9Fb/IdNLO1vgD0T46yYOTlXCvDgjsuY5J+3f5MKrwyShGIByD4a5J+4fzz
t6vK8VjxmksB+h2w4QkmlvTjYMdLF1378SZDU3WrMR4qrbmtLM3XBGXDJzQJIS56yBRB+Y+3sD+6
j3nEHOXqG/fsR1ZTGNpU5hNlbxOatebUvXyQS8xf6Bn6zuPzFvJJVNtsJbxB3f457vR7WRNhjPwO
RutOWj3N91s8nhdnElPEa14IgInZY2wZx3jnGY6sRKt2qCGXcqO+lLXN5dK9h7B0Y4GXpl+bsZ7Q
FDNYOgqEqg6DFU3N0e6FY7iA/21zlUJzoyJNndpeTk2+XnxW4OjH5G04BZPLCQmZPs6Vw56cbEIH
Ezq6vQytwlz+lsRwaG2jOruZZaHcBNEpoWKBPuElDUAmSVszGc0zGaIGDEYEGNqgm3M//S2/wPB9
Rj4yPfOUjovEx6P9cZjP0OV5d4uM3QsyF0xOzPhj2SzwOZtsejnWKTUxuZLWQjuxWKuNtnHTehaT
AvGF9RMmJzqECPPa1H60XzTEkIlAGZnBrfm3jplXbbEb34ijozbo3GpJJGTu8SPTwV0iHuc8MvvG
ResLdB+XZrgQCPeCUpllDJ5a6ynCzqJK1rYWMukHdvBOFAbbNXzCzSUtwMZK+3b1/OvSyA9CguMQ
4LClYSgTKIE810UPJcaBAhwcJ1BLwJ2kz268m7yOO3NdnSGye8qxxTb+OprnrIhaZ7YpxwYp9204
9MYbjR/3wELPTg8/vOLYj8o+NCdHH40Erbx6NvmkpsveuDxMIXy/VsGTMWPAkY6qGrea0bXH3IZZ
MAGX5A0e5YPaCy/4geoIQMtaCkwGZ8+tAPaGXR958udmlCBctK6yJiIBws2GY+kPgzmm1lgw8uLx
Jvyn874cSSD/L0FVHW76wwrMGycW8g7jWnmO2nrnfbmRw1bNUD2mZbD9pJqwm+eQjxPZ7ZfzhEb+
9lfSIhQ+hTxSg2XjXmZ3CWADa4iBQlOWjbfKQ1Dy9C5rvPwIIh0Xp8pltEampCeEYtFjTvlfDhXX
oK4wSKjkCNv5RtT4HL9jQ6SbzRIuPiCvFAB28PqzQ3726ePq7jED0C+FgufGqzOJ5YF/4Z0dB11Q
WIZBwKyv3LvNHQUjHROYN0YPspJxPTumi/Zh5LS8UZi4Ot4u+KkEsUoTwNeLfHGFd/w5ab4GBL+E
W4hnFyaCPua+2FkGRu97taTePlfhxC0H6h++fr9n/CWkctJgXmIT+wV/mKj68/H2TdWz87kDoSKZ
H/8XlKQkc9HlA35p6/0HG3XL6W5r/N8W5R4wEyJsWebZtbvBxjYAIE+TErOvtDDl9rmoLSRn6ecy
Q9bEaPzJi5XPWTs0EqN7VbTIFa+q1jWI5RHJt9pij8VN7SW/NK7E9ZtKbMrD4+GmfJ7T4loSOkNQ
JdegUfC2kaRQMLt3y99pSm/cHYtOMuQOtPErzWFfnWKRv9zGOH6n1bpDuSev1Nz6xCZCo6xTA+QX
YoPheOQYtE9H5d7YkZe2sERDHMZ8mG2GAgcYu2oI1vgD1CnkJgaAFv73FrQamwwX1n66svtBf0Ka
P/QZStYjxFbYdOsYdjlCAiJyyMG+Yu/yxpWnkOg98on6UcUx4ISlJGwTz4nYuwuodrdO8D8Lcmup
fdXR47sbNhXDsCN1hnZbAJ/k65pbAAS5oHm0gBeHrUD35jQqX+rhyrKvOURi4tY4427fD05jNLel
JcSTacWLIQhcAjraeYZgKkVrvqqFBwboyaKUqinDgg5jfk1Xk1wiFcvh6YX0sg+dlZlbisGgGKU7
ouiwNdnjrT7p+P1zfQ7zeMlfRooF2UAXCkUJFpgKNp1FWBj4z7/5alOgsFjfeknLozevKpS/IKGk
iWiy+rGEK79dXwUQRWJ3Sl6FzIq5VBUgCc2DBHIAa6jQ4hCslb0aCkTkfNf/vxnJtku31PXOS3rz
P1W2yjytgBtkYh5u11rrTVlp5s6c6F+wgmr9Ldw3IvPyBb7yYtC2hXEAFxiqFDRkODLOwIQPbnGX
Fey2WxQkuiRYz6lTQWUEYF28IC0eN2vSoDUWu78K0d/ke/4PSbQtKkXc75BFLTT66039kFz24daI
NGiuC9Z6/2ge+4VtQYYx7dReRGz8dXcIaSPgg6CDSEdmyVrAUtwmr4Cqo55q0T3a7jD4xsOds+Tt
kVGInOOHIOXBjlc7Biuw0vorGKYgHG4JvKUn+CX2SfbgAePwIk/Za/mz0P3JLI8y+aTjlQ2cEOY6
oBjCk7g5TRh8tiVPWaJDbqLzV29mybRqz4uMZJG1LfeQmiZ/uVgLqjqM9oQG9qHbM11FPTakB2bV
vXwx7ESlAR4ODPUTUa87UvRYwMP88C/04gI1HznV0PLes2TU+F4RMg9DN3PzksmK2Wo7Uxph/Bxq
Rlxq5XD/qxwjs7KG34B8SQCeLzxgNtiLRzPhcBg+hrCSaw30Sq4v4HXtQuQGy/FZw0951xcjzj5N
w+fEBIj2va9fZi4G7Zyi3m4Zbr6dBgeEEiuYVI4ixYVwlxWV0c7uk4wcKMTEWv3kMDYOnYSY5qqE
L4+CXEwGNLG6eyPXyYVvRzLY/FXGsOL/H4wcUmuYioyCevdH9A95Jq/I6gfFNOOQnvzacyV/WyUb
DdnLo07g4nQeWVllr3qDoYy7i6NpV1zW7hRb8xOQjtdKdsqgUWJeBwCkbY+QdYMw7JNQGYdwrkDD
gpfsb0JU1kQbbveqzkQR2Ro10ing4si4prwjFCH7Q7+JGJAUUiqbRk+gSC9iVjBTyB+z1rjYuPPi
srOSgf6T9Q7nJYn2s+QdSobm54bHVwlKxlgcHmJFss16ZDpPMTUg8iWXS6peXCv9gyiCN8SrSHoz
3FBFAX8NMpCUKC+WiAxn6Vc6e6vVayOZ/5m7kyrwdUNbnSgRBpOMBC5DMJuBUAW1B3cvQriI874E
HXPQOkYM2vW6vT/DGd13rFkXXZMGaD8bNVBnPHXUybNDX1VwFXJbIGu1wRjKMuCp8/Zqg5CX/HmR
q/LMWYjkYXPuyFkXK9feSuS55vvy0Wah/Bb9tGn/+RA7HoEzkfE8vBvicTgKc9NtkXsK9RmJbIv+
DerO/1LAOiwu9uJffBuIVlsPCbT46GE2VxjC8Zd5GmkqJO3V5P/j2L3RvUJWGHzQlB6Qyhzjacyx
oeF+K9VqFWq2nFr0fCj01o3vkpoI870h5Xzz5olIX6lfQYVb7zf+F1jGmSxPS4CnpXGB5bBUNNcx
omsy3mWO3uWTp1pGAbgE7P1+HLj3GoxuhcjJPVW31wH3e0ToqHKh/Nq2clDCqqwNvpFo4ZJEk6Fg
vZQbbaU+Cl7XryvIHVoNknu/0ZG9f2otT/UWIgX3ggj4QgOUwl9L1vquskAyY5uo3OZ38pWFFMzL
yM84K1AIslUsoL4LZh5i5Im38QfPyeDOKV9vnsIGJ7h++7XYkOKq7YF513u424/NasGxCJvKruWC
hO4gTJb2cu/n3LicJVmUNRk1uSJKdhFYQLu7ABWcFWU62FsRdMYnu+myWS9ZeUU9NGfZkD4l5uCA
1c4WDkdpFJoqrU+3+MbYgYD7Dz2G+7DyVIhXS9fv2h91OptIo9lM5ZV23C6IIDTgIyIGNEikSHsf
YeNlfSS/Fv6jG3IP0rD/ifWAZg6NRpMVSqdsHPAYqSc3iNaV9VAXXiOdDkYXyOL9XhcbhQT5fs+K
Io24Pp4CHHtIQtG0xvTmGuE1PSztiXQn7jv2Xejn/OCA1PuXli34beoe1KUMve9idIzfXEBaAX+8
uLLRwzTZD9W0FS2JJm3Io8M7SltQ5ByIYs99hSa/KbYMn1/GBJ++YVtI5K+mI+0zJvZKudTCQXuB
0dW9cswDdauk4wCtoh6a0DUdIcINEuq47JNZl9f8KU23eE8JBtrcIxhFgrJ01qUrKlY9fVhsWUPJ
NmhApZaXA1+TFR4KmGdcZbEQ+2V0d631pCpkO0ZDvSzh1O68XppWw5hkY0erKnAzsezmyLgy7yZO
fsIe3tJ6Anz/EFxiFPbd6h8gPH5gneQoe6dKinnjKcsnycrK80Cd3i/Mg3wvKyVYI5+JkVSSEBXF
ep/xrnIMLcVw3KFdmvjDR/MxNMWdL1Z2kUqQwqrU0BaXTKjNozvWrOc6qDV8AMdhC6hQacS3eMzW
ZApWeJe2C8hEVKmiNZ9wzaAxWzurcAiKhls5NymknCQXaJwNdxs3/fvai19aYNaBllJ7kd0TrlUB
2UcvsfSbqzvY0kx44nGB62aHjgNbX6ZBdxOWdBgjYvvMZm78VEVw4UQ+0X+G7NpSz+5o1lNdjTIv
4jtr958vlsg+BaqCy/NQn9ZFHA4D7Xot/e0VU615SlNWjxAlPjoa/K/BwihT4MNPKFcN8cZdll03
gWyGYgR1ulxgtDkg52wBjmqJxWRcnSjwAE3ZUqrQzXkM10TU8UC/xcgcFiJsRJIY5Cg1zzxkGjki
kIv6+d35YrBdIz2n90MLZwMEs349Rt/4RDmHwbJ+xMjHey88DDCbb70qi59xr0mQDxTdIyWAtbiR
uUqIpCRBgjxahW8gRV05mp8JrOArcM6OrQTTB7Q+AWTSsfmvLBxXEh+N83kszCXUzI/V+ToYcwu2
g7AcK7P9P9F28t2ObC2fzK6WGVafjUFx2dSHlKP/AW84eQxpbtm8ONDUKeNEygZNvzmUShMUh00s
/WOx/plQ/Aw+6o+nihQ4/AndMdrym4cKqGqvHk9rZgYjZy7L7jyyYOBThspNK8dNG2ieN5Y5l9d4
7nYSBrsij/yck+670wh6YVafr5f1azYjbU7hLxyP4r8RR2R10jEtpFtVlEmOI2HEb0TwMBnlRVHE
GEz8F2Nnm/yjyBvRw+JQKEcAYRP8YbHK3XcEQF6bvwzkOSR2v7Emb8k+anWjQ1TNveSg8xjyjcKS
UJN0S9nJv2FKaujjDAiO9OEChoF7vipVVgbxVfSua9MtgPfHpdfF49Ksa4aYFAwk+TVYEY68GGMO
47zLt/tCG7W7XM1RnP5WznXhQ5AacDdIMlXjAM0h3FKORFDcJR2cW/+5HRPSkf3SrIpYBHH0+/HF
X8tA6bnh2yxRQLMAp2PCr86RxaVbwsooDkSJNZ9dcgPsuff5FQtq+rgjjn7Dc4xU2L75V8a4NFIW
zfEQj/tpaD+JbRwqcRQf2tGhtjYtMQz2wCUy3Fk+3qBDSTFdm7i0b9SSLer9OFwNp/TPRCZZH3cK
zuWW31IC9yhVs6ZmlK5F6JRzbxK/bVPvhzF/hRdb/9iQ0V7xShdkRp/3JALpuElXim58jHUwSlBe
Pi0NT7r7iNykU/Tmii6g8MIz+hhAekHdVgxywXHSzjBHhUQ8UJ2zJb3Jpxex55yayFqXZyIsj16S
Bnyg36HpFnpoj34p6W4rxei51+pJknAcfAQtPxmFIBmbpMeuoJWyxgn/3B6GnjM2hd1Fh5le1LwC
gUIgwa7o+YhxWI8JQQwMY0WeZ8ZDXJbTUEy5vI/uSM9NuPbuwLi4Ebs5I4LT2Tnz6vYsdr8gTQTF
PXhV/gWPje/QhtOR4TIL8RCoRsaYvh9la31Dum8YEBvkD/d5GxE8WPKC/pT5Pwul+OZeBDl2vVam
D8ZSWVZxSeZbUsyQ6/evFZcU1dt7FuB7AIVSnlECdjbBsvzWsIqqMwrHvC2PcY4Vrtrp4oj7ytf8
WGvFM+pjYa6RMy05otDmOkMYLA/+X/Xc8+K30HbSnAGKi9HYqzmTZ5HiuxRIkjuSzLWOisj5lsPd
9JhcNoipz3jfB8N74gGy7873c/txo7HoafPHjLnvJvGxVoE4Q3C2BhZFMxwa0m/HmT980KvB3Yf4
kMKrCZOcxliuMJdw9YuX1k8Dii5DXCmw0NXfkHtAgYQtvAC748rVUuHW5BOhClAop3H48qO9Y/SJ
qi7K+lXszkTMg1B9EfAiXeVPJf7tuZM4zf7BhOW20Zgp0tsNJwZ9DBTHXC2gZfnpsCtPQ3szBTNB
0hS+ef7RAyRmaOckHKXQ2Pq1Go63XkNOihHUG8ZVgIG6842yF48FDtTLbS6CuUzH1VYf2vqTIUO4
TAiXxlBGcxeOUUviJzvGHY+fKzzge6La0RSIMiC0EgAH14JhP7Tfm1aIIu1j+VjOV/9GZMmV1aqr
X6AWf4czgh1siPQDLlEfRyas1W5C3hW0AdU0v0j6h+CHZ2DCnyAiheBa+1zdj0eEn95Oq26ZrFJ7
yaGuVYktjRDVCwFialWmZaDnO3VCpbOoSfxXier84vU3ArVBkx/0NPZWETizy41pBOCoAO2nwlay
UkedbpphW67bJtVIFYNzhwM/4czlKaF93hJmz0ubUIezT5VerMpLLX674/vDxn5a4YmEaKon49me
LP0eDHT2l/3gw4ywPU1xIjI6/xFveYCoSdZ38KH/8bxxcs5YgqKPBLYlzplHY4PunNpf88o/y5MX
b/rzuYZUQ5K5b/4Vq9aHgP8orPPm+wOTxyLPaB9P0E/yOLXYi6+ZAHYJWh1P4Y/oMn+SM8l2EUnb
7eiFlZvsydICrJLjmfm/ri4MNAGRr2u0rK7O6rxCNSAZ/qwXTLjEehpT1x02vUU6jZD8r0U/BYp9
rTGsHwIo0gzk89Lrs3H+oq0EJsHq6Xc8jgcIOPmbIpyoTDRRaEjrZcB0uYLnCgsxNBpc6Tbkg785
LQdZ7XxcnLrpg2HeUm/+5pl1JJpGwnCss2WHwwcw1oMlhGvHWKpt+SBteX6X7yacFEC+NXDo7fB3
c5D1PTazqnMKvyAmSGVHTr+Ms8peBEQVz+VDj+JieHTpyvjTwNnb3ChqmtcCa48CL1eMjcNMpmN7
CKSpSYWRqKebqogOtzbKomEMM4kGgOE6Bz8QFcR9EZQw4yVs6vn/5ZYP3laDxbjHWOEDiC7KxMLN
C6V4OeQkBIZTVAfSUYZUB2hczfuQl725HYXsFEz3cmaflWpp9ThRrBNGhG89O2El0p9VyQNzCPO0
9CHRx7OzMlTUwYUWL19Ioremkc60Qpx8AipIRZaCoNRGjGk/+FGO50Ofaz3wRGfuGxwVmV3O72iT
5Smjo/tmC918IVWAJ3v3rnlw6seaX0zr4h1NKxi6X3VAu7ill2qh++wVMz7nwsr1Qs42UUFuu1c6
9lTEUeyYcdeYMX9fFltzNh1KbakcEeJfjiL+/IVw5BoiTvs2gVFkR87VbDDqgeKM5KwbpZjOJVhn
HZGyPpdYmJiZvwHr1grsgam0zXeLPRO/CeepHMShroMjtF8TG1AXIHRMQLeW+GUkeoxWd0HddeU/
EZiixh/thswffdcL/M8PJl+LpgTbzjnE40O8FFCjyWBg6TOQm1jUVWhVWTDF4DbDeLIE3HCm8DJ4
QsNvSARN7yL0z/IY7d2Mze0SaoSZOTE1gxugE2l6Jz5/FmpJkQ6L1Pg9GaW5VDWBuoYPa9JyjR34
INT6ZFHpGz0EPh3thtgqqmMg9A08iqzZNk3PW1E3uTMdUADEJtuu6F9o67c57hx4yjEUFfvPq4JO
gE1vvmPukkRj8mMFFAOvqJgKoSDz8sobP5+r/heqmIyuWTI/ge2d/uJhBR6hfQsY5zEg6RSnmK+a
1eCICqaroWgFZmDtvyjC6A9JKOM0hEQtikwWSjYjaVxB9sO7j2k0btbqlcsOa7+njgtnGYwKGVAO
20nWKqOLyN00LzzZFX4Gg7jPbJw/N3YCTfMCxEh5ou9tK5LlYziudCV/jYdFClz8hvblq/nEtL50
jy4fQwOtvnvtFJektWogBNCKmwcQoV0Ye82sfaV8G4ZOVSToeLtYCQKISx5Qlu708QwOSlRHNcn2
LUHw3SYRFNlvWtNkOdgx0QEQ3tCUibUj41rZiSZgonY8c/nQ69nN7eA6hz4qdFWn1zXk6uozxRT9
Uiw7lT+3lQ6KNgaIO/qlTQG/ud1LDoR8HUWcnf6zZG+OHxff96mM26RI3WBg0gEJNVBWWhVoJy5x
G5xSixCMWM2lxUfvCLlk+y+z2J9o1bMLfi8iYQ4PI05CJYQ4yZA0QKBU6TMeQQvyfSw9A3DIGqKp
kRNXF4kg8Z0uWusjDNAhi14BU2Oxd2P2qkz/NMTCT0jeT7iIOJbvWltpzf+p+h8cBRIMUj9kdBCC
mgdGoKkXDBWaC//TxsBz/9VSDVnK/FHVM2yD/SDM4dBBat1zP8aLXhxzy7YsEPGF3ibChVWSQnj4
oGkEaOHVFewHtVzl+5PtrfYoyHS3cUz16r8B3vLRQozXgW7h92Pi+/2Iw52uQ4HIImQayEHFfj8i
6aRedUF0lWd+yc+tesLJ7FsiKCxPY2W22KIus1p/Cankhwc26mVEpA1IIhHU/FDzwaLlFWFEev0u
JSnUhtkcgu52MzFCXlkffP8IMX3nPUg4o0tY3f8apHLl8qvp9QfpIEnTOwcVyPc5M5KlYZd3uRUJ
xInXK0FxgvH+3CSHH54Agr9LAwHXerMt79e4/6mrp9guo8ZdwvNAQqiSm4XjEOw2eKXVpBMwWBqx
udX26jp67XlvU7Sy0FvxVNMW1IwjFb3wAcuSfA5uUCDrvfVLnHbQdz1018UGf4rtFaFdWG8bkr6Z
ubngCRKHcAo4aJlzXJSlxQ14v2ELwvAJFH6ABN531i2EJFtJv5qdQEfbZqwdTpvJwU4Gm1NHn3aI
dcpFwpNJTTETAvaK6rBPa6K4YdT55Gp8w4tydF9F8Tj1l17qcU2hKMr8ksAEuvzvtILGoq98Iak9
gkmTkel5J96eQQ/eNcD3c5gS3k9sNtbt/OdT4ghgnWo8L0TjbMyMk2UMHifYpN3IFRGjqJSt+qhv
R2wl1vE26FY2R+k9eMMVcPkT1uCzuAZ9o6dtWoDPOD3t3nOilqJD7Jo5zezoPdu+48GOCiwL1WS2
irOFlBO3jBaT3H5MAsF1QSdLMGJyC9cqWbmiGJlljmgbGkCSaNzv2hsS+HUn5mf1dEXq3SXS0txQ
0uBMg0yf/skXT0ahsPaBfSeigVrxCI2s/eublae6tIeNfCKHUAwiMAb/HfmFphcRt04PAm1BfcO+
0m1z1lTAZommb6ixozdXrKVMACuMy6SQ6B5RhEn95Uc7U88/lyCtC2+6Uqzaj1gKE5/ab649g7Ab
eKGxhoYQ1CDqxMaohO7cG1U2cQ2pVdEiv+IwUdgFvINKsYZp25qYXgs4QQGaS4chYX8AyIbdO8+x
rj3o875yRhk6Dek/IlPA/7mk1zQ71N18hQzPonyQMXGTMtrPCh+OwukggBDu9hwYuksAucvgJ4rA
1NOAPnCN1rUXs/Nk0eU05cGifSsHLhSqO0ubEgUvAqEdQ7+eU8Eaj2zIpsUtISbMRaKy34suVql4
0lmPiHs6Ma4lActgJO6xIDMJ+detuihcAUpgtfcI7uUcsu2afm+wpkYfeRPnGIzxS+h2w9snfzko
CpDxi59wvxOkTCsBhGrqbt/k3xmtJlOgGZPtc7Nf65/dRsubG1nFwVF5/0daHp7x+nmSs8I7pQmH
HekmoPFyKZrOnuvYuEMMyVKpY4AcxASvqwd7O4jwKS8rMUn1gOwkmdZejlWTSPqAre0dbNDupF1+
2U/y8XJwdnkFq3FQSR3uSj2/aOMqjYgFvDwe+oeBADwMEFFbHcomqhS6PU4dULbgcE0hPICadknA
aMszyqFX5GCjLN5bAp+1m76JU1G22i/5v2OeQMXcTk+6f0DqKIY1lVxWYF5vPTK/HFMzGJpxNY/A
OHi1lxbZJpcFMfpvZt0PbMONAW2F4pXMhRTRQ9ZyGD+3+rSqNh4RPwQ1+M5ptq9fadZlY2isUHuf
t6FSTkXPufZ3DxdWghlwmIKHGFzGLIwhvW9MuMXO2KoptYmN5b2ERbAcwrwW5tjDtlz5ZMhwoJsk
XzLA0FYCIB/Xp+oXYgMCHz+WzllGOUhOvN4Udo1tY7BkzsKPBHhs8gbiVTWhb/l1VEyN6TRcw0eh
RmTw6jBzWX/Moh78zOLlAtc8Hyxqy7tMgOknJPeQhPzBrapM/p5CwL9I5cIhDJh2VFuxpWY5aC/K
OIUgv+hqG1XYgurmPWzEcm5JV1HoUP0m1csvzfa6UMHgcH/o41eE2AuChH5c0AmfSEur9nerjcUs
UC9CYjEa8WTmhBlG5acnfVcwVp2r4stIBqeC+iZ4ghOPPNEdLHf3pn6EeBtaW7FXFCqsn3V3DpJl
TrUbn0BMjfx5v1yC3+OUFWZl+DVCunAnttGjbGK4mW8kDQi4sb4Bz1vkpSRADgTESuW+F/N56y2C
Eq2WTqgMpm3WN0ALAJVM6OgnA1GwFGifgttzw4WdNE/rLZqfn+LTaxb1fHWcAeek2I6sZ4sazeEG
XdRzfIQDOnB4gZmMwRU1xtxeqfcWeNESY8P/9UxydSYAU5Qv9PyBZrmKqBbWVd/DoBi3kJ/3Un+f
Dy2ixqJpNXJkoVFhKTALzBYzkhniL8PvrIQaO8orHGB0dWPV8m31wkK3nJ6Q6RK4O57/BqYAdTUu
QKXAypU0ekpLKEbcmQ4WsIOl1PrX5jILkr9If755RYqbf6IvsyIbc3pmazJVA9p/aVd2lBRmmNHm
Ph2JLNkJrAGJOrx3Kq8IGCJX0ApvGBEUAhE8mrnCAVow6pDZEeTuSBNBYKN48wmMIGFylfk7v55Y
Ua0x8h7vr3PblYDE2KNuoD3acx8R5IqvHM4eEEkKbMpzhF7gf2vuPCBrtN1z1DiGj+69N7CwvCJ1
4DmYkL1P0Ag5OLkB0omMCCDg61kBmX/liLtqmjpShzeK+a2RLN6BpxS4pmRTdAfi31tNGUtRsnvj
1qtNBh9aYaQkxI08/LdG32n3vVyeFRe6MbOG6JuaG5cpmdR8QU88V2cJK+pMVfprO+8TKL0A588C
R6Zsc2icx97+EgXFbCKEym7/Bn3vcuWgAccIrFpXdm6qBiNuJkigri80B4LMozbW84MaP2x2N5UL
JJVVrwMCeU9abSvN7N9MjWKPHXlblSfXNZDHT04/li8UTpWDkJwWYzvOkBzQPEZdfYI9f4pS5UyX
4+GHqY0ZURhN3pugBk8TdrThZCFg08KmNq2P4/YI9hRYqwD1huiM2Ts90vULLIJZCtKkITiwNTp/
GCizPxMrF7cmZsxhSFzZct7urcEeA2p9oo9iGAjGQ3TGDbB6UVyb8+biQhOMGN/LWtVd6dptJOn/
87TeOj+6B2bKRtwcf2ydQxvb3id2wfhjlhFKi3dUSkmbI9Jkoeb0XOOkWa5hSyEY/qIIFd9x5jVt
Yw7ZOq6Swm4dyLeRvTNpi71fyBBfeoCldstYT5R8XJSdTJ5J3OJ029+buXe3mHTNfo/+CxEyt9Sc
OIt2CNGpM4w+GTvvyoFr6F+zO5/FwNF2zxmQ+fL3GujRsbEq
`protect end_protected
