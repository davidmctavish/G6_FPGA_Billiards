`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KmBQFcd2QD+kNdok9pVSy+mGWrLkX1cfjcswOe7HQkAaL//+2eh9MyWA7iCeyf3d6lt9rsd77auE
ZHTB/Fk1dg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QEzlBt9msTE+rOcclHYmjKiZokGI/DjRL2yt3XgvDqGlPv64JOq2dg7pr5CbDR9qLFFLRNKC/Ave
HXTRb+K+eTpEPc7Ya4cYQ9g5+MXiwB7XQLPa/aEyjO3get5293ggZuzwkjZSHk+e9QqEk6Bt2c44
54ZWwitNxoUsEtZyS3w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TL0QuMHUSOmzGzMiljwv7rv+fdjjk1oxddi/yntmPUYv8VtZjSw6bnlL4bf8+q0960/PHsqwyv81
+G8ArGsFjA3CQMteKmkfl/GKlw/jFc2hhJ+hJn1EdTZ431Cju17vFLrxGbmfF2JpG6uCGt3WAMGu
G1fJ/VcvUYAU7TOa1hY2/jyUGZ+kSwhGTZ/4ly4fqsmslNZ3EEbYgLpFAp/bY89KPhWWSJnAqVdS
qCq9OYjG5kABfXiZN18ABG0VS1eWRKOZaodlce+Y/gZM8YZj2dctmqg94KhruUweeysu3c48Ck1S
AaLBgWKSuYgiZzrylr7qBC5Dl8oBgOPR5lyerw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dhihncQPuJXJisBMfg6qt1V0/kVXNX+63Zw3PO0eub9NsIOp9vBY+EvdwHq1kfbkAnPnkJp5g5dj
8jo4ZZkQ4/P6qlTLOl2VSHJYjdrirUyAOSEdGt3l160J7/RiV1QcAcFzPoLRIkYo/SrPrmAgOSjD
13RD+L4ONrHTFwpLC+M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p/aSq/rPYB4VskPGN3ZAnJ8z/CGp43GAjjH8Zzz77N5ByF29mwa2r5fYMj/F9VkgSkV8YsC9Tznw
lI4j6LMf9xzEX0HjWvWZ8pW4ITmEXtFV6uNX6FWbH1T9+SQOXk6jlchSOVmnkJTb28ykZodOoHXV
sHyYMhT/OBUCY+iWfh8BYWXEVyyUd5vsADHb3MkIuYdUTbUUFBhXMe9Efyrrd4jCrnlgHytJlFzc
HHZNJzS0lT/zBck+tKmXy9DwdLnPca6apjf9JkkmF7kUXw59bl0WfpuUVSCTVtnv4cgTqLL7Vr6F
wq7CBpoBFMhcwFp/IV8WLrlN0XiNXXNJSRga/A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
im0yA4YWXCc5wQFyCzlvx1+SU57E46sDOGpA9hkiZP53SMBT3GJ17XIBBbg+KlbM4PRkpLopDWwr
CbI7nH2O/1D9cGK/h61aKtTupijDDz6nkMhC7bcK+rpcdDKo8zbgwo8gNr9fjLfik1q7tIcX5Fv8
oAVjsvLmdfFzp2zw03b7SiUrvLfsGUFzid0cHMvLoaXIUrPsUUiz/Vrz8f1cYsnK9pFI9AhuzolQ
q+RF3ma/QzMRtNMVwI/8Z/E7WqsvlAD95qLZFTfjq+iZ02j+n+0rv6NBiNWXDLRWf5gASRNhs2TT
elqXQEbPBz7sXLgpqF5gtHp+zJNCf5P5oR4RUNqoujgn1afmDqYubys7fT188ShbgRVd+XS/1PxV
7+nRb6/0vtQI1i3Y/F1YeFMtnlrgqhC/+0bideWN+fd0XqMZgnGPJJwNhVi2ocMx19mULjjfBkO7
SEeTVOdc5I5HXWQn+EtdsbgKWp25Fc463+RfJWrky8gJW56BtvdtGXy3RHq6O+IAm3sCEh/GlGpr
Hi6GsS7C1b9d6ZCK7L0Ioh1psUc1jTGw843KjUUsVuxQIvajwX58mpo5NqV4Cxo8UDqtBEZjY07G
bVzpl4eusw8E4XT4Uw+B/Mb27jwNy6WVPTs32XKSU0EY4GHGeM0Q1GZGELFOJ+Ixj7J0bZYGHwr6
Rkon4ZnggnPhJ0+hAAboiUs6ydZVG3hEdbqg0q7MbWc5LTxWQpzZw1WTKaacEQXjmAqYniPOUKq2
QNeVhahR6cZxgTIwZQD0nT2Vu2p3A5wFgr99sbTvlS62gRpHXTS8T3WGmA/i8JXpqbSYvc+LLIu0
NkkV+hC/0/mcxW9xXrExc0j4V/g+xx8R7W1PbJZ3IVc9PSkKS+2dYgbXHKKY+MP6kZD65lGtDZ7w
1Dx1/5AzQEvqWZDC9xrmW5RBodczk+meMhmyliot48Fr5//QziWYgKMAK6KWUGKRToxjH8D9BglR
xHNf/AV58CT8T5OOxMEUiT1ofOk90ZMulgvf/0QOoDhpsZ8N0QlMa02VeVmD2ihWL89qWQrDcCFF
f3+mOkaKU7PclPW3rbSQ7yOCXNX6rSKsssg1akXzzQ6m44336msw2qFxuFgNrEIsQlJuBFdm46AX
szJcyp0Xcd1dWnrkmlkfSF/+qddqfkh5pCSvlTsgFzwmnD4Esb8ko2gSSZwYu0B8/LK01KEc/yQf
S4OFD2RzngUbjFUBgRCuvUr6PeQkPKjBB+dnx0dNA/MDVKI60jpOEoQ3Ue74C8RXOkyHbl6KAG81
cx4OnaFjzL0sBPo71J7LbB2xfayVgHl6Os6kbEZJPDsU+URla1LRkXOo91df+Vars89rAMmWNMJh
3miDDAeqaiMbLh5gauqqOrrfKRk07ySgxUB3e8JxDvRgAbhp3SmdVokS4muEXo9WuRY0+qBtZ8lx
lYc4ex7rGLjuJJOTyEpzXgtyijZI/w16hsd1SnhNwePCFIWK3Bz32Syo8wcJrXgypDMuj2KS9CRn
0edFqiyaH0fSRDZgj+JZ8XbucxJ5t6yxHMU2cDC6M3T5p6LC5MHwCzqPZ2DdnsJIO0SKf4pTY6dx
IfP9h48jKf+wKbLf30Q/jb7H3msbKEuyHMW2kJyGUQhbHoQ8JGo2Tq44L76R1Vtcff31QmYiuVWV
HG1e4lHTi1+IhjzEyjEWx6Kn892/SLDZ/sg07UoHm6wzeD/RG5pPVRnw2z7npY6BvMVXA6TQP8NE
eYBmNWrgKVK8weKEWS4HXvPXIwZmAESGeSYVAkEXb4516Qm2dg77nvD+BiPCEWkttU4NZhV+TWc4
TrtFh/6O3sPbhigBX8dK0XdCUJZHz/t2eTeYIJvHn4EFO3sNnkzsxOr+RwL/Yv8QleN63C7OTwaw
BIpOEnnLVLHUyo4HUIcyDCOfTqG5u2I1seTz+B3Bx3xucZ5h9LsyHKUEWSiaW2gC61zZ3gDcWG6H
tPPCh8L/LOjQS3XVpfibW1Dz5sQP24WMEqXx0rY3M1uNiFRHOWDkQIt5RtTpj6sbvb/d7JodS20/
SI4UwSVKBbaxl7I59AtSAUGo+J2xODzFPxKgMHDeSvRf6iPoG5Bo/ODZVRbq+L7GmAlEp076kf1/
ZD6WqYT4rXIWLurHH3wrR9/9gW/yMVgF76wqyEUa6BuRrZjcXVEOzA+A4VuiLg/zF9L9F1hrzj2I
0oFGO66Kdsj5B9rYRhQjYALK/vHUMOxJeKaRLB0QlCPwSpwsOL5OzV2UHxl4eK8oBr6pMgcXPC0P
Y6nynu0rF2Eii4YZ7+ULPbyflIrGlUaRaEO4bniBcA+xZAllt0K3fAvTYNbR5EscHBSw1fstVEQ4
I45eRgYCa66dtLDGlfj2WhSvCYSTEAM/ZbEh41OtdgRwgYr8MIa6my4Q0ZDWNHgBITB8AYrgUS9U
C95S4s3sSnU+orZOFICTvWRFOD+ZTfXUzCq6zCkQHGvfqLC1jFM3ybrHNJWC98mZvkiV54hPyED6
RnIt6VcJbpzi3r5ePQHWs8G5zEzkvj7bjYzNr2xMNk4co1hUbBEAqnfF8IY+nqOHysL3IBMTRWPk
fq95LbzTLM+YmszAoTlEqLQ7CmfB8h3nTkds7GYRaUDIvGK8+pMxdIOG0Nca4e77Z7wd2kHYhcC5
AE0ozkO2zoXHkvzxizngay/WI/zUGrrzqZqHqL0VI/+BSA4muTiofOCzFywEci52o93dGVuegd/R
KgX/Gtnr2aoLYjObcp/g2nuqfnTijLEcTskgjezgWx557uq3mOxOTsdLmWxzqyWKvyXuwHzfaCLn
3qU6OtNvCrA+Krsxx+x7xblEhxO5IjE/X5nW1aYt9yseGh7L9WOW9MvzKTaVyY4XjI1IRGcxQzQm
fQTf6XSQ+RMhSyaORR82kgIDQZ8FimbIcFV76tNphXvqqMaV8lp3I5SVcMb+LhQFK1I/ynQ007vv
XlX+HOyXuPw5xnRAEGx3ERuCt3dvYMTH6wt9k7YoNu9fVh22xfngDtKWY+rchx6Hf49CGt3HtN2U
1gAms4zj/lvjOJ8h7SFQhaT54jcNvDjWjahUktQRduFByQOcwaiN+kgvZQ69ez0hEXSjV4ljbi0Y
ACIbaI3PfqWwVWgUp7ZfV/de3VLsgzAGkAtPFu4bZePJDixd4CUOyvBzGyTWqnlARLXi9xY9N7Df
PKHCwBsML5ca2AeZOkvlcAkXJhFJqxBTyu3KJvG0o8L0wKtjAOS5qsqGRrYQ3hakz/bxcGmbmY9A
pOzCOqBKe73jlRGBbpMA5z8ZW4Ci67p3afIh5By2QK3iulxU3xQm8FlzyccceZup3SnfSwHPHoEt
zbERr69/GBNy/xy4sAi7jpRBPjQgPv7TuAUdmoYogiKA8SKVOQTEOfFpkER1MqsYSXF5WehW7Qk1
LAHc5feUGcgKS+Z1tOu4+vJKsxCes+FJBubJIAbIoECaLnfG1q7Mcbzb4d7JTNER8xouVQyEwjwq
69gq4CGOC96//CQMUxABXd+7cYftuyHQF6vbyTwFjfPBEulhJ+6HxuEYDejFCesOW+YSaxeOumZF
FpYi8W/ORz5ulNF+9vdYQXlMRWLaqzLFKa6OIBqrIYzuBd6qRKvDe7ehNOoWZQ9BKEJptXvCbBlX
Pq4y3k0quifbuftm4LWt6kEaMAnr3E/lFURe96xG9O1dWC14XjRFoGdUnAfcokZWFWU3d4BS4XGU
RIWZYTaRuoyX29LSL1mHm3GMFQMgd8xQ9P29LpDUoXxXG/Tae8TcC0/WEKOzwrauhyb/3gdWEBlE
ZwYg/QKF1fFY28Hss7CmMIcVJ0JXMH9TSJnNCE/U50YDtFIkeEV3q/0VomywliSDy93WXPEtUAKG
zfXDEScHIqDJ43PpwdZEymaxd+49xFvl/SaHdM1vwlyTkhy5QIWwLC6aClnUAtouqzb09Ra70tPQ
7ZuHXWvorRCUt720jnxEJHBQ1H1w0Zdd/hGOPAnG/v2ub3AdDQoX7/5W0ip9/TD7oiiW99xwnPoH
SdobCWk5Btmr4J1JkvNPwIMjFw3vvKgeU9fx8EVYHGbLXi09QIg58J2fieFGf3ZC25UlozoqFc7z
WvP4q3UC6dLMlyu0lR6FoaLRrj1k2l5P6u1T1uOUN87o/7+VV6Bzt4YNj9suZMlwBOu9Soq4gaKA
pXrLdaFwwChJ4f9h9XPIhNqM8/SBg1UYZRlWmwN4Y48sjzBmfDoOOkK9BUN2iW34jvagQZm4YYvU
DWXbq14liRPyMtUhRy4fXj1HFPrRpsoQv26M2Zn1CDsPV8XJl2T5vkVQ7GpFA9aGGIYmuu169str
Qps6G4GmPkaKn6wR96goZv+fA9qH15kH60VeI9c2IfC0t2kMfpcosDr4NIdCV3nojpvuHASpfCNQ
MegoTISzmj45QGQWjQFT7u7jL2L8A6m4m21Mhh/p1g3NnsHNCD2jZn+ksxI7OCAsnkafVG8VZwGb
3OeYMxvEz2hPLuaRW37aA38xHKEHc03OjFoFb9O5D5X6lw7lMN7SABru399VcFoP1hFNunwA06d9
ADc2Y7fhHuoWpuExmhTGSAgH5SyhNj0hTNKtBG4cujLsUC4gb3N2hwxVyjafQo/sOprAWXSfxG7x
Ul3CZU6T5nS+Teg6cjyIVy++I4l4OQqvg+ZDmf73JKdgqbl9cuk6Ss+4Ehu2MP+nGL6qXQCQH2Ps
OvB1mlS8U3pmpQeLaTvtf+4khKCxAwycpJqxYIKgHYCfDS0Lhjd/VLV6ygyTmwEf35oVHE8ypCPj
/GRFueV04BhiNNI5BZpI3sUOvF7CvbATkYwjPS54WEcxv2acVuvltBN0NqeQkqVCEkHe+hfSAOtI
Ukw2duN9sQbeyNCMhmOshyGWCpnHto/WKQFqi2vLvg2ct/fKeUGyogP/RoHgEX8g2+o57x4EXaaM
j+gnYDH52oo7zPD397Wj07SIhPHoDni3gI9N1L3MaEqlD2Nhb0hogNnUlPlXv1ni0QdKBQo6/hmg
MZae5Mytu88hHaKALzA5KbwJM6I1ozrRuPpWIgFC4JVupgKyaACpM6/H9uvBVru3YqHa5XH+z2dS
bJ8/29NXVkxRZh4u/9lQRKqy5dTyf4VzLsTgsnOl9RtmXqIyKSPbO5B1W5r8mWpKnlfZvCS/OcYT
hihk65V++iPyXtnrLaTmPazqedG+/zeZM74k5f4Xe1tkVjNXXj1JshMxb9OORC6U8Y4OOFc4Ci7l
sF/DiPE/W7KPIdLA7Tf7+hJrNtMpF2P6BkfcHZ7h34Kw2/y0Yv/DrYZ4QrYxUZME47l10L8Elrzj
0ipnB0GXKaLZgzlxroKU3HEmMtfRhCf2xKh/9TgaQdqK/Saxnfc1mR8pv0x4ibCHYnQAUzZvNzEk
qCltlk8moEopkvEYsBk61M3VUSK5MXvSOc82IjYjZyduPm+EaqaD3IrxkS6FNRZdkVokOVfuUrQd
vXb82UOl1Oa+lyCH3R1TeyPIhiBOdT6YD+suLNkOib2Km0E0DBTe9qvcMYuQve5dR3MEMb2cQVJD
OhNj5DTlxB35rFmgDrGfE2gRxE9KoiyNvosmhM9EbRFuweNNyilF7qgfxM/7UAVqIDS1HfebJLJY
QfF+WujqKS6D/5PT587h+APNaZuMoW7SDu04BrG/5RKX+1m5B04xCfP1JrLJKgTB7wbhlZCFhZGt
ezjJo30qlkdvi+vSjrQfTBpdbTP2TixYRfVtPyJe6A9DV3hBsUx4E6wW28BjmMYwk7MRKMBZ0Bl+
HWOzH8GKwXSFICN1OLkse2yv7Gcw7hM1xFIJlBSuVJLMQdkiMOroWW+xiqLpTkV5SVRHGz5fR1rm
/hfBWO21SLdBOzUXq2PPOLzGJqHgVbkwmrpLnaymozR66CvlAgAP2ELJLhRlN2NLYvgk9A/ZSpch
e7CfwBBwjHWxiiqoDS8ZX/YD+ZbF2W3Lc+4Lrf/HsjdyXVYouWmzZ4qieQL5OACkDYV+n/SMwfmz
p1Ih/reRiHnHh7ncuzkmpbXQQQzVeZnu6uHTMKTvhtMaa1yKZH+rkCUMNkSeRFqfoa7iZYtD0jQ5
PzSpD+O8mg6q5eP4JNjh7VUek7BUtuG8Oq1DLtPaTqtEeDCMtFVyxYHLNi86fprkXexvcKP+zU7Z
cv6Pa8GKxkHwCB5/0iQKYOHwrbs3TRDXYe68OfbLZjJ9MOSk6By2fV2Rg57ZuTJwfMMjLK4e618H
pS35hHZe60QhwNL7ZBlwWCuZo0WiFmXoIogoe7JxifyceVxeGFQvC8GcrYP44vsjPCjX+wBlRopp
K3S7ULBVcpuFVb+xkeqmafHXfrkphuFZudediVyyt4DGkJQ2PWmBgIah9Z09WoYYm6X0C+YTr67T
Z+eLyVW5IjDBPG0JA8/phhkvbBkk3ypUs+TUhtBBzD7a/trs2PUUsA1sRflnxlYcrH1zZfpsDweJ
U/40jvHRUyZXsqZxV4xmjtElMjaSdwqg+b3oyzNMqJGpkN2gm5yWLQbhUtBnEcawel+UANobieba
umKb/2bqBU37/8xe+7Wigac5U7mKBqAbjI0TIyTQoS491wJRWFdbjKT2EfFggqYbJBxkGKwsfxzm
AjCgHzCICPvmKW3JSZZwM6sKpFN7ON869EP/1mR8sS1aQOSbI67lzgGoTqHVd/sfiY5bAMRYJ7cx
ouVzQHBwe4NaS6vVO8RIKOEGK5SNEMGzhf8H6RsYkzqBlQtSyFQIHjko9N4vpANA13WQhc/2OPSD
xti7LccukdVvsAWNiwAKbRp03msvBRoYZeajrZlUEBHq7VxlT2EIFAD7/1YxZ/9eCuM4jP/yrzeU
h7ZgJGcSyuloTLE27RrVDiOLa8ROLW5/ovaxzdo3FmJyD0bV7ZG/w16vh4JxJHkT99La1/VhWeAJ
+25+AhCmPxflZUyX2mjSwPtt/avG0ru5TGbkQoQkXTKluqHzZjZgl/2fhI99isIZ6BrHPsaofyY3
qL4B3w==
`protect end_protected
