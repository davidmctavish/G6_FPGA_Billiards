`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F8rxxO4Ah0RXSVnAt9hRSGyY/zr+qnkyDl+TyYhUgsuQIVZKd7D6tzvDiNOGguh37ZiCMdzlS+iY
OHsAQlQrGQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Yc5xuxaUVExZXDua7pFR2tUz32UhxtpbUWJTIbJfPhB4En0QqCUcvvYv1KooPlrNX6JgsLwdqsX7
bEZhoOjusaup1X0FHY/TyHvEOtnrmxkvUbgz/AADykySrHfeBuy9o4w6mTwNtwt3pA89GcwboOkr
JkpQAt7nw4fkkhAyTfc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ofxo2qvOuM8WtK/fiB2hTWuapndArqRTfRLTYeUG9PQ6U+r1/hKQxDkrTBkrXE4Iq/bw6xF98BNP
ZMAPlt79bEWI6jP7RhW57CIJRm2Vl+B9CZn7BlHiT8PzV6t4uMiEY8sAHO6s52XvRSr9kI0uEl9f
/o2iVpj9dTv8qsWo8oohhX56VYLLgBCsDRL0lNsxfRHX1Dc+fKpBB/IzSWTaS/72QSauDUqv0CVD
bkGmJqFwbgRdYWpu2zqIKcszVI3pPfiuxD74nI6hplTyIsg215fUx5UrVNliwv7k1TYEgGq+L+aP
AM1ots6l23wy6+TedhXNPMZT3shd8Aqdd72tiQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
laGbLjwbjeJ1P3UPtdUe8LiEuGpWKHEVwa544tFk/WzaSeDZUP8esXw2yz3buTctc7mh1fzEY9+o
N97yXaK4J9AcDNwdHHYH2S4sBrwcfNTya/74ZgAv6uCuxGdE+mVkA3GrxAqqhpZNNxKraDRWyANg
Oy//2H3bg1BanfGhiKY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YA3+3LIscFTVnZVQYgOsy0z/8EI1v6llbJTY4+K+4uMKcgjoOQChRSbjSaPlytPIarA91jLeXkjn
AhS4WEvP9h3hba7q2LF0VFWgsq2r9NlTd2j0SVKTI5lBk+xTppM+K8Ho5OoKU3pPf2Bhk/g5T/bj
BNLUsdwgbL9r0PnP0Y3Pb5/oxFyemadbaY3YwhvmakPGWkBJ7ihQiJcRxjuNTNNBZmW/MI4htwSE
zzCcUSlxD2eLc240cQvjdoKa6FAji9AiT5jAr2EWdoJClUAVTFn9Mo+8UdJXjixOy0TOn0mK8dKs
opuVyTiKR9iScBaZqVCCWRvZHlAO49kzJot0eA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15616)
`protect data_block
tVJN0mqsaJQtcSi7HRQ8RaXJRAtd7f0c130GhPXO1Ps4u6E91TXIOQc/9uWMG2LeHtxZ63mbXRE7
Uxwllwh6kqnm4UOlY8SbT+W+Pgc2NfcnfilcTlCTYF0LNqTuZlGEWyGSU045RCBuNewELOdSjWQE
fU/b7XNpQMg7klxj+LsHQNEgsxp9l3ZEpgZAVOFA2G0tWd7R3dGQjCmUoET/XqvGiz60ikYxV0vy
w9rtJtMPr8d7mKQNBiR8Li3fj9WC3OPMd1PJV+me5braGYyv8RCTHL5L7ttWBdgw7n22z5iJ66GB
CZXgNHE8Ei9HSxye5K3Qy/OJjhQyP8l0BoYSmIwgu5P7geUS24yUWYpymePiYnSD/ZJYclvy1ULo
1Lp2xJHbrZLL7kiiQVSDCjpF39UGvYSi5c4Xmyh4IKviwLKDZTID+DJY6WzT19UU4l/7OP7t6n6m
GGf0nUmCUu6/qgfHFWf6NktG91Be+LfpQTlJgKecQW5P0ORkpPa3YXERuxd5RW/nT8yB9lD4spn8
ND+frRHi/wovwE4NBaEuFUuGdLSd+YXCCaVqS8Cg79K4kCofAF5c7w1AnRfDUyJqttcGTp+UUdFe
+5vBCTJlTOkktcW2aFm7/eKYqBeuPBRie5sxh1Mu2VIQa0hJBewXI9tOl7RMmLNXDjaLBcffHy4L
TjorH7sPHJYjg6eyHOI7Mak5HT6ZHaX6/Ssb4Lxo59KrzDjgXF/hqk/UVTzTqYJe8qZVvNRvX4yj
NF1oCixr5RgLRHRs9EMoNc01CdcZHSaIyVAoeppv0kHhNWYHVWduTP6mLBwI+AVZCicctUStD/wn
oIsvzKjnQ0kx6iQ9osWqeXBqcvsn5/85hzfz/d5nDkAdLj//kWfK6WMd3liO6hnIfVp7oJdVpzvb
4nRfLjdp+ynhFxGodtTeJWqTY0xwnu+rn+x8dI7lNX2LiEmslpExBsXutkY6Pb/4ksSmtyO01cZP
sOmTmAj65QR+fh/I7WpZRfhvsYJgpaB03VWMSb85VW9UdcCnAZfjH++EwyqBRcnDUNRts0mvWgrX
s3GvZHeLDjCUXTMyVipnULG10ucppqKE5j150r/Y3x4UZtD8BEHiC8rboOtFiu2ltdxhnujjUrwM
4u383FfHjk7aym4dgyoRDE/A8vM89KPer8ApBMbE2xZzJC4vpcfW1jyMWrf50CZrzhb+oWXNAe2f
ucOOgc1ZdGjFwyjW/pUVoJuUTyCZ9Dj/8VCt04ArjvqSBRVErVdL8WAnOEiJHiVbD1hYcKcz320l
9EDKkgTyojlFrUnk7XKZnFZcMW1bqrJusUP91/2UmEpwHmYC7IaeJ2hZvGWgxEOdtJdCgBK8KOS9
lwq4k0BaU8VsXnP2TEbZuzRh8ZFPQiCMdFcGPg7HVCbQEirShIVM+mcgS+go/aGbuvuARV8F5kss
4gl4Sr5wnD5WNvzXjS6r9Xw76Oo7lxcwMrDrUTEt52vhebhy427LibRh5QKu5ioFJfjA8SmD6xNQ
MdShq38M9aYqdSVE60qLzi6l0xD5xG085IVMehZKu3wYtBWFJ0Ot6OuL0gq5gFsQvIVWRCErF5/a
YHOctw1fwjzPdTPO899kPIo/TvSr580/oZfAW1tz7ELxQup2elqCaSYtjRjpO4aU9qMlKFgnM+k8
FJkUlE/tKnhaiXHxEOzk5OVLp1betQY28Ga8iIGKCMu/HmSxZJksZKFsbMGNC4n8Imp0UU51grrK
TTNi+z9QoU+d4wIwVgOqjgX2tBs3qSu8C3gk9skXYo8woR+wo9REowkIVzRH1jDdgRx/mTW9dRR3
XIWLZM7HuU8ux4odARLOAFlhoOHArCDnrVST+fNfchGW3kPIUGLeiFB4yhwgwX2qPfwIlSdwN0ms
oLBmOfC7AjuaIcA0247Wn2rutFAg7lJMRIVUzCQK2zuqrY2gDJrmYufJFIiii3IV3hLnwGTVUHmU
+IYrlTr6ESO/Uqllygk9DEhuzSaqVyx10bTzhCtubhNcuIu/43icMnq4Su0ZZrgoBVpeUQTtLjmt
V+rHVR0XxFXTaHwu0cJqloqdBnR3xHoiVaPI/gQR1HsSlERokDHTwzPsM/6P1zRPFnhOT1/P/Zu+
O+EhhyqPaTjUgHsZwk3tixdYI4dXlXgXGRzv4rTeHtaxsKZ75SrXqcxVRI+YMSKOAmnUakMW7lce
Vvg6CUD2nH8LR+xvzucB6JzYfS0PmYQxnPU1VCwPi8zt0q3uA1SLGI593tcmuzvKEsM3IxpSiDrL
T5JkvTA6oUh6VoFj5M315EAzI9S3ojpoDr7JxnupJg9n7XeMuNspPbLrpxoXiL6mhZTO/ummzEuQ
sIsJy4ZIeJD7gEj46uBorU7vgBlmgWpIqZF9r/v0yW46MHg0ulFQfAgAIVkbs/IRoiEpMTMUhAez
xVBVmR1vaWk+wFkuqlQ+EDCQuXu3qr2v9KgYzVyzfAfeIMf/PJ2D7K0h2GSnII/PxR9BqmW3k5GT
M/T+Q/i/qGyEzXX90GalluuZ+VgqZ98BirlfFdje5Kt/+JM6l02TyJk4/B6NTjEP2Za1q3taKq5i
d58gRCQ8NgNMRO+DQ5bvWk7a7uhdlxBoM2r2RFtQRVz2df9SIOLUN4VWUwLx3TmI3k99wY6jt0Jt
8nxrsM7rwWLUgQOgkca+gvDHwdsXPg5U8wFLjbLMlqvukAogIU28FQO32q/EGF8WqqkK/naLu69g
/KJ3xMb2YHJjR34EDAjZwqLonGTwEzP02dHEQJAadfKp1RF4dkuPpEUsyLU6MwFNOCSqQA8IXVzu
2QMBTYDJVfc04vaMkXGTR9CIsVCJOW4qHKJ3ROYEUIK5P1ES21taPMfku1yQpxTsw440ddwY24YW
p2Ft4t1CLYl/OCETGdqmu7rGKJUnzOokt90lrI1BIaaS41IBr9uTH7vFaN428ChmUDNfN3SLcweT
5j1UtiDu4LvcGf4Qd0qr38uqgRVMVEEDxHvGKuZhu3hUCB+Vu3pUjz9sGPEEvMctFjapH3x/SbI7
il0HUN/+lN2jFDIwSx3RtmnG6fzrzc5OjqW/nEec2S3qlq2TIljLXcr3YjzoXw6GQn6hoEB9D89G
uZoWEGiKgJCtp+7a/AeQSmVVS+CsAO7+5nl5CHMHEE4wJ1F5GCTPL5W5NakkeOUHDkchYkWGUyOL
8Z6l9d55VTY5mBwbZqg3GkF91xgbeYM++r/SRXTJ666GmhLmJKMUITSlwYfMRqnL4ESyqLhPq2fx
1dlTMUv6DXGEG5upClNgRYYIaCYS8A0GaI5XiJbiKDPhwbJXokfEJrhMiGnOlhyTCVZMPupWQRoP
wJVGVYFo03GmnWVrU0VH1hybYAOli2377+I5BOHfa2viyLRnxgZaEhe3LHGqWN25qmcQHIO7UKPY
/UHfeGFZViKxM6REe8e0kq9acIR6MuaGYCLhyZhiQBYlO8DjiMaFYCvkU7WYtE6wp0Ez1gusE4Fw
/ZZxrh0IXjTAgbRxmtqZfJBa/S0s471HPisObRI5YQoQKz2RojWme0/HqvO9piEWNkq1WPnvpt25
se4WISptGJkwDuoOQDRXWdWXSWo0hwJIq0yF73JO6MXjv92kewj0OZfJejpkd7+g3sfs+sa1R/ot
E26HvzKh5J2066rVInXyZOFNYSaL/ATMiJxRc+4/MsVw95ZW8qWtEfM1R2TmcngN4sS5PE8dXcrF
M12E3SLqbl16Donw9Lzzk2tlMWy98gvvNZrvMkF5Eodc0Xhi/XnS05SB6ZFZ9/36GSwiCYoxabeF
PukgABAIURd4I5fi809VdgoKBQ7sORD4J6MnyOTyqmKhKZD07WRCg/oZ0bUHMoa0S/McLnRtFFcn
y2HFSPJ2/fHeAJIc9q5FrjiBZ+h1Ij+i1HeRLoyzNjgslmvg1b+5n9kbYGOLb4GnGwX1ZYBbxqu4
LnQaQyx5g4IO/f8xmpN3cCfHQgHFV2zuIDgZjdyMNgFoHXbtpWjbw2yFuXcwIq10f3rdkA/02WXC
n4OzhXAvxo9WmILWB9XElaTHy/SPzs/E3A+JYPlZwO9Kc2iiJs/YhDAcybMuuOex5u+uJ4BpciXt
1BMn/fiG7PrJ6CuRXx0rDV9JYl3wXWQ19Unh2b+y3yKwtRKrEH/hXvTMUyyrXxVjCwhdtN/zXgv/
asFrsJrhty4iuOJf6GdH+TBWiSumav6e6NEpmXrFOzQ0PsvahWK4ZnVH8dit/n+3RGnkaVMroB8q
a/tcmWSEj/ROx2EMwBdrb+05zIUrWycs+U2yahNH5MJ6IkYmYHyP1pPG/wZf69vHFx7+0l+DRw+e
IOLNbMN/oyoceRHT3ymrgE4tuw7WwqJwTMzvnLfVpGvFrntDjFX60F8eKOlABn/Kvc8+V2lQOQ7P
8u87z10lcmqZYhkh5/qX6YxedUmAg1sMfPUlZ3aze3dd0JyB8xVaZiUJQYGnlufTmpsHJhFhUTwr
jKJxWZXUiawdeOUp7TbYOZAvMVGHIhYMxJ4Ep96t0bfnyKN0zyXIfoz23hr0pCiFESxI6jAjICSd
1L3UN715zuokGlXONfMbFohSZxQ8QAaUYSamqY9Jz2ledSpcW2kAiKwdyJ0Fo9tuf7WrwcBLXsZN
L8cayUR0r6A0LiIOHvPZE9IXnJE0XT03bgrQf4D2mIpa2r6ytGvX/nu0HHwNO8kEFdABQbiLWHu6
WSm5n1YDgpX2E9xBxd+u/pXUsz7KHhIKFmch04SlfCXBevLePGG7rLsWJtOhDrPRkDjG69W/9dlb
dvQmqbZQq3W7eShDsFFrwQW/2Qp0yauC9k9ALBnONi+s4iQiclriP/OnD/+ceK96+CUqQdhDM52F
OC0XMWgszwon76LFKxp4Vv4x316hrCjPsuE8AEjGVlLW0xDXI3M3T2tb8eT+hDCHwv5W/+HsHRH3
QRLmkUEU3v90chlbbgql8q39Oeldi6Dapa0DBFtxICI0KTMoyZGnXCBQLCqhTnFRGJU/YZyLHb77
1qxQG92/oyULiIDxJ9xfrZTq2Cp0+VR/opC7IjCPQ75IEArEhYioF3yW9rWJ2rApYNShEMCYC5sR
dXIxeT8TsOw7zRB30kpuk4eIjznKA0UmaxtssXDVFyBh0zKPkHW+OUsX10vnceX+rbIObFeIuYep
lUZPqAibj+LASG6VlqFGt0rl1FkvxTjLodTX/+33kcqDB5wJPYJnGhwxnMgiuZ8QYC77icFoQH0s
vRlMFmGT7na8RfYDWXSyBEj2US2P/bRexbOCy/REczb0LMTTJe18F9mKaUOsX46TZe2Yy9NgwwXv
+utcrOEQrpsshqs4kOELAUo510Awru9zOT1moF1E0MYw3MwqDz8AbLEAhFnZjLQg2mEzRmtVMTG+
xFKc1vU5s6JSkvl1jxNKBoRqZM9qM89BdlC/5kmazfqyDu5sJpVRGkzKt6P+Ely1EdtjRVGK/CdY
v4zK0TlVrFr1K7eFzsoP4aBT7cg/XCjv+Br0xA2trX2uBx7jXJOAS6Q99lvNIIhNNxtR/r8oyfGo
6f7NJaYKHT7o3JFCrfSVHBEcwz7tE0ESOna2R+3EtkBS3K0wl7wUu7VxDfsX/4GyXUTHVzv8s4MF
ytHLvvD4rt0P4fyci6bETg6GhI379rJ67MrwaIICv7iB2H9ghXssEKPEWiXjhnQyZXOxbslLrW8E
Y1JwuX/jefOcMrPcL+G75hBK6rI1efQRSpr65oxqyhpryQv3z89QVhxrj4W27R48vg2s0wjN4eTt
34EQElh2M3pLi5+B1Aih4frbFGqQet24DQ281Cp+7jZ9jVIOXPP2XvUO7zS4sq50jDXmHoG8wNI8
04V99br1R9dLhgEOhJN1Zis3Tig0XkSXn3DE/DhD9bKuSSSK2jfyJmRNhYkB8Qt7/F0FQOtVasv1
SRN6Cz3yuQZzC2MIMK6sxaJNbPVWfnz5RKN/Ocu1VCT5mtNhDQB/iyI2F2A//rMsBo9GoqUhXp9I
P4XJSchrmY45B36tV65N09xjGcGnJ44nez6YMhZ36qbmG1HOOCypA4/MxqGAZvcAVdviac83fszs
UqM2WRt7pYtrNebbwGRHIdIofW2bAA04vVW+bjli6i+Fd1LXmWfdOc7WMSXy3fb1K8ykztLkFmfB
uMDCZF+rO1RLlT4Zn2v+2MyD19r+FGFZuDU2ZNLtj5ZB6ydiAc6dsr/T0tD5FQ/erotvFrArpo7r
7CDv+5j6dwOoQh2j9yPQjPPA+yagk5ZCkp1YqnQPrv7DAuOYBCRt7jJbxB5XIubSTpGSUIH0ZLKa
DJUjNTuFrepKvSYd5UMJQxjapwKmihNqJhMmSQ+kAph+/A1KkWGcraIGFR2dhfPkEQ+M2Ibt/b2I
1kkYlHHPcbuKaj3mQFVZiAH85NPZN+ZR9ELz5rQQ3cDN+ZvsnBYIHlACGfofoN4pLq2K6dVeIvKD
i5yeE2iW5TzHF3bQo4EQqP6PCNLNDoFrMykHqHDGFHeDs/lPkgeat07bC9bLCeGB8aEGoGy3SmCO
968dS2xKCVjhrjYGRkwlGOsSAy4bE3iAk+UjEmIbGT7JPn5kVz9d90cxiP5YCOeGwy8ufAxJ/0Gx
GDQNLjZRLyrJBLn37E4b0flHci34x57/ikSchtSpvgDF3goBitkff0t0xGfX2ZaTOAAx/g8cjhld
7yKBbdJUpeT7oX97mtTDmExvDteHCwm1zwarJTB4TuNx8BUDD308OVay5c4UECkfdRnpT/JHZO49
84io1opcaqRJ/0X1JV1AkxTLFiyonOiRLTOMCxaIA6eq4Uaq55htgrPHbApUxhKNeDBdTTUpC2DX
qRbZoEBN5QvaQ/v3721/JjzK0rAlYYHabp6oZ+xLeJQSTBxJcdhyQh3g+HQMcVjIffAiJAEJqLZe
j2l84ARlJ+FhamjMKn2HuMNS+pOEpxqUTXBI3jnDTM7YRpXCWRgZ3b7bkFLMm77CgRpl75NRwB0p
UZ2DZu1BVa1dCiwe7rF40jGwRrelBSkDM9Bd/NVdo875C9U1lV7kKpKlci66povxLk3bTbKURYp4
mVfiKphBU1qFWuu4FkCuLzBzTbw8+7Wrs7HqWShw5WViv3xzyN2EAAr2Zo5ftsjRUo+WspERzGUz
8o8Lr9uajEmFjyneH/3n1huyHva3piYcMAbkEypeH5yzPD456HBJ/mqTaMjnt0bLZxwgMhXGICsf
QVLz0BL0x/jxIR85gOiwdC6u+ttfT83agBPeNE4Yk/Rb/S/ZSGHl26Q2sspjEibZcT/v1YjQxHjw
nkMDzJMRsjX4QOZwspZUvr2IcDXKu0TGkqBIGqrKu9MA4hluz+glpkCGEafk9UPyJEJuwcZQQ8El
3IIOIXIuOVnhQ0X4vEK3RwEwKG1kyo9fvqQkFrPob/uV2hs8nvmCOEFsJ+Et2eTgBN7jNee9Fh61
RXgISpGYx+YhF2aRWaeB6qEZXrS3JUFPtdZv/cF+uae0R7VTdAiP+RsB8oXP5Ffd9szQ/U27ZKas
iSkVs8M9L4ieEtO1roXO3CcR7KQleDvqLJ9QvPRQsk8hkRDd+ObC+1OL1BLVb0IyxqOLtjWKfqNH
LcKCFt011iNYvtDsRKrSbio42G19ut/vBzCKVa6l4lNXW09JZR8MDxCFsg4BkWht0mzVHN6EyFzC
z0Xty/5P8sGzBdw4zMGT3cKD0j0Tszb+YfZvQehHejyGsYIKAGuQVBu4ErowdxFkC+tKuWIP5Zvl
MwahbIPgQXkUwwbrSGZsJVQXzxqPzUqs7b/py7AzN0L9UtsdHXbaoMBonPkWfnhFmKBCrUCqVEYY
zmbGxjbHaWouZKoWqCe/mwe2yksful0knaN87tzyc9ARoJBuSbAUt1kh7eKZCDYXMaXamVpdQUMI
OEQxGBDIiLUbJXj0ocp/H+G+HNalwhWdoeNY+4wmAg9bpTWk4Xqqk6FbI15derZEwKwY1tdJ/Ngi
fRdsgQCS69Gyg7Ulqpd0Wt41g5arUW+JOnl+Dk48++aF96TQJVjBrzgU5uQkajwms79+If0s4HiU
P4D3eBukRnwGamtriuBh0d59F3sXHBBLxjNrCaruWeD0gKImBmAUTnBTMj0InPf9CeAWmab8EzB8
P3jKb3HFqAyH4oTJ8Lv24bmZ2p6Z8b7LqGqrp3VgZwAEIUNH/BNhvXBRT+Gn2ZYqQc8D/TATj04D
e+Y29PPfAUMbm9w0O1ofh0PV12aJMojcb84LaS+bKR2ObUBXYtLAYi//P2jV1Q6jYNjkG7Q4BSaZ
T77Ii8p69FPCx6B/GLVTayQhPcbwe1QvcHJVstM2Q/JQTSS8yQvkHevSHoMSonle6XHYokURg+y7
PcEutDeuf7lGXo4IynYrl5MB5/vWUpdJ3R+Acv9faSL4Ocy1LnSBLh2bdP0yoQ8p5d5kpCOksq1m
/IBIE1Srp9+fbxRi6oB8CEKnR2RWzIR6i5eDUa6TAUefFC6OB9/IiZcotdLcDtQzUVfKeRIbsCRn
M9sPReHMj0XEF0+LCRTvROh0lHj3g7XBGCOI7Y62lzvzfmlR5M0RzbrdSasessMKxdrV/X1un5pQ
eUuK6fx1fKq/4fR/7ZvllBcmIiv/sW7k9QgeipaamnlFJ6szf9OG6xt4WjQ4/a3FIeILK8gUWK4A
HBpgFtEVZ/ufg4B1sZ9TCZn0bhT4KMo95R7x36El2BimxPuiEPK1gw0wuEHQZ8E9K7HzHUSkmZrl
Jh4WXlZRBbSqQxy3oc9PYeGXJJX/4MgQCyIqkldiXWzNfak0TehHbRaRkvPzhYPrqp4RP02aL76U
9IwxNg61lJqljP04yzw1FKokcj7lapx2gFwyxJmrtd2Bgr7RCCQvEP+JA8kWBJaOzJlKUyvaYCp3
M8fKu+w5YphpBuQTdIMY/fBJ1x16nN0Jf2IiR1GU2z1/RJaK6igZRi001fDCYwe4qkhc+LFavGjX
U7TAW9Gs5Sm9WCKhtI8R7vbxWvPSpzcD/H5j75YBSM7RPu5Zg1hkvDTMxeCECuCRV8qBd17+X+m1
9ftUU18IMBPFckhwjNV+PkBwjlUN0hXO0o7CwkO1nBA8J0UlRNFgFgrbGs7hTLe/s0NXzlbWBggA
VVAI6RCjF1XgVIPZcMODZPGer3KoGKVdSE+kVMofCtRMHIjdkKBJ9ed+RIyyS/y5To4E5zdaGth4
LKdUO91NzLWpk0jHTqnEtBrGyVr6o1KMg6ggqOZQ/0Y+LYcPs4kQ6dMOf5rhk0aEzif7eBtbWuzb
e/6u4jayiXgYFFEEnVzaZ80oWkSWuYc1A2WwreZpJ5GSNeUvMrNZBsM5kBPCKfi4HrxnpJBiQiYo
+IANzPqUUJmPf1dNOfCDa/i2Phkw41cWYv5tXXX3jDmwNM+4cM1qxhjFgafvrjN2oHMHXq51dTGP
s37VZvC40NJC8vbbzKdBN5c8r8FJbe48hr0/Ze36lMnij92EoKQCRKCaIXmeGXK794ksZhLT5tfb
P/BRVAQD6BZmI1Gvo5wrX3qROdFcAbF55rP9EFqTBaZIClBUn99AF5V/S3kaazEwow8EPPRkmi4y
Nn7UiUIOodxozDy/7IGC38HALRtxqfnzEkMaVHpiGWrh2dDLmSkrohrkDxxhKdL0ySCU003UGVc9
vy1j6VgfHN3A5SN9Oi35xLpWu9Y4GL4JK2g+AOGfDoT7ticqTN0ds+IVWcOCwa7z6o7WtIFLUw5o
HjHSzdj+sqerqweAVg8IO2dwvtHAoHJILILAJ88R7Nr9DhCF7sQBKuH+G8eH+F7v4xq/YyFKdrJ2
zwH4SbCtE8eWSqfV7OC3iBg6VzROymYC+hdZMkNvYDZnD9FXzLB71SzfT5Xj1kDXBkAqk4RWbq9Z
VNW0V2wtwdV+4Qiv5OJqKMzBGXsGD3+Edn+Ex9hNXZPtvYT7xZC+0GOmQVbJIoP3E1FvxDCSrsPy
T6JOLmcUrnRVFPdK5OoKl/AuNxu0EZEaopVH8KZcU5i/undkRE4aTdVUBN+cYgo9aTx9LSL6VnuY
TnR+uxVd4bYaPOXdewuLulLHLimUYHOuauGsZDwBXvYAEk9P7hdqIraB0fzacD/L2gLMrCB84lzp
Hut1bO2RlOJ+K+94QWdsZITm1rOLQvgkO4kptW92OKho4ReqpaXdrHtQhyzUD08h+m4KpHPTwE9/
CJQiuVjwmbtt4UlTLraMHtyofD2OCzRXh5w9ld/bNi8cteMy1njpyEZlgmzCiH2Yc+VeHBaNCCPx
yGs4NoTH5OcA7PecEKR/fTJFBgpsepGLdPwozPYRNfGNzrkjcMSbJEYPDV2OeMcLOhfJ/eee7h7x
FlB9QHGtrcWYAd1KRj6b5ZiFPXKxwsIHDA/5imXjaHG/ohRF0vqBfW6qTypD5oPcokMDuiq+/2E/
CMmhzU0nj0AKAbLifENuwZwvFM8RneBGoseqi+3rhzj8oPbOvT59091/p0nTEO7PjL/zYU8n3Eys
rHolBnZ7QacORJPHiVYGkwvFvtxMPKzS2aUzmYeEdiYxU+pM8gAbftvqVs+9i/wryrBo2agD2bdM
XxHhEr5kl/psVfstf/jLSDLyjifiXP0pFxId+BIwAoj5Y5vP3dtQZSH6jwK+NGRVaXfYr0C9XP1M
CDTm5ZStXFFKI49ehpbEotz+r6AZosOzuUYKmnSfzdQfrY1ZW1LdAVGvxj9POgclatsbIKp5XDzM
kKA6i+KQoYAs2BMM9yk4g9tPhQWOd2ggLJkpiBrp0WjcPD12wksu0hMSjsFhaYpzZsRUDuxtzoNw
wHDl87ZAjjHlKSsGojPEWH2jP9OnE3fbQdfz6tjhxGdt7pCYp1MwjmdzXev7dVa7PSN607ySK17D
KLpdJg+AeCrAjvGvNnUnScwmVMU5r6FgmrSursdKamH9Ttsjzf98Jb0uvmRpQUKBjp5zOUd926zy
9faLJZMxn6KBQbf71x2XT+mich/XsI8njnCiQmRJmFm8cx0bp03KICkL2w3TQxG6EHzfSZJy364Y
4n5QwJ72ZxFpgwUMhCXaYTx0sc2RL8wrcq+rPHbyfHUmgtdiewhWqvrjyMU8fF8s2VZioexX05EA
0+kiqcFAnaptcKFPzEi/RXan8mQ/AId1DoQN+qDkDkACH5RzSZX+slpm0v+0w7SwRHMOeee5V5a/
zQZbCb4+xRbOajHRyOYBJMvSXyzpYghlh2lyqQw6ahAeKSXIWTsIC8NwvfgCkltAhVxDLN+cn6av
ahw2B70rjYPFhevtwh1mbFYmTmTGf6xby+aWlD06aENowCAXAThGDCdYyt1jKNzmsLAtB/TzP6HD
WVVFC/YyUwJB9o+8TVduJznVv3sfKng/SEK/tc2RfSqjF4NGlbey897IfIvzaTGYUG2ajRqdMDNX
xqpGFVwxQ0JOmfkgxhHqDSEvNj8XcUwRRA11soGzxyYnft1McHt7iPidS9dQ0cSfkEknKslRKrgr
hGuqoLMX29uGW7YzMf1YUJF9qigy9rtAL3bNtLtE7ioxP9VMS9bNLAbMQO/yMaEkfxz3BnlE3rfE
EC+MHMmTFJF8jpUMPJMPQcsTs3zVdWlAwR65JD3JysTw/8kqChNkbXuY+21cg0C6aebuJhSupDO9
coeMPd5ZqeaFXjkmg/WDJUdOGMI/QX/IJ0f20k6FIh4cQ9dDXH/JoZz46benNjEO06QJ6Buut0mx
9XXT9PfqBrJKHwauujtJg87Pyquyw2dI/vjSCyX7yKrfgeCvu/dtltJcP4AlUACnmyKP+Yz8JV83
v1gHXxGJaWTcO5476juPwR3qztsJz6uDfFqfqyp8+ZWv8yNGb23/nUiGkDwEVVsn9WF414PoZ/7h
LiC2QjEbOqRe/tVfsCx4/1Iu6SH/6pOhwJB+k8GXDtta2ZaQ287F8xBlAkp6gorUC1glXu9biu7u
OVHUrP2efHuatpbI3cmwEJr6abHzP3F33JVKqIWZIFoRkfnZkaS2FxEkCrRTLZfabMfRXbXut8P7
Yl25D6baWnAgrbksmHZt9C8wTdBaksD98611ORrhWMSEnfc38ykWOHlCLuMOP7XSkNQion/b8bAS
FGzec10mbW6x/TMnQUsrDyijn0LTBFLIHK2pI4OU3nJnuwqMGilvl0dYH9l4iKe1sqsQtIhuL+sm
DXH3DuCrD0pNz8dbF5VKy5lJQ/Ivne8ZivSynhmDvUwu0tBrDPG2Q64rbveZQFK2GgtFzTosoqTk
rtu80xlaVlN8BhC26qeIfBSrfZvINnhbGxZfXu9ZtwjIcIDjz11TQ8ta4slEYIHAcOQMi0XK99kv
kjm2wk4tCqKXVZWEu28RHxGny0hqcVJgucN1YzUq58mfojQTXNdFT9DOtj698eiDAB3lduz7bVb5
ihaUGCjEQcMA8LrH0i65/NyApT1eZVu6rFphbOZRPi1iUoW9PDbwT9XjREzaaNZ7+hbePxhhc0y+
TZWQ58TbmnR5WCfAIWlAc5B4DddDflOmvSGXAKlqu4Qa843i5825fxeOhUGZCQmH7DHtg5dwxwf7
pamsjIU/GZQN0c7yrfs5gO0EAZgX1xcaPydCLZ3islAR4dXqr2jzPo1eOdWrv75AZjFaY7GOglYY
FUrVHJNN6a8Or6vkmwMGoH2lu/rF5EbDjU0mOPZsZS1sX5TVod9t5J/p43y3eeC+Dq0r0Db/61kc
mmnMTkokSEe/bzmWNIf+gtSj+HYs4pJUwhJ0HAddkFCdRPp+T7mL/d4QA1Xe4A0DEg0gxUhf5CoX
QTu+ZZj+g5d5wwFUgMG60q1MLgeXchA1m8goSHWUNQzpekECxR6h+FnjHXBKwaPzcrSA2+/PhIz+
ICdlLMePyKy2UppxO3NG7/3nQdKOzkWY6IGo+xnDECgsZ94ildu5Q/gr0zgGLK62YGX2cJOsCtwg
JQD3SUNfGObtgn4RMixNQEiJUH7hk1bUFzK8qwDTT1h4ECHIB6y40rt1U78mCo67YLnZS2w74Z4J
eSCITbgXAJ19n0e7kr+a8pwl1KT2k5XqerTCcXyV9Az+uEiSBzaZ62LogN2m7GWtgdBtbE4FMpOZ
c3ZbnpatEoz6UTvoyUd1C/DLoTDShujxCiHPv2NGwv7MHB/YBjMia+DX/admulW9lqpdFgOAjpXr
GSDLzXkNQgaMQYlMA0VB77G8GmPvcO0V1WPvPCx7Fdtqv4TFdME2QxsvXRyDagb3TE0TWl9VgV84
RJ1vtwvmbqqJuIwQBOLkw2RKoHR93k0y7NFsc/ZMqYjJoaQTiZTWLqy7Z5uGZxKOWUNje6QUg6jM
7SiKkVuEkhYx9yvpr2molSoKv6Vh8I/ezR811p7/9fyhyigWpcW6mQ4VEHsr0ATgbmkqAGvisaFy
CLk//S9WTYqIcgMQ2snHfHRQ2gf0OV7mW2gjR1AyPYSDOr2STUh8pTh7kfEuRAaTyN2kX8HCak0x
eoyR8KloZudA6DFQ9QiZtkdX/GV3CFR2apupFmmxhKkT4PtmZyVD7p3Aq2rSTOEhR/hsGvlSfKH3
KUb17Xl0rCa0Ev1KaNEKHIX11RdS5ga3F0mO+x8Y9ZPHYx6dDlYiIAGZMb7iMdkgOXvVpcZ0MbgL
rngoNnweE9eiUrbXqf/8UO9E5PKMrBkzbRpb6e0/cUXyHP5QgQ8vjTCiiX7pQT5vSLknm5m/vbMa
hX65x/yclu1yh7IAlfMTaGApm3LD5j5Maoz6wLcD0t8+R9k3kiLR8CDIQr/mRsZ9mvOZhmm6S2Ok
awTB9Gy8k/ZxpcqaaijIH/xIVwj3K+o3HM3Cmn3zo9LQa10ukU1lyH806AmTdwuayJVFQG3Z82JV
uXNjQRz6+xqxXc1bkQ2W0Hs9Tk+rvznqEohJjfKGlyia+W6T6aWplt3Rl0gmmpWk+tqZHtmeHgji
aVBn+FC9iF13X1fpCJ8/7B7+eiPsFRcamGvoolyrUhzqf7XQZk91dqvNHhA+S/5C1730tpR8lbJi
5KmxbrRG5FJmuLNWo9ry1GO3RLPaRJuMdA+n3iwBo1OrKz4B0yWX6034fOfoc4suokDlZEwuhYP2
W+6GX7i+qqwJ6Uak2hMGPWbQzIa7lUf6gJTdw6DDH3fg3j80B0wrejV5AcMKzTEHj1cpX1sY+tuV
XXWSklw0PCIznQGOuRbDgS4CE6w/WigmJOP4v5HQc+pj+5tPMN4aheScHFOlz7i2O1b7dqsV3lQK
lnGmVJDjuqXcxBLuTmymcz5JHp0+4yWKfmFxfxKX9OsLY+3/3LwQnL8QfCZ2EaVuqeUESbIzKTMd
nEcjyvgQqtpeUfpjssEST7TIU4s1XdF074mjYQ+pYQTJMPvxytAd4lh9+xO1k9YPJOT0LOzhJDw2
2MYZr4FZrqX0oQRK+JyDZ3xXh1JzvzzwK4ftpNWs7cMwjAeDkcPZnde6XGkP8tR8sML52d3wV/T5
HdRlBkiajBssaMF0EyV6LkEt6RHfml6LA7mD+UXfnP27/IMDSkX8Nhnqxe7tTLXzPf3EXlIT1sh6
lfA9CE06tUVCW0NbptZA92CRzLvrtk2y6+iAEomgRxh0RtpGi/QaeHGRYEL8VywGN98Fos8vrhW4
Xicuml65i4cTirKIAp6zfYCUArVTT57ZYUlmy4YxLQmi2sTdIhFlYkhvTIhpgajb6IYqrJM2EXOM
xVZ2Kdc8WnnUxfSmmmFGj/RTjjGjkwZcSOJFWHPq1vjJRpmz/EJJS0OetGgdTDt68J7N0lleFzuk
uba2VitL4YaiGqtBuAR9gL+lHmXXcfmwjtgSryBINpD68hi41SZoKO0R3Nejh8WhQjHLrk7RJotP
IPa7WePregHrV1PoTqnZEZv5JtusTyPNaM+FcYS+p2vQZNDgsI736gisbNP4SEcuvWb1kGkAgWKj
k3dFYV7O01UQoPynF/GnEk8JyXLlpaP+k5UyFxda36nNQUmsRfX1abPc2QbX3fN3cfNhcsuWlGuT
WuJepCavFYoySB0G0jWwTey1ujn1XpHROcuVn14MbZ5vkHjKjrCokI3lB2hOEJBwiKuKBIqD2TJB
yTxzGbJDd3P8gPZRoxegHjUPcobBraJGg9W189ANYZmyYch2kZ0ryECHaZjjZAr/0dJ6yPljNGmR
80Tzbs/C+Rtyqdwf1y43EwG3P99baAijVdX9n71j7Aud4uOkWdPvxr0++YYlgWv6DDBdvBiZW9wb
8Z8fyUANxaufVeHi/eGUfFxA1H/T6GGHJ7evU/yUELIQVM/mGWJUA+zev086qf+VZwQ0iQRTRnSh
v4sw83XpDJ63G7SrnkL+kZvnfuZNUeIXH54/S4G/p+JbmEIXLP7n3P97e7Xqnmy+8YZCBSIBo3MU
0E1qKVqrxCRrWskGgpWvnjZUcKI/mG6BEct8mUHFuFe6V6t3molEGG5GQx8Gn8uVEn3rkbqVCBQq
GYwany4Q51nBEk2br/5SvDknP7CnpISF6vFEX8BMioWcq9aHLftg+uG8xUBi2PXuq++BTEdymvpZ
DNA4wtOei6Q1WCPNc1RU8OQLVF2jkBPe2l2MjfBD0eIewG5PCWoJJQw9ia+K5oAA4UPjKGM5LGyR
qaSmH6sSOHjjbzTBVlLktNGcpzT5+msEbtbRvinP1l2C2uW+vzfashSdRf6qCvZnyq2qBF9xc4ET
JB2x5IhrZ4WGqPeqS/gGJQnGEmIsaZVZSFeU3WyOuu/x1QhbwA8QMZ4X/NFw3rL21JRb7EoWiziz
7kRgO2PYk+t9PysVFKIZjgcGlvIzUVRklKIABWfmehtInbP2IfMK0WANWaHuHzjrdh3qv5gFY11o
VAj8yv6H07AJE2nidEqZHspoLUbvl6OwVklLhgdpzo8INCgqjh16Sx4AQDb5ZNZK98PCeSyHUQ/y
xyRtg426KoF+Wh586F9+y+WDNkP1NY6RyexOMhY+WcSC0EOf4L2MfPu4QYPztMguJfix5AugPva/
tM8eVKEr7aAiCK3eEF0jiVauEVSoJgO/XfN3uRPizjzruC2HOqPt785U/bw/ZBm5dFzGY7JZdui2
EXVc+eOjYtse1ZM30wW4V8puWYnGUXMOxxVjgwUpz7k1tiApbpcY1MFPV1CE5E2GenG+PfI1wlFA
UcqiBPPvZnM3pGYFe+PL55f2zwT5BVIhiLI+rTClxQiJK858fTLYP504AfTAdoH2KAyPHp2A2jz9
tDSoBhuxbPQrxce+8GKPRZ4VM/2aqLLv2Ci+GITGnwZSXAiE15lxuRHNuiEMfcFJaACydFDQS/E9
vHphc5FPOTYzkczwkrdlO2AogAv5svdvqMk9o7jBKmY/unbkNRBADK6WZzEoqPau1Af9+hWitOkM
d4KmWg0ERoSuBz54GGVHCHLa6Z3z66AxWx8l1QPGddphHyExDaDow3TBhwjBFlzR+3qazjecHfxS
VSIV9mStOJ1cP/y23egxUkZ4FgjlLof+g3NWiUR1wppsnGSGlNoXQ9HiVFsg2ibr6C+cOh+E26YM
ONzt7Sbalc76w++ZXE1SmcJD/lZZTBGwUeg0scbm6Up94iTvLVI0gTC+Me3elZ5fRotvNvInHCPh
Ru4B5q+qarVBCFO4QR9uwPfls9VCPY+jqU6D1Y16xVh95rVtP62F8ZIsKwK4gPJjuLqb9PdZXBrw
K03zxoT/fh8BY9sghdqq0taYNwBm1RAYFNWuKi+6cD2DNICDZBL4z2p66v1J+9i6d8s5L2Dhb+Em
DJPaUy68YrGvjzxlP7OBUm4MdPywwNPyjQWapxTnM4Td84UphG0qSf29+0NwPv3px1eTtqQoLu8c
MWct9DEHoQUFtdNR4SOUR9FaUrovKxED4WmAv6+kg5L1qoh+37DH4xrLdH3+M+aoHTXSH0cf6rWA
739ZDaRCONB/YB5vsMumMfMxbP2jRkIsE2WXbA8br/+kt7+1CzOMeH9qDPP/bBgSSvul/QwwB46i
VDm4307NqoPvcaX2GHenGRvVtsf249Sl5zlS915WFlW1oeW+B4sO2pm5I0GZWjbfV3MrNy6cllVZ
G5WntPTSpa2X0Rl+lULoAxD4ioEpiAFaATSrgetcJ6S9xswcDsxr71ilXaP1YhNFmOS1SMqDKJkx
9tMIkgHNJN64lnM6qHRUY0R+vAy8InMDVnhhK8KLdaYohzPpGV0yc7z6SBsq3i4RUtYAx541cvic
P48wobQmpk+l2P5bE1y1nnCAEgSaGV8fUHDxDC9yZMB4KWAMxH+5InNecjIW732oECGQdFtij1dN
XpJuAOTqUIC3vTYqoylOifOvJRA7OjCXVZ0yORGcsRKuLYkpuWSena1lEnj1ab9uuekkc0aAEzSt
kPx1GQQBJ1P/zQJWoSDe+vzA/zwcBdSzUz2VvbeNc8PUdtb68JqC51/RcTGIY3iqORBh0NBHKT4W
cmLzaThOPiDusx9+k1OTxgYgtVLDdl4Aq8+L2nFUiN9TwiV6dnGbkt1auK6+c3vAFXmfLC8UoExa
v4p1q1JA0tG7WKm+CJLxZlf6tyCw73oqUQjgBWPh0Z1pAPY6/583GoFpN6K0IeVkLTC5yTkoBbdA
ZJlqnAZ12f9U2iCGps0MsHN9wmXs/QEFJ1BMEup4IggYDg1MoQ/+yLAxa+i+2X9lkXsNWL7irY7F
2jOnBF0I60jysDNQZ4hgssGf/8neGW8W6bu+HOEC42RvhzC2/MAObDDm898Oc1FoJVFgfXbZ86yI
g1/Gtik2jAor9kYetFCNJ7tJP63jDFaqh1xiCe5yg8a07w/3yTEP+Xa5kFEewSXETH8mFuE1lUa8
awZzXKXjF05UdTicFi5rNvdiotSywWmp70QPulbiAvQMsjBP2n+LiNy1qTi00qHQBfDCCq5sxGSL
1c3IyZBFXWBU/D6oKPPJkBeuT6o3leqYasVZBKGKEXMWOsI7ky+5pNZGhLV65dd68csquES8D3z9
MNrwO9qvy/FiwoT4RxbiCSh9qVzuXMFAzgKPjfxx0mhowi9p/KODPNpyjJCCKF9bCOG/K06Kh6aS
XOpC0dTtBMha+hZnpTIS+a6OnWQS6cqig3Basi8s/0/94PvBb7VURYokfw6ws3ITNfKmjiNBem3T
jhY8zDVo3jO3H/H4/tj8jT37E3BQswQnT/AOAKxR0/MdEwhfh0HqvK4DO6D4u+yTTyjKW9wSvy25
aHNXZUP+oMZuatZVHtDVcy+pcIspCj51SUZZgP2VHjmx8OQ4l8eaBNXSBJ/9jRd8mbhEvdYoH72E
UOHJha4yh5E/aWvMQdifpH+JLZHVunqvLaODZeZIxR/ZhGC8vH3C3J6AP3IryrEGrl8InLdlTTpg
zwmgM7PkXfluPJcLuxqiSI2HZ9BJ+k//GIs57bijwoP6INPaNeLV8awPGXP+vZbc8nqqzHyDQ6a3
WilWk3SC2VyqW3VWmGvvnBnF5ksZWmrN3SXmod6WWhD86fC+08iWNVn3fQk8wQiqnDA9PhUzZ+9+
9Q0OuC7N3/ihD/SoQ4hzlVHgH6wXb9uGA3WR4KFrONq5yDU/Ly8UandsPR08QGbJACxoPIicrp9L
xRKyDMz1y4yCUXJD4RCMig4nNDbsEvpTTLioU1doMJNmA5mZgZcXYU2hvIXLSFs02j8GHeMhxc66
PMo4WrEM6cNs/up5TgalHWABITjRKU50N4MRV+nTosWHAA8NBBR5YLkKTFZPwP9/flsMfRTttcoX
0R1ewl2EFGrJEqLprDeZbYG9zfNmgWZ/LuRG3GMISpmqBXTQzfzZ1oNvuYQx5dktWuZDZuHd7WcB
70o0K9va8bNGM4bDb/uWxJ+wBtytR1JKsBjCRMOp5WE/pHNGLggvppXFfNMm8rsJDx1/8yCuJO5F
5mzX/RKfo5muFZsMLd4CyciU9PQsn4h2dWIMFjEUS3/QU+TbNn/I8+pH9T6sLkyiwU0taa93vsAi
XWxKFjidpNt52mJpeSI7oxIog7ozu0KErpaf9Oc1/aKemTETdawPorGprudUINxllkoIObYIPdMQ
EWeAXa/lRkaDes+ZNuT/M7s6qhEz1Q7Cr8e08coqNyH049ZI2ynAWDRsH+mQ3Grt4dckEs2/qJ+s
84fTHIScw2Rjhtvfq4UFYR2Cw82mMUe6Ogzz9el6DvS1LFyfMX69mxXm8eKtY8+gR28h5jbWnCzR
TjMRu7mKdjSvcgxJsfz8OWINzurUawpISvDfp+ZwTgpEA3SRhM6iVM9PSTbptuRhiHvYrL+POif5
ehui2ATnqmxSv9oHNQMS9bNrRBn2N9PjQklV9IYaBB1IaNo03tnNhFi264ezpfW+QWlY6kd+fx3P
LmmPECEnmUc0j9ESS2+/mJkwoo/7Huqbi9V5ILH/xDSPbxZFfT030N0n5roQwlAcktZ8oWTydCWl
mCU67OoVeQ6+QPpm3K5ui6Cwe2aSf+W66ds7unJhWpUL3+A8AJ0W2zSD3S25sK/92HttfBGwm4+D
brlDje2WaCRPnW/y80BeS7OFUuaeEhzQWVH4Pa7WbVCGvqFHnMz+1O/9v/ZTTuz2womhDM1kEE44
3pK2JOQr5OKpAhepZy2maG0MEcM0mJq/rChXGdJXLbegZ93bIYr5/4IZwNj4aVV8vbWraFiFYDok
Kc197Xg36DxwHrQfZWG24V4CYs05qR0v56bNixir435/+dBMx3ezpUGjJqiPWDr/+yq0z26AbScp
JCiErM/xCafnb6EozSnlXZydS6eMfj19HtAStczr+1cturHxFiquGe6qXOB1F8NwGLuqJ4ipeohG
i+zq5bfRF2pkYH2TbUy4BevvYYM/+e3d5aKQi/hpIkUvu4pG1S9vTcaAe8X5GFknnWNVf98gr6ir
P76UquVC8rkesEi52XQ4DvltvVs7W/6o9/VCaw9agWV1ncV9iNGPyjhKpkVikPGJEB8evwOCCeRl
d7x4llxi8QWpEsUS9z0/Qli5KRbH2OR0FZQgUHSkK/OrNCADzyB33FGlswqlTjG8nySChhTl/ibv
yWlIvmcm7+gis/dklUA2iujwy47+5jKd5ZSmFk+uE1wOYoneHkIiULZAYoF5ZFMoucQiQulqQYwO
T/Bhc2lx6WHcQ2i+swWPEKRuk/Loh/IzISWVl8NfOV/Kb4o6fNo7nF3gkccGF9WmK0GLHynj3zHy
NHMjrgJqx0v08s36/8qrDyMhVnFoyq5vVUkW2ROiq5JppiSvXIGl1f2loaZnMpxXRhVx6YDWoMZp
LYlf1wET2oBDVRLZ1BthG50T6sxNjHUJsdQZV4eXQT8zRb9Z+8WWvkBy9cZiU3wmSfO4stKpOOtK
8x7Ohur4e7Kpxo8tNCIrLhh49khFkoRWdnB9eHVoSaQE2TMPln5Zsl89L7Jo3Hr1NCaOBkez0jMw
As4Ow3X1/j/NELHv2VX9BmQ5kUYT6uG3ty0dmYKDKXMFkJFWMIIIYs3z6Fl8njSgvW8UshAMXMgd
szJ+jhiDGLtfEuH0e95vpsHWzpKU4AJIuzw1gjGjLyoIJOC7S7q1I2F+/XU1sBEOxSTJ4ze+leiq
f9SuDeeVP5y2nUY0Wu7+GqOO6iPz8/DSJZ7VGeR8YPUicdV5BdWMLhP8jD4BZGjpVuIbdmcfQl6a
8MpvdBlYYQhViXAzb7LQkTyx1vq5XMyI5eNx+hGMeVlnQE147w6B6H834WxFoLvIX/hfwDeuhpBJ
JyyI+jG5sux/O24U4oPRen9tdETDtJ4EzkLWwtCnOUjZjOZNmBuJWCG17uVLnx8N6vnEIdkQgNRb
PSMfD+WtW50tJ0ly11OzWkC2SEMfodmYwohcSi7BurV3cFpDQO9pHk6ZmxzpocQVgAvq2O+tpQ==
`protect end_protected
