`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
o8aPZVQ0BxSqgbNenLKYaM8OG9BuMpMLjosc4pM/4XokwsnXiWNYPCiIqtdZXduYAFKSLbO/JcIy
ely4DWOpVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X7RLnFiGs7YNLCpniO3IFa8dL0LL6kXh2JuOv3Q+ks9pDRtxM0hyteUB9OxaSXAs3et0laoVU732
S7YBeuKMdcbMKG1glHY+nTQSwcAg5ySd1uCpGFnLiryeciaLwPlqMbkaoCztY4MU/5udJj92CsaD
5m4tdotJuY7BJtFbmnY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Iq1KtT1oizXJuvWScrUC8AGDrBQHT2l66zYfHcN2c1dKrLCgBcwpXtcpqfrBjAKa9Fe2nXVUNBxP
xiLw7RCN81PI9GX5KfofCPQ8S7gih+kSZuf9SExNS934twFM9YoL96eVPCCNzUinYkhZ3eO2oPIV
M2RLffKZio7oTkGAPsuk7msJ6uYugOVmQmyyEala7nWDXYOF1DN7ISVltpaVsfXdceXx0ISW/puh
aSRVtoE0JmOLo1sNPp6Ds1gu1J1XRtCJv/vO0gssiv7Sn30aK37tj2dPYZ19kT/ZGmJRhfBm16yv
Q1uEUrkGZIucqC4bZd+kbO9THqy1FEmpWhs4+Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vXBQkDW8IPd+SAbz+VT0oLGc8e5BDDXxreZAHG0Mbk+5edp4Jrjv4wHf7LfYiubYwrNzWKQpWCVF
j3Z5BAXsqTJIuASxy/xBV89q8TtlsQNQkbVdJXd8Zaw3qcZAJHkBLHeHlhEnbboIgmug1ePbJ6pq
9eNKMHh3jipZj/Oqo8k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lrse2qNm+82AMBhVltdLqPRTQzgawu35mrgainArfeF6W+wGJyR2qr2UjVe16wi8IsprVcTQL7yF
tIE9NL1gWdowgTDZQs791L2vVykzuw1cw1lquy8wZIoYlLv/OiLXeTUE/fnh6DAnQBPNY9j5HNRz
GVuikrNp725qYKLHHpFAErYyrMAHZQKl+ObE35GfgGvaoS80yqt8EPAofkFitjinvBRuGMMcT3Ba
UPiK06uKMdQ1VD/WiJafbjSLysUWJJZJ4lu/IH567yv2ULIqcgCWt94wcmL9xJr/oBuidZYpvIDi
UNymE7sBRnQrfldWcWVuBmHxr+j9GYjGqyNh+w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19696)
`protect data_block
lVITVv2PQktlr5bJRJ6IkI8Mqgu4fGWZcNiXYQaufRkI/TNyfCP+eReUfefdooGTU29cHA6fHqxk
0PaZdrMXMwlpoSMoMx0Gqzxk4WzSq84QabYTOHF+x4Iw5tviqPF9eIB/6KxJGeX4R8MdCyQaPPaA
6lJqMX7CPZWutljESd5YAeno2IRT9ErROJiF3Jd//6cknRtDRdUJ2oiGKkgyYmvf0XmWU8Hfwi/v
eTTRKI4TgtAyO6eh5aUTaC6+KhFKsrMm3165cKb3DNhpdmYgN3D22BVLErwjLDXEi5CIAzCZovpt
sF15rl9XCjs4jUlSiNfgESD5oEOuXb2zTjfSaZvKYnMwuang4ECfOs7zMRrD3B5pEEVLk7kjHnkH
4R3cv4r6BKAVcA0mzPz2EoUhNnmsqMO30u7/SSVNcVM8pT2hfNS4jIv17UiS6teYjoGMPOSXIibf
ZD+D+o7d77hyVAXQWqhaRzWTv/P1ESr7oCjPjPsqvGwiywCbiFa4b8/HiSZAT6156LvrorF7hmby
B9Qh1xpCIrl5a49HW7bZ+Gwywyt4DQ72RhtC9WisPfSpFt+Pplt+0kz6yYD7lws5XAMb7tFYu7aI
ek6T+cJB5OHwEnCu03DpRig083SUL+L4sQLMNxwqSaEywo3Bj/yoJh9Mqa2xV37cjPqrL2nraGMj
BYCiKgctNWqp15FVVXLEyx/CiPHAvp29YJW6BCGdhzS+IfgZiIcfborUvD/yOx6R3tyjkN8Y6u4r
0DHt1OCPPOsAob7GjMalX5NhocWbCP20XGktPZJrueeQG9l7imyun8dLh6HLensJsxg6QRhfxYCH
BIR/MMt7ftu4A5bYfOUGH1dTU3QvX2LFSLTGl0r95e1m47ygpyeQFG672jmtVKzKNIja+D4/CFFI
VlWR8Cm6tEFumZJuCLwdUEY+qOyYO1aUU300s77BIjruz46niC0ZOhphCan5pcm5Qcar83F6IsQA
A16se5t1Q0WmPyTvxsX6IvE2U14GhbP7OOZdMOr2eV1jN2Dk1az6DE0zMrtQebZlRAio9RprhMsF
q2uWnhvdbJnqxGwluvjfA+NidqvePyQqSjIuCeGVVS0XSDNIdJGSt2+cx/pLs3kQIFlNKgBsXW2w
sfeTl81kk4I6W2GRfJRsS6HBRbQl4XxcCMrQqhYirEMZKOOBg8rqsFszyMDK5VLXqOaL3QonmoNF
2o+vMXeE/3A+NLO+NIhno1uEZxhMJhzxqGanqvEpAANtzF5FEU083ESM/Zig0c0d4IcVJUTay/xX
gBX9BflBYofzLGfTaSvzmNuJRupEtwGaQfVhM4IV9Nuc0c5zaTubzdxWSPnU00l38xgHgA9Dp+3C
R0B/JeW4G2B2r5RDbbpIKAdD+JXARV2B9YQM5T5kU3GX95bkjW0WarOnfX7aGeY/26mrgAWA8pnZ
LrlwG0n0ojd8YKwDClVK6R+47m3bDaiT9K06FD4dKrKEnISu8aK1pAXk8m/qJaya2rGiKHO/G2uG
v7DDXsrEN0xtz0PmDUgl7v5NJlqbPkzNhsO40M524s+WzeI5WuHu7xX54+/uut8OmGusYNk1jUir
rekvK1EAYfoZ0uCj3bGv5deAgVK/ZwVMiDned6E85487OfFuBINFyb1gtwoxgd4ReD7py6W2EjxY
v59bowfgLi6JVCBn7wNEYnfSzzALk/Pb5eXWZuA4QBXnfvsnjHBw2z3/RHLcQWNPwG/CHIQk+FJf
P7yDi2sryzzSsjmqJ39S2WHv3OPt1CK5FNuTizHGx4Re4Tf2zEe0onc0WssCkh4rrRbb2RLDDIQU
n3yPXVUVuVHI5YmnzMSmFrP6cJHEpT4lSV3sWboPc9pJ1Le30pQavwZvDoUu92agYCf/fXYmafLY
OrfsFoP6vtS9KmOixnnWw3sPaXA8OG7wGn3+GK7wch56sAF+3YH/EE7rJk/7pgCpxFY5PzG0a+Ck
vFUqjoAvcaD+8+Bidn8l4/PvDAqys/lE+aFaJX6t7J7DcxSMnb7yPgTr4mwT0894tBh6264Bnwb9
QaUkCMqAsD9M75irOSGv//phpm3y3X3WkBgJIniGyq2pzGrp2HM0Uh/PGAMXB0PCfLUO6GbWivJI
Gt8I+Ua0aBc6sVG1BjzMwMq2f0Od6hANgr0VLJId/7k9PZ8ebpAINL+BOYpCnaHd7FJyWdENeC9Q
DFjPYZ8uwFeOXsw7SaenyphQdTLi0Tp10170yBDdDC7yuJYsZvyD4vWyxZygjE0uggFSxHL0l697
KyXwf7+dg3cU3tmsKualCkhijLwbyGNmEsr43SccQN7/gA9nAUpmawfi0q1DdkRcBRwFNufer4Y1
31Eu/lRHME0XI8wEOuv3QBxQyd1mfjxGhd051siuCpwTlcxcrPoK9zH9agQ97fb7zPWYa8dHE5yB
Ls9jARscx7yePW5OojrTR1I24Q566jcu8muW2ldfKxNVhraPlltQFEwYuA6RUfzqugWEjsR2PCpd
1K+3T/AP4bTTRqH22LEPWeD0XG9pQNcg/0b8IzX43Iv3HSRNgRt4JnWcdIHhl7T/D4VbU3nUhNti
B06UOKnfdywWKrUJVgi1D+Iixx1/K74UYnDkRFg+b+fIhcfjCjSNbFTB+Gzjoi+3PJefApLwjfxi
EUAWtIENoXmXrFS1AS1qA+xmife0N6BeANjtFMQHlfNVrQs/EY3nOS7cruWh1tZZgEYy0YF+5D66
rwIaQc5HmYW89D292dTN9o7MsnUgonibkaMovWsYF98te0BnqcKdUprySyl0M/KQnHXU4l5AFzkU
Yv9kAzqnfgTD6vHCwruCndJ7UpGVFa8m8j5gCXIv7SyxakvIuBL9EcCl3Af7uhzbc1Fs15bLcdIg
IxpUuoES2kK9fpX69LxpPQ6IvmHGzvIxjh3MmVLJtqoyUahcCt8y4f/yWc1mCSadomK/CY5lzdaw
+GM052R5wvzXla8G1pmV2jXLHjl26yKkICbOigtpdlFXM5Of2t44Pdv8gsd4ZZambH5EaFVj3k5l
2qkpALAHAkG5CU1ryEh5MIrwjDvfKjucdtlod3TzbFHSo+boBpe5t7GzFdN/Q4yiktS8cif+h3kB
UKAmLZNqbYSBrmJvYlSAY6v/7hLkJr2EcCOwfPnGQ2bcPG0nLKK50nk/K5Ox0KrCzwjKPc76M9V1
sI2/bwMYV0q+fxTZON01hYTtUwH7FAWSj4TZCUqIOKkLTACqOgVHcEMDrdAUVRcGmp/9EP0U/pZd
aKjfBGd2mAhjmKcrbv24PhJ5OZILo2Rr3sll0bd0jOb8nbRaM6mlHG4J54EioAkXOPi59j31LUNx
exyB3DhfGKyECoLq6SD5lOU/u3shOhE3g3TdqKReyzXHAKEv0vKSxh86LFFyNzzIcuaUPIXzwgdJ
hEf0U1gPqBMarKdLg8OWELSijLx00pX4+jopRigZQZ8/7KhwWQeq880ilSxUPDmZhQNiJxJrvpvq
P8I529+OK3zan+xLND9sHgZHWJhT7fjxBTNrnV/rNl1CXxoUV7XqHJ9qy6s1vV/uU5bP58pp7Pzr
YKulzf6bcOzkUn2418Ej5k/v7xlHypHAAJWUlZftOljBVgB88MLSPp+XEkBRL0q/+Xfj9Ij884sj
EZ2AJ6CIZslCVNSPfFbKSIkF4UaVAzqV2wp9lwu0nGsyMi6Gpb6Htals8TgLMD/E6peWd9o5EMdX
SksSsIDRBNDHZZhbN0VpeMUSnewoqI9BX7dUb5zvvV1tfcIeshkdYLD5f4HnrKR3vJvdRtdg9bWX
itDJaW5qGbZBjijdJqSv2iGwDQvUuqoA82Y6hIA6HBd2fxp3u6sopkdZRjsPgwUq+ndUYejtzCGT
+tl/ripJMBLtdWmDCwBMiLdsQFNb017luBKscgZ0Ah8vUHbyshuqa4g93xZIczu/UzjchT+IgA9g
lRXOjlHg3RmkGeXISphHmIvyBKIGH949BcTy0uf02n/BmcLct8c2pOUhi97daUPJ+nT+/wNmYY/9
ZkDva972AX54EmlKh66G7gf9dzB4rAnQVnUlUgBmfsicA7ilyOd2ycXzOU1e/70S3jpUblVCAOUX
O+/l300A3j9dD+DfHyu84Craf0jhqqeGl5wVjA39PiIpP7ofsh/rRpX+XYWeV4Zvdup0D1JVOMjN
IZBSPg84QkNOCh7x1R3L9cVk4IhLpf8mffsPksSduiqdjAkfeM0KqaiLK3uixFnnWfhEgxYZtDvw
XvG+ZgdWvg0EXTPN1f+hVZ/rnqq+sk9n5IHpmk/iCWlWoZ+cHgqFztvInzm0YEQOX3FN5Rn4JbiP
Ph4a349XvzAvII97ELrdAdTSq6H1yzGM/X7wJhzx6Ysq/N1DGjSN60vU6mya8QeFc6utSFVICtcs
hJzalHtO3wOF0a3lPrw5dctl9+zqRRE8e8CyoYy8/uaiXnJsZ/As66003n2QGKk35Yi/5kQ0iCH6
ZrPtb89udU3C1x5hw4n4wl3tdloFbV3ylX3z0WsbXLA1v85yVWTQEIdILpKmO3lTR1WAqfyef+Pr
tF895S7VIJwYpH+zbenfPOZxF49FLa1TTUq+9gilarLf76LSnxdTruVVQpHuM087CnxoQLcFSXZo
wQ5eTkrx0ZPmfkZ62A7RIbOKxlbnm3T84aK2Z/eyB25oEYa+nGJPv4BLNs529cdG1QBGUtBOyl/x
EU36hO2DWGtkCIeF3Iw0cKXo1rkteAv5xwSg10tI09wj7u0DGn+tlmTi3ruiZ4HD94Jtgyrw101R
2g+owViMzUS5F0AJs8dAIsRiuHMmtLDezPYkPTKlodM7YPgpFrEfFGsbZOnppQYc3j7w65g7TfMi
sdJKPo46hzBSPqyHYobmbAKft1Nz3hJ7zK/MPKYiZB1N2vHJFJaiQjF844VVgwX7t/IR6OGKkf99
XBkw3WzEn/SOxc700QfOM2R8mM2V+LUFk6FgguJdLVBIweHaZLGUZy3quO1v/Op/PqvIYoEuWOtV
Cu6US7LTCWm+OYXr7t7CxQCjxinXU9EfVWeLVFwIj4/7leAUACHG5iIZAVCaNVJdMIrUSaxMDNzp
N6dGo0lHGTkb8rLFEYdkiDyAwsf/yj3nNQJd4mBMg9wxz7TCfbKj47W21/kOlCk0Gh7l+3MAyc0Q
k4xrpHXQ6VILn9SUzaNiuu3ZRDLli/XEwvusnHXwETsydppJ1+N3yVhrTJ202ctlHC15/zGGM2/I
sFI/y9JqvTTCSnIE2POqBVZZzroVI0EHa5NHA7Bb8yuyBc97JZBpxe+UzKolP5uoiKOk1d7xEm3X
tzqHNdzLd0ngDyQM9dMBnzeOcgHLNl0skcGJ0X5pUloLFRISJR0wFncT1/6WRVCcdPU/IqbyRjXp
1PF9z8A80fgiEDFbgHGtA9e6h8HEzNQskkzmTa/fLu6ruD8wfk+BHekB+14KqMJt/04PMQJIvNPp
cKuIlLqxQZqoq+KKqvADDrwj1MY6+Wgh/2zFRBePZJUALuAZecKTHFIOELO+JO+pgLwQup5H/96c
4HIg/WvF1E79gzk7cDgyWDio/9Q5dfMNtmLN5M1og9oqLOMxkEgQZ53dupQFw4R8YEUxZYeifDg6
XMJSRH9weecvVEUEtEY3FlBJVoE3cg5Wx1Wmagvjz57Dgkd+Aj2oZgR73SD7eO3HDkYQm3CYCZGS
NzfkiWVhZE2CzOUX9A8g48AnYxvbi6VdHbxZFl9lbofkNTuuLSUs8xxa1GJ6GssVnVbyPqBGjEnV
HIFjTMnqTqMIO+KRQwX+HS6nWcYH06sfGO4MV2p/TbPfh9BNpqP1fch/7DEW5W86bEhvS509EUdL
yQtHfRXpDGXnI8EFnrG6MOgarFBke3Tq6bu0YWDBo1K61xpzk4UMtrn0QtOJW9L8AyKjqjeWuF1r
DX7DVOP7abv+AiSCIDLo/hwFP46jcHFSpNmICgZ9NSgL+Vhuhvg2NRuupMbVzfrkq7QHoOyguoDR
msHP35fZj7gspQHdyaOl6Oul8n9oBQL1ZAVwzLDLIzmDpwKj/3S8J9FP9BhTwHCa1whe9KmKlcXZ
eWMyw34sE9qSlvUVFV/Xr6/iXcwTJTuLd1fXj2EnDJd8mh0ohB4Sd0BqCJ4dga6Ai3ATEiYX5Vv1
2f4cQHe6js9YbATVkuNf90NklFbHoR6VZ2wCuUjZRcXzaiuz7TdKWnNfs4tba4VWNqKgEVQUnal6
U8lqQ0YioQupbri32EjqKSNj4PhjCPInNlCZ19kdbeOV1AnqogWSCkoBfOuC9MMuftJ/rePCO4OW
SPb4aQNaKstwtbaIyBMYXp+ei9/bt2bCyYB+QjkEyqFABh4gHzd9sje0BZZ7fdR6l5Fo3W3lyA0v
FGud4lBAnSfaO0XhxHot+0kgjOjbnd+sh1cOqewPFvTRnKs8J3fVX5/plHm2oflEVmOW0BJ21LZw
1Rb9HbNS42zNvO8k/EA1uDY2InH0TLJPpCCsIbLUzJe9v0e4yjCrRcQoSU9a7gatsv4xHyPnoku4
z1LMmNiQcvXPLdSxrkg+dQ3ogrtzJQGzRHr+ExJF/+FUH1zwtWkql8+fzlJD/+eZCEO0GF/TSxcU
phBxQ780KSxl1xzCd8JHww6QJ2yTv2xtM2NpPzhCWe92mT3WNAE+56z2UUijxz6mm6z/5sHeR1BJ
6Xzt56OBhTDAKaNxijZXrFE4R3UHlipPSZjV9B13OLiFF407KbFDrHz6i1v9IDFW8pq4HZ41TRtO
sBSgfxUpn1xDSJZSQxBhDe7iZJir5F9O4mCaL/jQPK7xqaw3OtsZ5Rz+yIAFeFP+td9CIOhoDxlW
Lhzv8vuzb208JsGlfVhyrDb7ByB8kHmpjuAtPrSmWiAfr4d6Q8WhyeZa03Lf1ELPJG22dlsPD/Ju
o6FTvz0Z769fJCQehCPws5daxBbaUnE6epavL9uLm7h8kQ2XBWYtqWWa/OUa4kSu4XJxFuJIJ3+5
vPe+AC8t+sp5Qg/db0NScdHnPMAufhaN1qQ4rlIv6GEjD2sFuHka84yP++MPYGVgKxnFEsSE12Ct
pAQecidjzW+UZ4I21VS2irhpY6t16QlCeg2B0xGD9QMX0ETEgkIEN+1knHneHSQZ2NqO8BOjCsx9
j/yAhJoZ6gpaI7tREIUMAw9cribC1Z/ghIAox4Ub6wwOQBSB7yvNwztgTecmBpGnA0gZWzLk/riW
PBBaIKN7otcnJNwiFnh0hY/uFlSDErUcdEwLEgmrY6cytsFw1K/3whHInpgS1ke5nC6jnqYoJO0h
/ZkfOrYAyJXREYRPI7v+dn7H2O7LDespIll2/6jihP1/J85bLN6h00PYQp7SKbacCFupLjNjebf7
X++F2/R/pnIwlIraUzqAOzm6NX5XKrsPbCG+coQknTUCWDGLNLa2362neyWbQpGmGoxNWsTQSMTj
efb1O1XC99Tlt61e1HWql4DXdb52E+bbPX1WI4y0uNq5Uy1iy3vlWZGrevrTgTNmsUwjLm+86Dob
+N4XBdaRWmBCBn8jl9Opy5S0e0HjaxTWnTIXffLbsslKIEU8DxZl6NNh92tDXwbHbQJiagLv4r1n
wVXqqFpbBaVxRw+UXWltR1NIW9HPQ3P62Mxwh5h7Rs6dVcP4usGwrWCsIFwUbemA0jveVDbx66u6
LWzWR6UmvhC8MgVZY1MZPZrHNxgsyjZPxrlx7vz0Oz/jsJ2bmsZb0WiqSDCR2C0Ovh9puJZs1K1t
3G8r1Cv10frr52dqV+Uz1DXKFCDRxYNkAzYfrAphKGOen8Y56fp6UWWqDbv+sCtNMTDMp2eQPg1Q
WMBZE1+LWR2YuKHXMVW3nat6HLDcw5axZ7Aj+JkFfMfTbcYDN2y/z+d+6xIW3gA35V3nvncVSJU9
4QU0KoAqnigtNkv9FyDs2S42ElMKV3WRj5xyvn7FOYBKE+9OaLGFdx6Hpss6x8GTn890+6FGw45g
dtMmW4bP/lxr5Q49leOJgog2XEp6+TLaj+Vod6w7KPlN39wBjVmtdDouKuk2Bj+PqFYDDe6whJAg
eFU5xHPNZJLYYmkFGGlVeT4w9+4uiygCy1V3pc67AQXQLDuPeZvvy+n7wUNvsXBAYOqnT9YOtv4O
AFmWY6Lq0xnLcmJNCbG+0XMy/VE11EKc5ZM9qVpCP8iJFgnm578m1HurBT+wG9lgrdDURoaHNe6s
+89rdZiFbdJGjnyJYQLzjn+83UBmnP/LPyc/AnSPWFslFW8UKvSq3u+X1bfTK3R7bUnaZCYTmjwD
/duJctz/1+hl5b2dObnaMEDdip2/KJcjyLAltzkR5bucmNQE932Za+so03LZ9NfsEhSaSi2PIHcD
bHdlfLZZNacgoumN+FxT9bBYrgA3k71miNjKOHI1CJ/OKiZxSxAn40FU4ZRSZDS5w4dJUtAmsPhR
AzNzfQhmrBvg0aGR7ExyzWcOnwUZBw2tDCLxG2p3crsgmklKoWCYWxxWzgAp3jYR5CYtbxCXawL0
SMTpCzwo3/+kmAkr1yRpkOvlqgJkEptH4WC2c5+WJ761OxWWnbOuI2zGgj6OXxZlG9G7nMQSN89n
v8GYttx4N0dd200TWH/UUjGRfpP3xzZQebnSOQEEo1oqHlMC4/Z/BuKobom66LYJ9cDS90BXnpRV
9EOZ5GkuXYGfiirNjU/XGyxWxUXMr0lhJIJOGgnlCcWyV4ksuLmglOXZahLS0WmN235O3/h4PQZH
a5n4svnp9Bx2z7dhHs8f7WU+Zl1/lefhK6Ylmnx/851Sq9mxKoN4VGyWWKiTJm2wv9XxBDSKOYKN
y2M00i9bL+ddC8tOf+xtsJ7YpVChDUr/1pIXmQH/RMcYGkqgwOo5Hcbd2JC2NlauQilCeLek3wmj
cAPPV5S7JOg/WjD+5Gf1La6I48qnToQS6Y6xqC72O2tQRIcvxPt4RlgTviBzvFdW1qd0NdPPe9UV
CDiC3DCBHur4qJxk9RJiikp4h8mMPW7l8ra72xb8THzUwMu7o/fk4Ydax0h39HNLcw43M6ZNyFBN
45L/r++eqqjw3chYnMaR6KqFQs3no0FGR2mEyPCI88+X6T1m6/igJC4LK3/0xyZg8QWC1/Y2srab
f4qyIyFF27r8VKdx/LUh/Vejs6SjtgFxhooTqk4CBJ7mXrxEnQ4NXZ8upDFRgBj60pK/TMth3mZZ
0l+9W1RjY18ckZ6QWytg7UgF9DSS8PApM3mxUOTkwiA4tVnqD0VBvEEWyb2YgGoQGvyYh6ZC+1ak
NG/IrUsCtaf9vYiOrY48bmB2kHpShowGwJDTwZlL/Xtg0qEXI3OZ0Q309rfZMTMYg4ssv4ZivN7A
w96fMZryZHs/XMu2EXjr65lls678kX78nPdi9tN/RaoZALYC7RD4kXy20xkUiaIrJ4wBajW+NzIM
oJvhQjMRPPeAMOBZ0sci9Yc0LGFcB1Hw57YfzkXwWbI/jPvJOPWTrSWHcFvC9FU+UJVOkJME3Oqw
utSh5O9iKjHkWcH1HQJ/GEiDNRHWiWi8ZlylN8pinCJBvg5crM/t6uBft9HNt0ncIxNizd4ZlQeI
ViJSMVNl07XAXmB4TYZKZLHM3d6tFRqD/o4S3j6LTmWoAW4JyR5VGSgrxU4YJtOLSmHlesjc09Ux
W0zC0qADFKZM+mdm6ofkNaDZx1PdZ6Nzjixu+gSz27Xv5rfh9i3JTBM5Cc4DKtFpYAhtEAKpvgo1
pyPN+K1N4utX33I2iRhTKIxgEcBvFJiccskGpW7ypbojrP9/zTS+TifwaRb9clWAZ1Yv+RfDp4VO
EWcYQNGqgMcOPq7d/lBHZAoauxuCNfdwQkM8XiOryIqdk10MHOSVUFDbAjes/DkYMtOKUTokLftt
qsBrcRX+EBSTa4kNe9UMkhyHJQ/Z8EEEMCaIbhsrx8Lsk8sGho1Bl1dTheBPu14AE0nD6kUDejHA
+m+LVi+JYp/BXRmBSv7YQhooGlAYQYEcH+KyAeky96xv/ueR29DoVaVWDV6xqhTc7DBwTYqDlTwT
rwNYboiqpJoTTCecVmDsWp+R0FL6mA0xv0VfGJXlnEB/vwINsxy//eHa1D8VYOH6IDKITQjm1jCx
B6eE3JRE09Txpzd75a7ngO9edsmZgVSIgLDx5/yC0AU3RGRmTQdFxibahXGcULbtjDp3W6IpUpz/
zLXFRpczeyQk2RQH4HaCLOamPSppwiCZGmFCR/2AFZ0VPZlTOIuBv2hi7b9AgXV0fK6Jyy2PxeOM
YLUuOaA0k3GkBfD75dEzC6QHbYignx22ZzblI9CSmlXRWvu0P32mlUN0+zlf+SgwP2kb/oTjaTrC
0nzHhQvL+9drgzGNPIYlJsZA93cLrQ5cSvTV8S34VjH6CEqh4K5yrg5kcz7tsoxEhXewA9YEb2Mn
cWTEnohSqMEL4rwLAw3uHliu1CewkQclIj07yCp1QKaYKbJP9wbDCgfU0Qw7QMAQVxV0sXU2Ivmj
YZBCVa3ivtafWIaORUtMX2sUBkJyiTJiJEpR/onHBXruLF5Nz/BazzwadkKbxaS4Fs1lIyXnpck/
AcFH4j7LBk9I/HmiVBRC2OlX0feDH2eD2j6elvDAjGf69rid6qXag+DYlCxVC1ZVyJT+P3PkWVO7
RWNGxTQJ5spBU96lZUOQPLzSNCec4Rc68eDTjPwWG9TKFPUTsX4byZ29ZdpgYUbK1PiUe/I8KKXN
UBBWeFFOVytDJW1hjlNy9W/U4ca3W43R/sKCAkDdbvvjjybhxCWk5qOorSIozzv3O5BnslT8R25b
kS0uB6MTeJMHu3DbMEydUO/NFwB6qmoGLsfVN8nJDD0pqEmEP/PyEtOchp/qiA8oWYgDSmhdbfpI
jx1IJupVjssORVwT6h50/a8EdobUvTk9ZCX23Nfy03UUfqaO9NR7OuvvgHN5QMYKZBJtYH5/uTcW
DpKK9Ttrc1dVQ1iJUdnlYxZNsuIKuo2WFyxN892usWN7GseL9AssRtKe+dr5GrFcxTG1DUZQ9S4p
ag0nPVV6j0JOX4bn/CBSqgFybJBTTJ4TnXDNl83HHNsne2nYHyiEC31ChwrvoXQhkynHmZ1xGFbQ
e+YVY2tpyVvTMewBP65k/td0OONTIOmj7guSImIGoOndsWq98pEaSlzgJ5iA9QuGrs/1mCdmzCE9
TKqeR7kxllytnGwGBa1n+0KCtmtpUZ8o1DYHxr44oEdOcWhp+0epDWuG1YYlRLnujzIJIlmQNY1L
p5gpub++qQ4NXJRY/Igx8I4x+8mnXfN1J6fQuWsVxfpKGri28iH8ACpP4HE+PHWctdjGgSXIY0Fr
F4MhnzCykHAI8apjFEp8tObIjw8qJaPyyqCR94U7jlgZrJOtOGbJNS3LqvWIGeO9phS7S12gpOqR
C5vdS4Thy31FnSPjf55+oaigFFOEkrq1h1D0DngEKa2KL2rc+i8ZpVtQyI1eDQXHiEBVu747AY0N
QSS5NEorW4zcAYb2uZQTuxgS4ltX8DQAlsf1xBZ9DzCBtkosjOoIIdn7vwFruy4AF1kz15FhPv8y
9BwjIPPYLbMIKIxQCXyf5AjIDJGtyyEUw5lvAWuHyklUWWGzb7yb5ClsjkDx9av6bopyF13Re9XE
5iduD/i/hBC6MvlQ+iI6Javg9LE+9pPSf6yd0wyX8A66fM4QhWrDtAFIr/ZaXQsG1DAXf2VqVOXz
30gm1zXBFhooZYOOTEjjAHf9Mwow2c17q6VeT+0vtnGP0pV2cepTMMhSZ87cfr993Q8v56EqSbfv
3dDnNHUxHJq1F3Ui4d9PCMF9IErf1En2Gi0IlaTqCyVZwYPwMNVlHEYJGn6oNsF886c1/fwexo9g
9C3T9QlhTUsJbL/mNHiEsgNNewuldnpvRB5s+wA3XxYhyRyzmRUNUjf0Hsl+JphHa10aWvqaZZra
baidSEAx5cs/Jc6DUfyXeg1XjuQgjzbPTDOgOyS70YP1LL/N1awGRvtK73eKEUOw6rL+G2yizQUp
FtxaORjEzxyZLedf0ysYA3Za67EufrZHNrLRkp5RzVI/zFf+ifiBV15V4XJwv9ygou4IP4bVG/Zw
e1pj0FCUsHHdEGzu/hBX96K11GJA9HBam4Xk833O6ExuUAulSktTF2+qBXymJ7SqcEuduv0LEFzA
iB2bZQMQ+PYwC2fR0UlEN5h6j5iPvjGpE0GSRqK3VOgZTRHIdgpJY6bBV3ByEsE5mFQ7XqoXlRQE
9t7wNfuNnySDmdWPq7sLcjKSHZf3CAih+Aod5PDZwqzTuw4vBXQlBSr/rQnksX0aHX/wQHbyJJDb
5ZVOL9vL0PiYk5+qKPAxkoRHA8hAB79BjIxA690W/nRzAG/XZy1gp+5K9HqhcdVsOXpBKxTUq0kI
po1Dnp138jyXElFcZIiOCa0gh6gL/oQoS9OJfR4C+nHa3x2qei1aM5B47yfMiCjfrRzfwxIEQWT/
t0wmB14Ico1rsluOHC70YInKnz/COf3ie5HT35JDF7hLDRIhgE/e+mIYW3UjAEN+uthUTtwNKIKb
V8rsZ0DnvA1D1iL9xlOBLl57qUCgI0eK3hUOXY5vRNs4eNgv8+JHfyR9vAFh5RFPoK/x7UWgsQyc
LsEgxda7bhmXiOQyiip/3piV03nSEDXqZeR4j7X7yzYVJm32pHqN6M8eXJKVE0gcB/wfHp4kPHaR
httKhkxy3d+QjLDm2c1lqnru7HIdowSFH/DvXmubtYhz+4Z7CNx+rVVibTnBl9R30c6hjwT1SAQm
LR0Tc8Q+wSoI3cPDwdNimz2rjoJgHff7JtOXad4tE0ezZ8p/s3JLYlgKm+flDJfc7ZFYmF8Wajb9
blRC5LhkMMxSGzYZ/1PcP9mJR6N+/2U7Qq7AUKNiSLgVgjkiNruR14qCnF6pFA5pglz/TN1DS93I
YK2umcPww1xpHKVAdIKLl9KCqqOdMyqbB9utXZ/3J3FfHBcb2g/zn2gF1g/bcdMXbtpI3VI4tGha
l2iHfflV73r5uvh+QSD1750C+JUsEKO1RfMmXrPuKuZPZoauvnHDUuOYC/NPYPbO+p9FY2UvIUme
UAJo/H0vKuMh1xI6+XObid+3cm0At6BqWyS3ddhRSEEgEQnN/0V7Om4G1Nm4FLDFrCCdzcfe/Qb2
YGPAQEHeGJ+vo4ByuxEFSlVB82f+C8GSORmE5IklXqxUAjjnvXE1MtbHRRTbePMBOe72ZBymhfjd
Z9UA968wN4GNNG/uUDOUVa/wfYCT2F6D2WSARaGguwbOl9U6gTq7CbXX8sfNBTizzBodTSc8ekTn
AqWilxrxLmbM5tdUkw/cKZrNoiUyXHSMpHuFBpjWeHQrgj5xK5ugoa+98AMKUY0phar7oMVh+4SV
6SPZbh315KUqvXI5lndcBTHQCpx6KMHzvPuDZBdTylXepB3wDLt5n2RZvE80SEceNJVXqb6pn8D7
mwsRbWHwde6SqvorokkXrOIoYqz6HpPGCUebznouTAX5VAqV2pQOZavqt6KCcZe+8yYF+JOHZ5s4
gCT5f1izgcEG1ZCtDAhBqE6uxaNX4kI1EQPz3+dA3NDr96K3JfePEV9YJKniK8VBeIElIQSai6Bd
GzUf+m2aIl0xqYUK3jsuQSLWRgmgsN1eqWHM/sREjTazgMzN7v4j9pqMsoAuDbFtzCKLJMk9YAS3
Zuq0t64h795bi6sBXcc1j2q3hVYxzTzayk70VQTjJvoW6flFEz3Yp/2MG1lS9ic9mAiCYCc7RtQ9
1yauBqMYazh5D3w089H+bzgo5kFIJxnte3w9yUe2PH3DL2Qc1rZJRrk8t440+cgZSgEPV2gc9Z6S
XIV9yOg7bRhy9Z3mkf0jx9Lfmsg/g+v4XXpyGWOKTWx0/JeubBQeg+kTcbvRiZxDIfToewa0QE77
3HqfNSmXsM1oMwXPyHdyyLcNMAA10OXcRxAo3Uv4Baghk8Ki72L0aBlxyW2m9xJVQEuLICoUMNy0
uIS3uCFvXCtmL2nVKOMjM59pNUh3ppXFUQ7LU4soinZXCUnoglS0m8m2Sa4eZ3GOhAj7Xp+UGp8b
VFOg3n5JwMm7xgOdk3rtfEB/X+K5TTl1FP/am5jWOe6lMn+x8bsrTCAnKJAme+lpioufOGydH2RE
XON2BPQ2eUqnQY8NQcCjDhVm3WCtGWM3p+atEFIM7aL/8mRbVe7+UYyyxdyq1HeaUujcz7C8BBTj
py6w+og3XJS4zeTQa03bXbuzf+afQaa70w2La5krIuEQTwbPuKgAR3bvzFXVRPja1c3T028oTspX
wEVoQVYrsDuWQ9ajX21H5SUF8GauPNjPrBmWggVFZF1aBIt7wJkO6KvL3MialTWfaEC1BaCQP+4v
jI/cmVs2UBUyhDlbxeftj7slbmJH9wviOwPvMXF82t98X0QJH5Rb2Z2ru/52qDnl907zyqHgNviY
eJWtMBqCSVXWonBf+Cuc5m1f09C5E/dzGPVIRBjopfBv7laznSsi1lmn0nYay4jctGrHSOWnPf6V
ua7Didi8MlENCPkJQ7dBjetJEBraiOSjOT9Htft7vJqUIlF1S/Z/36SyU1z2x6tsQk6SVs87cqV3
Nc40VX8mosI/FhsErybP4BEHrvw2QkyfXUpn1y35Yr9Zxv0G2pf6RS0zexoX5tl732ta20Ht3a7U
SIBeJbgMRtsedk2bgsLznniwa83/eEOXDHJDL4yzUjcB/Olc7bigIbHgETfXwZThurQ6kZHkyq27
Iopb0K2HjX1ZreyJrx6z4rI7951srNmdOHkxaYxOHyVFKvaySY15NUc1WaZM39nBeaL7dWCDPCSB
VYYRnEyzDwTAadpIJFIANS3HjEugDStBumyjUNjXB1hxvz+tvzZbVyWBOSjFUgxzQFinfA0SWA9q
NPmgc8m+Gd5/Xp4xi7PdCk9E2PURHVZkba8qo5L2JdQVZnnpthqlwVFRHhOfCg01zx7wuuiV/+Qe
yzCaS76GqC62RRKC9923xldeHY4Sgx/DngI7cC+pFWcjm3YCr71O6mFdHDob68bMr77uhjR11mIf
cpaqpKU1gHQ8uvykpa/bT0Yl3UgNYoPEYN7SbQGIySgdDMDabGD/qTFBYv3fu+agYduNvGoimRET
zatmRSxVnEhz/ResM4+0QqXoD9we/9r+kjG7xaq0tnUgQv+INsF0s5cwvWXNK4kXnDHMtFlXjCBE
yUxRoWy5kfoOdBe7ZsL2lx46ORPiF34z5VMbPjEZYwgwnmyCDoQWpPxqQ0b57vwmZzjTMSACOY+q
lu1tyyvkRQmKLDe9aKlqDlcpnhvMg07ofTjJsMR3xqUn/8KRQ6e7B0Gx6TrWy5KGo7s26gZuEVII
YyhShjhvrezMjWbGsug3WOQiGEMk6ZSWfh38AzhhaDL0qkcUiLD5ksSdaGnvpcUnZ0JycL+uZ7XA
0YAHysllQb2vMz1nAOX2yG7toz2Og6gF7wmAA9tN4G2/t1cWisyMwq4FC9o/seogXqPqbFA2PRMc
R+JVdomdAteK0N81usxp3GL8bntZVPUyP7zD/szu2BNT3hlQ5R+IiYw79pjujgWLVGLw5GsIgjJZ
kJxjxpMtJY9TewqtC2V7BUpn9BpXhCY9O006oXmoXboYwX73nHdDnXoIESmI5N3GPXpbYQ6m3Vpe
6L5glFnCEZ5aLnMi4tjvsC7B7LxotaSfcZLdNRtdM+6OCnsAGcwIUwn1sFU+4Yp12UyotYqUgb6A
+YPsS36+DqRQ6oosHXPAFUacjqAFW4uZSxMnfH6VZSrEa8H0uhvEwRJsY0Sc+lyQLid+cWVnwR+W
37KHc7d476tgQj0YccVBEvmWKjo1BdlpWwtp38/EV0YdoW8LHsdwWpdvUdWGrn3dMWrDyOwxJKPL
8IXaZ+hqbXaPQlgrbH0N5JPZayeXs0eHdHjmp9EVI53bKrc0RnLnzuPGZHkq5BGqC0AR4jwD2p/r
QUpwYeldk9sDAa6klzKNVlocAJfcpGuURhgkOjjm65v/0gxViokVqFyF1pqOJv7kk1RRDttkTrKf
eG3YDOKArOHpM+W74jSgQsEI1YxNrcosrQKyHfYXmka1U687Gr6d9kc0KZiSxGhhWasO5gJlHv5z
zGrfX0rvBlV3GAWOrRfvZYHzEHjJR5I4cV9nwoCtSKmFxPKvR6QAXKr0nOYEv5t9EyEWHiD09t+p
c/0MQ+sImjijpiYKns8cnDJ1EBTS8TxPMTfH5fn+t/LZ/+eZvanU8M0fE+719vi7RkhFBcFp3wr6
wjyaA1iLtRPnlri4nyUvB/eGcwFBAaU16NMCShVVojyC7/jj8vCD+1A9JfwLa3yrgDJT6m+B8Zmr
hQGkEok/PUz9NQNik6EE+N2oR/vIa0ZZdpd4I+9ymAK3HgcMr+TmVx+j0nboSgIVHevvrZGYPRvy
tWbY0CmV/TVjXT9dVub8pSDD9nudkzl+yj+L+Wr3C9JEtKRth4ePL6L8i87Z4Z8/rUeyk9noNY1T
/sCGuXyEpgGmR8zccbjBXpI5nmR1VJzgWBrcqI1Av7VwYxGZQXXH0bXZTmeiT+VUbOyvXGhmlfHa
tnj6O15tEJf8uNqmXrUyCzZGoA81ah8bs7FVclP/Q4Yc311hX212HuSP5k5ViwczaqA5vfSOSz/m
pLXZ0i6KM5VCNFoaVsYC6DOe3O5T410RF4RBN4MvuSGoOIIjyy4TuIYp9Ri1h1zyrvvAkLI/LjUN
rmfownK6ZYwkaqTXZsrjWKiBLsfQqBCXdp+fIbR+0ZZjTu8m7DqqH44xfbE4MqwuUoA0usVrnbmQ
jimC45jIIociabt9fwJqNY4gPukKUVrY2TjPEYu06kBXSMwa3KTaRLIgHiEAdMVyedz0lF26f9nX
37p1recaIlH7vIghnc4LfrIdqrTfYi5SSb1UMJJldvtPKagkXfLMHREDUb/xAA+BIdcDcN2whNKF
c6np2FcGvgLAss8BsZA54b2NazZ+j2tVdu+EEH6Y+6ox0BiCGrkYN1bIbhovOpxMO0BNsyrob4Ne
P21Y84G+GXRMHEGGfEhngQ/SHyDqo+UtmwWi5LniDtnDhbcD0ELg3PHLh6aPqroZDJpcxOaHLckd
GiRNkmPA0cjz0Wy7OiosKhw5qIqXL2yuScaTm6puoqBkxHsw++1IF8Z8WsD1aWCg40FnjxJNZIef
3tyLq3RG+P9etEQ2G2XYSRU2QVmPLeuDTGkvzDvA6BVtHaKtT6o8PL9PD54v2BSp4sSMltbpB3Z0
D8UMU3EulhjzzRQDvQHxRK5lGTCmqQ42eeYfD/63VEz5294tzNLC7nwf/HbBKABQbqQeEh7qpoWK
ekLyV8zhrNJw4NdPqVIMHT/BXTuvCTGoPgMNuAIKFo8DqkmT8D4ZeOnHAyCfBMttW9NOnhkmdHt9
EfNVUqrQCKPzjJYWQJ2U86MgQkh4F2rwVlWq51ZcwdACcqek+pjdHQJGsQR/jDjFIaVjR/u8QbIM
gRnf59B4/93H5AwleWAzDiI+YSCpoauSHUmwfrn0nOwHot3lxv2NXhz4rHSazED9l5TVUYuKyMCd
TxbhTdcDYHe3geIEfk/X+sfQbMFy9LiKNa/gZL2AYLAh28wRxBKV67cISCpL3//0e3sqiIYvfi9q
fFaX2tnxwgwNwoKXIUFyvPWiqssejfRIlGWdA+JGycpp6QLkpFS8m9vW7P2JbBCdA++zEs7UdW3J
C8C6rpkd3+gKoF9eOfQQrehsZcz8fTU/0GN3LYtvt6J2IpgvjoMNzNGqNn2+/S6cuVLNM6IZnWec
P2uyxuW/ERUCET5LOshjJ1Ekh1TnYWYQnvRDXEOf3gpXP2WSGWHNELZ63vt88D8ICGYuyQOt008q
fsbFuW0ZchzQerCjsB7etSb28MTXDPPA/qwnN92qo89/lmaPJU06f+pLi+ulVI4kwBij6Oc0G9fv
nN9j97dZYF3NBF8K7gichhPzics99SwdwJA9Erw0u2erwk4LcS4O5j/IiU1YqWZJBllI8oXWpF+s
NgmwjS+k9iA0QhkkjUWOx+o1CoMCNiX0+F93jmvq+/uDlpJujEy2AHHFiOzRo3HO/BI8otpEE0N0
cv8xmS5P0Q0WXUwd7tjgb5NCVZcWDAV2wZeKH+X7YG+e+lm7DEFUcE4ZsUFbLBzfl45+uyg8Kw62
cA+n+AXjrjtzObl4GIXSH9Z9BNb/Rp+5Jb4sK07Bk69VbtEiPTxpPTFw0xEwFs/ZYpSgfRb9cp2p
eG4B/yJHfT/Yf09bFdN8uXeNeZUCbTaXHmK8Xkc0K9fGPb2OsjTJKSZkMSwa+/jrJmhZIpp3/XzB
PeAWlB6J1W22HNdg2VfQQEU08R9kz5/nfANoSjENU3FvMU2plCNpgogrJ5u9h4bB3GZKF+dPWNWy
X9LlVOhpjMJyRSm19XNy1VROHwYeQbSc8d96++coHo3sqtFxwk1u5Ect6i7OgmxJFyRpwfd545d9
WGtxAxz6KSSDJKLXiYoZ1qapRkbYVH/5OSpg+alpiy7IyTU85MTUiApZe7r79uIs0HFAPxyrrjK7
FsCCbjh/qyLcnk356hQKcxk9m77MZGOQbk4sDwrDYJkTC+0PJqhnAZxohX59WYjW3r2Lg7rDglMv
iy+xW8WYm2dGxfbyXz0J+B8/UcpTvfs92UYrBBLMTzlHPaiuuiIYQPC4pvr28gvQTLhtSLG38Fmp
urIwifNVq4B8zcJzXvrXfHNqSQWGG/SWonOqmPyXy97RrbK/YoOOfInPgGyBWwxiBUW9TTL/eD73
FMM5921Yq25U++9w4Ixc6l1Ab63fmdBF2Xgt6EPMp68+Axj9xBU8V74r/g8m0QMiD1bqsiUMPL81
J4XoApJexjc6xiBN1whAiU6qzAcerpS7b+5umS8VKLDCwYL3q1KcHtc8MxQS0pt8yWauYkVxUWOI
Uit1+Cu6YAIuxEPy6SOZEnYgLBYYryQaFFz8cQuuKZtsKcxT32WESrnjJZDLQCT0f5yqi7CpuUcb
u+CeyYRya0woS//x3bcTWBkc93gfnvCpL5utrIFi7rx9YO9N+AYhyZ7e9U1yBSn8qIpsBjGir16Q
0dy2JyBFaIAoJaqrnSP5pXvB1z0wl/DhwZ96n4Av7uCt3V2BdDa16f/jD6VwAhIChAT+m/vqfGId
hLRmy1OBbCuSvWaRHc/bB14vb1qt2+BoHiVN5rBcARLUd1Wenu8J+iGQ8uSyX+nGSVlz7GnkB6dP
Ra6UHS5EE6dyIAK6EG3SlDgeCvlQE54Uit1dTsiJ7KRjUToHch3I35Uc5O8vQeapEQcUb3fmNEUn
nMl9V8sHPe8Xy32Y9fOUiuYmpPBqv8/US1Ua1eoPG5mbs5kLj8k+aeTTLV57zZGNmfy71FTo0f8A
+9OKPhieFzD9hexOQLvXbp/OlLrZDJBgDZ/0LceDcs1Zf5c3PJb95p8tVgY7XNAQsfPgUMeEepCX
l9FH43iZ4uFesexJeIcA2P+75TSLfCA6HvEpfZuCMl8n/q1tCVjWmcnzkhz9RXqMFJbJXdipyqAb
yim1+5BWo1A4lXLNEr98lp0OMkz+FiZGqLFVNj60U5rwpGLZxezXZunjCX5WU1u5nJT2H5IBQwgB
rDNDxUDOoM1mCYfIeemba8+zY1+7s2gc81JJBGkn3KdBadU6+aLL832C/xhLM13VXUXF138cIzxN
WtM8T9ksWZxbioLHjgNnYtDx/zERALzj2xofyx9AkR+XDiHu1pZnnie88JxSquWjZm0C7s89gypn
M/XdvHRX+nZhjR/q7ncOJ1vQTsJwZKTPc0/wnw4mAtAkUMwtCw0asrawmeEn0v2RK/KpuP02vNpr
At51IsSsOYdDiE7g31FTCdhDY05uUM3EhE3xrMK3oit4P6Am1sfHX9DiVIJnBbZcXB7o9qmHNYkF
E9vPIHPputSGQVxmyVBvGjDqUrBvh0W/rxH57NP3fiNsRPWRAyUNHdOE6xNtOyRewbdAkN0CZ53D
cpAeJM7NJt/cmJXl5vvocTZkR1vYp/EuyE0v6p9VwQ6/cXgh13ia+D3YhwThwveqa05nAUlYXpR7
8v/AWpc0SJn+5nx0CLyoqQry4GHzNp8S2bbffsAdZn/f6SPgYOZSWRk4gZ2UnTw1gIb0xRCmndkx
QdI9I0iDOLwMMg3bC5SJ687FLAMz6IRdObHLsFA/e3hFCi42vgU42bdPxj75iWejmp4GSdt+NeyB
1gkvcPgTSc3/K3So3dFKhJAA7WOHTzigRxdKMgcs//kms2whplc5PJr18rQ94MRBnTxzaYyDadFL
2OCZT4WvYiUgTe2T10Dvxc1jCbjr4qXjDdjtv/T6xuj4ATUkIlueBT9PFeZccNr7lTF1yyjssQ8e
7Odh6nMYNDI2o/jOiOCF8EzL6sBzFL5UAXR/BN6h6kUApxfvHgZvLI1SbZJHBK0bjSnmoKeNhc8K
iq6mzQi/5wsPLwGie10nWXt87S24j7UBsSf95mQ5cn3AtEMzOwJ7cuVwQAvDWqFaBXNFDjP9DOSL
BhsvLS6tuaZ//GT1ZW0OgKPBylDasUIPjDLs/b1tstVxkN7P4zwDxt9zUm7nuqO/xZzRY66/cnE7
F6435+Fwox9yrfU4IccLnXw1JwICMuEqapDx0LmetThD808piay4oeBm/FlQYBaGlgWLCELKMYmk
Os1k537Mqar8LkntaVpZj3fQQuNNorW9sk7S/IUfIW4o2xG6OaI/dxjeSVKh3EACNbwhthpCwnjB
UOiYv7hbErKwEsy9iYQOfvYxGDr+g9XXYHol+i/h1ukLu6kIITAZxjxPqEm/T+J+i0FCPon/TjRk
3TNZW5m0dyhFyMPPXH+JNcboBMBxO0eiPXvk9qGga2QS7Mna14h4PWgCuCP4Td6IMOsxXQlSxDtc
ShmbmtdW+d486jVUScFDsTwBI6iMWVn+ew6NM5f3LYvYWo44/RqyuBfoUeqIpQKOOmJU2TZMQSqq
0x0qNv8Pi3BDSmQtAvZkqlA/42xFee671YgHH6hmqZ6564G190NzyR+45TIQPy+7kJgDLMiXPq+i
XP9+OjlVp598vXPxS5OU3suZuiLou5pqSSXFT7ogz++HNHeVIHxtU1ToItof1F5AiP7//DBQt3Qg
X5oyolhDcgjAHKhPxOiTB7OglybB3Sri2T9b4anzsnDuYJipPv8jpouJqnoYbJnB+nrxAnR7kYs/
lZdDcqKzn3h6c5DsAgIEtUWfCqVCZBwk+cG7K+2q/+t+dUPB61nSFPCJzVnNgO0n4hwdykun8BRY
3V9mMxZ+3UPc4TQfsBXYbqytWGfyVAhuymwQaXBDMOrstbn7HWGdymvX1ULB55ERTnyp4/D4dUQp
ZAKmACOI+GIF6vmb7RG+CraPh8QDmt6jVIAAlzPBYEvFt04pnWhkxa1oHNJeec1EnyejcvrXWA9M
f+RZy1EUwxe/QtzKFk7BIVPCXDu+ebUVLlrnRgLnZq9b7bsUtKKwKopTizd6v4jFgK4IMiJMPKbT
c3iYp+YTWk31/pFmVsJ+eIHz/tXFwfffc+SphRSglUsAVrJBgpqUz7UPY6ltgpkAzi5rdmlGH7VH
BFi9iO2h96qwM9M+dvjTNE4V+wv4P/t9/DIT/fMOFdjmKX+7EZOl2AmeC8pixjEmraiO4EB69SxE
P2l6Vd+XVppkxVuwyezK64QqyYPrNCMyC/DBc0ryZrw3T0QBlyd6bsg3wWAZt3JmxsOgyDjTrS6G
g+rBTA92w72V9+Ho6oTkhhumf/XDTSz85HHuBY+K6zBlkDRgR5APFrdB3qZRafkg/emp9O98ev/b
J+Ag4EXszBULXJH5ObcSCO9t28Ip2g3ozWsA6okyQXd8W64ZQvHwelnwOaf/SHOutU0fDUNK5y8v
Z/7TLMiPo2NBeyRKgUx6gfsetd6BKle+HJt9YE7zyjMUryzQIVid4IP4Kgz9Z2yWgBKgoIn/TQBl
yU0oPn+L+yFnuSiK1w33L4N37KeHYaWiKYhzyrVotEoLNKGGsSQP/xYbzmiBvnfKSH2lbsigqTYX
BkGBFUxPdMA1+eGY+dTGWN07hoT3VqAwz5O4dUyEZ6MaoPn5pZyBBzOMjIN5ulZP8S3modaPhJQF
0k2G7ShU4FivupmQojCm4TDsxq4XsNXQUoH2FjdPlFC5DS4Wwlr/RHT6F+YuFNE6ESxUj43QPzu+
9cHVqwu3oAOiQ+1aZ5421Z8cNu/WWblsoJPignnVWIEMIEYSZsQXvG0PaNUMTQlT7E9HbBQfEd53
Qsnb+Xy77vRlSILrw554c4F3rHLYa6Eqd6sMOrXP5lUZRuGp64o4x75gH+eA/zm2zDH9nHKugUw8
/xflWmW5UFBdp/1QqDlAQTcOtOIntawJSODsNFNfAvPp+aTGbDQyfi7b5ukDGCLQCCACb+b6VHWB
SQMtkVK/t7HOZopX9B5fOCg4L0AXzBfkbwloTvgzVxjrAYNf1J85S9XXZGat/srkQSUUSoPdOv/s
fNRa3LSwFzWHQDgAFjS/yBFq04UHxUwdfsoWdutqycDUWRUHYqOe4J04ZJ8AwWlI1y46pwYREyVI
DxS7V5lQsr+U6WcLAWw3GEyOUd4GPMvOPIyTmSHhEJgPHefCeJkuBKLftZb9xbuNTbRHNRA+s7Tb
0aV/c/XyJxcNmY0gbPgMjKbTHm6HF3RR+bPV+Pvwabvq/5DvSYuqUvDWppiWSDr4459TsFmOYsze
MX6PKAthHdK+t9RXIwZP0ERFGrfqR1VHGU+XiVvGp4eDlWgPVE5PTf2UljAzCF7WmQ9iF7q2v8Gr
+MLmd9AORSq3YjeNi0Sd/QI5Ico/XoFN2/hNz5c0MfULC2JfdYN8p6XBjfcuuTT4KTRcJcSdPh8b
WUAC/bpPjI+lMKHF7Eeuf9I/0dTAPOoLiRpjmuIpEU6EpXbMQW1GKQuC3VxvJFpnpBRg+tFgzaOG
qBG1RArogrqEUAn1yPCU7UQ8A+nRJpk+0b1b3FpsrsO5qY2dXCSzR8vs61ID4hiG1FmOY+uHqf2b
LPFjpLNtjCmZPxId1FXYQFJaT5nDTDJwHPkzoeioBUV/+vZpg4uLQvssXa+YsJVrmsxKGW5YBSwu
pfDevDmmlCN4Z5Kt18irj98E8bh8uurQCLKKGjwiQcRqBXy76wh6NcWdS4lJ9cGKSV4j/hoWGRTd
quCcsSV2O/U8Tsc6eQ+QIqnKvVYayOs9L3NzcliJinYaQV4R04ITFlZcFFZr7xpoiMX8SxS0obiu
Cdkt2u6jZHoanl3nf5jkZYutIACS39Gqfs309pO1ZKwL5U3FTIv/qhVX6yV3VZRoCkh7yipe3PcJ
+3yoSvdZHN14G6uqZ9P0xPHnPmrf+SnEhJx1ri+9sMWC2E2gYAKJt4oqd4OEuJcy+9w6WY874eLT
g8INFWbXfVLJRDyegJy7mSG/UNQhucuPVFtSHqJRTX8bETLRGlUf4WNJee5WUo1jRxxTkAuVOW3+
qBHq2oPBStHsvyz4aBKwAWeNHn5WGgCLyU5F3I8b5efp5ySzULbLRlehIfE2YL+xPG/QqqCyWgPw
acBVtO9ANEOb+lAzgUNLBKG3kC9ori0xd5JJFJuZD+tUul2V7oaiRiH57Qn+wrVaTfRyrM1DJHIQ
LqSCyL6N7oIyfHMDdZV80zmtSb1BmhWvll+UhAOFwZ9deOIq+yV0LePi9MsFiWtbt7/zpz4WDx+c
tgcC6zRVNnAL5N3bEXAWH9+XIavi2L41q/8DbMxGKNud9My3ykW8jyp2Rsimrj/qzB+bmGTRUpd7
bY1FK2Z/6icuBwCSu+13vJ7h0Ag6V2WSTCcP6w72xSTtxKpkqur24eiWwJNLIYEwfZ7bzx+wIt8C
8/G8Fb0QAh0Z55O+7uRHm9aI1nH6PnPQFVVNPE6+CuWoy+bI7w44T9dBiza2folIIX6a/UWOgPyv
GZpWklsI4Q7ZQakMyEU+llqaG2/u8R9uK6WpMhklgfnKAU7XXlMXHBGj+KOf+j0kuJ4BvxG1Wm4u
O3dRFISDznu87yZ3byaUn55WKz4S5YSIzczlHqvU0rT5La+TwO2nIR1mTARJO8ZhFDUq9Jziz1Kq
5ZgpbgT00O1WmHmkz0bkw7P3LtfOo16ybThWY89rsTZbCwd9beLO/ha5Y0dNlZMT01tTZ46bpuzP
7pZ3HcW9PoMyhN6laon6YnV2mBmShXWNlITMqlm+PoU3rEapUkLo62ducFdu+YHbLy4Yu9jZrvhb
KW9Knbgu4UT/1QRLWJqPPE5b/tZGHLLHZAfvYAgRsGem00R8IYNy8y8bCXyfrWLc3Dx0peb1RXt+
74Dz+h+xo8XMQz9MBRa3kIWS41slekfjnDMbUUod0ZHRjFiwrOvesHr8nEUNLrttt/s85tOqs7u+
OZ3WiOHf661DR8BcIb4X5Bt/CiawPDWWcU7X97t3L0wcJd2M/GbQodte8B7P9b7g9VbT+GA7TbPS
YeCQssj1/EPAKhlJHwuKRNB2BYFbEKIMIedUXyey9YJ/Gb5QM8LjwXak0T4hEkMKwUyaGKswiueq
L2ST41SxTJVk0nPGaQaUbxjadiRhuFmOFUtB0HrHcjxlUaIYPbig8ypvTWpMSiOpFywCBM3DdJLG
orjYasURmhMNpcgalGK12XWNIgCet0FIOOp2g5qPbeKX51LLDhxYXShyTbzzHjj4LM4p0pcsJcyB
BmEBY1FHscJEAdtjAtuCE8gvuljqFf/WfvoTWMJ69xSxYSeyZfRlMmyKDv3YsvWF4XoZebZuap0a
tYPHca4TrZ/HT2NpNdPtcWdn6MxOvL1YnEARbeBV1IpuIWyAiY0+BE1P75CT8SZ5HawSx+/2HDaI
cSJgqiBVc++dRpXR/8u8vBT6rUGOvq+9SnrdGBGHmRCT+HwNWvLLPXVcBMqR772NZ6xNrwt5aOX3
+rbUmvoS9kUUztOxG4Cns6MwXxMtevV0oqVjLgqPhJO84XG9CIcE/XfRihMDxARQj9hFaBgteTmN
LLWXz1KxRxHohpajOxw4Fp40bLbDn5ofm+qUMfzxMjpD0EhIBNb5k4QVaVjZNNMkA+ovwNK4J6Ad
XR7jGwfCMi2NjATPqtGkYiZ2BIb6H5gcdJI7iFCN+kIdGUXP5BCtNOhIB8j2eue+hxanpmLAKZ6M
cq6CM3XnkF24XfzIpkEnGB9MGjm2bSH1Ny9JP7xsYPrWrWxsj2PxT+Bm6cPa0eu0+XxARhYyD6R7
a3GAXfQsWvdwM5kwfmrVshnM55ho/dcwZemrcgThl7M4Jf6o2Tdpi+DNoHpINFoc8RJJg1vM65Sp
nYYyd+z7GE7Bk3scr8RtrprrbZElG+Yc6JfiPD8ze4SlzTnuxA+JK44JIXXSIntOY/vFfMbKAHZr
bLPOMPYagtvihtttaNasIXKpGfuicS/X4vZAMwOwDRpr7uR+VMoiLR4bQMPsTXZdtgjGUexwl6pC
lGqLejCNkrBFGreuoyVV524CUa2mSnPBjceI4Pc0AXTBqi0yWaPSMBFr3+uD94m8LXhia41rqqI8
T7KD17mGz2QkdF/DjZUXCRDGoKjlCemiV4ROmlNn7BvBx8S/qkXId4LiJePKbUo1DJAW/VS349fK
aMuqS8Uu/9bjd3pKQRdb8dYCPCOHFiNgvaQKUDpf8vJMF1ZTGu2cbNyywhng3VOUDIowfw3slOLn
UzwgXT6rTGQy8+YXotidNI/XE769fWfPtTg9Fz+hY6nB/kgG6Rg/O0/uvtfjHSI3sjVzVPVMgKtL
bQnRU7xMx0TIBH1T7gErg/77AJ64nxqDsrKa4DecfGy2fZbX+3xRC3/O5Xj4r0QoXr4gR9atnhCn
u5i+EcPcAwaeLvxemwZNXOlKKMVwR5q/Mh6EAJTJvvNyeGKjabEnO+0jcM+iHLKJ1gQsgC44e7We
WbKOqlJRo29CzBqqml90zDlkXCfPLE+dkRK+Ir6w6Pkxebr+d4jmvLB4V3ztNae02SJI6ALwqZtN
W28uT1xlZWfE20n3DvwA3S+TV1L3cJTUoff0c6m4zHYXiphZTin6nUpH/KIgv/cC00pnRLVbBtpj
DG6TBnoMl/oXr4mCoaWi2kT3RWO2JBanVyNwOnYrv2YMkcxkepG5z+iQqQ0FTxMr/OfNZM4Ffeu2
KzVJUxGazLeAvVNmE92mQKHEeUJLh9Q/TEUSVmqALaKZBeainANUIedh83dpyH5sWtur/p/VFlSP
bRXqrarTfZlZLLdfH7YtBG8ilMm/TPe9oWcTuaOgdw==
`protect end_protected
