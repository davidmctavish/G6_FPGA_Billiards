`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iu3+/C9XFn2DzcgNebxbu1rMESdiphYvYrViUXuKf99RbureDRcnEvXlp/c0w61/why9HzjvDtj9
i+J+I2bWfA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iZJ6PcS/rbEHLoVa7dfypE92VEH4VT0HpU1pGzdMR2COPCnTEdPYxisLrH1Im3lMaF7fk5ZyosHD
jfOfNndXaHQCKrdVlDk5fiLF1BW3qw2qehoNKuD56U4BEA5IQWFoDrpyXislex/cukh71E/1uelC
Krm8cVaK7cdI1/o06ok=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ajt9nMj72Oun9RAn43YtatA8v59S5pMe94jQyebAFq8UVar+hrHcUmn2xBgjxNVJBSG5QQ6pFv6+
z4rYFA2u3Nq3F4LkJtShYtOyXbfZ92+rWupTLXiGl6xvHae/4hhSl0EPp8Nf1SWl7GPKM16POrCD
+wkqOAr1HXgwv5hVOv+ArhnvnOc1EgUm3WSv42XXbIRZU031B706dcgfyrO5ImThC4r691/FSD4w
oSvuMuLBc/MsDAVvo88/+vderX3tybwHMvlcXc+osfUvRoTH6HWfYSOvAZeRsiQKBWLlrx2kFcjR
vPakWCpU2J5mwQvIJgiwdoA/giBDYH4S26SNAg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Iecvoah9HxZqCYIm+DPWv6gJYLYdGKAIbpKC6+g1+tQAzZui8+AaMLuxr6Arq+NOnuslirKLdc6L
3z9AfnHPKdlOwHLUs8XkG2bpQLJKCf2qaqItJDTgRf/xLOcFAh7K0laURp88bcNMxVdfUj5k22Sl
xVctAods0oeO1RAR164=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NAz7Saohu/eLeL533aMzaMhAMAq7PDCeAJg5gpxHQyFAUgdH3uJnV0NH/md697hPG1Qg5ndYeHey
Mu5GaWxek6F5Cw1ZX6wD+AQco5LqCqAqjP9cnFEiSaoLmIZlOM+J/KiTCb7duwrdIar/0yKiTBUF
py3fX0T2JE0qsJxnaGpgXMYqI6goxaDdb2uGkwPS7gXF2jtcfWdQzqfAJck9+Fq76QJg7o7Ugg8t
2xFlrxgyn2ftFbVgR5UVJRbM/E7FNV+Uuilaf0U2ef5qdpW4bOCt+Mu23fPxtAA6bM3PyBf47yYF
7xHBsH36ACBYTkDQh6U8g6e4bgcDdVB9NLQpFQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11552)
`protect data_block
DLgpWg2hjJ02rUrNzO6olEJ/xSD80ixrx6SArUU+ku3jLi8K0MTTdmLqVWstTZeXGqTIP6QgWrVw
ncKdqOr0j/zD+vNltPGbVmi3BgqOgCox+UbBdN62rJ22shD1rQZvX/js9h5JxBNaXnJYoJ9BBVpV
kgjuIHe4V2yuvZOnaoTTNOcyjEuUbpee1xmS3pLuBg9CubpQXP00Jzju3Az5U0iYW3xiRCAJf6yc
/wLi0i+XSHR8vCoV24yN04JRIBlZ60+YjsA/1bO1JS9ggPrFKnilFIoCKPpf405XDBdHnfb+847x
XZlFI1Z4jzjwV+AOjaEEHDtI16jMmQZgDWIPMo/XxHjXkcPVDm8hCm3UjamUrsTmzYquAT9qxeAO
OC4gpW2AgX5laA7/eT4xZj9VQRQdcosjBMjYyRg9Qbp5BLEctE+eaQ0gpXtPfF+4wzI7hk6OpoiM
XVDTCMPe5C3y2zFNbOpLEN5Dfj4uRk2JpeZ3pXUw+QCO0oH17oPqrQ3AxxOk0PfV8eGS2GLrOTfF
ffBrYYjfT+boFFz4W1tjfnKI9pGh0Tx5ohpQC072XapLRi0TIZ4fJErYdgAmDokXvdHulfVQmz/U
Hl8IHgoZlE98lmvDesoS4Ehs/6uFX9uL9SrmA+gSXLWfMi7By2NFDw1OHjjnEIMtH5bYrTpTkchx
pGyvHvbVD2SEL2otLVnqfGQtVWvBZY68SV9938PmIKoxSC2YuZqruyU43Hn5Wqa/3kQIM4Hpapja
K2rY8aV2rf8eXVr/+EtRRlDluKabAmL+l7gbt3T6VnoZPcFWKbGsaOpYbpyIvPp42QYa/e2w4fa7
5nPrnaa+M5JhI2u0weLTWeh8A0indzm1sRsonWSSgfq3bhJ+l0FCG8YZ1lg6fcFgRBM/bRrWRijr
uZjReqya5NPylzL4azN+9SZEsRNxjwRwbWnPfSOUzmjeQhfOHGuNNuFUto4qEDrBOkJgEK/l7DpH
/aUbEj0y2tYSO+2H+GHmaIhj3OtBsmT6q14NUdWqUjrUCaZ+Gp9wfP+2yQaEuUEQycil2SwSXO0w
T1SNddEhDKTy11S460nxEazme/rHRPw4P+c501d0Iq4q8gkeT4YWakbgDMU2JcyMaf8oM0RmAK8b
eHnks9Dhx+ySpIPgk7ZIc0zfbUiAbAaSAm8V+rDBgatDUHxZbvGrwKgUJK5GVECnxUIczg3SfffJ
nH8zvjQJK6+dy+uctw9KB7g03TswwVVFeGV/rVyFLXKq4AExf5O996qM1ORYFtMejuXDI5bBgUr+
iUB/nTDYW9gPmh0Or4FHT4xLQR1vdW/W9FQIxz5i/Q01Qh0Hywk9If7mbf3mQRg0tzG6GxNxQ3+d
pJYtRIM4RlPs0qJmRUSqhSlE42pozhXc5NoHWYScb5QdDlakM3j1BbcRRO3ODcHKIg34cg6DnhS6
AmB2ba0gv1OHTm3/NyxzYlJc/VX1+Pc04MBSVYCgt2huttpvuty6Yl+Gg3nEDxjXeePB8hk97wcw
bK0MmZnRr5DlEw8kVsuOGAUk5IXiQZHAanbjmNYwZvLxd93GHJiwvS/yuomqAX9mkBcreAHMJBnQ
1ZQ4YK4nY6zVqZboORajRZjjcP3ZCPF31R9y8UGPXpQup1uGa0DX/1OBmjUINBFrO9eGNhsvm5PX
JMuLZLDCRVw3khn6HkGPiomnAx48HOQjCo5afJacH/+wYnN5GwFE36t8qZu4uUL4r7dDds2GnNRs
v53eBXGFioLFsP6szTsvOsCs0g0UqejDYivauG7RiMANOZz/pzKMLrxKJ44I7vbYAm7mUq14u54g
DRp/JmutCEkcQ4cZ3wwfgaPVe8nXMb60PwzNWQ5VI6TpLGRfu/JTsRK3yyMFhvQYq4opdfuVzzBa
+lk/vwjaDnSghBPOgEmYdLAv9jviQfK4NSZYtaN503yvIIJaExW1Cm4kfseDtvn99KRMj7dEIGB2
PXgZT3gzGRh7wIhYmy3WXfmr2QhpDVTkTLerD2QZOmeLkACk1BANwdWL/1+KinBz0VlwHUoEtv8w
6b0bELjzFEVPqO0aKD0OfO2fDu+sK+P7z4KSI5E+YDWVlD6YCizBTPEVG/n5MK+PqdcoO8oognf2
ra++H7nNuKVbpMox8T5yohBkPExajjrmhPl33MT32wbiF6+nc2EA8ATRl3ofyFv4gLpfD3nscGTe
tEkbSoFKMZgqr+O2exsRFgrmFQKbsiMmwIYj8SX7pZ3ws8I3DtU+1ko8WDMSJaf4rk/tn/B8X5IT
u5gKsHb/flYBe+7Ugl6an9qgfEMk74agtZMPWsbTzgian3LkARdS4LyGlKDRdr8qItGxpbZu+H/z
eV8BW2Nyt/n55JCN9rEOAe19cIA7Sp5r/B/ryXfb7/M0Ze/HOv9uJ69vgZooyhjVVVPfHoinvUuY
aqy0guqhzMHqtqkgWRkrOIuW2PLkJiI9u7GKTgOIcV/pTydibVjFcGw7c9KY9LNqZAUcIOH0TstA
BJ1shGT6b1oaXgh12c8D80i/OuGcoDfZGHPnZb/6H+JjMVIsFdRsMKbT5jR/I5hpttzOgP1tlz1a
LArOv8cg6eeC4pWlXROtK5v5zf43m5JFFRs1sUfdRHJ5SeV0XQM6DY4nHPyKDqjDU0x3ghTWtygF
xvucghv+Q1AGtQ/P4Wllti8ygtK7WC0Mi4EhrN9OsRTkfro934fOWq5Y618Id7vDpLLn1+0lEw0A
JWesdPmCdZTlsTDSLvffFFa78obd7FufwwGS8drPL1VH2yH4Wppczz3SZVqHT4++n4PNhkkd3xns
cG9iFi12DYqaSO0y4XRQgO3O+u0yoeT4XxjWD1MbidMbfrZf0htD1UfmfC7QT9lbZSqla6VCDzSO
x6AGTMY3y2U/zVaEkUThiQuUbDZ6QQ+jF7iP2nJvfcSWCi+JuQYy7gAKzTPpfA5xLxQDXF2EPWNl
ASpycWL5AerLrWSk7fhu47xUQRGnSgi1ZBCOdmmHqY6vLsp5FWIeBlZo5tNYzzQbbH++jpXxad+B
6u9e9zfHUJO7Bfnh+OCpCWuF8Z5mSaC0hHPA8NgF2zcB/2gQWao5a7U82i1nNNnX0tJ3iLeNE9dx
e2I9eGTubtLOY5cMVYM514LMCZpcqgCPjfMndhFyZ4gcvqogOaGLMOU+KCEs98+/+K6avCriaLmT
BuWSgsmORlWkqKeKfVyMSjhoZqSnfzAVJisbf2AzCqyZU+mVn9Nza0sDi9zI5ZsG2FjV81rNXTw5
0oN+tQ72q3DkCHZjVqbQY8yPJDWUO8Z/PnuzQcXmEG2DVMoT/W6/PF1rxhNuQe98Fc7dsBxcCDwH
S8S9CBlq41+zen9MyCDXNYVYdgytnBdvvNYHNkVQcdtf3mk7CSRz9HwUhEuMuC6wi/7iJyp05xi3
cXMhGMwFrPBRVlObv4caaJSCn+fetptPaXI2LX9MkOXkffmiuLQgvRpcCwZmFpPhD+iAXmRgSGwT
eeTD3rL98Ao+fY3f8AZsczpSX43uLdvUwCJrR0wpBEu5UjfAwSXr6vEQkEdTLRcdQdUYgKinbMlH
XiKNNcwmq0UlVJlMWDNhXyYWnkwkyFCYFOfis6mJZm2LPzeSgIpL3OednCl9LxSG5Svp9y7v26XJ
lS7+uvAJFQDse9/KAzlg5YGtX3pDHAG6E625QcUCLXglJ4mnp0sE/eVZUUazvGX2L00IvOQdQBO7
pUoZsN4F7mFVSNggzClAnh/4Wf5P/vx0+useEgLEDX7bwgql6UmFyk9NsrAgmtiO3XrWS6ILhfiz
sHxy/tU/i3bTktLLjNTVUIGKLqOrWzyL/q5ElDffj7TSJtl78m8EIudSRn/zp25wQU7+tY4G69ci
77VDCv2bVEyNRfUjygmx7pkmqtzBRzWXcbWRxl+gHDKVdZJ+fQ+6dF1CkknesYKO1PNRfs48Eyls
DboPW2oOaCfAHW7hfpNpLXwbAftjmPKSMG7oNFGm+qnXCCEyq61k10CRG6TctxZSirX2bsBMc3Qj
kmG5bsmlcj8ntoUb91Y5S8eRPouA7aV2nrteRrQLHM9fx44Hy4VCjaYArCRb70dQcMgkdzsQDj8S
nbJTz7OHCRgEMqLDpZiu9zGjMkNxhLCw+VJayKMPk1Q1rPfHHJdlYiU/3wl53KypGy3HHT7gHcur
EhkmhmKCt0Meg0VfYfjl5Y3CZF9FFeH9lckeN+2K0r2Avx3D1fkeXO2R0Gk2JSFXCDOaO1sfAfkk
V1X0a80WsUXk2/bO+ijqHgbu7lhFQZ50MLucDC55MTITIJS2vLuhrDP8xEdLrJv6RG9+sjw4rb6m
2n5+p4uf6cIOWEnNdcg3whLMudTyv1YjPotupRZT+wTErFIckQSjzpQgQsP06p2hRjPGsjJaZUQw
9WirsrMbt+KDVgnhNhqtxYxGAPBQj/Jz6YShJmOkL5V2UQcTK/WyQVaG9eJaIuaBmYa+9ef8MgNS
Znt56iS/6RSX9JXPJig88eebfpYtzNd3bK14TtbKJajqnRF+IW6Wg7TcVFJ1vn9Zv7rWRG2NQbWj
yz/qcQmirzt9CODm3nHkzoKCj7H3IrKYBfb4POKnNN2/ebjSSw9b/WlUw6MAIMYft0y3rjwoddNq
hxT6/mutBbIHUbiTxLm8+3Y9jDlF6kPJz5UvpsZ/bMldee8kQ4nbRJDC8qyLT19ojcMuRprlbMWu
8c7MMnyj3fQzkHxIiC6RAEdu4z4RUCLw4jwwRkAQ3nSBeElbdSkpdAnf/4mlOWJ0RCMjVSag1c4n
HU/AeLj3PcLnRWIpl8x23LcbXJBXSe3YFVyRnFXjxLkvFrJsgsu/svXn8FMKPFNp7uM2tVMF2mur
Wl/YFRH5Yl+w1Op28+mc4Cp7mTp+G/pEp3hzgpW0oGbmWZwyi1cIJK1VTg6zHdlUniESbP/6woU4
LEoYNnw9DUIcfSwqCtcuvf88xiWJEpmPNAlRHzDS++qkTi1pr9UhDzyt2ZN9a2bMzpGFlvdVXKEs
LJNxTN9ED/2S3eCevPUhzXy8jJG/cSovSNPQAZi6g4PQ3NwnTAXUTCbZw/hksJ8e+oEFv1x9Up2u
2Jo9rc+A8K9W5BRQ4B+Y0s9O9mR19Ku2zDCwZUm0PYqCkcp06SaMhNzVpwbGcSgM5BMF0kZ1c34Q
6SW+c4eBnvzKzwf/jt+nRf9U08J7u5e1B6dpR3VVU6QYoMHa9ddUuc886TzHkvS6jqPEpMRLu7iZ
rnfMD0W3DgW/SZ/BGd4u/nRPHF4hkrpLaFrkBKJdtaKOMZezbdbwspp3qy2vgpv9meheuGqsQagF
BIjyCXu1dRQmHkjUShsVqpZuB3JlRhuvnWdNq2AhNVmibh3NZfMQuU9u4I6G6kjc8+Xnb3sMOY/V
uChC4l05rz7JUiIitHc35O/LCFMeQIc7R6cimcMkkfhh7qhvzE3MO3SEceV1BSp9NtglVfv7ZYy6
rhM1n7OBMk70Ts6sEgemeO+9O++EnBbH91Q9Fl3xMpyR7hfcfIOytgWXWvBgqZN7r8q9BmrgrfRW
WMKgV1t33ZB3qO9pEtHeh2hLVBLVjB6pKAVmf33D6uNPNI/jpPv3EHGidBEftzPNT3t/hzRAEWwP
Yet7bEvUM3A6Ie/9YADTV6Sb5MTROuztWkYNzNBeNyo5N2jxmQs0cfFdOMkoXBmWWAwXx0jVaxSK
7bgR4kAp2274rtCbG5edflEuiwK+ZhoiGzSUK/aarNHPic6703oeoiUrMPmWg9is3QkCphjnCcJi
IN9XLSaTIAVQ8MOGmQcKVyjzXCL0IudHONpQcNL+Fm1qJ8fKucK7i/9uCHcQWgXAcWIbMGxHfWWd
Y7iEpx3aRdfU2+BivUjVAxALEQF6EN5xUV7n3BrAAC5qWmodUbQpzZQJeOSdpZNSRc9oQW0EChgW
diGuIIAgFI12VBB94wvqVGdwrl7Y0/ofbZAUZ2aEDEuuSyxmkJFweT19yLh/WxV9lZgv5oiqz1ud
w8h7p3IFuKYFINWau6+6Hgi/U722WGd8GItteIVq+AG77IG7hSZ0e7Vf/TD3SuN36y78NhKHjmM2
35SNlnZ0JAX2F4MAHltF/qfuTSTZAF0+AD94xKzclCkjbKX4NJmmisJN7hf2/i5M5+PHACqSPWic
uT+p6MfVjkMX11je6p7iY66bsS9BZiYjgaGX2xlKkPLSegC0bTaTSSMo8ukGL5iNO5InVHRJ4nFC
a9YaggJK8joQAPPqAYmZcRhw7MF+PFReSDO5zOHfKayCN/IqLGckNOfC7CYqCpLtwzzTZY6ET0FA
53t8SPDu7SnHpe7SShMaOnCk5ktvZU0zzlilY7Lc8CyobeTWkPoQ7HAz1oALoDxV30axspMF6Nqw
kzvPcFVK4z2flWfFXSPcvjqWTXY8tLQ+EffumbZHgfOdmtO3MF+0aKmkudCYcpokqfbiGwUBouqf
4gfPgBouP2XQ3aRxEvqiiISifr2SHuv5yGiva+xabzVMvsKTzFnEECbSyhAi9TPDOXLEiaxABWAt
mJeQLtwespaj9rbxtX8ODBawK4wT8mZx7ZYOX0fMxylRwiBIIdBPe171bIOawGsqFGKfamtKMDjJ
nlmuzE2Tib2dXfq6cxI2Bnb0Cosi1XZEJZ+aBSJ0GbxBHQ7cCPzAsCczvpNOXQjGaMTawX5I57ro
avW+q2x1eZs96A8JiNTR0LTmT1ypTQ9O2B2cuK0jjLJbeqPkDr5jyW1p25lnRAML+SU0HyR00I7m
80o5luA04LXuawxJazikdHsFyfxUZCvG5UBiK5NkiNlymoAnawzx/N7LOr+I7Jqgg1g3mZmiKiu2
j3Svjn+MvSJafljj021jokOOigWfpbK0kGIiX/WOgpBnbIrKYsrpxSvR8nN/Z/ZB0meOrpxE025J
LoqPEiiDolb3t6eMS4jdUiwPGpljPDy4K5Oqt3k5J3hcOtGIuPtptS43szqmkfyEYOMLX+2p4U8N
dkbs/Iclln9K7BuX5tUVBU+UOeRCShbjyoWObBefsiYlvOsqDpAq9RWLsRl7qwPS9LIYm8zmnmAy
FWeYoh2fKWLx4OG6p/a3y6FybTZt6fO6KHzyWMQrURtU/kqRBBqvtJ6x/k9R04JfWGxlPPwqKf68
Mcn3/93vmLcioCIarKit+e2vSL4pmp68FQA8g2gRp9zyFfA9aXFG5AishhDgBYigXApTl/Yl7Y8d
is6wlkfnS8oV8pg+/hhE76JfXQ57fn80ZzRwSu/9rPpgNxEyPUQl1URqEwPvp6KwC9qtZiggA3Mw
zqMunh9vTbP8dwa4/oKvDcmGq0vidmOUkm1PRDc1wW0SP0zGAkntnyV9ng+OAqb29YjO8t36O4QG
0/chSFwA8wxqObkn6qUpFciFNymumy1RUwrvxmhDgmg3uCmFhsN37tfqZV7ugM/udUCytG7VbuMj
WJqVcyBBZhd4IdK/Fd0xJazwkQ1gWlVI/Ge7kVyTPlJ+fdGqn1o1CdSDO23Jd+cr8jGDRScDclFL
Mo2O71gJNKjs4EOM+8xgvXHjriAPVGA58R2udPmbDEt9j5XLq+KLknA0jdiIP+7NDq3PUMOLYPyO
RCNTshYchRYDDeDMaYFqxz/TO3G7/PKh2e8aL4lvJUovCsAw2idPUk4ILWB2A/w3/2XtzDZg58Wb
rhorDA5IInblSbZZMxl5FWLKKeY5HELkwcUO4QQooxuj//tUqLoH+Cqh1H1GmEipgmHYN7ZvBMn8
EalpY9haTgL31rECHUg3cbK9B3Au/oL5aDoifRYGnsdH68h6hClhCzYFONh8wf5HJ2rQ8zARbgGm
GRvfQzr0aQcvga4qJGeRWi6uyBWyDrUxi1cXlenjuqQVeGI2qm5l0IIExWJoJfzRPLxkX0IvCudQ
NV11U7ewuG7y4dLPkzKP816mk3JVQyifvywYdo21uugQK4iLRnYrk93xzFAFer9eOSATfDAnYTrs
4KnnG7ZpVEkmbRUTWDJcRfvU7keWjt/igrrquU4NmZWOeplS+C1yOClb5FGjS0jG918RGY2kLL8G
S6wULpFsw6EgnPNJzNLBDMx2wfFW7EqN2IL9iqlJlnOckelS8xJYk7Q9AYHGt6pKs4qX4jUbi2Oh
rI7WU4nPBAfk7ck68WFQcb5UWjqIPL8GHRvaQgNlQT8Z6MtGRiQOMAe2uv7qikuKH5un5+lKs6xc
Ju2qTqkpHHTYeMI9sHTGZ7Hmmf70qnYV8+a8HJ+LUS2paEex6T0dy7kVrpPh4RaNqO86pKqupOeE
fTt/kFWoASXYWF+bemjaZFfkmALXzGYNBd8oM8DEyJ8u+D+4uq7X72zC49IwCBSGzeDV9Gf4Zsg0
8oFOCPnHWgt2NV9/PNvg1cPx3t45EQ2MTo546nBnYgIG/eR4p6EsOOiYB8ee/frd2RCgA3CVrprZ
B0j+iGfHOOGvvpBazPkRh0attfxCkDr8hmxewzwLZg3aA3znb4rmVam2Xwx8INiW5JRQ6ismFQLI
8xfVnE/6dJINXQDTmIyscHf4k0BgFI9rsT1bXvJ6Gobb/wCSZzVGusyB85YlmYnhqHoSa6xIfXzz
rJL+oo7V8yTjEHAPXnZ4TueBu/z6mrkO830/W/yLWdfyWSIePqA/uX6IJ/WX1H/iNyE6aBQLSfK6
eBBNa9KhxToD4LPMFCxwsvW5coNKPKKAoXeQbLMMxVZC+CL1tFUph5Fz2WunZfUKLl5a3jDMqRjR
5AAY9fHqeDPI9VbAyqSnbamYO+lc/BstqHWjtjUeD6csG71gGVnbF84LqZKtey1Yl3qpC7a/JIve
lX3EKml+mwjDMndXZEPkGPH0escYbGZaIeRnWN1mXusfOCy2AJQWs3r6W/12/USxD2B5dDMUYXzS
+aS8ptvU+W7hTVHYjoEESnsYaPkSndFzKdM/ikwmvtdYPZYT9C0s3Qb3fX2sGAJLNMe8LVl/vU73
J9CMTuoL7PkiVPeGc80rEKPBmix8iLikVHQTvWEMe4/95nej03IXwayphmO1Do0KWPKPVXsPgvxp
TMxvZCuIMLDDFMVN/46HPZbT2O+7acZEWHSRP8JpnW7RroGecgdv5ui+Qi31gc+2DM0Y9QYgBNMw
q4pBfgI+yEf+8jveTR8u96F8Sokp5kJlt0BCBbve0WiiQIiLy/RU0EpODpKPl0oDVaUZ4882gtTm
22FA2yrDnhm81ojfez3QXt+eqU+/3PCIlGuadMAmX8LyQJmWn3DqN2Xlg/Zv34CAi65zjGYv2VsA
0BFCNWpRIJbi5jRVv01yZ1pZCpdDgD1og3nRKqBswoNuZOLieauwwbejO1jus6jOCwMbO/Z4UJs/
+AjxGldp+NpM2wGzMTkTm/jPuzH9wPd7rl2Q6OxfQo/HoAmhqyJeOgICrjEfc6llTCkafltLyHte
MSmXt9JkAt2sgOMyqTjAsrMsRd+NdJXVe1OdVa+I++3J7lwvD70QKJp53jwHFgOKX/jb2LlFMwUz
V5POqXf5HOiZg6mERHeZ0QiCTE6P+we3CzTvLROjT3CgrnIrDdXKbng184+JLSOK042scQZ4tDj/
oj8lrq2WGk92LFsDE2ZrSrrYrxlcZVex0rJ8fY89vyJ6y5yOJ/XWOW73FzSXCJpph9kAOTB2CagR
j/QRD9yEFRbRi5oEUEUj2b4+UIx/2nBDmgER1HoB6iLtpRVltWV0UbSw+azqLjRObuarw4s3BBNe
wWFvEmdI2hB/lJyflCF1zWyv4TzJErwcjMyHiaT7edXR5jbJTXu6tQiUgCq4mlGs4e50uebakjMq
lmVrWfkzu6BEwGyyqpoq+XLtA6NJmIo2BFQ+Ttm8Oza9LXouzzorPi9Rm5jQtQf7jW5oiSxb1dNl
kUbjxswS6Zgd7yyKFpISwnPf284EaA3hjg5LbdhkNnkqzj5VvvHXrS9udsLiXUDEuqH71iDERpYU
Odt3umCwuZOd7eoT4Ja5zpeSsr1lkx2JaNx44cd9lh4BFMJhX3z4Nzrg1ht2Anzmc5cu4hH43KEH
skjuo4wNhOBFkJT0vzW3TeuVGXkW3c/Q3oeloQLJGdoC2oTxEv6a3lFtBY7WcJ3YPi/+QNU942KQ
jRbr3UGjpYwaobVlLp3eL7cbD5JfuK3w4HyoSGLgzX+qjOxGMENAFdWaetuS9Zda2DB22N+afuhR
45aBlyaHV0//pj4QneWe6zMJHXttLPgL8/JBerSJraQPhD2aS63pju5uNVjABsH6Z/5ch83H623B
4+eFKJoUExEoDx8k+Vv7oZTidR8YjtTdKmtcde3UkE7pnDLnAHrkEhAtoTsLnVOHsXm/hfJV9+Dx
x7xoYZ5CN4/WqaRmDvip9TOjW/ueLQh86Z8MCpJeZxbac0oC2Rl19IQn36d5pEj3TUPPgrzVlsz8
znUyWR5+BZdK4rFO+uhMj3nw4mXcOAzD+QyA8O1E5OPfcr+0vPN/AOLtuytDPsASj3wQ04Dc6ze2
chOVt9UzrFRL7atjQilqajXVJmh9Nb5ZIQ4aPmdD8vpHcdB52sg/SjivxKP1REdof2qmVFVy7O0H
XJ11V5+q5vsZUBvsrusx3S2/ZBDgxfKoXc0oiSMWbp8lguRIKJRAFmV+CRNmEaKvwQ0ZgLb3DVDH
SGgqQqc8adI2mykPqn52b+wDaSjpFhn7vfA6l8skZZXz5uIy5Al7APUF6BAlGguclWNM78QENQ7a
IescYad9yKyhu5iA6iL9Gh1YHZ4oB7ePT8/hb5t6cTrWYg4fhtfrRG7AKnpfWJJMRIR9xsurQgtT
mYX5pCOZ5ljC4/Hr6E7bM15O0uKNpwAYOolwsS+VMZOnaaDXSIIUpIkmMQPLJ/Ja9PIHjlZRg/s7
uljAFfAqHSqRRKz+m1wWpjUvNHYpy2n7PRUrLaVkT8BgQcV61mshSIMD/gWjHPxcGZB+bPrz3woj
3w/bvetGa9rNn18Ccocw/07Q9rSK901ABQI+GIluI2a89DSsBTtS6Pnov8lkckHg4GZK/gC5lMbT
Rz3Tyb54IKVehDTNmplbDRmd4U4FAvqws3MDRzxBLDuYpmnGaosbM8sDx6Fvm7PjQjAitjfi1Spp
U9g7f4NqugxJbNYawYBjIf2fv+o9TnV+FsycZxVgIsXJ7ju2G7nkXVkAjz5sz7kNE/pYkQKJOjVW
EALhHhiZ1XL6Lt1iBYYLMyWdXAOGR3ixY32M/ymeOG+9uOEtTPlwmyXLpx3xf1MHx3me2WHm0i6Q
TcX8ToCJ7/8qjxqxOZ5F8FnOqwDF+2IKShHdM0Xu+4vHf3iYgFJFXcNuwlQQtTHx7idJqqqorEdE
XehzxmRpdciTqIButCACf7OspXdNPYSjQ2E7j/kwSF66Zf3i9HrVGexxizxwaoyhTV56GmPsJJb2
8ymsleyDGqZuKAaYWWiFZwwfxkztFx/XphrW9tPcguLUh+0BKEsRHGI+BsZISCAIFz8zGNIIQTRP
E05e7GINA36Nx62kIVGXYFPJMH9wjA7ckX1HccaTRjE5xCTvpeceG2nhLWcL9nmOD7u0nWUjEBHv
PH9QkdEt61yn/ECT53O+1jCeYNH7v27FkVfR1wt+AiTZoqB+a9TFPC9oDDvFAazfbWtwUaBxlawC
a3ye178qp55/41cFoLZoofMmAeck3lBgH1opwmjrbarnlm6Fck//l5Znzvw+QNhDQXFUCHcQplwQ
jHvI7nIe9BZOEfbAsNqIALAQYwSjqLP9bweDtTdcc39G+zBtMDJwQw/6QnOwtauSnG4MWOBsdTDQ
FEkfpEHwIPnKTwTKxVRK68yYK52kIoyOtwnHbZk+ExE8kvunzB/k4M3FVTEDrDJ2gclyf5gZwexg
qXMX3dgbdAL4UBATsnpj3u5+472SZJkqqyotpqYPxn2QBDRwTCao3QfnX49Pb+85BNKl6N7HYQ13
De1whsxseMOFY0j/G6hypmcq+mGZqQX9wOHDA0iYpiacMsu8W3x4mW4UFq1l6/6aPSPfO6tK95A2
ejJnAP/oFskmRQS/86zujqfgWBujyAGQpxRm+IsyUPviltVRkin3ffkTXZN+gIRE5Q0R2OLcVJ8J
+N1lsgNM/gnVg/T8Dk9g5aSkqQ/jLNcqW8KFoesB0K3tUt/Xmf54Iw22p8SghX5x9dBuEgSpwFEV
41SPU0eB1zS07+o8VNnQf0wLC1tUqwTP5P7nn+1NxFJzwy6QAAcXhkfC2t2rgYQso301gXSgJRmY
pV0Sq3IDUlSRoNUB2teQeVRzaxr6cuUpgUpfm89NKa8Orh+zay/wetRWDU+fEGoATiQuyvJJ9Joj
/WjlVmEGpgkv3n7xyw2+CBKhAMKE9gErSdzeQ8It8tHklEOSIHIs+ycaAX2/gtixnXwxGE7iXzdY
yf5umQbJz2ToRX8VNtiwyBxaiscDZ+i56Q/DJa3LETPlj8YJwtFYjho0YIV2hl1KbUSjhKu9JUu8
+d4KwTktZCJr31FOcGsBBD0pES2SHE897aaoL6+7mzDvS78z3ufp+p1qxGBXwxP0deGmi92ZDFpT
nY9Fhy0tWVohW034f2AZSCyy1WCVLubQrBZMQDt1mGwsZ9OvkHraoLG+SqyCDfkeq7R0JZj2+rGe
MDgZIS/VHXEVMTJ3ut6of1k9RCx+szE3bpCrDeDNbxDuXU9YYG7YV8ukQPv9ug8gKLLKlDQ9VuQH
hUKNxisSE0XcN101cYvpvJhh0zQNjBiFZBMpmFex/T+dc6YAJgoQjeJtx/qxlHJ6cFmNsjTzGgDu
eEK9iVRFlAqrTW5r8kEm1tYrK9KtYA4uXE9v2kP1pkqND4N13/dXIkmcywdFUXJCJdNYEs9Ge3bU
2ShuxYTwrEQ2HmCeM8y0l0Gu2hpLNkk7ABcpHLa+9m/wFDIMynnAm9mxwl0nQ+UPtIPDukIdqcP+
GxBPGP/37GjiEjVlTgnrDF4yP9ruv2HM3yDD4TwVdE4+hEmvuJODLPEc+3LIqSlQwX+4QeSYuCSz
JKLokhdPbFUuBgiK95r8xK5rPRS1zj8AbAY8mmr47nC5hb/fNnls733H6tjaTIwBuWMxs5ma5tE+
DSs+0KppJC1Isaw1mYrgmMabqCMXqH1as97t5l/PCj0Du3thQjHUkPcdggYEB4HYQ4921+DjLlj4
oHmealJ+YJ8SjScem0ZnFKcqNhJacHtcnEOvoIXuYC4WyIA6kZuD/sIq76xmeET19x4fe2u+IIQ0
ODv2ykSvyKGVBghGHUstbI+rijVjO7KW9AC5Ko4gjE2PYe891ta8WHHVwZHWN7Tq3GYi2bNN5nO3
wUKIsRR48aorzG0CKTWvG5fUUSEUVvkvmLP5vigRPMujuvWaizB2N9Rabqqu0L7kximS+Rvk0Dok
FEHqYx29+zAD2XX8+IEI59AD45iFhM09yp4SANJF/PnOSKmpyrcm8mvkoHrCDwAysJzuTgUrg7QB
7aG6HEIJxRiriEfoRiYsDKtVplzHzPREI0cTJUkgHJ66Z886z2Ky/DLOwBHWAx9j53YmAypSsz9L
CODqzRbpFc0BRz8eaT+S3ThDRK0UBbrf9DuAhpm1pAaNiEC8Rrw/M9Vt7IZbZnkVItCb/cqAOBrF
O/sCD7kzni6ivQKNy2YnvR/l02uyI7KgDX7QYgYtf7hPstt9qrNIpJ7uTZZJFJLFc6asVzOsHqIn
sOMr1fInt4uBa88AhUxX3eeRMiD7agkX4rYO9ejQhIXnihCT/0IeaGvVB5eUlRoS7IOpA0q440BQ
ryA5BIQNWU6bVwWp3G0SHR0GPbT1o+a+++UFcEbHm4pIOj+UhYVOyymEG3Hk/SsXm3T1rZ3xnfrd
wE5AFwY3rdj/lHi//Gy8aSNKiAogVuPh3oFNOfobEEankjL+g82KU7A3XOFh9NOKB7cZDWDZ9mf5
My8PZAzK4T0NDn52bCCj09mYzSrhFvTHmBVB2z18QHFrVvdgPWOuW6mkIZVdM337eMN0tEXPfqEy
tUI0qTKnUmSsB0kgt4Th4peXb64hQdxZ4CUErkFFOoPWwLp5SIQT9RkORb1in/EQ+0JWHlJNlLf4
fi9kjelfNUciwcUnNtOOi/wbJGkHWe79tBObSyIv0egt6kcKfmOv4/DO/3KkMxJlNBMIWTA18PLX
RbERukUprVb0DqUs/wjHwH8LGzmCyAW2GmqA77/5jy5/tBGXG0pBhIC5vzJLpu1szW/O8+S8Rfoy
DO4xtsWN2T1La9b8mwD0aOWZONjgZvhemQ9xwgdXG6kmBl1jmf2L5lB7lRBKcVf9Tq28FT6ofXLl
iTfVuaS9luHf3k9yJ72CX7H8Wy31/vfGFGj8fR4ApCKE5KwPBurOHwppGmVNNI2qEAo8JuGLrxnv
t4ADBoMAs05ABaXJeuFRw2ELoCNZNPJ2rrW3gSzG83xeHsGCeXgbea6Gt7IxHPgF1YrxaOne+fFJ
6o4c4myAsdeBBfAU4YS7XZxKjRW1JXeaR0Wlt2GzAJmhbcFJOVQxtJy//Gz4FzWyYpCWZUUGYey7
uxtn7U/6OksXl2JMyzktefEDh0hxMS1AKeeuN+NpwcDTTkgI2QAP9Wh/FGbkbKXuRsQwrulEQR7u
AiGVFWRaH0D6q6lJWSlC/4eHTuR0mXF+fvmNvxXjWk4MxiB2WhW066aNbh4Ab7kEmpE/OftXeSh/
1dYNTrS/OXOOzPVbQ+LgQLJK5oCZVm21zBiBf8Jwtb8uSIPxmM4yWRoq2Um5RbhrQcLZmLrGAqQj
hj1fYHwczs0sOe8hSci5t0ccDXhulhdG86TUSBiXFefoTNjZwHBlwuc7+AzGLZbuLJzpmi2KHkjZ
5qCOzltlfvwoXGH2pc5Zfff7VlYGlLeNvAxZwmhS4ejtGKjbcydytYI/sNR3aqg4KKQZy8IXrnZ6
LYpsX7NJiTCmEzFVFJs1xsEgRD8l0253iEnnCrAh5N42wladbIuFJgowWWOl51kqUscNrBEtHiKA
ft37ufyAs0ru4Ywyc+7OT4a5+eEtUKxHasCBV9zmhUZ7bHrQFivHD9TeFAokF0SfS0Pi3aMkEs+0
tTD5Cajjjiy0+uZWUT4+RI0FnAKOFYOfuVxJi+HnL/viBIpYLeCtsdP77wp1Xazw+N00KnbUivzx
SCEwUP1CuKm6UWCd3rScS4uG81xZvM8UBkN0DxeaWNXF3bvaQXkgnO+tmWEdKQqrzI+wVibHb6wL
5Px545SXIEfANCRYZomm3SNzN6D2RpjNJ52fxhEiVrcQWjGTM8Jwc7x9vdgFjZrMzjvZ1uw1qmI1
M3zP3GPAth0XZ7dTD/QLNYeJEfjhZ/RZkLhAse251H6ZJkHzRq45JGPQ8rRTD2rg1U7tvu7oChYL
Z4yVEnvr+gmvL6uFD28nTFRxJE18guSXZhT53VwbekJeGeGfdZ0=
`protect end_protected
