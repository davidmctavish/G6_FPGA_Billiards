`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dRPyPKIotlmxhYMz81rVSAdtdHlNVfc6dPI0wUOlA/0fsImqArsCYqsRQVFrfdLLYClSf4nvhujs
MeSx8CMIpA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FLY4tYYoOXm7BBAVrydNeUvulYTBaJU3tEKVwzI6Ls7rsvFii88AqR6fmXsDOxpjxiy6De0KX1vN
NUUnSjDUvjO060tVufULge24MY+Hzwbj2AvPwmzUIKEaTBn77LHOOipABrx/mwE5qJ3tKhoQfe4q
4bG5Z/Uni/09jp70A/Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CyyXcBVJ357hGP5I7+JdONSQCA48iZ5g3oYq4wcXL0C5/MGI+8dxnSi/tBYIP78Tg95/bPJdXnPV
9wXGYo7UnnpMcOuTj7bjhxqDWj2sbkJHXSIPW/TkljIqXrZUmlOsiSuNXZELXeaEvR1aZwfV511+
Oj+7zPL2AtwVm7pUgGIsjJ+KGNOr5N3W7ahYR+MM91dsxcgxTntT7pJu2r1HZdcthcv2kfqmSViR
UyIW/qjDhpAsFqU0x/hAVYVS2QX8BnZlNmtUN+4iHDXyqVy/grUexR5N8lRQ7gpEIfybMkBcICO5
gO92tuQa5zaaZTDrpPAx31kPdTJr1bE9OgYouw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BDXiNBUuAX5aJjIB4q+UgX025MyvVgGXDo8jdQHlx/IugIpQ6QtT9Mb+ZY3H1ZGzrrNV5MOp7ZEb
EHtjD7VnsJq/h4/qNCQrTTjpraSdnOn3jUuPdoqF2HDjaoOI48piIsdS0nvsfGPDgrG+7CVStygL
mH+B4ecIuVyXo0jJ/+M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XX/tLKdqlgockldwi6lD6b6sEX49oOSDHrVNKL21uU5o68mAYzcenXPPYZgfGemnageSaunbZLLk
/Qf3GE7ViE1VFNjBZBL+lBdt7RtPLc5+ccpD4UZEtW0iejqjtKIP8+CX2sqvp1MTuQmDvfXviZs+
UrRSRWiNFU+WmncjEeTkIc0kDDTwyOw87Zd1nGlDz4jvCu3lGm2l/cgaXa5sFKFiClK2glWGidjU
j6AbWjrAzYU4Kay/859TYFg1ogGRoKOdTYaKMRmFg2rHIpiBmjy092TSifin4uy3dFF8RXF1eyW2
E62EsOhlmrA9e87Chom2L0uXYmZb2KiPmrsCmw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31072)
`protect data_block
GdAkXmS1zhVrET+Qp53/KHnxlmAHKXR6spvcqWmk2NGLm43Bs7iCYHhkihwEGApqRMdD3udFjjEY
N4NdjaBSgG+8Ajs7vhWF2ZHgS6IzOvhK7n8L1birWz+0pAMi/LXJMGnw3+Ud7csCRGnCz8CaDfsi
DrX4AAdDNWzU/4J0V+7SBChkHcPeuP47EZOZPNPd6Kp+A4pIghawB490+80um4duyM2dNauxD+Rc
RW+A5UJ2DgDlA1/WZHiJ3Hj9cJLXSoTC4LkdRH59BG/ZS12lz2ms4WX8FZd/Lsf7QH5zVH/N4o/2
bjqpg3xp63E5a6rJI/4LXD3VKY/mGlN6Lu2AABEhRb2Mn3js9C/1DGmdgFuIUw43DKDMMt+0E8mP
suyk8Gtj5w1ZKhCH7IsvEO/DwxgoWpQsBOiAIrXaWMxagxwJq8+uIme+76wXmCBBaHQhwo2H3Uvj
PN9Go5Fi59IwJbN0akA8A2Venud8laTuUSw/cAS4Vtuy9dQq3tTEwLxNRI9h2AQ7+ndbi6p1jMIq
j2LQD9Qs/+HdHFjFR4f16J/tdCTdd5A2dDZ96VLfeG2AuCXBzmGD1MUlXTN0VtmRV42++8qXg8KN
HK+7jgaOGvAfLBK+ak0h9OS/UgaJnqmFTAL7hCRmqwIV/WuJ/P46W47aDqmyVwdoF0tfnNQCXPj2
jO9+d2V4X7ejbkSOJifn7tsIjhtmJ324dbf0KZ0ZzYmjXooGIEMEusfIx7NUCxEzxhpnXXYTx6fp
YeNcNGgMjwcA5kL1BkRlvB04p1sEcYLDcpFJSIBwB1NhA2bJDIAJnd8HfWiHqNjURpc9XkJkeJAh
KvmEMi6qYSQxUocfnZ/dCWQQZkuSoQuPDrBVC2AMd9P5W594CoEec/Z4pSbZgKhtEZhJBcphoJzY
okp2oBaQjkAZQ/Eaylr0hd05nJP27TVxO3Oiai85beYv8gHrc0k1I0tTscHUQ7MR4v7S3r7n/bWq
0aMnnNe+I5rYYWgBzjjKa20Mma/cLTs1f0Q5AstbjqeuqUKvO2WMdxH03muJnGZp2+K0l2Df1QD4
tl02jUu/YEyw92I+8JG/z3RmAxNBuJLeiXrF+6M3nF5v/VTzWamujkrunEJRcoietfwOIujSyV4d
7M80WAD3oSascXd0Lx5aijoCGaLIVreDtZkI+DD/VOQwq9GXivgnpOFs0dfEsxEKlhACsV6ooopf
w+tY7xqej70YF3jGRAOwTgsW6c6cg/IcfOYKZN1tEnFBkp0poOKCFFt8Y7UXEvivQp4KdYE7So4L
lKxzdwa37V+/M0uHaQT6S84e6Yujx6c0WLgEkhw4GFTZyEJCVyq0qanQ66BaY2VmpLH/b7S4zkTF
ALolp2QBjO6vU5pZmKhXeUFUmRZqvJE5u6ONkhSQXC7lanC+H48DWDCAYOM0OCpe+cf33WJ0luHN
ZVtkBM6BsTKr5fdWTXZoFWfG06AX8r3WbEdOVPsz9jIYWh5sYMxt54RlEkgHZ4Otjs7rJ0XOJAbt
Ox82qX35jXLK0al86XRtvhdkNbF6dAUdR6BfQ5OpiD7CB9UmjR4vyc51iJVzSGNGJURp9F9SGimn
hEUc/g5vP+FdSMm9HR6CacllWdRMHt8fq9W64rVvRfQCAmlXKRCrjHg2F5dJd6qYBQSturaddIAg
JkTk1oeeDpln4f84h/g5K18HFjd9TRzqYBV9gm3ooy+aXNA2yy8GqNQT3bDlph8IrtZzcE3RwzKj
Paww5Tw1s4kwcAaFugg55Kj4PJKmpA4Vqgoiy8SbixWZJ7tTsCdroSwscWD6abnAtkdJFR7vCWgV
lsWdgDajbx7lUzWFUKO1rk0WqZUhwk/F3fB4Rzvdsd5JQirCdRbwr9zGkUyrtNiX2lyy6Arec7B8
GeobhOrnvj8R4NSZMKm4AVdLOe6y0RQNl+cjJwGas/8pRUhR+S0SWVAPEqILR4TafI5fesXPulK0
cEKbbCFFT+nixHe7EggsL/x1JUftKwOlqf3aWgPPmSK0+4lPY8Y2VdYAQ0NOoo8eibA7J3eVDoNG
ssWl5GO9cCF8nQYLS5v697Zqt96lrweMJDD9PkHNekhrN7P1n7jkhTBzhkuMDcB2NngQu8rea0CW
c6A2SQ3ErLyZYoM4st9JQSiD9KxnybdwO6Y+9MT6Z/G6R3fiucyW5Lt7I5fv/vS3pNK1NUWNsD0F
u+q+SxdICW07Gt3RYHE5Tjoh9yAsUlTI0IljZsGT7AVy9QYBAFFQxkSTR5tOID6aK9pbhms0ZOuK
3FuTK6HQvcUaCqHKC0p7O1rKO75Bf2BHqP2KTWdeBOXiLVgZVRIYOrunYSZjwFQ+BmRPid2pv4T2
OiyD7JzvK6roYH7Gucvf46LR6BO+1GxCv58VBiOvSQMwVtoCC2ZZh01zRGudQy3DVI/g8leP4v9y
CdKs+6OK7ynZAx0hjeR79VaGKp6xZQB7OP1E/6a0CfsWLC75CPhZUlFCiKv9d4GZYyYNNTrK/pRP
pnAKSZvDsI7uma8Hn787GtlCVONZI31ua9PLlumfTR2if5HLjrwLM/lyMS+EH/Lr7hUfuzAEwlzV
EHp3fmkKnadtfWi8KcqMTmAlAJiz6huooA+FUmKwMR72uOjYenLVlHUUbIotNlih8uzc/QIqJZyY
OOPh2liRzxk9qczI4ezm2+lZGd7fix9n9hi8YpAYml/r84ffWB0J6fmTZZldySixxYaf4SdWUdg9
23159bQzzsafpBmD1j3EeSNw7FYrLl7srxKMKnXl5yA3Xm6kKwvrFq7vJ+1ycM3ze5z28Q/d+EnV
3Cc7JIYFCShkJUDxG7Ewf1lF+EaCpSgJiUnmUzj3Pgv5FnXuKQuUlApEb18PreZ+fqmnt4YNgLEj
CJLdkZLtwfVlkBsWAGBtH96UxKRBb3LL6GOscMwgjMYaqRCuoeUkfUaJ9pe5izPDKxBySQ715g2n
jPFMSmvPMzQlf3RKp0f72ergo/5jaxOO6275HEfG79IvVhoSuZ1P/FhQuNgSJs5H/5SmXvAZ8/CL
7eBOD+vxoQSQU74PG3Bum7akYo7xVWPy/A6t0yGrjqsSEwTzjEH7fDOrv0DLAk+h9UKCAhrl06V1
+usX1X3hHk+69fD9OYNM+bNRcA1LLeq/kn0u9INfljkFebEyCxwx00W+7ZUNW6zDoXSwDL8yaUnV
9Tqz6uf219qCmcLz9Ik5SISX/xRLtPduL4LdGDNEfuhzkWUPC3gdqGV3uXPbNpEs9EiUZDh3cTzr
WjN39VuPpPQ+MWj+SToYGI012aWNm8tAuxDRIkVAp/FpipXAaVyd2M6zlF6X4ekSjYGmYBHSxm43
pz4hc+cBdsxN0swg8gEfkmSW4rjoSVNi8kOiR65iIecAbUhVjfyy0gUCNWaNtLah3hI0JnA2Hanq
3GNi0qInOpeG1/1b1zs1yIe5MXag38oTpeMFlWY4IaXg/V2LvVfnQHY5BE1VpUsD4VIxfewK6aIg
kbM+nv+Xrbq5unpYKtCdG8Zn5eeuEY9N1aiPVl5oPf2P/RixPwXAwck1PEmqmWJJP2akdpFHrr44
4RNyFyR77fFINIQdOpRBAsZFyDPtoV1kDJTSxIZGTl/k2AQmX6cASWn/opVxCbnvhP8bFgQXM2w8
gucBRMBHj+P8K4RZcmAfHZ2dL1Lk+buRESbEGzS2tQZENRXB7E5umS7Fnwg7t4Vw3+ynI9ucrseM
q+0JMBIQbdJjo8cePraX3phojSUqTgOqqCNu4quoubscnamT+NdZWbiAaFlChHrYGCniQwasZ1RF
aGMWzLIpz9Qd8kZYx9I0CDj6dsfg96XOdxBjwcXORmNIexmSJIvIY7HiRiDbsdLIk8uoZTDJbs17
f3KTXgoJhearM2bQI8n5uybWngg711GkvMFcVipXTQturnNkpJZ74ZVTr4V2Qw4R2EDXJ+/Vzfod
EsAvHD6wWAmOiPIDeOv4ChrkRV7biRvjN4GYlNcRxzwrqjHnh/5FdHlW9N3ZzDqHKydLiqwVb4hy
yZhb8edj/Ja8j0A0T5KNXyszdFpRW0M5479WOzmjsJXInFow9sBFRbAG3KjYqoSBIS04H8IIIQ9/
Nen+dXr2Uqqpf5zNbw56ey9BwMDuH/fORX3vk9LZJX9tuXoFTXx1HHxeHeKfB4lU9ZSGVxYsFn0l
FHBMwcZ3l0iJhR+FN07zM6YzCWJr+lNOj+OpPoygKLrTxtU6WArpLqX9wMN4LZmqrYfJzuFZvRy9
dZuyUO9c/C51a0EYyyDibvB5SBbgB9PjuYNCU4fdzyDSYK14PfRHfMFED+ooHLk07JJUIpASH4V6
ucQA3vPQyzzB/1QWsrKwjrcfd8GSF5O7Aqkal+777NiuHAQLNg5VtOdPMmS6kauLlL22W8ZsI4eS
MazZO4eGlns/lM4KOyknRv9axm+jrT44JmNv6DcaARlV5O331AnjkLNNRL1ap+cWB+LBgx34V2VP
ICFFW87XFSdL1OpauF1Ey5uBnKU3AK0Yl0jkQc2crMSxSVZ8qsxJgnN7VK31xnFFZX2+Md1UGa5x
KKdoD/lipQxconpRMLybpXwNs6CARUvhcEkh6NA22uWeFrIHcIWuKjHtA4lskNvSsedw6burFpRi
5RFZcGYkaW+c2+49brAkCcdnZOV0PodWKkPNB8pewwynIIMkmHUsKcDBaIdxT5dSaT5YOxnFC+PF
j49TNiMeRqe/z/TiXErKL+EvAx5fIM7T7AF/NiQyuJUl+FATXs3BE26MRrco5pN1scn8ix3RjD2u
7wV0bC/WWhQRD41yduCMQfOVnbM6gM/575ubWV7ozYj+6DIMfROioD1xnqxziTSBa88Mkba8VIoe
t7l+6cZ5ksWyrU9kXsIMILiyRaGvUYSwbiDFCM+L5gzdO+BO6uUF+/RMW3yyIPSNTkWpF4Xkpauh
DYB/N6z8K7zP4hDXqiHKvGqbxrCLxYWOjmR4RJGe5KErASHbuYlmh5LzxTepWCwl1TZ6GVQAosHn
HkIgXhSp6tjq6rdVIibm8tF6Q2PJbfO6T17eJKGNxef0rKiP1bMMe0YgH8G+RHG1Q7jaT16qllhy
y5rLfTkQ8EH8egixSyHYjppaiCCPVqwCotlqmjnRu+Y7Q/95QmqpB4zz9g5LccZDVW/HA3eXU53O
iY/y+RuUwRC2W7KaYn5zAZ6Scrix0Lp0+fWRxYVtw6nc+R1cwm+a0+igWlFhb41MUiL8J+bwhJYV
C2BcGbUPOCxHfFg0tQyc51IQGkqvsBjeOpQ9r+tWWnK+tp4VMAsMSFlWoya9JR9DAPcP6f1mloVi
JTXDzzfbxhGsqky/+cIyj05VqfWclQxHMByxqVc/R73IOOcHWPwjXaMDuarXc09IsHq1m5DyY/Yl
KgIHDzTLxqoJTWejA+6hm8nwOibUFetAVKpSyWbO+T3r9UG93+YIw8kG8oC+YNNRxq/rHvmwNBOS
NUN0pWlVFTqOcaA0BgdHNCIGgenVPqWI4DT+cmNoT9j1zd3DK4NQG9RE6GoYgl6+3vCKNErQFX8K
uwSvuklB3XUyi0/mZIqn85L/yNC2SLEReoRRsZ/BGj3lr49J1aar+0yDGJmGg81fEc4lm9F4G4/N
BVhAZ3d8/VBEuyrETPIUYnCv/orb7irGjT0QPgI41kj1L6n9PSViIHl82T8L0wnX0ioCER4SaSwJ
j1RETC25N1GWkRn4hX8t0veQvNdkmWz/r+2HQfZRlhA9fcejcXgDQ3OgWz7AtaTKCahfhJ0+ViE9
RRPTwPL1W46uEWnz31OPpgxbt1kza+ZTzpk1jhXPUqUwdYgou+F31JFZIVL7BAF5MYtK6Ta1VHSO
naNSbHPskJ3jByMKPsfqeyjlrFodofasmIYbwtWOKQ5TjOswZnOS3UnHjQ+f+Fd3rbWqkNrnCCT2
hqDTqcvpSkS652lw1up13Uw2dMW7zinzVSSxF8+5YrwHSrvL8NfoauoOco2JgVxKymm4AWOc/9+t
O6PSACbKXiOIvvBnDUez5tilRcR8jH2TXLDKgxOZP+3BUB2T8aFqwSFU91AaU/B6TOBtUgBcwopx
Qr0Ynjg7mZmmLVtjmRKc2BlX4T+yuHcPfQqDuWDSVCVpUa+bk8ox5lT9Mb6x7gRv1X9Mrz34eMEv
q+frA8hwLMJQuonaz5xkyz/uTdCyUIZLYhITQd4zBzdXfgl0LyTwbZvN3rXpPmYEig/WSVniUlj2
STIa0m7HFijSfhByB/5/9qA9CbQehBdKhj5zIOFSxZOpYnttTe17PRCMvfRFOmYvX5iUT5UTHIN+
EXkiXlBOlUAizsdBtwJTGgwLDIEaBRXCAcqltRaxgwARtf5yElBIZJll1ilmkfxY2mqa54DaCCN8
ab0XgTiIsH6NZtkQ2nAhNg6YczukmokOpz4yL5hnoBirLMs1duPOOFI60Pm9YHeXQuvjmWaCIa3W
hhc47n2DlDuVI2bHb600o4dNicMqZjf2PaIaHdBddFaen3ArcfQmgJgGjr+XmuOM34JhEqm4oGKo
CdznWzCsLVksq8sIDhEyCUUX/rM8hjJN13dipLYRSI4sUsUAYerclgmsHS55D202j3JXqhP8CFcD
OpmPU9m50hyJsRooXNYM/g0lmJ1OzHgsDtS1uXPasTwhiZE18kTJBl3HlxpYcG4Brax5r48TgUZs
Bbhb2ZXbrCk0Rf7FlKicDRHhHK5M9BLqm5ey/H12ySJDLyYHABaH0ovVgNtuzvHGDmV2buueCykk
T6DI4yg33AFChHUyFIsJBPGpJI3WlVPNJQZUphpRhcFiwLIOCpxSBGwIRyJw8yeuS37IpI3DuQPm
1/imNtXPcrl+4X/Q64aj9e6rerz/ce3wesOmqWq2jTy6E+n6e/+lIK69/gf/+6eBSoCUh5YCL2b1
D5LSi203eeyNFogb9/tF7Km9UJoiVmM8hRgsIxg9onv5TVVIjiVHpjLMtmIFIJxPCf6KR2+iqAoY
IKEuX2q1gPS9kIsVCW6D8TIcZve29CknpE1lj/hF3aYpeD6bFfpDr/DKadSh8ujYGFvE/Ds210gr
u2OxNVGi6vTfLB9fpbJUgTQeRsHYlKS5kcXzMYEiu0zHpPBc7enm9GSlJZ3YI8o88sit0KIZ4Ml7
hTLP2uPtg55scPubpdKo8MqoxI1ksaa36vG6vmOePjSORFQh+qPufaHgjmqWUoL/FO5wXwMMHnqa
Py5fERqxgRpYNj/2xHkDFXAE04Hmh0WXM3LZOUHIBe/Nq7UzXG6y6iDscibbg1XCfgElAtinTa2B
AunO38dWVcXU4yWn/GVj9xfgjYQ0kUqm0PPnvsr1TjNXYkZucd7GNvhglLQclbj3Jj/MZ+O5ih1F
IOZZeixi+Nu6qwnvzHGd3qFQGiHc/7GPB5oS+b6MHk8gdmYpOIqntS9+lhz65/pBxwRN/w9Ab1la
0gtuOk0cfY6GgcI/Mv/jyaxtYeCNcM0ms96F7zEiKj7iKhxH1R6xE80AhvGKteUYl5lcU9aG0JwE
XllTdEKDW+in8vzUHH3anzULFvm64BguAFc6jQ+cCzX+aut84xdAAMUKTvRQNk1gAb0MFIPseQkD
KolJLHZn7oty7aWyTpijH/5jqoWKHzlTj/qlUfPirBwliLkV8DzAeoL4DsGxeeQmfVsOS4KAfxvX
ssE4kGdckjhsNSh4y9uEFO/mFcxommfXGGtSJ6p95DnM4AflmW/AZs0g8GgO8h7nCsmduZpHuokl
biuNApfqk5bzy/fwPO7HO+qWSyjklQuhemAN5iC4SqAB9C4VR2CQIyoXTPqE+tENa+Z7Sj36rq7D
IsX5E39/toifIiLd6qtOa0utDNyqd0E1cQiYMge8v9h10a2bBxNjwFJ684LyYa20zOkuWUUdJAOy
yoPy+UnCGIleS6ITlh5X6awo1K8ruLK3ChpDo1S/0WC/cxg+dh4xaQKO3GU6fyMmjBIg+VBXnlyw
mwIIdNkU8lNZxTe360AAJpm98djxVzhScXI9wCJJQOjxRhwRPbDrzJd3ZbovhTDivZLhXaPignGs
sK5xV0rcSM0F7piAPk/yyjMuiH+aBckhh3w8FjzfdC4zfzV3+FWTHo5h3BIw2PRHnbqwCmYC54Cw
fKCF7lQBZDhl540jBaSrUpuN6ARNsfKb+/mF9SnVtyZ9yN3rOGqtMVj2h/MLEErz30nq9USPmH77
3Y+J7ZJbmAglMgM8K7FI/65BwAckb4dcgjioKnBJvNHqCjtqQ6hfmdAVqwOJFdi5W7u6ZIyCmXzS
QR6QK/7OTPrnxJg899TYDkiaR47B/qbYuqasLhpNKFhBZLUs2cO49YlAWIKbd0U0Xodu08uyPx2c
N7lF0hQY/8wLt0cRgetuFnB+AYPJL2P+0aVG6Op30hnGfnYyZlD5aeohCkljkMDHd4n2bbKArMGB
W9kYUarx6X4U/Qwfj8KnXLHeBkPFfdvFPD1rmVlURKm3eTtCm5I/2NFnrnpOa1RDeZ/K0PwjRAzz
Wm0qx6BqqE7mgK0vNooa1fSN1SMeZ7WOKYk6j/TZailTvnfAFFGKG/jTtGPh4FDl/Pt6W41E0TWq
AsAVmj544br2dwrjDVclYndtuDp9ni5uMwi8XHk0HcdcGBIJ7qpViaP6rbTFL6c6zvp+opvxFUW2
F6qcvvBdM7wux09llhKzCxqQLpaIXM86I1xVha72wiA3yQp6Krk9Apo8P+oMBIE/tzNX8wZ2I6i5
tMsTOgEpNQy7Eld/o0TJIuPsCUFeRHvju7uqanpvZaLcnE2GBHfdCr2FWCu/jAUPl1q8w1Vo3vot
k/7u4KT8tZIG+BEphyIwF6umj+bIIQpEpZ6uZOIy52egZOEz5vcYH+EAsoWe4MwbMRiEZypP6WIR
1h4daHtRNyDc81hUUpHtd+WdDFhvVgrVgwfcxogTWuN1f1chbNANxBlH0T6Scmn4qQkB7Iuj5Z6a
ZjNL5IldkzA0v4b9Slee8EyAG7Mjx/DIuBhbzWV2IAUYhXoiAvPV9h3xtwSXN7he2mgcQE9g/ch+
OuGK4SM9kdbd9q97VTK1k3zqQCnzKOgvtU4jgPCp3A/4+0Ez0Lt+L8JAVA84iEQMKCSdWITwVNkt
4NwBuz4nqeEWpQ1clzt2LXwaohrrl+3CnT6ySt7kVZpvNIaMCBKdrAwIQB18i9hmf+yiQqBOuApI
JZq5UNdQ5+WszH+8Bj0Ql8+Gs1KHII+JeLNSu9AunTdfqIgHaMz1IRP7cXiZ3IGidA2O+yRf6S1t
jahP8ZcrEgDSi7TCHfhf2vGKWJSoc1zY2H1t7fcuuz0/bIQEM0gJDviFbbg2ZmI2R4p2VAdjoeSm
I93KtcdTQKu2k2j2tgIa1nSzBAyQLejW26W4HnvHxPAesgkJk+pRwS7pl8rp5iy0UhlwGQJ25A18
jB/1b345wOpRvNfmhHYbu+Vym2uM6LBv5r/LnwG2/qsSRawP5GyvJChYnfQvfx2ARNV4K0vg6pyJ
4eOaXlJFflhLQVZvzOOXfaAn0TjeNDXBmwOrSvlQfgPMtAUXfgy2iOsnng9uUTK2PCIzrZHYdBX+
bdTeeUL1QGdBIVt1y+kd1rB1zeMhc+PXDVJZ/z01f10oAW14X+BqJR3uRtilG+w6rYfVOpZ67tB+
+jEfiIarKEFCWrNcqnOMoHUUOMgHYGg90HEPqHJrU53kb7YuyaiRwdIk96RU6KdJf+FuGViI8n7y
YfxJuDg0fjWgReEELd1KJUKHaMHnqPHtoTUenvv8EJLXIrBoF+Ce0910fHeHLdWCrkSY1Guy+dwK
vjQ0dZ6CD+0KVSzJ6NOrGJ1QNRV+HKN6cdqvpAw+f2f+p4z1bmbUgQFEJhF/xPofMLTTTMucNQUf
76pNFpOi5z2Zy+oeujueL+BMUk6DCyP1UuyxXiUEBbRZed1K+O143RmdtAxAvZVTGMQ+CLGEIY7L
0vJ822dyIySLjzYiaooznZdR2IQBpCMgOZVloACNeD6jpC/ImEy6lPVARr8sioJobuARa3W6ySob
Gx4WMjpYRCFLs5TitOMHqjRD2jO4hOgX472215aem1GdD1wf2NJMcDVaKyx6tiO7d1IF1KW5F67b
jG7PMkXVtHLBC9oPpYg+MlCDAb61ZUtvwjZMPQzb1a1ER8RvAhO2rrBwMl6s9Y0QvCb95q5HWV+J
v0Zhn2Q2UgR94QJ7k4PjoySun5p2Zb3UMGrqbekmG1Jt01S+y1Tn1AcVVNhDXtdCTLedQadfiptI
sWd4B5lQgXTwVkjC867DPtXyY6qJ/t3CG+KfLF3IIsRTcfzq1brgL6qUkI4u/w48IlVqrHrbW6EV
psLw/4265JVRb6p6NEJkPoW7ih9A2p9AuKWgg6e3QNWYxI/peHPYFdtOXCNMO3utehQIeCiNHbRR
DUyvKit169z5wjVcfKQioGQMzjhEiS5BXMJgetMv28iHztOc6y1lpcldULbTWtwwkc8q3fRy7z9l
xoyvpYZcnZyKDKDHMNkNqwTf1aMgKtgsjzDT7wHFOHRud7I76OZD2p3dngyG3WUMSk1wauqrEPLj
mN+UtNVfAIzORTANiuJygCmQYyWmXK/c2reC5IDefD9FXgszHFiBrZ2p1Vtl4hzoFdR9aCLzn5qK
iHzvv3ts233Sq7wAhIfpfxCbLrDNq+YDiywOWD4X3qrIhAyZPt3uZWD9suG4q3uPJwqWn3ITeprE
TqDB0LeA7ayYlJ5R9TqQq3nyhPaNp3SRfZqHYMEqbgxzOC7sS+FCvA4MQH2yhIgHiIe+Ed8beNZV
+VfSTjOUW/4ina1kLQLCHBo07iha7kQelaqgPhIvpwQou16Ozgl7RSPZCVy4JrI3L2LB/Gnrkiyd
LJH0j19Govs3Nd0QqU/LRwRdeCKYNXEYMzDvxcXfVwxEEu9shPDdpH0ej+rXUPXAzvqydXKjjLX0
HLVXTRib7Ka9O/ULxlrzaks4sAXdP4xrQ64aeEK6WxEA+fnvGWfHt4RrChGB7Ic36tQQl/DGX4F0
eHytxi8OTmkJQ+j6YbMKsP9wvyKJqHapKRV+LM3xDEX7jaQpQ+A6IV7wwb82RUeVgvVADGCUva4k
bsIbag3JpByvUvAPXW1ktqGwwsO5ERUMTNx5HDSmfkQGBlwVgxXKX1770alq6CivdZVE2qOkqhJL
CI2rR38NTIaTHMCQpGuFIMD6in39J8XgRgHgQX4pPv0j7ucFFbMOcdIUzpabmHnssHK4OCeFDsfK
yhX7L7tE5wx+iuQY1p4GoZMHm++sKf5DXBmPVDVrEVjCtkXq2PFCQEO3kzwyF4fwtos3r2Rp3OZC
FUfPi979uu4fSUn2VzrLfmVgF5uyL38V4hQ2HlkDPFJ0wtnY/20yVS96TfHOeLNLSmiB6sJsJQ2s
R/gAZ1zOb/TjSVKLCfbXogAlSkNEde9CoIoNHueBz3d0Iz5wczrCgRDsoh7FmMrcVV/f/44bNyoZ
z4zJ0e/NT6sn+DA+RYyMEZMzySRy1500Ima0Er8DXWU7tW+ITDwF2kEOtMLOWcElsJShUmwrWkrx
MndZvGsISvYSyBZuJ8gzMvGcj2b7C2csDLgm/oUWxrSYd3UVO5/lD3hpXhH28AqPCvmQoTd6PYvx
t2UFM0lHT6gOfTrWSKE9rTm3fUSSRwSzC96/0B+NwkkJUrQCPKirGd1PVNz1Cws+o5Z1RDUrRaJv
YhSdV+/3kbDfYUkrfqoYUOl++9T1uyFB8qOublRVpmPFcb4HIgU5KhLn+jeb35gyTQV4B1fdLEN0
NO1TXlOxhRhTh2DQtW/XMFCODxOmzmJ01bNPiJGQHhjC/hbStgMMzQehsC2HHxlC0zr9D9SfIaAB
kyb70D0cy2RDA8qmDW7BYW6XA3LYitNxfJVt6O3eHhKWI+ced1jnrgZ0hjZdi9ZC4k4CyzX7sQCR
IDrtQMMC2cRtQeBFjwDtkS1NwACB92PsUcf4MDXdKfHtw9W5vEkw4dzw59LuwSPSMKQos4aIR4SE
PHndVt1Flq79LnzTFl1S87GqFx8xp6UEoUGHnwX+s5IBqEe73pe8AroqaVXqdDeTnGK7lhvr+Gng
PC6ybPvIl++oiD86JmL6tcQpWgHfXRZeBKZsW3/lP4H+AjdITpYqmvCiMIaeCuCUZ+H041BfTc8I
RVBS5GGxQiTuMfBZG8VEA6+Ik52gQRjug7Iw5cQETkILol9QuhNHFxV7GZNF26eWt+rBla/gY1NO
L2aG1tm8ttm8lhXuoOWxJFM9nE65KZowVPJQOfJXaywzLVANa3UtCXM7UqNqP5rfL1aMdZzu8BXu
xLl2KmIbD2BDTiCY+BJJ4ct+jS1WQGEomH736gSCjXXMaPkh723AVOC7i1dL8V/JpwJwG0DY4eKl
mxF0/j4Z37xEVr/3rdwbDhdIPHHBSiS42KRZ7Rx86YnBdiYPBK632EdgRlAyWxOjVUFKLIpBaP6T
tIpbAHzRzCIGU5kKVw6upqpzHDjbDgi+1HP0il7FPKh+thgSa1PvMjhz4/k2BwaVhsja2tXLM8sl
99pCFpj3lq0CEbbVxtCXNKnb5CSSelKtOjqYoI3J9y5rLIu8HTOdJvi1AsSRG9tDadGOMnHkw85W
Oy88X3A2QVkMkQURh4zkHQpTY++YR9JiVwOrkrn4mVJ/oFxp/Ce9DE2oL1aiqQvXao99Gt0RcU+r
UdXEtBmY2uBPY5ka9POHyjnv9UIRrgTMQ4+Wq8ZkV3TqlLGmTSckhLa2OnTb8BmC1raGGSDWMJzt
NKOXKOC72CrLGqMR20RkHYOR8ejortJwWFEY9V61zlI+PAckLvGxnxk2bdgjCGWNietXXCqeFiDv
CQWeJTlr0LFBTHboFra0LP57s/Ex5OFfz2Al1cvN93AKrsxTbjdB1z/5n1kuQO3lwHqd7r+cVgEC
iT9DGWbsiVhVtPNq81ZG3+PgQyLSZFVU8s/FCZpnDyIKXZ937s6KVaYBgzq3LYIQW1VV6RszVUlA
Fre8FE2sxSoYYMHflFKpTzcS9GplXk44Z228w2vGR3QTOdqF+vWzg+58A2JIcGn55wNpWA/rgavu
0I2JOY7yspTebHFu0pRtCi4R6BpBVNA/I/F3YW1fStQ6B9IdZ2mOWInPgEy9aBHvv4oYBPHWdEqE
JVhZzRJtZgdcGcoN4Er10xtU4p2XPNTMc0l0Ac9g0yGVN1CXc3QxXNj3zpZLddopNBy02y14mflH
yGn+ED/NO26nMrxgWBSAu3S1TXdlgj5zncrxPHdRt9YN8vcf6jyNsv60SXLPiUWWl9Mjrc/WmnMR
9aFnCDrN2Fmfed5+pVRh7lINd8XqRK/qlO4G8qcokcBWgMFTHpwDo6Xub5gATLrvbRLFhJFCT0cL
Th0vhnk+WRoxA1BD+FRv79tfuQYw2DP+tfg/zQ8SMUy/9LYdWjPxFneScUHPqPPF8mD6VDcV74s4
B+gGLCmda6RAfjQRIXsltgXwDP55yLqio8T2W+tC8hYRXJWKJUHFRgFMUgmpXyvDRfsmJH0a1zjB
AovlBML4ObEO4c0H4GlXuluuE6a8DemKUpGI62Nvcn0RA8Dk2cfDgQImmi0xgo36e8W/Q9QWp8Lg
FmRHToU+OgH/tu6gEX0tGBH/8bMYCArU1Q9sepW5wFjLUNKA0gOR69wpz4znxRm8Xq7KQjHYofck
sIlpRRwIDl/a+4xf9zoRz98x1gyS4QiVIgw0LoHRiWQDQqVtOYoXL7KwlLxgZihPlbAMzp9vIeqK
qiz2qcpBuXcpb5DRd4ag/2NafbvuedmsrqXkeDNvVn/WOQqHkvk6XROte8/BMy3WFNwwPk3M5kC6
dKpeLH1YdyVC6lspQE2jz8CjviNzlT/xrBwqngCf8gW7DfIW4B+cRlYNgfBRcTLLhT4L5DYd+LAn
7/k6hK2atm036zUF7ZYQ9R8h2qEH0OzjNziFsOumOJY3OxQBKf4PhUrNLiDVcT2bQAtWLhyM7AJ3
x5LVUo9ch+KN+hDSv8czhXsVed1W5D1hrs3zNwvPHoeQ6qYRPqazeCjHvfLE3SLVao2TOeus6HhP
n5neeaGB9AvhStev5BjcvkF7aqO5blcEOWmfwbLuJwOMcUQFpn91lNMZ6fXYCxWwWTKI1wnwN2as
qFmYfq0i0lajwsCySRFVrHW1x9+nJsJpI3MeUkYoCAHUWmnCNwoFh3bdVLU618KwNW5h+Crq5NLL
HI3hU3CNjeGuzMACor35fKrwn6YGtfTaEPPVWqeh4Vh8D9gWs7V0hU8FOYmB5RovbiNFK9QXIRWf
3ENlj1iHV8evKPtwTyfaFEiIL/2W4I0UojxCqOsB+iK6JpyU8Kb8EnlYTkiqo4hFnNMqcPjBrWEB
HxlwDQdOB7Y2Hgi2ulT8npFfG7ZDmNJXOcrHRWovh9JDaavtjTGAeJlWlGOi0kyr2dNBrQ8S5C3S
k5vHsbbbm9Zg45V+R+DPNeXJuXfT3SQK7lGGEyxZ5u2WKqvH5lGB4zk7aR2O2gFVwoYpc2eKFO+N
zPpwZrARrRnmfbGHVKSHyLJhYiLajIs46yPeN8hPKm82n0xyO/4zGih62CFb0mUv+0H204PxIWhr
gsVkBmHIAZ7q/xxhVu/u1vTBAU6mt5k/7gqZvStfuinph+yv8EZIWAcsGqbPe1QG9Z9JjTEt/cY1
uWS5dUVkaAXUvKtfjTv9LJGzIibsO6EmniTDpP0J3/iY76OVEfXLCb3qra/gg/sQXezmJAUVsfM5
tbhgr6ocDlvHSyosbCVgk5jnHPzWp925XgB4Vlrq8JS4JjZJL2vXsmY/OaxAF5mWU/xtjrRUWP59
KHsAyehj50bcyNrkVpuDwgScs6JN9uE2wefNZrLE/fUjsSucTKezmiBlx41fcT88LBwiWelPGJ7s
b2cgN8w/EA6/vF+zFvJ9QtoLjt/U5VE9EDBRG58mlC+Vo0+qZxauCMLD6uI3uWcWOerQrQh7vWI2
rVYHrY+jIZc+QdvZtpyWBTsyu9uNUayKNWziEgRlI3ieYvEELQ4FFPNRvA9CdZUYAmtdbJ9g4oPZ
piGsvbnZDbZItuPLEdmsqm59dSlvkgn4AyRfxRV58iDnfSe4ZtA97rNHnk7KDFrqKLduoDo48nEp
ytfURadbYyKFMCG1gzeRqJN7/P0/lzZyzZ7k4JcDs6EktiBKoyvTLluwbHy7CxP6JqvFKm7BZdlB
Y6PBlR5q9/g7bgPdcXHGH23sSpl+F29Gq14/8pP980syqdz18/iU2QItlHjZNDQbyy5i0HWwyF40
Jkom2/jRkhMz6LUu8S67fdqqjalRWdmjPXFRyNkFEDOwbVMJcZIQxlhvZpp54pZxAZn6C4nj1v/q
jtnwjj77j9CwBnWm+ZgQc40RgEoD/+sbHlH7tS+ZEGDzMLL6Z0tBIKeWfpfMTGHJ+0qzQgvs+mwG
kT7bwAt3xGu3xxMGbBn9W+t9xNaC9iIq5v8uJorGGKFIA0VAWPVtgVpkCpys5/oiN2yu1SkCFZb4
qapBMOcvwLshCUqdrJeIe17EPy6DZt23ggFNZbeuN5rpGHMQMsnLDcl9amh0vHNJ2IdZXCubjgHy
O2B1go1ofBB6zdruftcf86VxBlhYSWdBgwM+eKWy1L/sILs4Y8mXET7tIeITh0Qph6dG0YEASazC
Rnt1WC0FAaWCchvOaw5Arusg/yrzSsM2GHKY0NcbcmjlZtlGl+U0S3xsRy6wuMmSvdHVGRDRdgwW
7vJOaMGEDbM/m309+dblS1/dp1fC+NhyRQvB6emm5NwRB7ypWlOPabEtECTFOrE8Z6tE/IY30LE1
uyothDR+1yvL1CRamJwK0+5HNKKhfonHxCLKb0+Nz+9OLsIAZutkSS2QWQFgoDScz7ysGG7H45vc
UIgbL4cd1iBYW/K5Rg/ez7HL8nUS08taTeD1eJngXGi9qldolYOlHxel3ebuYJZ/IzPb3/yRxrkf
gjx129ZPtTr9uSzJxBetF5l8HsjOh5lHiGMFOQ+s+5e9w3Khb6eQr/EPrj/S2aE3eFAxWbMTis8F
4JmLmQYITF9DM3NGKnqsDISJkEJL3J55qMrkpFKnSMJKeuLVSn2SL50LXrqLmout8PFMsx+8+cD3
y833pjYrwko29u3FJ9kiib0f6zn7h/+V4zOSlzwtt+zYze18KHXLy0AXxFbLhsRNI40kwfFg8Zx0
6vzJA3v6dNnImZUS0hq4SfvT6/ownMOQb7tdHirWkCpF77a0BAX1gZkiQJ6iE1C6rts/6O+PuYL1
x5vsrBrENAOwpvtFfGzLbjYYLkGHtIjyKcUv4sth1E/lofU+Cr2cHwlO5bLuSl6aZhOwDvoiqGDY
AiufSepo52fphWkTDzINXU8CKMnFtxsEz3x+xCnSHlfP/8jQ+1AF0C7Y2hEp6xhKIhIQLUttQw1m
q95xdNKYStdqzDpC2xONWrRKqpUclhu7ezg+lwTejTaoQaIiWjqdqUNwk6JxrmVwzXOEIxMs+KZG
r5MTRkalCUSrZ+oza0J+t52TLio2gkFrwfGauNek9yozzGdG7KFpHDNKo4l/ZdNGXPfg9Rc9DOV4
gEYki1NxgLkTSGsGpl4fkDkqFYLjNrhma6w9egt47efGD48D/HXo/S1KC5OhdmXy3f26xxPliCA3
QPRpH4kAbrw3bJJS5Xso/APGqF/csJ1VDh7qpuAK0td4kwecPDMBb609oBKt7UQGtv6XNRutxldG
cmUTGJDTNOJF3p+nPjgoNmbu059nNbkNzeIyh98V7ACXC+LibKUJ6Buhz2dr/Tfm4sx+HAajLldk
k9FHAxem0VPlLQkP8MhFN+Xe/XxcJqdeiX4yvvk2a427mfTiTcHyWENwS9Iv/FEfXxJuvmzGC1eT
zTWhgpuAkgwvNxoAQnoax6nW7YEHLWWv2qq3+ryjMM+agNASJ3/lvxvx+tv7f/ucsAaHqWBl59ti
CQZuU98LN/OQEGqk6hXGvTAQ2I4DGjxKpH0vHppIfhhDcP1s8oIYsvTi0XQk6YvrHymYKBhXu6QW
qVS/ppswlzIhJjKaF9QP+ikix5sgzYszU7eGHMANgcHBL9rZfGpi1yw72b/91mCaut7F5G3M8bdB
A+BuM546Wr1dnQiUxQJQbMDhajgXdlPB5/pO5KpBJLzV6bLY6TNwThx6rDNkpj3wWnF6RlMCyIu0
b1ZdQlCHRMxvzAN/6bIGsXGpAcXyZ19DzcRVjyN/jH93HCaa1YXlfiw8lDjfpui4Uqdg9dWPo4cq
ZlrxEOa4jFloiHV0xJwL3fnvkpJa5eSlkwDYm7ermM536EFXawjvsesyCIMYUDqzEKZj/n0S4iM4
07+a7UNO6z6mWm0Hkx756rkfuF3ZQeGyOyaeXQz1vMk0/UNJrykWAtckyKIqZRUp4kFID7MOGHuG
8LHCzWJbJU0A8eupPddyu5nZKA9Oip2FzrMjpnRfGyYscObAccApmzvBAmFeZuLVeNqoiTnIB6nt
J6PCbW27LpKG3KZ5X+fYERt6p0XURO4LVhxs+cRfdkh4E+1l+qpMJT9l+b6CNeqPD+8aRw39tv6E
ZpmhBvTNOL3h5o8q99Knsnj3pOiYFAD2it5xu1z63sJC/zXL6Z5nbT309YGJ/4QMulcQyF2WHuk7
+EPgcqL25bGC0bF7KrBvIgCYktPtGc4E9Rmf4oRCxfIv9FBlAJOAsmWZMyv381e+PF4123OWjV3K
ALLBQq7Vlx/uNHkzr8Jb0DGWjGxm2T9XG43BwKcNTbTHZxYXTz7UzEKWYesJSqhtng4cFOvWYr9a
9dbxPogCtm6f3KQp5UdBywbKWQLgUtWwdxtrvsOWlCvn4nzuhXs+RVTdfYCuGcVHd3HrR/AynRct
dBqVTw6/TVMPJkNOZh5PVUyg/VOeEFMvMc1ohG1A1G3C/jkX4Kauz3zZiva/8jMVhJfvgJ//YPSk
j6vLN6WC3/WB283XNZ+CR97tVK4ZGdbbfJRtolFAQi6SJBQxVGtqJv5axXehGdaebNYipKVJVI/y
AruK3KP0tj3zyRpZVS/BR8v0zjF80lwy8WRxPYQubtmnydsgGklyLfBRrXT0jSD6Rt+fwAJJh2MS
x/oXdnbBvCo2H8mJzQAPsHeQBDhFY+QkHCfRBRE7ASKnP0FaayxiNTnSqETFCisvisAdGPf0Yw+q
xh8oWYaFOgn9oHNVGiuZoZl+EAW4vING6nIErhoxp968omrK2WztvGoWdZ3a2CHXGVRr9poOcbpq
Jkkz6I/dhRLKzM2lURslxJfvNA46ruqRrKzuUqLFybiE5AdOMA7rz5VZbmoZnPl9J0dXahhUZfEs
vFCtYqtdYImSj9EDy8Lj1s3wRSNfx3jcfBqpePbUKirJO7WJ61wXfUrgdAgsiUrztT78fEelGs7W
V67r8pLbFBiEJ/JMnBsCYX90NCZC+TqlcM0+uYlPTXAq9vKmbXGkgp+wZMIwn+NUihh0BZkzUCVf
iX7nmOK4m+MXjkRS75ZyU5G9zSRUerTXB40lAyqON26+7WYi1HLHq0wOMr+0HgnxZONDga9HUt4o
3vJ2O9zn5MNDsZrafcR2+cHoHi9RKN7gE8HP65T4Q6Z0pbTrK974fg9gmyuBF5+HLt1U/Z6L9vQD
JBTXgp4gGjVZAdGtGacutNSQELpmd1XHTlDGkR/sN6h5FZ0lpfm2jVnX92YlFeSsYcnokkx8jPtJ
opeoo7GK+VyOMZWwp161eKCz/GWRFWX1ivXcMu0cnrodQ+TY4qZ3PjDG4jujfDziJPtRxeSzVnsZ
of8YDNhIVtwRgZ2aOMmdVFUHcBh0Fau8Soku3Spb/IDYVg0m/56L8h7Nf2WW9LCX03gLa2+4oIgW
FrOKL1U4BrAUOcWtcxtRPnKzHBCeshJG1ZavN+dFocyXT0mOw8IMpSLQSf4Gg77I/dS4hpe/ITox
3Y9QVeusp0uoKL3Nnoz1poot+zQkdaOM5WaCTgBp8EpLFg0Dnb8I7FW/5gLsrHOhksY7sVOVWfUN
8nvm2WXYi+dDvmqr433fYj/SpkR8TymwjtlEoz9yObbJY0nr/l6+jq0ZyMxZFYlCTXlzvbUSFRNm
wPobzXKoC5SNos2d/om/0K9/XAWr+9KfVDvMi6Z5WbzsJWy/5hg5wHOQ6RcNOUSKCjIew+cuwvY8
tPM/dOreHdstqHZrqClMuh4mD7kV8yH+FdwYoLXtiFQUFi79yB8fbzisFFB89RfvlS+tT8Ihae2r
B8FNJWhK+oKi9ggVnmsdhs1j6HxFLUgeF3TKfFJMHpVEk3C05YD9lU8nSGJXjSHyZDtYkpWm7Gr7
qvjd+IG4QMTpC04bDxUS5el4YD+TG0s0cIxG3gmrD+DRm6w2IxptXXjUPkB2aGjdOslwoTDhvd+o
Krk8UlfIpYau3OOcSUOmuztixoPzTUSjqDRNpvQ96NxSW+i82mk52NkSj0LAJFL2RSTxG4y+KOt/
HPbG1IbpV1bukbcMArMlacUhjkHDS53QkdOeHH57cmzFLIekeHQXQsITh57cY2qu5FOo7jLpvOc0
96ZKQQb5HZDtrzOlS5k8uewn4ZiiBSxrN6jdMUNnR/K83s6rcrPvkHijT2Q6M28IIhGOBymo1xzm
NPnFsVJgsUYDKlyHXkqPRGX1JDBaqiToHCypNVhaSHpXoCyTwKOaU7flvwJzJhWP0R7kZvtd2g9D
ME/FgLD24D12S8RUiwssDEdcasbT/E4k0bYmku89XePRDloRymtBw71lItt+IbC7orSDuHhqJf+a
rJo3asLvJzwbPApWt1jsHckT11TEPdHCZWF0nWpwE9X+WofwtkTtsDgQigWD8p0oEJGjOHMVOleb
yYrF1gitYaPrPZa8BgQ+Ns/t6xM332Kvz95Qyot7qc6WqlYCX/Soiu7xk5lG1AsiDc2x9PnwGTNY
THWx4PSiqNm0bfxCfHwyWgDfXWaeafA+17eI61O0B398Sla9KwDZ6M/eZtVd9s5WVmwYC+U+WMen
LYqaXlr+4fulCEruoQmYeGqnGff5aUYfAqio945mCX2iHHX43L3RnROHAylBttq8XGeELbOm1StR
doRC655cpVv1V7mSnvq7+KjlcgobkNU4xVnxhscsS9B6ftUaOS4H5TdXEB16ZGVp8+GOzhH05eMY
QpeS1oIsjkUzKz9Q2htYTwY+a3rPbMN2eGyK2aBIW8fE7A/IfxKEaqh6EZsUV64WxeGzdfUQ4nYp
ewra0HJpWkDbpVQeO+uxDBN+QUgl8yO3C9bBvAHWGZaFtEOOndvwWO+N1SyvirIA3Bs5HIqH55Ce
QyD1oKjT/0Y1VLqGYWiYPps4+GPCbt/AFudaMXhzJZT8PpFKGAZe1He63dPddFWbcvUSne1wsGY6
OY6y01bShG6P4IKBa32q+Jw50PQn6pNzFK4lc9BXfJFHse7OjlYtXWi0Zs7YLnAhXtu9+qQS4Yq0
lFeRTjTlVUjpHOKdq7LIxd2GI+viHFvoRTGT78BTVXrrBWL4fT3jGkFzqKzfsSEdnSfxjsBxB3L7
f6XSeMlacEVhAkcwRgu0UXe+ijJzBeiGIVPFfLS0wkxT7I+ytPUR5TEeMXrumG3PHmXYZJmYj2qh
i6AggNWEuW0Wd6Z03bDgN4YduPXjUAJFaVKzla9QIsbeLrYjpNtAMeOy6T22kaXCzrOeJkrWHzlg
l3AnJQWv86Ee+MjgtMcZJRPRcx9ck/v0qo4DOwI0Vprs5niHGaVylqM593kPYYPYhq/UQmJE5UpW
HNS6CcJw4xr0GqgBv1Yp+AwnPG2wUOfQvWQ/XIn5utCzT+FysSfmeA6XvckYBPs2vHupNoTLx2ah
piEDXcAJzBreC4gJhc31wqcgChfAqDu0kjfO5KtnqxIiZ+ev2lF82S0ryi94g2QZVtUUTfNgbTgE
2xkIB80A8wX7CobYSML49psSgGgUX80HjtJxgLkQpuDMImPp60FVhb4L9BKqcxHkq4xEmb6t5IIm
Os5oCN3xhn/5fV7xMK801JHxHhl3z08ZIsGnEz5JhoH3dTEuHKOMPH3cxOthcAuBo6v6w4uUQxNS
GF78pu9mRwVqAIWgs6MWQsEFSri6lKLCct8L18NGuAoE7BP9o2IDWH8lwxfxYkfnhf7bSoUYiyd4
ZM8xknZFwveLvwoyGFluTNA+uHTrz8C1ux9D41E7coEsp9RNq1I56+QY6h4yHGOORWXXlpRGOuZm
YTycUQp0+0cjZLqyvbHYuDGa8m5LDgoJC34wGlXu5IJPZqE9UQ4oKuPFRjX7p6Sfx6aqvjPX/94T
T/vR0uyhbnpSgpd0NmSnZ4P5PiVZWOIPZkuCas7qNq5syg00eRnrEwiHD4VBFvOULywUw7heNGh0
a+ri3AhoGYqt9pw4gM0BBd5reoERayAIjtmNtFWEKgLSWhvSGAr166wK31mENcetn9KTOrnHq5fh
ay7+SoPpnIFg/buoFuzS8JbfTub1LiZawKWPcDYYmGUB6/auNCyA029NKP9Rc6yZhvKPSYItFHOp
ee2rKyp17tAApDLPPu0jfGkJ4gegIU5rlY3QWduMbB8xSJLeafonyHSSEbakTeH4Zos7r5Y7rBCQ
7cRCLlTfHtSgJaUXskvRIZNw4A/LCpJgmRUnE5Fv+KqlEetSqoCXGlTz8TAl9Q5mmYX+51YVmqRS
n7yuPQ3Yn3QjXnGe3W48HpF+rOsxK5u49oZMVeH1y07g8CfQGttIt+l4eTZEe/7GMgK2k0BJUZvc
+wLZ6En8NZ2mB9SZqGbMmmTV/6/8HCiK+rEt9eqkUDw2in8pbF1WpKvIiImXB5IxQGH62nUEcyVd
fzJC5h5SVHUBMeqPhZJ8I+ef6D8VFS9u8WoB4be5rIVogf/3Bfsf24BknytjxcbIIG1pcViMDPo4
YXdEYZ761SHpcHdgdPq6Xau308qXya1lctKpZNuSvV+WDxaif55DQuf6J5lG+1qmpkNV2M2RVpRw
EWA3lat17ARnxYdxgF/ufFGfQR0iBSMcMTEroguVXaYPG+H1VVe77iDyp+AKyMqjz4Rn1AfvZ1ro
dEug8zLs6uFgZpQcreKU3/LCr2gNXDLYzGvBMyqes+hYVvfxq0uoM0Odj99JcLSSthzt8GeJ8071
oX2g9Z4iUdHWCcU+0c8BEjBLbBC295+vs5rRm4vcpFmWUFFRyr+q3Hn5czqm0xQ4PJqGl8o/OHmF
bSipEWThmu+budSUjSs+ev7drC+Y9riJ9JUV1Y+k2SLFTPesNYMxZTXY37+TidAJyQAUlalVBFle
PHWF5mpXK/YLDEF4Eg8nAjiKh0fnryteEgBz7VjWl4NRYPUgc0i+fSOVCug9uUpvz4AIbik3eE2g
+Tyzo6rAeuKE9uUVacJnKiZJQwdc1eH2KUhA2AuBzcRqdqGXv5xX0S7yXSLdvI7vfcIIbU8503Li
uzD8Q0mEqGMmGvHgzibjAb0hfDU2kKR+BaQZx+7OcQ1d5K4MBCM/8ALvkp+9cTMeDs+A3mTSAMmb
SOyLDbpjTkO7guQ4CNplwlpWxit+EjQ66+G2DKv4PFtPGWmG/USPtYrbsDE1RkU5NGbGrTk4HXV/
9qYP3RJy22OxYxscVRp8RGsTdVpGLYgAT4aTrKNvC0FRjL5zQ7HcmnEGWmJ22lV3d1FZ/ZRxYWJ7
d6WTC+LL1bvRKMD8618rhF+9cA16nL3FTIvTwtKKfJjyF7fHcXytSjoE4oGsINRpmSBWyN5HaAnT
y4DAAe5GyjXJFd+MxeWfEfj6P5dStgN0Jg/CkfZ5IVhbhJg5J6wNr4U/YqxQ+TNCahDsoyIPSAXm
Uggqsan+cGanjphxP7Hm1HaCFUZoiqS4vKjWoxQG7v3sKtOu8J/U2VXuHrWeS/02voYXJBxNYe56
RcJRIcgCmg1hzB3k2JnS0FkLQpXXkti2+WWeg/NgVkyyBLimRJo3Hwhuu067PKJKbyzbYB/SyoVz
G+xFxmCmFjcsgtmePnmI/jby8UOKoXugXpgKkFe8SYrap+nhgW1KPRpx+Oj2yErJZlv3IGu6POZd
kQIG/TmgLpoJTFkW5cpS6gLbZo1J/+uhXe/FI+T5LQXSrhfFDnutcad0fnJITkBrgL3M6yQb9cuZ
c0kPs/ncu0U6gwgBBdrniHfGZsyNd2ubdFs5q7/ihE8MLa3A6TcbEhANu9tZ/cwYJ+gpdZEq4th7
hLC2b4sc1zHZGtEW0aGMBAcin4pjgI5lr4TbKlSxFUJSPaOONiANibxp2kT9ys7dqwCmcJE6Z4qC
fww4lQhq9lyNOwVJJq1U/FrM10f2/T0vzPkqrKT8ejT5h9DG6A9ZiBMhWjmH2x1GwQHpxnz5ELgn
X79mmYuZ3ZUQBG1tLz/ULL01XMTkquOj20+eByPGULEF+ykqTRZ1+k5o4Hp3tqsyF1550wrK7bRW
FbSq10ArsptqZQf2L1l31Iunk1C+h/NdxNfzJe09oqrm/Y/ha1vVbzQAvmjgl9t5PmzzhCze/MyR
rYIAnkOPAIWTZB7rOylLiq+ytkKLY68+qZYWmnowoucg4A6rNQdEc2q5NLh5ujj37efQa4jeZ4dO
JR911ynXsoaz391yk7PNsg0u78yBrl27sDasWTvHDP8Lxka8LbEeIQr3N9OAQJfQ1zEXgrTfOCcq
ol1SjlAfghWOnqbxr2MIal0Fr/NfwIC/fc59B1i9wiYSswsOms4ysfblqc4MWeS44ZY+Xz8fuSaJ
y2Os/k1MkL0mtryEP/Ttlc/xU5oCWMMqHwYVFPU6W00DeOkJgNHI6ITCFQtByWnClbKK/AjqULtB
5r6H7U4XtMGJQB+MFU6b5fqWKDkeYyryqS/HWBxHJKoCIQhviQngx8Xzc3FjtHF1nIiXo/qRuwdX
TsOTSk+sgAhLwcihtsZbINqcwfEL2v8o5c/8fDWwVVhudccWU7DGr75kBsZ3XeOZBGkiM5QxfdRx
0oIE3LOVtWIh94ROQdqZjNKGlYTo6r+ABiqneZexNBVsWn5TMP5wrbFeiAheagMHis6LRlr7yi6S
Rb4OTafG2d9AS0J0esMShYSd6/z05OpHIGWJY0nTBa4yv89qdfp2rpxbeOl/4zhZHhs1hFdVU0R6
N9J6WLp3qFoLCOf+UHDQ46wTxWhBvDpHh/faqy7SonAUVXCHU1iyI/g/kjrYXbdd+kifDyV+P9+w
dx/dJ0SjRID/N/uhlXlcZ/4HegozM81XXDO/2OpQFRmbHghSReuUUyAGUPuObJBoxJYw5X9oyFrD
+pVWxYLJk7AO9Ri2JzB7f5xFAYkeX30rXGCpKOfpvBsJ+phVpiuopn6XSlZdFJS3mDp5AwWFSWJS
zQLX9qUQpYo8igtvmC5nIYA1mJvmK1jFJkTU4Nilbp3UMFeG1DeJGWmvHbDFkTo59IW85cePnE9+
KqKsP4MvNI3S6RMmnfJgXJm5ESlmOeXs3NHaWynvfWD7CBSDOk2HzqW8sXhrr6ooyPdP17cbo9Ve
ONt3krFL+7NLYq3pzYuQbVAmsknlSkOJWDEMLKHVOHrfRjXIh4hVCe82AjkvurfFTmibVdyb4f90
1Z8a6B4VYhasAYcYm3Ih7y7wv5efI5YjRlepXYhCha4/56jOpu2lGuv/u8exDqp7I+0JziGkPFtw
aS3kvrUvE1fQkd8qsW1zV3HFP03aA+ClPy+WoJt0/FeTm+uWKIdoML0si2ifqCuqQoYf3cgWMy5I
w6MvcKz+21YJkpOICzJbzCCaSQf4jMZayvYNKpEGrI3aIqs3obNlGTRAIu8E60YwcIaO/oAU/p30
iSHu6Uf6pkLTrhkGzGWFYBx234/Bj+JTh09YT9sxamxEoY8bBioC6ez3AW7VynvHoVVKuK0eClh2
Gg8iqQDMOpFBVY/6qbISDHP0Dn3p07IfXmyE9btG+fQyEbdYMQAOpy3iFf+0DRB5ICI1cuaMm6Xd
HufYgdAjgjz5Mp90U5xG0UByCLFefmUmXlkJVvzeS49q51iEBN9yPBhGIjSDZs4RHIUm8kB8o1FC
7k3wLzCpo16fgwsf8cZgFOkP+x/8wL8oN+d1G5KqSZo/XIigUi8ruEXZse5AXZLllHIpYSrsvxgz
Xd2WGX45V0xSGLJnfVqWN11Rcn6iLsM7av7zABxy1nWXXmBPElcS/FnHupMon3bekPTHuDP5bKWD
HcKp10/rIeDUrZPYIG/y0KaO4PEf4qIl4jcpsplRCU8w2cDbm5VdDxGQNOiBQd/HSCiAO4vf+Fhz
JcPNv4A+G21EGpkEzmDpIkJPgK61mtj8wPvBPxEPpydka/SYODFYr0pWtIpwCBWSp+xWzjLp59YR
TLW6iReDNt9rcCEIaIbiNeFUowaVNBrnvMVBx4QIoWswYAsT0T1QQH6/H9ABlFIl+T/eBQbkX3Ck
zlHTMZyIedoux/3Y4xzsSddUUY3alwtTN/R2c7JOzNtnrqCxy7ZpeOlsdn6WL6KBusOCKvVYqwW/
MQ5fcSegJE8l8/EdXU9ybuJ/cZ34ZqgKP1t7vfEM9/z/DcSumI+haEfEQOqXgwzb2UiSFtVIVxbm
RTIH13THHCLhCVJHIID4HX4DU7ILZbJXQaow3FKN9ejxtngNh0YMWa3B5wpAWdSwApJ7KLqcXuMz
0zIXJpvCd9On4BOD55RMUYijBf6USEHDn8+U5db0IDd5Z3qqZi6btqDJbDdXBayFLBV7ZagyAnfo
xuJmM6I9zRNIW3e8bMIUivsXUqTx0e4ZKxnrk/3WhPfj3xMoQoryTlleNqcswDAaPmdozatEfmUT
SwIrT6yOjM6spRSm5NnkweMTUrNzTRSXZfOp9B+TgcVcJvNyHT2wbzyEwUfhI2F7fkhpaoV74grR
BIIpSfpfCeuDlp7duoNeqlDaWJiDP+wlJxGUA0SXnO0xPG8hy30DZvDJJb5kZDiTmfsbws1e9KHm
+BkVwHV05byWLO5edfNTjNZlEJN7gkfOMLq6somoisaodOcpSkwHexk2EGAF66opH9TgzCkb+oUO
dUkd9N2Dp3deLTWBPpGg8uGQGELbm5RN3OWi+8U2ISmWS1Xi6y3ynPX1ywL1k6VqeKBNHOaiUaYs
ZCvQsxTP+vLHuOpbgWRzmmfdYrbeebqmqGJInTWl9/N5rviAsCU/n+q+drH0Xz9RyHBLvpnVEvz+
jMYBQzQfMOraHhbxlJ6BIEEVwimovUdbrJ0KUZJvsn5WFnQD/jwaVt8zO0ML3ENVsUVOhL3YF8sE
mIgjf9i+it8dBYINOTcFPAWUfWAV0IKUG434dn2M3rzpw7BpbZYjY4gc0jvz8U6BMQ+0KGDRtBBm
Q0CDGRxcSEyycpIGhhhiFg8/GKWMUcYLY6ab5/ThutVhuJu+SlV5lrF+I/1QQevguy7U0Ccx5vKT
iu0LTPN1C4xGA7wTA3Ehe20KK2MynlOMduCTgbAQjVYueknYeqGNSGR/8BsDXf4DEyrXjaNwGVaj
/NglgbErrt31oeSnqQK7KFcEpgDzc0pkB5PY1o+FdlNSa+WyQBBPYtXNqlEuWtBdDBt9/AG0n33P
6xGubg++5qyy9XvgjpMlFL5NpDJAesCSJV2dKGfHmT4y/Sxtj9pLsqA9nAZa1tsds0T3uKOwZxQc
I4mGPsiQoD4RcjDCI56Uv0/NuP1gCVZY4urNv3SKRhOQ+tptgKBIHP6Wf9xLzq8qd+F49nDWU/h8
AB8RqAvZ7FM2IMlXq/o7UlQDGHfiEkgXb00dBsDa7nd7KcmVl5QtRv3Tcgda77NB3mhGCGloVD7Y
Y8FsHfbbWiafBy9US2283JtnjNu0Tl7Od16Q8ZvfYkV43mF4OClEHRascGF2gD60amtHHVYARd6R
G/zU3rvnGT9GZTc9N+cIF4hG0TAwixqQ7b7CMm/0IDJ2fRoSagb9e501zyyBlXwwbPF6m9NxfCkh
vaaN0aFArZ49+gYs525PFng3r7P/0FmLKmLVJ4p+X+44f/etH4iPWuePyqcSi2tajk9RqQtkKNkO
DZBOogR3opygZ6v7AzsC1IWF3aayfZ/TLJenVGM1pQ4fzUE3//VLZU4xVAi+SGMCcNLVWBqPQj0K
98gDRxyjs5ERCkaOdQ02D2MLXA6QmDuI4JgxmhxFDkxKPsHI050xLub0kzygtRdZIW5Q0AeDABtw
1piLHDELJIWv7JQnYRuWCH4KGuhy2zMjpjqz8hMQHe62kBBR59/Kxdk2fo0j1KqidaSe390Fmq5x
HeCg0wkJrmyU0l/UZi7fbLW65lklo6BrNDmInpGPfyDnLYBh6lEQXMggiaSIagrk9UU4EQTgb+Bp
gbA+rfsp84G0aR9crT+U0IrjzyzCSVBGIVQd3pTKJHBmE/0ivlS7Inxg5c4S3wP7TebtLcAnqYmg
LalJUsJEiaDI82V83N+cwQ8bDpzTbuVmQs37cSADMBeJ7YzgNe1RT80MxScplH9+k/QrBqrr30i1
XoOdJ4z4bgvc9zRGr7mbgdr9R07mJJ7YjCOP4PPBiLaROAopFMXq2nnN9FZo4NG5Lz2Lu+Sl4n0n
zv5h8/XqM4kx7Afuu8lMHhwVoy3t58wLsZRZmX5n4Sl4E91aa7WcETJQ7av6yO43QkW+T4FqjSig
uUAV7Qtd7X1qTCaK2uA0XnDCy7UKkHYKE5BJvb6KBIBiGXxbiRYOvPVzdehgZrdcNPYrdJkeYi2h
NSQe34DKfZjiILFBrAUZPbnlRhaZ/Tg4frumtlywlPuNxPA+7cis1kfhSnX52pyYRLuSU65ur/oo
ejdteEQNk6KjKyWyZmQtNsSH/G7doLfoGBzDDcPdHEBrS6fjAI7ltIGTPci146WfePvjzaPd6Yvl
kfFP0q0xQ3wy9g3hGJwuWkFo55yLj8MggkrBkVTnvR2WetG9iN59nT0RgknDFoqn/rYvHARwFtWt
edu0HMjETnORpG9hdBro/IK4cnM/9RsiLmqwPVcB6gAzdn+3P+LKvr+KxbjmLAatiPxukKYhaOu0
bNZhsZFfLMTep0RHwzmu461I6ncK7W6jISetMdbNAJYKmDzgM+Eng/WoDletvVMvhogkJb+YhBl5
fH/wQKm2Al9zAR4W5FwGbQgo3ZGjQVWTsYb4VsOwx9OJmhV86cymD1u66El2oNkmEedsdWu+hQs7
fgn+4FsMHHMzA//TLbiWFgntF7QC2wNUvevYL/JkaCWT9rF2620wPEQaipyzNFWXTe89JiCxXz66
aLrFZ4Gz3n7njgMjZTOMi51NAANmXCtXmU+WhVbIhY22cXRxnLHS2TxGmLhp8g4tiq4mJuVWZOCT
a6tZXflVNKF3Br/ZQgA8opyECdaf8GkFCupVaOojH+Hr1T5bK9lhBrVjxFKcnDUvXJHaK1dNHL05
hUyWxczBSs0kSOi0GPAdBlXm5B1xuQZ744QB8pMdDBGpMUfoL2i31YigeJLld+6JSKqntc0dP1Rr
+k7evDNLN8gnah5Sx7EtB51Grczp7agM0do/DrrycO27t4t09KHhKMii6bXJClQudsFcGppuqgM6
W5gJVsP4GAILObOtkhQcbjBqUTQapBvlUBZfVCpVvhgi03RnVEQpoQSe3Ns8pKqPg9iATNQ1aJYH
t1v56FEMDq4Aw6D8KPkSRmK4hFag/IXgoEZ9NaWkQjCfrL3XVq8xsXOWw49rwsIrxU3Hek24OqK3
EXgPCjbnZI//RHTXZISL7DkYmuWM/zu03dRS8m0nkIXsSH7Zs5TWz3IVHYXuNOha9AeeH6sop/wi
+YTCHxNVz1LbR/4r7A+cwWHsnZai9GLWrdrAlH0+sRNFRh68O++oNva4gaRr+pqt8t7AExJvOv/O
UHGoEYSvrFfiua2XRvlJSuobfkMnGNBbmZTZ0RLQx9Z0VwdVIUSO9xHOWzKhVVFNSt7gJK/3sFM7
KpThZINBU9jKxr+AZTERPfCuZFGrfqflfRYw8dferKFh2qFwBZE8AmnzLYiBFoU0uT7LY72VkCJA
VKO24yCshF0L8Luwa4SV6qyo1KhBRFvNCwXmEfllDuVvCs4JyVSeHIK8hLrynmrPHrgqOK9rMF1K
j71gQbEglxisC2PkUETAmzLqr/KSFLRVrlF1MqASrAs848u3F6eedHNqrP7JRn2QISRCxrPM5x0Y
0WeixbPaXTfzGpijgXE0kuifwz7a9PJrd/cCpcbm/+TwVZm6Q1j3AjGHcRq7S0r6vcSvJDhm+ijZ
iI+xcgl478JzDOMHCZnxq/kyLrVsqlIrwE0fjT09PQSR0FId3wCVxzb2xWLXVV37rWsMg3xwJYr5
T20UG+TMzw/1V8e4CdyMHLqKcact8eLsZDXqJUNp3u/fFb8cq8ERXUtcbmkmIp7+Kpx66rwWueRd
DNrQMVfRcvYboQ/tzUvOhJ9n59ZJPn4cJnV1pMvs+4qzhUGUt5riF2E5UuznDwJAUSeXP6g9mtZD
8bMkMRk5SA/5oh8yA0YfFAlU5DTW/llBar9zssfoFNHSpvVOO8V/ikL2I9R0xmbGqiKcJKPiydcb
psiF+yCjqpK1S8XknCMfxSr7oLA0LDm+cJISdbJ/W32GmS5zV3/6WX64dKSLD1KhUyB4bB9UkM4t
8BQS+6oWfF/cFkkM2NQAEL59frKYyzMmd4xUQLmS5BhdTtOkc6spyb/+IgxCwnLJDBWFvZTLb2Gg
8MRXbXDt1a/e9NJ9XrxWLfQSuD2Ra3CYK8Ct1fMkRWsZIZphnGb3qiX9dLwVvFTKp7RSQJm4gsHh
UZu7fhgGYEDyp5ttCo6Zm/ojfMUHq1R9Ymqm5YqaH4f0SL9CUu0dqMTWj86SfR3+xUGtkIFkluH5
FvqfxRIEJTeyn008Y4HC+NKlr0CMX15wHx0sumAp13VrIGpZux+R1DwuWev0VcF2bDoo9UwCvfbU
8gOtdIj+1fHaTYsCEJk1uDaeV8yKnKEJC2ML5OqC17lScHtIzFXXEljGQ0BMv87Bpgp0odGY/QiY
lmukynRq95a+TfTreuLojP3iPhPfy08zp9wh9SI2T/FwtScfH82+ucu8+RNAx4U0Atwlb49fiGTc
xlgNFyWlI4J0VVTMC2TQifnKnh9ir3vAYtEkKtzHaSgDGsqe3ONwGYmFYPJESZEjgvw9aC+W/qD1
TwknNtV8RsTKFsQch9K4+ntsyv6sYpnRt3+jD5R1HMx9Jw2SlKY1HD8YwPyUJYm4CSEC5xxD/Q5F
bwZAEtq+6cLbx175Y3w49jMtdfnPjrPmqFJOYfMNuBYOyPEv3PyrINORUUS9VaxZXRPIVaKDELnF
YOvlkZgz47ytSm4gKJyRZWiQ6q/fgFlAbh7tmJBSI/2aQJmlFq/sEEo4W2csQ8JkcN0r4y62sTg1
wDxk20m8Wmd+pTmBX9HBbg8oqxALJQJuFPt27WhUUw43AAwutQUqBWWdeAI6/lNk1LHIS0L6MBZI
B0XBrAUd1xQfAp2F3wCrTgXiB9Z8eO6KXtb+ihXuu1qtcwvnlEbXzk7FT4SrYHUQcq72DL0pdsV4
OJKaxA/9NO7VT2s9z0yp6P09G2HXYkv7qCsy7pKtJJmBbFJ5zhONyhmozT7HvO2l5QUg1JzB15g3
L6DgFNbsjnVboVEaFgIA+IDRnlTEfiXqNM3mzVHbbybFH3MNVi6UoPc/sW5R6BWq2w3VxfE6yGrt
d5h62ihBKpxCeRnf/aL0IXYXFJ5VH3nKO+MHEa/Mb1PCLTmrMHrNoJ2YEUrRPWS1u3HmCiOIi4CS
YJvaE3mn3n2Ly8RwaVsUPCMqCb/kNDDVzjG9ZA1AtSEbUmoKZa+xg6sn+iaTvBCjCOTz5tlKtf8N
oqHIcnQI+Y5P8kutuP3dXWbZgMfQ0MtKtaYRRqrmQVPl3uDpP5fSt3KOLmLaedimAFvzkjYR1ZM4
EbeEm249dbPAFIuIRis8w4Z7Ngi/gGLeTLZSPHG5vguYijtz1K5FcNfttwDV2zSnPFYdNADWEnTi
CNKtT+cl5N3mssxWu6gqbcsSKoBSVEICycyUCuKZYpGy4zSa7TFHYTcZ4Jba+29qwRDHMlra5/nM
Hoq2oe/K4c+aFSZdDvErEEpoDlZIpp7cE+GVT326Zj1zwTp+6jxREXyxXVQdgYnasEpkAwLdcCni
a2YuCqDtcMz0hiiZzxNahgVzk7AycINkpzCy+q2sSrEGiVSd9VXWh5Z+nShVeyNmhWhygegK+IjF
E3K1RZWQ8Ang5rgtMJc9wliOSN7Z9p8Fn9j/1ZtbFzF/eTtzlLQTXbOilYt1uCJyqYRHhWEyVgIK
V+ZXeM9n9wH9Qz3nNUY8uGa6TkiANzB/nmXHS/0fW1l3bR7HBohD6gUbep1SA9jrAr3XdXcPl30D
WkhMLAgvf9/lUZGi9y3xXFh6FpjrMg/QcgULMLcR3Tml4UfAQSljsih0m7t1BThF5iRGnldVE9K9
80ASztvnYglfPzvzo2Or1tG3tYlM55xvxG3M5vxBoTU19hSfQYBIt/dA5poB7kt2ay5Ianc/Zicq
zAFhppALx7r5MuVZ+JYdNm04CXhvPY102H6MCo66tJAR/0RU0N/INS0fTXgt6yYBm0mF7oLj4Xk0
PwDcBUapu48zq5Fb/WQf0E/6Jm5QiK1VTU4CLj8YbmBo3AvGLHmR7KBceU5uy92svHvIpMK2SbWS
XJuzeh1YD17XaJh4njCzMnY4M43FSIe2m+LYLXpZOumsj5WNq03lvPehlzddeMYWc54VqObfqmA9
Ii8DzXLh83k7jlOmkqFb/1rxgzOOBpFKnDysEsuxELeyvQQzBPqoppftuY6Jw44wX9lMWweGln+s
OKAiTZX5LKtQyNeySlHMx8in+pURZdfzpHOIjEgjy8yrAyezQyizDZzkTXOpRgyeKE76hhTW4Tu9
9dC0kmBe4nJ/p9eI7tciB72035g09AyLaih6rEIcqKXy1RO78GafcwakjkQwDENiLR4pWfc1+EQe
Jinfj5QG59dtA+2cw/hr/11xm3HgvmJsY+JbrmYu6ZmSsrv/F7yMVoBSALbaGm6EmUksYocFZS6k
hFGlTbGgf31z+5K1f1X+4SQhcC1p+tV/N6w8rjH/2hhmUo6VZkGV2mmBLoRE+sL5UYJc4MV8ULUg
kJagq9bFpEGC+UhKfXuUUU4JIX1jflXOawV1thjOwXRwXcP6YPWYqq11RXMZUyCGBk3yCFoF4sBV
LLxqS5m+WPtbYjTeeuZZioA5DuknJpPSY6kFbVeVrW9KPzn9mU5Kdm3v5WEgsrgwHJjRkQ2UHMRT
F6NwvAIMeWEXFogwUbVW3/fGS4PHlktQhJ3ojcLgqYc4KIJgYDSvaosg9QxsH1aqt/ilfsQ2rYYY
fZ3T0RHyBj0FwA63IL/3aWW7FWJ+3srJHJj4RJ+l9p1NDtQ1vpspP4dqr2t/zns0pwe8ypF78qN4
VIcKc+kq4FqTp8QgEwntXMNDZSzH0CjJ2RKSP8uNP3IiTm2+Wq/0i2SvZlDJCJbaa3hczJ4hiO9B
PcSyaTV1rO7fVml2ZQKvr1t36FF0np5UdrdBW4LpmKJ8OYtrwTO7DZnb0rtIMYs8yH1+cV6vbVlp
+T83T8MeKF/fOgh+tdWo8fA9hEi6AEZJKr+BxmJBI5Opgd6FndG04Vv0n3mipaoUMgt2ncKcznrJ
1/apWpog3wM5hwQzG+rbq7itqgx9rf1IHvFBuGA0a864s5qKVwiCxNCmK3ckob/lMbEH4Kd5E19V
w5Tt4o0+KV9196CPBTipe8Di0DXysKDOXXo63TtTAPI6DRZ1JHgk0wMKYHmDrw68rItsRgAqr1o6
hJV3B6DtcTOTJ2BjYfYY45gndClrjNRE9oHgpJgNrgGybyI0VynvTSDT0JrLsvooSrMJkMLD6v1v
Iv5rIro12TBd29oAuJh7KV0CJU2l7D0zSIV58OaPMozg/JkneBIHWv1yW3cXEA02f/7vGZ+nxJqm
xkDz7q7pUVfwIhFSgkkRg37Jvnn++xMQw42bnxV2RZ16P9Fl+QbaauFndoOhyeNGeD/SFPkuvN+f
a7vgko3AAdKliVeSb+hB5poh0S/FfPVL+yIrB7y4IwmP2tLU8yVNJnk3ntnTQrn/tmm8UWuyI3Br
qdAsdIkBM4obfHFANxbWPglVAyCoGVmSOPR/j0CzCg9vBR0/D2mHe18zWlPC5AKMJt1HGIJ5tjcb
a87lJCfn9GZiOTqfrNHiZwcmFVMMOd5vpNX13MpN9adHmS8dMePAxlMBuc0daCQO3opphibd4P6v
OgXaSTi66zU3Ji7Q8TNuLwOud9vEntAt1kXJUkBYCRdydC3jybwTEWBcX5mbiYiGLWOSh5Y7WY0r
53PstgV/D7/ZZZer909XTdHBt+lsIjyWO343fu1ZzFD377DaKOq/MLv6AcWt4ynTeOAuMSkswMlj
Aqz/DBY5/9R+dVJXk7TZpdDcSnU4P6lbFZt3HQsiU13NZ+vS+gvqDZ5eHZLSRqMJ8WmHl8cgwe1v
ZcSF1HbiNwomj+klZLvz4GCiNTuA4+/pz802q6nNgZ65vlcAdPvWn7j7R3ifR60hoO4dc+gYtov1
ADtkjsSj6Kkpc1Avwo88V1qVS8Rlkb5Pobmw/Wdf00wmTBLF7/sjz3QBl0Sp86nIlAWr1ZbPEz8+
K/nyq7x1PyFzHVvwTaEqk15Xp/h3Q06Ad8KBuC2VBtieOFXFmdttMUL6yOzTQlBp1F5hBy171K+w
55pPuVPIgJ0q2KWZFIp/AjAmJL46zcLk1Xu218xLhGwWFUqPMMhwb6XpK5qSOyRovTj+WJEpVMe+
dJ1Ak8WtLFKDNDs803nrwdupxmGAjFhBTge0kxtIw/3t3Qd6eWMNIj6DHZZn9nDSTvywFGy/4wAG
y9OnZneUZCRuQ+rLkt1l1GlN7V0CA44n+bysOc8rMCdSKgDv1W0pexRDn0kPynf/6797OZrd2Osx
fxV5YJtBRRuWgsArA5lX7tvq89T11FAArSMXje7Exc7r6m92f7YAMFnUSMhgjvm87ocnU4nN8M1Z
vCVOft1DzbJJfEXJZDm9f71GR//IPEy3+jDXSbZqTYdGP3ADi88vcT42J66WdAJjMKBpt2Us0/Tm
3oquun9FaY991hzsQ6YnSVEqaNaEaQ7bskNZvAUSb1/9vwP6KSO1nHZbCZ5Cj3yqNLUjhAxk82AH
VOQpHkEoeeJQ+c08CMjT87qQEoIVxmfApg7sJ+HXoMEJOBrBgla0yDIMm8Tl7MkBSfytjiV3KoDE
aS+zhHD1c/9o505/8b9xhI8lA7W56nMPIHYVpus/Su2umaJwtBpC/YDqdRxzh/Ks4876c++2ZL9P
+hNhD10VZqiM+oGA1OrRIO0jxoAPHctUfXjst4yf/cCU41Q6qUm1lGZM5DfbG86edfBGDqfiyYLC
WDGQiaqqMgO2tmTdfaRpPovMLhePydt5RMDfZA2IhKAb4fvQRtxZBQ52cNUXLDyOYmPhtkY2ghkl
MUTLDv//9oCFdMQs0hipDPQW45bbuOt0Mwsj+WwMZ3CjovDjSHw5tki9l9QAGJpXD4U0xfoMtiz/
UJFK/n6RxxhLTwIHlqLq9heTG6NcEppjd9TtWi+GTc4m/sk9MLtgmuRPY87TCMnA61K/0zDmv99B
Ykh897Sp4tnQ5BVGp45HwhZ4ndw5x3OkWzWO7ZyWjWVgJR3pcMZMv+n89Vp6oHC4BXZRlsL3VkDx
2Yi+FYntncRLfSd4VdEnvat8gQJDGlOVBiuY2FBwK8slPKRv8U/MnUHYALLfShy3ObNRqAGSRx8s
a7IPN807pKPjq+1p+Q+vjlw1Ksh/5jBNzI2cs84iX93ago0sMKm/ZBCaifkLcPYiLrXAMjfGivoB
KA8px40FNk+Dqfg6POUnBosswsLiqyMNFPye6LpEVosq8oQkkTxnELMs9g8AJe6F5y4TJKP2qzyp
qqy54wI5ZKI6xNQQR5SH0qqnunlPoiuelFcbwwK7CjWg3HKTQVHbwiuGBIqirnTuvu7waVIO7LsP
jrBxtquSnpg1ZMFQY5TASox2wtvyIqVq62Qtvs8WovxFBsbDLmzgUR73g+8dVNJrIDwulk4lglav
a+/yWekOVlz8UewWlsI58eoRj40v7tSouWxFlEJ+ZXifjCZhHrL9LTJLJ6x3y1CmETccENfdqHuk
Bp4od01MEu5Wvo60T4jFoBDE0i3lTRucY5KDnPIFZdt5ftZ4EisOBPamca72v3AMm85LC6TAbCaU
NWQ4B4M2QF/cQ+ETLwXouJ6L9kdLJvjrGkl3FgRotuAxL6ABi3ObG+1lVLo9SkifGdysy7WCmPZk
QBgbo/DmRpZ7ZYQQ9yPHh5C3VnTxBvpRsOI5viFwHTCxn3ZIciQlrKu4uXbW0JVSj+0XLB4vsh65
UsYLP+SPO4nuUVHa5u1tcrLcHatjBj1a3llJ+li6YS1HvICF57iFg2M56EZReDXD9hlmtZ8LmXYh
/uZDAohGRiIYcZy/5+v4Z+dvohFPiHITD/8BlGmKEOSygcoAXdzux97L43ay6OB4ZVfrkxQzbZVV
t9UEGvlihqgPp5GV6xoc38Ie52HgzPENTaErRvqTCKHq4aAWKMs5qwgJjXHet2BA6Jeiw9UzqVpN
jVGMrLlFA/VduCoOzVTuW58QPfRy1Sy20qDnsGTDRHd1tRKNSk+m2RRkewvk3ORXQUx/sNmGHeFD
Y48L7lG5LxNJ0TULiDTJrRF8//lrCvpdWcGinIHE2u6VH1fBBnsnGLuz+ApPMDg03UiP+iF6tmza
3mG8N9etlMeQr9MHYjJZYWDRKEvy0pvUoWcaEwpf4mPOcS6f+0LtiIvAqAxoMAvdfCe1KvTAgQ3K
0NhpDpKEYi6UaBycIt+G4W59Cg0s/qFRby1VmtPV8ASETDpgQ2OeeSBOyKXgvWsBZ9KZu9x7VPc/
ZyNW+9bs+KXUBscoeqoa+Pcaa9f8THBJzhIGFSsildopckNrwmnSTVTytzeN5aA5wZETep1W4+a2
OGo7S2LmYEG/A85IBwPJO8P5dq3B96TLZADeesrLzWqavivWLDpYB5j9a42IfyifKSH6yFJIAaY3
GiaBSuNWH+KQbl4yiH3UhEujSRj2FsY4y3cz0EoWXToIJiC5W9256vAJMZRkFwv2mgHxhZFwqi7v
pIkIYZxryl0MAMRrecRgvrVq6Okbol1Aj6hmQV6ql4UfbpdkdOXtVad0R5ZONR2FJZ/dp94rwtXH
cqxXGNBxF/JiO3Gkt1WNZRYCKXUsFt9LfSOxgZtu4tre729dv/R2XiiVesEU/eX7iYC0y2cYeixE
JNpSWslfPeZv4bqDK+eTcoM38cXcS/aS1sARUIR7ADJQAtBhKQ1cCDta/d1tarj8QKTxAvUB4lTL
5cEl3OqVPMAnW89jkzgZQZi30KD93tnbZA/QoQEwKe1D4ZBYzNwyJuhKzCaWYcHmpqdbLGgkCa74
tx0xE+9fHisJGU4kBmj+AQLw/ks9Thrkj4FiWhDgstKJg1NXQbcWAsXGSv6eMbOHjJx3N2TZSGoG
+kXnCp9V1H70DIxIFHZgLczbG3jyNusVDefWP6Oc9QCrVdll3N/VQaWmarcf1L8Ta2qIpQF7/Ivg
lepuJrIARJYJjdwwqqDGWawUP4g2H+rvmPcOu+z3alguUsjiz4v5sOOuir8ggVolSvRuLjXHiWXK
w5eVNxU7suZyhIotCBZD1NkZRDTdyrdD98NWSjHANTR49HMBmkkZWXSnLH/u6cCAXW9E7xLbulPV
jppLlGHaG9oXk4RE8spV7n4go/H6WN+s4Cj0Cq0g66q6Rg9ZBKMzdQmdoGdQdVFjZv0g0QlUV022
SKHlER0x7U9MefswkGfh+drdy7R/py1AbkEKaKMl018qpsa4mw2gl7H0CfU624QhWidwMaEU3jpB
vBSvPPW9H6iO/ZlgmkAXZBr4SA69aX/Ce2aDgolpYnQLdAQbE0TBzfhJKvkpXcxWB6f3tL7HCt5U
EJNGW4uYF96wK0pM9efQ72/2UUprUbHPYxG583oSm96Mo/YnZx0SxkxYLRWLJhnee5OkKGch2Vxe
HhFKES9FbPY3w54sM3BinZ60ODmJtkWpSR1SNGtDpWOtKnvo21gQh///ZgQLTLLaxUo03cLiIuBx
c4Sjaoblf1wQntCL/RLkV2tN2q3Yo1AkVoHquntBvIKIrtfb0MmUGFjljvakAR5LYncKrParzrxY
2sOTV8IxfqJ6n3Aw2nDcc631RwmN1W13A1IooEPZdgxM5vy18VMFWot2pCetrVsLmWRbMmeNsIec
6aT2Xo4mMagAu/bCScNtncVjEr7ugynQudB6vIxkfO4GTdOVe+MIAkBQZRanBz2amk6gZIUJBaUH
XQIAS5h0Izl92i6hRsQbkfLK7q954PEmiYsENU0uUm+esfW8pMoJON5O2MPM/WW6Vk3JRArmTLVg
sOTHv22HSABXyp/lqkhx1g6EVO/GqztW7GN7o7wJw/Bf9l5DlLkZvOpLy35Mg9WYRiPViwQiTuBn
FSic+LKeJHKtz0XqBPTlHPZIEt7ZFQuSmRwh7qBlzKDtD704W1H1A3vv9FjG2Zysamg3Ik74xlIK
411afAwJoW6otcA0Z7oRu/vgblGlNkp4jtpRWYgRBb17zv10UE+PoP3hKkQp5WD/GzgKxjzu2pjU
vtG/qF8Y8W8TfJ/HybYVX4y370jQylA6zf6AUlFMnEVzg5zyBt0LlxdsQXm1DAmC1KvGJJvHgNnE
e/tP9k+M6eBLhHKvKBtGG/XshlL7wrr4FAm6nfQd0SRw/y945jGh4X3wAXu3/lPx3nW9pdvFw7LC
hLNaEFbYPVIChWkefq8l6he7Em68qoimr0BFmWQs7C0S8Mk2pKZywPUn27RMqEqX8KmO2prNG7o5
ROEZ4VRy0ZbKiaPnIhvqVcmsbHzrxNS47JvxBpn72LeK/GLs0SQiy/HhRKafM7KXgkLgqeumBjjD
4B8S8ExsCvhadxQ/L0Y1quyKsk2ihy1z4M6PaGVEDF+3LCJsQyBPvsGa6tFlMUhzZkz4M0JkHE/G
Q02L1w3BoG1EWy1F6Q8blKs7jceSQu87gtsvsPMfGQePWGPdDWVy0EIu8nNZOSxw9NkxrQGQzRGq
9nHpKJ9wnvV602/Y9ZXIkwGk9ZDUXXzhxFWvOLPSJ9GujLPXDFhDjsVpKk+szuN/0Pm7oD/k+uQ+
DjBkSnqhssqT2Le+FGH5YrCprb2BfkaMhlmPbBkCP0dwxpAkVej8GxJBkYdhY+HLxeXP5tIlgGvB
+obRS18Tia7wEtho+lwBKlBAkKy5v9H3SXVxMhxjtyjMf+dQKJk1QHQmy6gtnZ3UsFddnC5ZSm2B
qcK5VLrSNIWH1H4oVpMXa+0KvNegXAqfXyGGQihlsq3lW7BGHLzpqzMTl3qyXMEYlVWS2LQicjzi
MU2wih7/zuIWsX1fvjLNGwXBN9+HpbvW2pVxF6pqM2Poqgj6wQXkxNgyUp5bp3uczw2HrXsOK6jo
f4Hw6ofOWdCuAQFRg9+awkJ65JsDOBaa+tmTRDnCyNMqxtkfsrQRaw1jh3R6nW8d5TJjfuuzJCw1
qVz5525HVoB9ob/C2zMMj/TgCc7JCXapA7KvQFof2ww3OAJIbhHZf2ImANtWqhYmuwq8xA0a45w2
cH+J+TazrKvaSLsw4icdlJA+FMkyIDCDESnfBICRCuWVOixZu7pd+i6eifuPcbmZoQJZnMGHDmgH
WwnDrrOYNMKx9exIYRCfP4beTG5+s/a0s8fTdu8+5UxUr6INbqRShN7tPekMt2WN5BlIkW9RXh8G
WdCjHnbCO7AE2yBkypP2tsUSSqC89WCPa5d/8wBkM+byeujMZg1Fp4wdjtxv1cZXNMCevZomGYnW
Ayd0+tnYrI8ezk/mVQa8fqKqm7HOK4Aenev0wKCxs2PlbVRfTMxfJ6lwRItuWVz1fvIt2Zntf2SQ
p3p+BcKOef3rj4nsqw6201nOnFZOrYOSg1u4EWrMdWIjS+7hvIlToShVrAVeXsQJMfnwG79uoGgy
Zx7p4kimhOgykCEzb81ItXKrWMSEM9n/6Z6bt9itszrwBmlZwwohOUEsZqYFRgo5VnLTywQ3nI2j
uziNITgfHktzes7NYp8NMiBeHvf2NI8fzoUw+t+RbnCJoMNEmrnvbLscnyhfPKNXiXMGdLJ9oUmQ
EiT9CkdELbG0dzCIdyU5Tx4XyIFCYnrYAJeuGc3QX8AvngZHSn0xsm0nxhy/EpyqYcfE7taAVh+o
6y3BOiNDW3ZN+ZUgRmh3TwwmzfdHgA1KY59qSp6PONHyT0x5QmeFqC7M5bJW8y3LilN+8o76BhHt
EAoIQq//rrxUOquYTzYmMwGcHztMz7zw0iRCJD5BMatTJNICXuWAPA2Y4KrDacA21E3Nu055n+Z5
Xwx1ODgcsddca8ZMikyuhGTXwjmNd6j6z4ZRV9vyPK1s1XIUHBFKZTm1/bIzSdZUsim2dtkEA+fU
HArthR3FuQ5zhGYgcBT0Nkvnh/dYncdWp5jkm6ZAg/T/DoGEjvTiLQT8CKRHXjT36CX0P5A+/sOr
sSRbklR1GqcGo5okDHTm6jb18TjQtX/6PMTMIrEyf4FiC00buQhNUlw/tSwR8IgDXjdahighwbM5
Fg8Ud0Sjbaoh86AD4BfOsc3WrzDL3a09gPE4yi/nZInuBFFPosRWCC5hiwvlzrdDTtYsmVNeK8MA
ixVa7ycCXGAQ59tfrE7SuAFrK/N0AXR8Mbp+A4FcpFIYiQ6TeDeTaeW7+G/9+weF5Zpfe233vjut
JLLwcTTPnE9fIdr7EH/cD34pnJ4t8YvOAxvi0vI/J2nDluuaHBBRJLbg1rON6YEeqxNInG4cPxFp
KJ5JKELFleCj4+FIrMfOtqJRZoiAZJTs2LmpHwQvvsjKZSUXIg3vjHinA6TX6XBzmoRVLp+D3Kk+
mmRUw6JFAAJZxMoyoZot7A/YsUjdp9V+AN+9YP5VvZ26RfvDleFH22Za71j2ZMDgfueaPSmErW4E
2FaITucWUX2CAyR3YLRdIk6ofBjKBHc0WOK70uDGirGINISACcF7LB1ovBuo06nKdiVYzAjke/38
9TYttzrQ7y/nsYZNgII/xsZ9cKCBay/wR+wyH9fN282wPregiwU+fGM0XolVOTJXIdja/Ja1qOqS
HSvSBLeZif2C/2nxaeMFnIPl3NRf5Shb8NRnKQdq3h1QLGMtZSioZlNpUGollFz/N0txlnGi2ZGW
goblgs3ckFOG8dtAOe1CicqkkspxuHoUm30zWMuYZ8wcnbIeEwmjLTlWD0PnjqR22LdutznW3I6e
d1Tuo4H7MS9Cr72RWd3iZ61wUf38Rn9shcQm2vFFNLrmLp1XULZ3HOBOeBBt9gnz1J8IXryFfXkI
yjXnvl9ZurHwizrKdlLJFv/d+JkXFXyx+++bizmVUBLqwtfut+0S/974WYOywH2HdejszhLtzTUx
erv1hwPs00EQNySNajnWiHe9zTcjGBZpXjG6Q/O3IR+soOi89YH3bhEN9hB/DqZkaaWCADYTz6wN
wDpQ5+VB3/q9nT4RBg/81lMBZbP0gTuU2pfGjgcSxAn0RLGiXfFdc/2OMZpH4kiZ9Qq8sWcxOYVa
e5WEO1v9zFgh1SiHPLSDXfkEuhaFhU8+38RwWsjMh6NBtGxqxSSwRbGgxu868SlQ5P/KFHIuNqnX
+Uhc07EHseiv9bggSGZsujqeGQmssj1nI8Ma2JdEWjNp5HT++H50vDZZZb0rDPGcbmFZfCnG28hL
Ei4Ls2RC63n+lcB+51EN7I38NULuYKQfKOhzS3EULQlbC8gy24fW3NPuVmf34UYVV+LqN2y/I7KB
LqJj0apxoaLySj1EA2QlGdsJW9TlT/ZliL3XAuF1M57JtlL7Av7z0uKWz12sHl0jIVRrqqoUsgtb
LVYepUPWyiTVbM1AwN0rlCzthFzw/FUdGuzd0CW5Vb7DI1kpiCaz19ZzQtBpQisCauXVuAkFyo20
aPZpkr4MeDK2QrspdUjhjPrxFm1ZDmvsbQMB4cUkJ9R4bVP+DSi8iqH6YbpPcdPq8DeKhgCo672J
Ty1V7J/7BKKYNq277E/lIN3XSZkpXvIw3IYP5PQpOi0j5zviBU3j/JR+sJj2s8mwpDgHvkiTtNOa
wy4rM+N3AocwSNoKaUyWD7XQNgGh2i11D55pUS4xr/2zHNuLkdQC/V3+LRU0fwjld4hm2XPB05hl
XYObOZHz2Eulvb5nrEUsWp5kaKhuAO37t0n64xFFSvbpfwKJfnsVhDtc/zqqbud07EIl5HQzfQzV
92NYJX5EWiwYbnM64IOTj/xZxkNaxHqTPDHwIr9t/nkWj+Lhy5jZZHvzgUkuWwv//430KgGDcoPE
kAo9xfy7lSVFKpacNqOV45tUis4DueyAoeULWPWYyteCvY/h7JbJgAUrJtfJDKdaFLB61Eg99IU4
EiuzLaEO7w==
`protect end_protected
