`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BumwjKwgynLUhacTS4vb+0b9403BmW4VMNuYGlqISXP4bHDu9oNGPA5musld7KjvTtBeB9gGoHkK
AcySYT0PJQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g6tt6KmbRdBXCzU/P6DWrgU0p6EllTgbpxudZlztJiVsPXvpU+QlPwTF25rGm+z2oO4cMSKzJQUh
IzbM2xY/2+K4e1IP6DsW0dzPaA6VnYkGoa+qCXNRe5f6eW78a5eOVPjFAQhC92irj0sX4OF9ZGwH
ZxPKoyqM6IpbUF/a8yA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ftP1GTVKBNQTWoQAaJUcERKmQ7iHAMlvf5sCSX7ULb0adMAtQ1JhHoIKrxmyvXFdFtC5J0dKWFHt
DykYiZNxemuNRMvKLFT0eUOEhcfe3PewgRTO0Ngibrm+UomrPRTCy5n6Ehg7Ee5560mfyZHFX+mH
+yMlfI8kbCnRtFFc0igmC2nh4u42WoeS5ulV08WbOkaRXn17JQBIGguELaP7I4Y8vCPCm3W0+rOr
94M8bGOy7VEH+REU0+2WA6YBTTeFP8JRGr1Nc3+R4TL2TQvCtuSa8LvyxA1ILKJiOdtsIXzrrNN5
nnZzQfT7LprMmhBYjmLeMCe6z2BZKW+TfTPYzA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T48dwGGSrrh9RGcmQscpOin4tOn9vVSUip19MyrdeKAtZT4nU++z5V8KhrJO4rJ3vPgQTnvioUD3
ZdhuhkHmRKt7mvIPjz1n79KZuuKkclVEzeXwJp9F70hvXPb9AEiFT6NZwW/pf6hwpWsJI95Dbkiv
4hvgUY52W8s84zaGLQI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L2G+8KcTk+T8rvtsyeYAUTOSN7D/VZ+AIxK1ze95FB3Q+5m7zks8/cV/fMi9sAuVxsHsL88yhYLs
xcK0YKWwVjEWrxpqqokuNw+TJzONGbv0zEtd7gsz9e21aPuhIQ5XVbTI9dObdJ/ehBrLh4jroVUs
bW+ClUnI5Li0V4pcpEQ2oaF4k+GgwQaQLJ0FeSKTU+sNQRTS9U1y2WRJNXorIZQcGnjmHAbqr1v/
QSULdWUjHpcWGdUmjm5now4GWKK0C/s1lWNAkYnrDZzMGM5BGj2owWx35K5OYu0dhgFsCpxpt6uH
Zl0xAZqCTiEpvxDP+vgwhKI2AhKIgPG7qhGBRA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10416)
`protect data_block
lwRGukOVJmlXlmti0awYC784bNzRZ5gQ2Eyaq/idyvOMtiJ0Rg2ayvmNSEV9DTAMW9RI0vWxac03
uFNngVIfMDuO0qPY2yB1NC9/VJ4OWBBITG5OrkeNF5KhkrdHHwDzNgjcTD1wvGEYhpY1l/OZWpLW
bgLWM3JsH4j6DKUIWk3C55mST+IyTg6Ju3vYvpgI7plJ5/trwOiINMpHg5spoHZtswN2lRxZ+uXI
/zvdFVMaOQ3ZALK+9sLQyj9wrNEoim4MPxPv1tJJrTkBFCaBSkfVX7T8+H/lvQcOm3Y+TE5m15GV
2dPB0JCwS5a8tUVmQRMmbpR1YG1AlbOiwTlgJksatDcxvvzzwaEfQ5EPI6g8wd99GoHojL5jfV0R
R9C+ji43g2hxXAbfnY+21PAus5PtEh3tVikn1y7G91wY6WMviu/nO6Ob9oXHZzcxHEHBQ+I8CfZG
dNWf/aP6pV6q1rbRJEUmizsj1L1o8LyGGMPG1mQD13MJcOyikBx+ityjO675VJZgv6H1oyOSEaem
YBksx9Mej6wUC8ooliSZqLj3sD7dIiJKIpzO/ztKMgAfZg1gAVAV37wjck+E2eW/JPV5ssMi9SGJ
iBPb8iKP+cnbuC57fg4zsNTsvwGJUrViU6RxtkOyPHdE2S3P0Ipa1h0ZQKs9CxvkLhZrPt5q19We
yAHOGJ+5F3w+6y71vBN/WMRcqTfFMivZIfLmdGc6elklJDX3DR9SH7Aw1bJVCuSj44IhjOMfb9dY
44i8YjZs8QO2zMtiwPPQ/yJlaXChdEWoGgPucdk0EKEe9IwLdEVqWrGR/eWwP6f4Y8QF2nJlFpYH
dTf9L87tMffEHNOeoAEeiCViFN971xOPrGeB94Bi405KkMq7BkYmIJ0Ob6wbxTI4ya24bVPE4c9m
cald7a+jCRKJawuTAci7OYNwOsEejzP+PzjBNo6ZjbTILv2PATS8EYBVxBSh0Lfathkt9H8mKhar
Hu1q2qUBuwwAQ8KslQtj22fiXx+xUqe1PAZ3+PuoNfDnnpqxbNk9mTRsRPXuE3MP5Dzqq+4NQSTX
vr6eZO6DQEEvJv7bHrr59wdetchyjPpOo28nuKt7e6Kxvj/QHGtvd4A2yHPCTBGRRMBlWQeLuiSE
x4+F2ZKmZkKsgwYmu2WBxnEgPg+Kw//SO0LsGZUYobswIApJ3T0F3BWpu7fN/VhA+uQugdvtTRXM
BDY39jU9hEH0kd156g+3pY+k3I9P3eQyAKHqHINQ/HeVtZ3KQjie2xpES/Fx/bE722S013Q8oYFa
LyQcZ6/3AZvYwpIQynMgBX0sA2CVAdQtsvAsLQwYiS3G6F+C7cXcBBG40EdoK5XgF/JxZAMGiyrv
FVmpGYfBm+vpxSdxJgupnwQAfahCM2SbyE6B6D4GqL6DLg/94pnODhx/GjSpJCofQN4h2Oj5B/Ea
C0KUNqp7uHLmHW6lt36Fc0N0LwzLxnQZhPJc9PC0/ErncEbAWpSbXYUXXUMZbNzRRbD3q6acy4Rh
zFkbe8ZfFp81qMNsZDXQSG/bmAfEmOwrHUeVST3/0me1gJbDqtzv+BQzSkqpnwE/2vC3ad4OCc+N
YTn5B4E7MFKMgTXXsuDSdNps5r+WeWTGTh4Et7rBRSFby98Ui69pLhSjA89xqANL8L2Z4m9yC2m5
OJZ9o0NkabIGrLVBQZjJgdfC4dQVFlkrdFkj51dMOdC86I2urvrj2nQCwN9CSx9SpemjSyJ6UNea
SoL8ZFaSfcGDY7RV/EyFMeHGUMc2/P+k+9PCEJH8GmXOVBCAfmFfe1il9vFpZu7K6Vcp7r2wHcxK
+ZGTsvmMTXj7r3m0qfkFbBF57s4uP7zjChAuChgy9E/LrnZO6sA7VP0FsBaw0/U0cTrJDc2n1m7i
RpepPVVazDY52z7dx3l3c9ILfEsTp1gNadGcz1Eumxdak3ZoSZhqTLk2kj9pIVtK4ZJeMXXWcBPk
5Ypn1WxgNqYHeSBspn16hREyjU6I70u9Jygmk4vHrgg92B360sd4/LEMkTJiFW1giyISFIahYq03
WE1LG4eHWtZIWAnVfMw+VhgrKAwoc9/OnFQorSrB+sVo9cJUEn9w5FZEfW1oX75A7HJtGIiOuZGl
+BAwn8WUqp4WbCvk68pLRIqP9dmSZMlmJjK4t/CUiOVdTwa4qZcDHBJQvYv67tZT/mCJI72EJfp3
tPz2mUwvVbhEItwcuaomQ2CAlsyl7YciDKumdZ72VTdEJdoQ/gAABWp7+SA3c9FSERnODTS16ZeW
Fkvk5HOhPUPH7klcXEtn9+hRZNWUrSOFc5T9B7NbZxBttcVkZ+g3cRPVIKig+PUpdfj7X7DPFV6n
zfr3XgBVZUmfeH2SLr4e+ias4NqM9U9XPVgUhOqJnz19Scf2pmtR3yXfu4SvGow5400VGVe1dhVZ
gJUNmT99ER+7mrK4Ein8l9bY8ikAvdm9UtE5/y6+Feo0XRX4D1rxI7RSMG2WAXbHfjhLS/A1DAra
sVxbS7DzUbw/1tlaqPdZ1wBMkfiFYYNldwOd35Y4nK/V5QEbtoy34gnXHeXBsFdPVY8ph1aV/4cj
/QmxkQHoqQLbumEB12DADJP6dPuaP5wcVMAdHlgOKTeuqKR9o5BiXTo/PcDhVHW9/1WSS1zoFeE5
njZKWqRu7JvfeGzrQTYgy9xG5IlAH4mBoZS8g0VEW+y0IozqvmJ0F0o+6cWfORCzLpTGwHAO+wuX
nevDshm1zIc/wlW9P3fi8SXXHJqugV6NdJLg69KzQ03KOhQFFW8r+5MytxcwQpSsXMCSrCa5E10s
9lBbib+Gt16isu+FJ29UnWB2mO0gmPPUpjug4qvKcwDPKunFlKYoPu9WFouEWKdeq906cftiy0AS
5JBFrqkEyyEbf+nA5MbBijEuOpvm2WbVQ/y8rnvz9JObocdu+paVHHrt6iW9Uq3UpMg9zxPqLVMA
qrSE9IxdkECpkBjT9FeX85yHmLS//jAnPIfJ0bcqIy7v5FOXAdTXrtynw0NA6IUHS4rBMqm0ytpA
2THRDEi38ypFfzZPTQsQRQWNYGuQFj5YygOug8Dfrk/ffz9sJTGVLPdC2NYOpmhuWRcXRJVe8pQx
e1SaNgq3rpGKclroaCWhl4XWmMl9KJ4Ic58voJobrmFf7faeAqf6CCvSllEtYtn2NWxYzCzB6/4p
XctI+2+fWCPO6KSyuBg7tE+wWmzwM1W6smooHBJIPK8XnyWSE5vUTZb90/OrZem8EnhI69AYtN/a
Jy+2jvEFioZMcZC9ANtfiFqJKZ1El/i4cbRAJ8EtUVsBR6+keEeybP+P/O1Y4BPpSH4T5PCKTHPx
VkwI/7AQQpw5GpT7twyx/jC8hjk1Td7KptUBDLmPgXNZEeXSVvv3+Zve7rKITKjKqwB+fBjGLWjL
+FF6gPw6ZPaWlgrQgJDyGlcStNrrGKTZwOhKF/edKhplboCA4rO5Pb8gkI6zGynwxML75YEZf1Iu
G+T7Jr8rOP+m/njBIn7YYEKa/hMLvoEdUyK7JpI7wHM2keBSHf6rZPyXHp+tNmIFt/dBgPQk+qlS
CVpoQ3lYl9eiAb1rJn/u37L2hk9cRS7uKsh+JON1b78O1m7Q0Jc6IozbOsnTJZp3Mxav2ivEVg16
69m+EpEdNG5ryTGwoiFUIbgsDNEZ4I5nXrsVrnjwGO2RnUCeWERSZweth8EpDj+Iqs979j0hNqNI
Ls8U/BihPEG9vkvpbOWiFNB3M9RFO946fW02mGxXCrn81wB40+uQUZIFD1Xsv61AtjSZTyCYiyC0
Pd4B3DFAa5JUPZxjg6p8FiDybLv7/6IUsgtAtj8R7CnSAMYL/8tllcQKZgTU4KnEGeNLnVjHLLMk
TStA77s0OLcsg9Zpsl62VvK4ZKdE1brx/Vf0FshXoaLJis89o05NDst9RlBt8es1C6dIkqLjD/fa
2ZxiXA1HnM4m2GBcHMqXDqCFMaqXBNpUBzV0NJhe4AjUrmZ+i2VjYc1VbANZClSeQ0S0z/vthNvo
7Xxy7UjqnuHIdIGTqoOWuNcSrro1J4vUSdLIkCzCEhPfp354AYXQpUYR79L5Jo63NlRwgRGylZbe
g5ZDvvkVufANNxnA6KcoDFlo/YIFTqYEpnKjesAf+nH0owh/l+6RXIdkLscQpU3/KkoTzB8Hflgm
EanOSzQCerzND7pXzqBco50HmNy/Y9ehVsF4BXBpreOaBf8r9j1dwVhqFmJdl8UKi9k1GqaJSCk4
iE89ijc46zpll1vDiZ0Rb7qyv8/dtZdSSc3Buu+SPtAf9cscvcdGRRLjS4e/pVj6GRn4co9mF/3D
dajc5VEEWISaN+/W1QQuuaBl5Uxo+KSGi7puRMkDZq87Zw35fa6pEuiberoGzpf3GnmyWcyD+7fZ
041g7S00sgaIAudXY8fv6BpP8WFagiNtHpZIH3Wg0OSM38E8wDXdIWb/RWAp5VqOSDpK1PUhbplt
BH9aMMN51zdkdWCcB3iI3h3VfvlbroCCLH+O8C54lBm13MIau62k7jn2On5aVouGshnKUZYtcYGc
3RiFnAu2RbrOX9oBN7g17FqMAKJSHmCV28p4AEQTXz21pWEgLt1apgcRberQcJSn1r6hDtM3LGw/
5oDmLBE/BMaaUCYssV2U7mBwT47yDgapL9ZvKWdXsTz2D1X5+WuzCN3an45j5Gqs6Euw7twjRZ8a
DLau+kQqmIqMQxu33a13RUcJ4LGbxVsFaH0XK/SCdm6oYAThWlvNcL/Idh5qWArtB7GgXvMF7qz6
86jkrYmgmzs9U7rJYvq+hBw+Z5efONpieZ1ts5PQxGRC1JI9oUqDChN7hr6WeUeObx3EJcTrn1cr
AsaZ2rw4HD0/Hbal1FFCXh9uONfZRGxsg7Mp/sKUbSVHcrIUTkFRjUqJIlStnJozW+wvDPkeEpOf
fsDowhan/TWJRWfMrM5BTzMBqL/ZMAfyz2ndMbaqs01coazAWolqIfTJWtXR5CoZEvF9Sb+uZwW9
XwRduRrVMV99Ph4NZjmRw/706uF4C2D423FaUWvko5oa7vcQDkb0mNr4RNu4KwtnVLTIwyX7TxoY
w8k5s6s4O2trBAGcqce27td40fvRN/W9GuZD9ekzLUX8sCC1zKWm5BVBvB/oE/2DCFMo9IU6exT6
9KS6qrK6ovfGF2FqR8wBPDguifnFEzHy8jwLldjujEUiQIA+pQCll/wfz9Q7HjZEFY0joJlVD5n8
lI1X24bucpiOxRVPla6+U5OkZixpKn5tP5DLfV9rydc1sIykRwpU1C3KsY8Hq6jz+w27wou+HUAS
8Vw1Fw3UXZTvt/4JpiYRRiIP0anpTqYJZWipL9j+mmLSvJ+MuUf6gi9dbBo0DxahyQ4/RAnvJyNH
+0P1IHjcp/6SwNx9xf/uZLM1HHcoTm5lm/rcMhqKCnWm04IByW94PA/rb1JIC6gVa4ZcjixL4Yyx
uw7wNto7nN+ZYKg5LK6xAXdw6Q5gc+d4B0O9dk+rHHSEei4xSN1lz1Q3iAEmW1YxtS4hCilC82sq
kgpjCoL681dfplglBrU+tYcTlxGu8Jkj33JHVx+7cvZeQ8/FuwNziM2FWAtzoVZmxe6UOjOpgTHh
fdOGu+TnNbPF6+iUB2IgsCiM1U0srE8MibPpAtzjnTFurdCPYJTYCu88GuoNVDzvtAzZ1tQFnY1d
e1chem+yqiWOClM2I8hTY0lWT/m9xS1VHxTdPOj92YjErdbWAjEdVkEEfWonceywR907hpAu4YZj
jSv8Oy3VlQRcutmhrZ5iVg5XSfyk2qzpdf33ouqpXaLoxTZFhDv+uaxMhEbDVSmi1rcLYmpIKGuG
G9o2r0X/lPLFNnU7ZgKd8c4spMM1fQU97MjC2k4xmYrSjsmtnosao4JmojYPojS1cx3TsuXaH8q0
QZhzTJD65ZIxjfnkeK9/aUO0ahFvS0J0YkZce43WcXKQHfyvbBLWbF/39xOkXEm0L9XVmNP3UHaV
zxlSEVMcFubduhV/4n8YG3QHf2nIBB7fLqjMS2Jkt8w5n382pAUkGcTpawy7ShnYQlxIXIgoZ1MH
47SPK6wI/p8jr4A6rLu9h3N6y7+hQ9dXxLeifigD6bdF8saRECST6vfrTXrwngqFPbu9oeNexzyu
9ZQGAFxkYAtjDCERhFkghzfGqjZENypNrVFDM0mFa9TI/QKULvTaxBgUwSnpu5dbbQxseZt4QqjG
Aiy0TAMfthogOdQmh3z0UlSkyPGB6PJjWVpFrf/BzKsnwzQv79TR6fRfeZaD6eGJbNuQDd16QbYu
hqA8eKMHV9OZZoFiA8khrsWBCkHd+tMn5SZHNH1+2tINXp9NfaR4L52O/93aGQTvNvAbsEZabqF/
MUUYqSpi5m+JDfzxhCDAJwgPuLK0sZbXZLh8yjUbxZYHw5fg+vsOPsNMwuDoiL70vNqFFFa7Orr5
zhNjb+j5dndi11L/9BUNnA0xlKUVCGeOTcU5PFsmH06QoRgD3MHnoCgQSisaSlRh4lehNC9lExJ+
b1Ad6AWgVbNyQvSOqeNLVgGtqSzwCkDeNgxc+HfPAI5w9GkA3Rm2yxn3oQNnuNG9WkNVIMb3YXBQ
CbmuMgQeE2eyqFADoaiEZ5DmQjIQfcIhmFXJhdHthXFe3Hlb8carAHqw/791QbWY5dqovK4JObEE
SUhTs4Hz24SiC9mCRIbb48NTWNHOMZtaNYFT/GEieHM42/90q+rgUs8keaTuGdDCvk2Xj4+3g9rr
dl/DWwj83ut3HCtDhA2Ct8pAoX1XO9f+Hycyi4dNKX4LoWM/jO3ArE+LBITxHNNJ6Jz6kDXoCsh9
o1sVS8D5/44T9t20Ef0QgS6dQbO7osQbSz0qIhGyEU8aLN3ZM0yyjGtZH4hxwBKc+f0/W6GHDms3
pdyNbI+XOTaQqJDULuisfHdSgKzYo8ZUr1qWWyv3DA6Ctk7lNb4my7XYyHr5ldoNty+bvcYFNS1T
S5Nf7AityRyhrYZNtxSxH9XVQqe6ti9JPKjlc5bGwQDl2RyHBNxy8ACfbShFr0judqzJQIntIgRp
5H+xwr0QLW0arzsQf9OcNNa0BzaClzgn+z152HuQ6q/b4t2YOmasKTPMa8Csb044VJ32zAX5YEzW
jAnFYK1TMPBMFkwNo5WUfVBKci1dk9TQF8F9C2G5ffBxx3QLOTFqpeAspngCl5ADLEq7p4dTyEDJ
Yeis2xR1ULEQPubbiCKJWwMkdKV4yV1N+RRcDrL0Iod/NKOsaWiQPq/Rc7cJq0xdbQyQ/1sCRW0i
RUlwj5qkgpON+m0t15FN64C/HNGhatYpDpoGbTlji3rzrRYDNWVELNQHv0f4wMB0NPW5Hv0MvEdf
rp/MJZX0DvzdfbHs7S0vtFq+P2LLXKeoz5rcpGdXToVQGaqb35DvCsHDKYle52UT8AjWOBHRJ7T8
SoE7RRA/DBim5iRDZV1vQYoDx+mz3pUk9E3ekD/ZMt2TMnCGhsagJOE+fkg5gNVZAI23A/yv/mEC
w49vej5J7X5qqn5hK6tQR+NhqW8WUzR1TRhyEkrxp4Kd4E3pKODLovS431fdMsK5GQvUd+ofKLHW
OJXdxcm4r2r9DoPmXkptdgrIO36QY58b8NfMmKGQPQgkJ6ScKroC8hEulSnWtWAGtMf7pLzM+Cwf
4Y0quROmROouhL+e63rmT4s6CP5gvXuQmcca9AeWt4DkrwYDy/U+4cXaLH4yCyrpSwHIe3DJJv7p
mgnQVmwa4S5uHBheG4/kXgwvInI93QC/mI6lU4z2W2UsWZZc8Wg4s7vrooyLXurZFAFFAQ83e5SG
XcJX0VqUeZzEnDO+EuQWA4XE92A7hQa3Yvqvqj7P4j8+h4rvklWgUeQKEo+LO5xMXIpDQe4s70EW
Ev7WAf/B9RFt/ORQLZqRmA2xZLesk8wsOR+ckY+kLy15y71VyDDH95pFK9Q2UfB+AotVHz3A3CMQ
lmgjRRIsHhAbusPY9O/lyDRnIMpxkIHW48lPthkHCE1vVoO9tvqhVrg5Zu+UrELSwuNsTsaGYThz
TwJdAagFopOZmw3pUm7q57Oq1h0UE7teBR4QL1xRfTTZ0yRRNrePLW9nIyrgB2PVLoJ7vCp1IH+r
XdJtu1RXdfMLBoDZVATjrfIIYOLtQogCsd2ef6QxB3oAlcuE/NUNZTq5qXYTkgB+eVkKH29ye0Cy
Y/wiYZp4Dsg+Giw8G9qw1MNuqpdRpPD2qW9XNp3SEgD1b5uulZPzyCoKfAVa+4+ygWRdzxCEhT/K
2O7UbZTfNBtVhUxB1y8GsO2FvpAm9Zo/nED6MHzBB1qJ8EPUG/vRrDQSeNe809d/5rtgMlsn9I4J
5SJ9DeLIiJ4RobzlZ4IMLTfpABJFx315EUDRXMul3G66p8NR3AcbLjZ0Ccb32xWhntYmFq8bxPi1
9gD4NJaZXNCxgosKu9yyKUBkAUjuSZqIY8Br8PXAGMqcycluJCocSIiP/Doc9qtmhsepVwrApr0V
pIK74ohUPH5LnvEHHr3WOk+xu6ct15tCrPf1NYvRBwVEUdSW2jBUGQYqMaU1TOKwPW7EPMLsDFQ0
PTswW9MqlpHy0J/7jvRwADBMSwsp6mObAlvNFy1E1idjKZ931g1z5yiOns+gtGDZYBW+Edn1AQDV
wWVhvG7wnoQv0FAgIqiRdPNqCszxFUO7wBcA1j0FcLU8FZY58w54gcPUkw6RAO96WaVol5nXnY59
3R6R0XvzWEiKdJqEoLC4hb6NvCYyXuGonLvIzRvEERCIDaDgXNkUSQ/f/2Cb+WZpmcktayCL6qiB
RJR8z54Na6ni2VqMAwMoDWnf5Bzg2WtAd6o2jKTEiCVWPC6fm2zR6yWjWkfwUP0SHCF8QfQnorlL
lQ7rR1xD8HdqoTwvzN5UO9Yuf+n+sn6T9mNraQHyguFEDrEZA5ZbU6+bMdx9W5yDQfz0mdDq2PG1
LY7y02JGh5dWYSbcr121OKKMoCehwNW3+nTea5+w6c1m4NWE5l3IHKU2WP0rXmMFswK6n2q8pnKp
iyGyA+TgX7HAR9OyECS9wADIzEZMaGVtghvoYTdYtytsQ8Hzy5H6Zby8hXQ0JYNYQdFOUrkxPID/
G0L0eiChbQjPTMVsQsiMTHeZYK+XIw9qJtDJhUWX+vcfHy2O0q+OF61l2QnktVBHlMHwfjGHYT7T
gSVv8Lp6la0ASmAVt36g4n5VYa6BMa+a4Tp79qZJH373+qjet9ZPEur/RP7Mz/7fbvke2gTSv34j
Fa3Hg+wyx4oW9SPd8MdFmgdy3A6QviS3QqCJWFvekPoWpYOuhQJpDeC53RQQofcP7OIdBLRLZXwL
FVOl9tRTIlMDc/Z1UT/XlpdErINwLVCPC7K07Pcsk++QyGfUUEN8CrDjrMqOREzCUyEuHCEpbTmm
nnq54OawqJ/9aAPxAXcsTUoKSCM49FuN+Rm9jyl3sDcW9iiZmIBd2yU4B9Q9AlmB2IPVHCbv91GI
BHmwPni/8Rsdpp6zSTAQda6nKGRh7ytIecyupOhYM6iLwsHGM3hfBQ/TfNvFqh7K4bqAYv/zKkio
uvnTzh2FYNDaeDL0D9NUXFmkyowvueJL3Bg1BR8ExxWe/PHvyegBXh9xFr5Pjlx7Huasj7A1CfHH
81ATb0edetjv1MNmVBpQtRQ0opKiXB1xurzAZ2xVFXMGTHwl4nU1EkwWZQ+G37C/NON3yrkiXwy+
3zU16zkGX7+c72BzXrMuzsEstcHRFbMzO1+vfwb8R2rq9FsIGDVTJ8FW/0kYf97FPDtAw9yfIJ/H
Pr5yOypoODVca34lyDCUR6/BCNBPqXS6uK7bG4gvONnTg/yoKpHEiyLXhmZAQCjNvWSX7ibovKqW
TIWxkmxJFLHEUaxAhcW1M2iomyiPMg/NFh6HCD7puN3rjGjV3OnLkVLmVvUcE65VqtdlpGzmjEZy
Eq11wnjPW/2d23Xxy9Skf36mzoiK/JI4lqqvsBEMNiWVv6OuaAzupiabI4FP5syRw3d0+Q0I/htg
cfz8W+eGovKYRCavZV4lyR0YrdTtzLJIq3edCvUuy8ZJFTolpJy22P4r3Ic5JnqaiV00MFKrrjp5
mzf2VzsjE3B/3exuo4t59dat5fbODa2P7yqjwlBp7meYHFoIPg4MmC4AjFs4Xn1N5/PwCEg/4JJK
4l5v1p7cy1ISphhph3P1L9sdMIrMH00t1vjSKqznCT8YCeixN3aRfb06nllvHt0cZsSCLaHy145Q
CVEZd3IaiZqWaRZ5ISXjT/FF3HTvKf/3GqAmY4GXV8ZgrgnwdTcfj8L0p2aZ7pSLB44b4+qeI0FP
R0v/c/W+P5d5XD0oJvdU43bDDK9gfUqtbgNCQNbo7fSNp79mq+0OMA6c+IkkTDQKhs9PJkwkQfTS
zRd6w6xbDHA+ECiGKPyG+wPFumH/dGduVhd7VsRB4Nxs8ZWDUKSqU9eCwbeXJlIE8Of6zl3Z/H+i
0jfatCtr4HipT6DzLjH4OHqzP9AVo1z6Cday08xnmITD67NQArD9FYXS4yv1cRvlMtpvXLIIuQFc
rSbPMIGhKUx8x79m18Pk3GXfZWDbcuxck6HIYhM2MUOGWT00JHk7Ow/J2qQk6zP2raKKk9u/wFWL
+sWUvGIfOY0kMmfQpVGpsKpNmhXIfQeDaKZ9jL++OwpN6OJXdTV92X2trsGUzRzZjbmdUYp39So3
0pyLJcmp3xfVTqI6SMNmTyu0OpbkCsLJJ+ApO3FlvxPr7+497fWV7YG7AxSKJaWX5j5Aq4JhblD7
TxT5wahnOuzDdOddXNp01hcI5dfFxzjFBP3cTj4ZoTRWegO89xn0N7BFdnfykrCD4YWQyUxnF7/n
rylIsQGZu1xGzO+oP4s75159xP5sFcGp7dGwF91yurVdzEU6NdVJgIhPMovELcazPRqdQqjcDcRk
0MOasjg8zL9LcUvcqtZVWHnFoh+aI8eocTTLlBHl3Ayi50K1LyNiOzuLtIC03tXakq8tlzgZ22P7
lGmWTGCfUlhLzcUUI8nJ/G3UPIpd7LQqwUE3R4OqikosLYq6VJPssk3gjZlAGHm0T+gqXnfLJUBN
VDxeO0oJHxG2KhkCQPJp8G2u89Tgh3kw1foe8g/Ox18VPi4v7JWqXRsqnrIslxVCabsP+rBUJAjw
EphkomXeGt9u5dtyVJ8HGVUhNP3rrZIuLF9S2j9SWEisbtc3r2/HdLhqvt3ePK8cu0SpphHjJojN
Bm2n10FGmW5QeMNFQws+EEmT6pITPf7BMqe73/8bjDBwa6oh2HTmmHZlnwsG8k80txFsPv+Zzkag
qJN7TH1PUegwFNj4fJzemY41z23PdCyAZ5I9CVJ6zfLyiGKfnU7hyCXG0RVdLQuB+nsp20QlN9Ma
HX9F6lW4mF5qFxF1O+BHMc7XSIiLKsk7ZJlhzRKH7U7tYOc9S0W1CAv/BQB8GlGzYPsIwZvGxM/f
ZgQuL/KOrFeY5b/vbJIj3qLP+hVXG3Sw9slOKlhjaBBREsbPLi0F+APuOIf0YpnljYeT97CIwwk7
Shq9VytcsusAci7tCA52New3sCHpYdplQo4ED8vUfyMYLDn8pJ9rfYFpxJ1o3LqxcQfWjKUequwX
qG4FwWDkBTcwPV5Ja3MM4P55xXbVYqAyWN3rHU8Wf3KgK+TbkVKpb3T/ok+dz3Rn0ZAETYJDDJCd
hh7HFkFNfhEnPcAgJtHTQTuHkDe4BwL8UJ7CPDZp2rXKUvlrMBs0I/S2A4NruL2YgY2ORTmPtbn1
kdOFIhRYly8UnL2fAWFDJw7fr5APpuP9/GPu5urhGjjOFisEv/TCRihxOvmKi/ICL14ICb5w9LUl
CjFwdSaGYzXYyXr82mhWVBobrHebD02O3eoX3LN+mrHkeEA8O4Ff/lXWReqLkQIdd6B6mYX5kUkk
ZxlVzY4AVtOlQb/x1Q8GG1H9xsxKaL+DynINxqCuNFIqGaKndqT0kRVTI1v4HSHogC9IFci0yyrb
UoDWfWsha2Ey4Pv05s6M5r6v+9NvZAidfh7Oc36uA5BSEn/bug6lfA6SNdm0mbmUdeXChkyt9A7O
9W5r7X9rbb9ft4d6nCX4yvS+0p12ut4AkAE7iyCVjETNlCv3Bqq6oMPUcgNU0jqqKNKc+CQnFwGu
+AYgYr6Pwu3ePzlCwzRtvf0uTOYUjXqoUNhG/4E1+dH2tzHXcy0nihoPr/WS/VI5cJjibkcLUFwp
U3y9U0kABisocLqgZUtCp4SHeLVN5e47G8rFheRg0m9Ese62ILCORyelVfLOlHev+7ybRTy+dxfk
QOMbs9DdCbGNhhO6kpGO0nDxan0eCUGW/ku5l/BiF7LmkUC7WdfvE8K2F65R2trjL2bIb+QRy/yZ
rL/ARSZwn77CussX2sP+IwGL5M9X3Z3sCG8v89jzW6sOvmZW2y+uXlsjVYAbHZWmh/8Y+vtAZ4bn
rBn1kRCdkvU1PZZx/3QNxq0azjkq4EC0pZiP8V9FcUvIDi9j7vvDi+YVs69V9HngH4z39azItLKp
WY29EL0wwGzv6S7uiuE85uLo7vYDpsbFcrT8a1Z5wi7yApIV6z1E2u/5+X7QVPafli1EdcOJMwIv
eCQ7/MMQ2CcMWdbSGRVpR8SBIKupa3KZ/obzwE6Gyg2NdJW3i5Qc4LG843A+9/RxsRlwkvUzzPE5
JqK3L4ogNKDj1k3bhgpCB+e8un6QTfw/AI1W43CxV+oHTftZsbsCy1+M1WfwD5RaLvrm+UGgiV2t
BRholUfstswXjYTAU3PiH+d/m1EqRSyMqLcRFh9eJYvBGnhSJYmCwALR6/p74HYwB35YwrP379WA
aIuuKpkYFLhwiLa6Jv44PNgTqyeWJ4CpRY1hjibyeB6yOtUUSqmMQIy26/7S6DoMM93G595P5d4w
gS4fsA5A5SNvBCQArrcsMF71B7o/CVuBrOwDNPGBmukXuYSz0cbJG61mCcJMxivFpfqkiFFMq7aU
MDXplkdSj4F/Iee3aUZsq6KNN8HCLTZ/SwEP20m9u/+b/VFD65VqwjjPdkYM9wOXSkGEpEWxMDQN
TZm2HsOjW2s+3sZi1r8SE04O2vnkXsrzvbpZhiXMV0q5WpZxsqjhuqBm7gpCb9fJ1VDe8K8RJpMe
scBRQi44m1hU+1RuP6kolml/0Xi+bmBJu7VgA+255iSX5nTXYWDe8CIdRSaecxqw7221B1ohKByt
Gu+P8lc5K5f3cv+wkgq9afi2PCE7V3hGv+aOgZgG2vt+OCL9BdvFRGrG7FoTb8Gx876s5DRpnhbX
wm6AXn5N2xopa5xVsmpq5WY/Z5A+0OmUw3ruHhmrdKmvwKJSZ1Fht4t870yn/wvJZ928pmTfoAba
mWOTh1Y0G21outCNKlXoTG9ioSricXfLhJmpB9/YbajpJDDtTbIaK7HEMsiNzddot0CySHI4ESaz
XhDPSaLY7U4FLpZLc6h3EaBjGbMNxYTX/ZnF4tCbI2H1BIGUNyAodOodjIp0+cSJNFfpekctK5YF
fjhqlNoja+BApwDMezo5+T73FqK3OS5DCO3F/580OnyCHAMLkqS4Rje3DlgpAWi0P0GzbfAQi3Fi
scBD8wpi9uyvkD201YU3ab9QbQcdicMUhh8mylTe6lkpYONjLgy1YIAqtFtzio0AnW2pt0W0YOZz
h91utAUIZyDZjBCPwGyAzha9vqDY5FAw9ak+rNHx0LEPc0GETJdge1NF+cm8muFx99O+PvkkiUrv
uLK3vigMVefsVE1ymVfaIahsF6g8aMHG305419qQ/WjAWTL3/IKF/LkQxFTf4O/oxLIDlK/eLNm9
zKlxF9Hp84cdTNY6KrA5q9aWuh+k+XRFaw6pGH9jIyLWw9L1ydMu5Lv7
`protect end_protected
