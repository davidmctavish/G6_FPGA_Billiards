`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HgA2IYn7DDAg50ZQXIF+3uF9LGQQ7iRnh9rRjI9Qf5gANpcevgVL1MizfVT7NKiRIjR25gpd/frh
i5ioFrwX9g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jGWna+ri4Ln5Ol4O2XYl54WWXvApiw4AQvHKyG5WPA/wG5gdYxJB5TsVgAEnuuZW8XaNRVTjEJ1g
xQEQ0pfMwvMIi5U6dbR13ZZNcJ6K5RD352bkLqoevz9cM6sx0mdobkv90Db/JxIGmA4NxmsNFJU5
OprkhndD6iP9cSc6xF8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dE09sW8rfEVKAE8tJxbijIBoKg5aImi/bwGIqMNMo00RGPg+oZMfI/MapbgagkM8cCe8OcVtZRES
JNvPFDz9zirNP3oDs2Tt5klGXNXOmV0H9wo8twnF8t+v2V0VOksCnwflqXn3kNmZ7gktK4yiZrUo
GVG9bpriTIEerq9osaZ9zFU4gNqRGXMTqOCkqnVKc+guoVUqmu68nXogrnzzpdA9iZQhEHM4eRqL
2cZbraX6UijVKuKZ98sS+y0q40tEseAiD9qQj5m/TTizJ8N+QVgEEUTB7YndGZ2+7nWBRj5upize
jwxV2AwuUJL/ohewELTaCEAH54sauhn3IsA9mQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vJFMkpaFUDrnI4gxuqkHmRkcal6RLTHDB5pKdGHAIKJW9lwXqRph65+R46SI7MCZBwm9XXsphpzY
tUBz6PT7VpCSG2rrI2JAPI4Gi8YMyRIIIhcBRcUACFKwtU5BGWGL1kQl2dGkVReJoHz5rMC08XIr
8lHI7RXdVL0RJLoKln4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jz3Mt6krjLr0CAySESYUYpmpNSb2dzpouEL8gBb7U15BOyU5048hkAwGgdP61H9LcXSnDSLG06Eb
YLCo2Mq+Be79txxWDS5LuqgwrpUmspI0vd0x/0SPc2pTWWU4sSPsuw3OSHlXP83bjxUgZLwrFEE+
CZ9S5e26tFirr7RDMOQrjTM9ngvsabDng0ByxKwSSG6141sLFDk3/PcDxlJX63JCw4W+o6cTzXn3
/EfJownOkIBmT3+tYE1QHW4CylG4rnSmq5s9IIoayec7Lhih22HyCiw0LXNg8055ZFcHBfuVlvHm
nNiN81PGoBCrXSWTmw5QGIQtLWxsuW4jfy/Ibg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
qx3N9tvAjRHZsKRahdsaaAsrBR9ILJH4cDbAr2QPBYz9ar1wVfVApd9CX5T4Xcly9H6zm2jFLK5s
zFHpgkhaTuyiuQUzdTc2Xp87TBrVKrRQbDqlaBl0xxP+vhgXMOhfCqg9vwvFxxdj3oh+5H3ncHUM
+yAXe7dPJJrQXPoJfoOsy0sClO2vKT07R6tqrRR+ois0uAL6jl3Z3v1GZpA4eD4cfk84fYMUSR+r
j995xf6ctXX+BaWn9T2emCGMgyMcJseKYIPcAZnB3SLJmdC555mbeST9HTakwLHA7VU0C2K4LbRh
dRZ1maxiq2kIe80DZoB4WL+7rg4Gs1DI9uoQ0J+alSQhuOGrytswPXLvKed4TwJWJIJYq+BP/nfb
7qNNugNySJNhctmGP/IcDt6zG7fT8tvb1myqJMfvWlum9ntarZPYRdfrdjHxfvDf4hdxIxANZucn
6CwA+6eFWaPh8wracLt2yiTcaP5jK30hoVg8SAWSNdmFu8tLvsBnLP8NUbi4AJFOXi2fMX3/SMjP
kA9k8u1JZriJc0Y/5l8lAdSBRo17i7JjWdrrHeOtbMn1KvhrV6Q0jK9gewbUWFmmFaFeTdd+BvlB
vywJBVwSWCcxTxST4ycKz2K2qruu38WzQ+m+cijgwpj5V6o0NY//607R0VfDnXmRpaPSKIDojzwp
2tGW8fY/z9MhdUoEbpau06E93SxAXSMwvM6E2Fxq5X7H6kktW/tvAtDBIRYAbzxx6hKU0F/+sSi7
pBFztVDBgD79ViTIwQbWirR/isUVRl3cu854XZO263UJGlvOQ3OqWFqzGX/LgTKV9BjYZi8mbH4X
UtgjjOZcADhBLA12ADpBhHS6i2uMogMFfljh4kLerMv3RT3MhVxJt+doOPEsi4PCMiXAAxHbXI/t
cNavdlsBr1NjmyHVVzQWtI9Mp8w8F10IRZzGZ+d3/Ife0OiIV/PZHu19RMX1z2pN+8Me+wMQ25NF
1l6a+tiBze8av7EmVT8An/65NkYjOz5TLevuCYkSu4NFxK+7FobMEwXa4R1nLX1fxCltWwzh7MAg
dAaH95yOU/hs3uEI7dVAc0QTiZDQpBTe6dF1EktO4WpC21E5IOw6jPTE9xkpGrj2DHyQe/e5CGD5
QcOk9lK/cfmS8NS5bkphR3kqgNZuk/GY8Wec344Glr3d9AdjYlH6c/T1sjpu1xcgrN7Gi1j6R22l
Gr2wnS8RwidzNs46uQY1otJe7B0GhRKWeOadkuP+SA/OeDC2DKG+N5FXArx0P8m3rnbCy6sm7M6+
QFtxqcwOUnsyzlie8xLWatAwGynqXWrcDeXNHfETPBxg1LN9dDZV12zsIw26u7KRmdAyp9OVI5Cb
4x4XcxVK/Bk7eK0951ZWUPtYzsYrd0ViPNiIvl2PmNUhTF7UbAjGAqP0zpBe/GjTC3wQmA0kmaQY
7jvufdWBeHAlm3LW4doeO3hLcjUzIIfzf5F5FyFUoJiH9LQNqU/WfJd4PS0TQfl86zU925bIl6jR
6LWF9IDDRwF/qdu3/BlhqerZIkPow8TXi9KeiSXvDHX5KrBbOfWKAnvsa/Dvcm+Pf24VU220X+PQ
JKM1H3bkzaXnjNkskkWcF7iUEzsMvRLomouZdj74bB7Kvj0XuxvHDK4wZzcv5GdmBxBno9PRwAT0
fW26m3GRUbZuGzipg38DxBuTeDajTAD67CWMYm5hJ8Ok8F/7jiVV70zOgNDNxrO0Xb/lTCABourS
6ZjsitiTXJwpLmuH27GHK2+4t2W5zK9hPRlwrU/UwwV6yINS0B0i1aeUH5g1Dc8Lj9HXcqfjuF3e
8D/TxFyhyntNAhKfQK5vpi6NrhVj1E6BuSLeImbmWV0xbLzxkuwMJm6Vo61WHqIrj36ynxwKojw8
3zg8p3uqbkvdI8YExhYjlwq1Yeggn8kuaB8VuptDLquyABupRIMExDkVJuv79cNX8iDFFBMMD7aA
uAJIPAjO5Hk9KBD8sVB1XTgiO4DlM7RbT4n1otzZCrb42m1IpgxVsClswHemCVrFgEAmSNcHFTVF
1rMRLJ4EYYBmJCjFn3EXV/8e7NpgVGB6ZVIthnBTBsY+Dxx84ZD4lTUhXFmBub08nsYT4O78F719
yKStNfkpkVw+nLxgtyGyT6GB19AoAdBJ27azqhqa64+OXZVcK3qTDVAuG4V3Bv3qXvrgo105jgNW
sS57R7hsUqZrJvXxCMmwyYhICMnOlboYIi1z6HBVclu6QbsrmMNbCAx0l6Ijgp5PewrIdqiSO7MX
B6YgUTL6KOmTyOw83z3A1a9aJRfU6Lbb9Ng9qBS1ZEWgsyTtMchKsu436AwUv33QRZONhYTT+XB/
Jugqpyu32kBkEHe+PnlmFS1W7TZBUkWvemqE7wpGFel9P83DNjM85/S3ovcdBmZbt66OhnWeAkCk
LA2Sa5FITIv25iqO8GeBuk/XxrOpr20kp1h1FBfmNxYU/kZDlxXyW/JQ/5FMIoTzBvIa8jwqYNX3
jXwlAEfS1IQsJzuC2StTvRegQ1VZC8S1TtKKdswKuXMavVxpCsrLeewJuA2h/zF95atBy8nthscZ
nqxmJNEF8FO2dhHzjZzjySU1I587znlsd9A3JJxB2k8ORU4td3tRQDJUWl9s1CaglGFhoHU9p5yE
o4K57dEiDaTO0ZQQRnqogyz4gYeJ+/zjKZ4Q/CKhbhSnfzcB2ATk8f4DOlx1uzaPXdE45x718F7t
nhZSOXATvMUjf4l6fGKwvN8GbJtrKt03lz5VpY7ZnSiM7S8c/DlX4UOEn/vCxzsJ1DWDOLf40G5Q
hawM/e941GwUn/Uxt4bM9qBwJFcuBHcgi20dfzde+uQzMJlw6zQvDG8blwfaBov+1cCh9VZo7VC5
ujfEnaaJ1zB0HGGIMV1iF+eqmsrQksZslz1gv+7BuX+WKCu8nW5aYTHMb3V9F95K39bjA0AnnXIV
tR0uC8U7ex3c82tOQIVink69EtV8b1EXTE1sumyGSk6j/NfKK3OXOzSHa9WR5OVSPyinfj48AUa6
fj6QUjnvBt3qWnLlWQjgMPF+M7yjTrcdpMrGY6OWwYQPHl1Lh4aqX3b3K9VG4z9/aI0K606p+asQ
A2o52LZOpPsmJwhgA4kO7rYLCTIhzTCY4drExrkX8kJHWhBGv+elymJiwtvyyugyiER3NcT+gTcQ
go73Hy6jC0k5c5xRROxYt+Kd3t43/O37+yYBQGf3LBSh7tor5Iw9ungx1Fmw6JWpEeC6UKy10rC2
uE7Ni6g5yubOhs5ND+N8mpzJrQlmz0gqxR/nnxHMgJZgVXTvdbHerw1qQc+zz0fYJED73mgiizHj
au4Z/ac4/mgHHsv5RO/9oIdbDWA9oj9jqAZHuYacGrmVoPIiK7VkHlXI89IKHpVO+Ymbdk/EEJMm
ShpICNyrkbnFrV+oR5hWNOblbSQyyIm0eCZpaVK3iZtAyAHqDtsHKjSiUAge/tDTv7kAhMn18I7V
Hh9eoE5UFzlKyZ79OkSeiIJUuizbV5LlwB0CArKBZnGjnH2EW0wkToINdMAy/gbBEwb3wXHhech2
z1lTkjsfjCSAOWYwjU7vZgHlERLx05GajOu+7EXxBdwwnov1qmoyyMxbzhQfFDF9WeOiaABukyJk
0gSSzMSS1RHarf3qBDB2cdu/1CBS6HF8gYzqbB3iuxd51wmRPRaiEQK7YOlzsxeZUAojyv0hhVA3
qIh32KYJqwHSNkYWAnmSYK7ZDnJ1on2yrdqjGmH3bHbNGHelIt5ipkG2gJkhG+32gPbE972WFfe9
fxYjnR8DmhBEhBmqU9pPTJc7sewe1OuQbZGDw/kQhjaJetG/MKiA1uuKGAheY2bQNFLUTX1quRTy
UcYeoZDXOaUDhX+Py0EIVcWk1GhwJSUmHT5XC9H6CKAMr6rerpi0Son9/vmlqEaoxlCibtfbwMBX
DIu4/YxIBG5bFUsoQNR+KCJxCsIlukY+b0he/I5dDbf9HiTwgMikTZkzwxyFcR9WaBphG9o4N70m
RmuMNExx3/ImyftwJu9QPE0cZdSQ5FLvpe+nSAsaSHmfEZhovm3LIsupgETHKr2fIrEvbvD5JUVX
bi9TRssIVgTGe4L3dK4J5Is668V2KWy3rsWfs0Sk7dICUYyE17xTcnLlgXWMQkuHWk48yLSmU8JH
1S8UF2Hx0LBwEV7jiT2W+8m57U4k7exetyR3XIYp5uAecH/V2mLc8LT5quiQvCkBu0nYxNlh1C/r
YHln+IGXqL5i04VGJH4NUYk8B2AwmhBEGYSEAViQXsFwTXrijddOct8fT7i+ygLGZGjauGZnoPgh
ISKw4UQALyetbeDMQxb9k3nIrCr+Vi9rO/PMpL8Ul8Tma4QynCHzQwTbqv20U904wuSHjoNsnDXK
+zcS69vi2gROb0qPkadk2T11+SqAx2rvVkDj/SH37+GfDcagmLViKEjtiig9kqBrVDhrbCVx3FR/
80TT6KUAgpkgnhJGylJwkF/dmjXsiD/0P+MM24j8+XpI0Gd4i1eLWSt6SZU4xOHjABzQnpqOM9bS
rp8OnPdvPIsbs5+fUCDaAjUD8RwAXTb1L3TOb+PA4bkQkH7jYk/LD7PZ32/PSinankQraKFiJVpx
MB77nX6EVbbYLGqlAi+VmDrdMiLWysmYIwPZvTgVhdm1d8ZT4si08BSuO8A2+i5cQMoFBj/d47j0
bO2kntewUIHHKupVH/aNxtw7fAU/MhSeessMVP62SY1zeqhZU3kWEVpqzZZ43rF8PFMAFb43nvBv
0FSuElOk+7u6K5MHO0u09Q6/2g/wO/kft4S0XchSIFmSpa0zr1PU2y14NoD0oFDoaFydsx4vmovk
nx0O4dQUmf9BeI9lUncv1lQ1F+jTfGQk1g7K2DhT0gQtlhTgP9sSXcXvwaWhJa/v+gYoTa7RgpVH
TLIn08F8ubz0aMNL4X51ol060eeLB2HxdAn0+STX3XBm5uME4Jj4Xp19wxCSlbGbochRi4DrJ72E
gb5z2kpFnKItUgjXdlL9nFddhJfp6ZqfiAvcCcGX40CkA+WnXsAJIad8QnOnI3ARvdSMIzZqd0nb
GIwblfVkBwD0tQs/2+8r8Ovw++squNWADndy11Ks/9qosFC72N5BToO5s88PukW7lmCvkUz2jDv5
v7HBJ5Gulv1YIvqu9/T3IvwZRVII90uilUbsjvOOrOvoBJ3ajE2rRUZ6SM5FfCy5k0M838cCCsiA
UK1mr7pO4CjKtpuHD+ScAdowzb21Li/cranMT5RPolPAbesD9/z2NgSwMGSLJnrcxlr2XQUSFcWh
Sj1yhSGqJvoo2Jx6S2bgFKO6tBSNoWTpxB0=
`protect end_protected
