`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TesOEhveIGXmLY9MB6Nd356LpcutXfRax0YWtsFjcHaBAdMTItbmZYXbhtjUdYTyqU/g/cLu0zrs
CjD6kNv14w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MOKL/vvi6+byokG8VdTkvaq0n0RXaRoGpLhgL3Er9X6ZUQBbcu1UNq492dtEtCzLHhEd7zAE0rcL
QMm/nHgVwWvfyr6vbRq6uK4OeGJCsRJ+R8ql+CzN+BQuSR4aKLciKEgW/Lt56XJvpYWV+esSlN0z
sQGhs2zQTaR5zVqpEsk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q35NfcTJ5Rfa9Nwlen86X4Qu5qPti8pQm1uZCccb3/R1R59dckaqUrP6OHVgzDWJwVmA/jq7/aZ7
ED7w3Na7gQg7AkwP+FocBv1HMBU33Fjwji6pUNb1715H4bIMIObcmZCi4R7NW4sBiNGbYBe32rLx
l56QVlTBpZUyh/Qs7R6EEWgsVjCC6zVcqsl8ROs8lTHcUGG+bJMWBzBHx94W4iC8a78sRUCyxy4U
LocZbOD85Klu9fRPT4ZQSbLgJ6+z9F/gYO6SXXU4oizDR+D9TT+qT0X2TzsO/U0caX60WI5hsLfv
Gapla0a420FvLl81b9pFvO5AzpyCYfT1uszOXQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
r4Rc2odin9JujFSAKz9V5+dxfMS+GZULOeBqUgWDUJ+fWwQmCeWKDrNsUpR2rdWOCaG4D74oiBzw
muXiYRkbgyCU4o9sNzDvVTXcUiI2qOV3dB9Zc753JdABcYjxP5+IcpgOYN3XeYJQ6bCuFB94ytJq
ILYOpZTYnwtL0xg1gXU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NavOPafGh+rDhmrBhO9Qq6OgTYiCpjkCMSWXPdlAzEcx5FPUA3vjWT/H3MWKlpBc9Gp8/lKAcBHm
FoH/+QXFytsnAw8PTM7Ti0KjV4v0OHCwYkds9ch1QW0EM/ujx+4+eOXHHA+LZ8Rojx74i/V4MpPD
AXK/2In9qqSDxsOCv7MSPI1c/LPSWURscvA7NPEeyEPBvykLrQ/FssHCCuI015ac0C1jCRH7dARy
qrfl9T/+WDHPYjHW9c3tXrRrV4wdRBqMmLmIXkpwe5Y0hd4ULbfpMwrnzcfoKQ8AVDC+zwzU7DPQ
pyLoOtkLZKBqfBKePe0DhaAqYdWVyNykKKICdw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16848)
`protect data_block
/g7fTg2AyPuZMGv6mvyp6x4+cVcvKAMZmSh0r1UwTefni+MUdlBJ5hWiuIjLoaMdhzt7x5KzTnGZ
RP/GP1CCIYtjQNYagbv8g+XakUVlhoL+yNwQQ+b3I2fT/9s/mYBnL5wvSVxO7VnWX2xogJgUY26k
PE2ErZAW4ov8LgpAGWEY88fbDYk11ybrFTJ4ch2Ya4IkeOLAz+LXqyUNt/JbP+tBxA3t/sdb6KMC
VV6CQK3Lx22o1vxSGtmQ507nPbi0lOYsEXSpBb0ahFg/xi8zGNOUk8HhpQuwIH0bju3k2Ag/beSH
ShrNroeZwr0tiIgDkLLL9TtUqPAKLJEvsMAL9RVkmBlwG08hrv412Itwo850NUUltBpuauB5nKYN
m+VupoA2QXfYTw/lrTUNs1aev8WOLo1LHhjZWfQQ5XyDRDkOH5o1LIIybmhEbnqGyz17H9YkY65U
ZWhRlDAc+UA3tSpBa8y1ZRwCJlEcZZX1K3NQ2rp8bU4b/WedCjobM8Gbq5WQswsnHeWgDGckxFeJ
7iAf4eUbNvPMu6VvWhk0FNMsE8ut0czsTo7G/jchX6JF9yuvnaNe8Il58BAhxrbuIew8KAFWq69A
AkoJP1mumlqYuiX56HW5nV5fv6cih2UqHBRDiuKid5PwDylhHXxvIIjdkCz73c1i8w6TzazBqtFW
aidogjxDLQB1yREfoSOqvmfH67qW4mD6TvsASCmx+w86Td1c03GztDB2O4ucv3io1+gTonatUSb4
nbN9h3kdDFn/KSCz4CyDwZ93HZYhVgDrZjEmcTGFEdKQASqSgSyTto9ug2d2vux2W064TWvNvtud
ORe4GvaMP/vJJvMlsDdaag1xfNS9SCEzA34PWuE3/2cxut68XX0YYzBSGjs89E9ZsIYqtzSo5JdU
uHYbmOqoYaGMImNCYLdmu0HpfSmpV9osiS/ALfuWDWbPjAr7wriWcvXKWs0Kwv9XK6IemVgzsIHC
Q8O01rYLtrnRrdZHVNfFRi9YOPafQfNDhYzZ8lFJArBAe6gaj8TBV6rrHGAqxwx0+/f67rrZQ7hz
HwkM54BSJ9/mB+pFTQL9D/ybSK0/1uLl6Vm0hBU83v1KXgWIaNags+n8VZ64EBcfwkYljvOW8Dye
wdoVAi2eylK7jNvqcFsDqwbp03wqE3hHeqxelYAyCtdpTYGUoP4OUWVzq7wVYv2MNPDhXRbXgxHx
2T1FGDsK0xLHNSU+FEgMc7B6+9zvEhqJAH4WU01XJluEh3J0w6iT+M4Aw1LnlvlZtyJy3GaMj3aV
EGIR/7Th+FHQSZa4KDjIz5RiDcTfGIzBEPVnlnP6n3M9y9CFgsbQwE5bl+lC82HHBZKyjdjSYkOZ
a6fTDhCmQ8S1p6YY5+hoKTgWw6Aho8WoPfkCrXgvjrSPyNWQuijIwEuUpcHmtoB/oqzMs3cG+NjD
9RH6pFm1LARV9Bba2IfvXtwAGtGT0U5P8KSUZJzi4NMgffDt0M+PE+UItDhwSY9SpiG9hQ9Yj8AP
gw5oVM8Uk5oUCpBWz3nS6gvJ/iJkU8Ex/prAXcfxNuC3ars2XexnUDXdEg05cTXo9+1U7AL5kA7k
PljtRD4uRNqjlhix7EOYp0nC0VvWsGXhloEnmtcPr7sjIuhX25EtNYbl8s36EI23qGO69rgKYgRj
yxdQLoOkrEYanCNzQbAR7NlPSYROpwbwh1e9niqoLWzW2LyM6hK/i3+fFAIs3veKLdNRltlxV5O1
RcEHENXVPmLWcl9BdxC2/+mBuTIC7JtD1FkE4frawpDZ9RVMn7srrCVSCRmugAeqvTgUmsTY5ABv
w8yqXam9NhK9V8TMmCC1Z/AdrL+X0JgSx/uHTEmfPKx9MxHCcugtbQ/4HPWPSUdL3lrzdaej5wXm
BEPX961yGA6AEOz/SXVJSg3X8q1NcPnMljSf40f6ktuQJWB7yrkT5J9rTdj1ijEfzfjKR0/AlLX/
wJASt/EkYeQjJzfFkcYuD7UCtk0h65nX9+bocbhmuwi2FyNtFnwf+zr2FeKfcdb4qPk5qjDgmTWL
DfvR6qCEXX+OuXr+4Oi4fdHd6yKMk5yZHj7pgGxBFx5WMQ/Vuv5Me4IDOsrH3rnrLOWt6G/Qwh19
Y3NkZVD2pFNL23fxd2JAQ6kASZ0RqBkl/OmMMGF00wozHPeALS3Y+oPsxZ4atMpjni2Zsf3RF+bK
oWQnBVv5YhCfcETn6sjKDqgQkHnLjyu85YasOWnsd6NxXM4a6XNKHtqCN1llOLrpnloMizILtSUb
mTqziII5L0uT4swczPglCdzFSF1LSN+c0TRokiMNJgwed1tpUTo2sYj3AKtzddhjDpssLfqVJi/q
nO8wpEToSxj/zsb3CRfKBywmm/1KsHoGqCqUte+PMRJ6Mjz9DFyIcqLjgPRqsRicdrh7inNUt8ej
lsXj98MWwrIuhcB/0oypRSED9qpwvxExsqQZUhnFSb+AJDPR4DyNInW5kPLV5G9XgYFVGNaW7wzB
d3vWlvZykflPXflx9L3WJO0VpGO7WYt/gkwLso0b6qt3Jq1nKfkm00Exz6YYST8eSfLtmXmPu+3O
fvTmxQ5XvYImwnqSZLCclMA4yUUGzakmqjT9OkCXIHsCUjkPrZ3bZzabkT1i2O0bt7IdySx/lLMI
nbEXUhqQi0ciewlcax7NbV9slmjOfW+0soxx7VFHUAEmtuB4nwsPsbGOp4/gb2SkrAzTOlEnbmKY
DATp7w6GurI7jur0hXOETn+2pXra6no5w4YGHSsTQhpKEgl76ysy/heahjMQ6S/pbhpBvDp5QN2l
XuFUeD4yV/1PXPsjflLwQn+HTnunRK1evV0Pb2/Vx7ZTHevUfaTXrooJ+V10aRxONvmFg09V62QB
KS7eC00RQH+s/zdurd92XQr4ngAL8MPoPdUC1/iFdPT0IqCte0mPYjxVRwT7QA57x2CcEJc3Oh1r
kkgXaMNggD1DkZarLsm+BLwwOruT+Her35TA/0A6n/KhFcagaVaWId7iEf6FCfHp2uSCI1WEdzAg
5aThy2ValprM3Ymcf5GIDuy8uRK7W7pwXoz2MgOEgDNyAlUhWIXd9Cgtd3KAwI3mZrM/N+HeiOBd
LwlARf5A7s6v4DLeO2BgHrb6Ccu2uwATYXB7cADBYIX0uYRxANdoRNZEuys7c+n0AEyIxQqwOJmu
UaX+pSrND0w9THVDcOOo9iH1JV846LeX2upcKBY9rlyZJ1r6Kl442evwOhT7QA0aphZsP6S6fp3u
gVr67dZYnE4k8IVLO8L1GhHoa6Jpqwr9+AX5Rtra4N12proRkD387fgfCVkTh0x0EoNACahEvAF1
tgZJHrdkI6hd4wHnKGR+9pI/GU4zCaBK4W5VnvY8eZ0H6cL3Ib1L22EElZCQROtn32vjuQ8bQoYw
vCEg4F1Gpo11MBIyFXi7w70N1SoYdrDUUAQshgQAzWjoAXjQ1LLPJZDmwkp9i+I7fwHr0FZf1HMr
hVnLnhqtMyJDCjjbOOQep2jzvu/uK2Odmrcq1FLHeuODoNU7gbjbHL3qg7K7VjaWmTpt60WT9tqz
fAnIoTgK7aeY6wu3VZwjPllS9sowO8Q7feQv1IPQI6hlJ9CIJmWruVoDhxH5b6K/Ml+4j+vb0C3u
GGlTd/RSWdJcREOAK+7vRlo77bqw8FSHkhjyw8Nrb+qKIiQTm2PeueXI/5EZhRvFHZO03LB0BIXf
uWHBFMNrZDZevoy1yKsmdmeYOca8mXBwXXoPuHEfwl2XJZqseMkoBLWmdreaXfrPvsFAapkhfduP
5mTHFA9OiGFmfsPkESP5mavltNHj0UTupnnOIfyTBJJ2nWta2cc5NWc7h37aFVMLk6Nljh2O2glS
2I1/8SPjz8WklAoKaYTMGnKYF/xXXsEd5TGRhjQxoEFKuz38rBSitqujeJpCrqdDkhBgDsO3Yd8c
adWc2qHRS7ThZf1PYxAEPIR1jnv1oQA3cwboVDxJBSXej8nrM9KVw6oqmJqRglv4pZXbpdSYRGKq
rnxcApPSUY6BwUM8UkeBzh1KfHGFdymlb1O0wW/bsQYcdGbwMGTrvmKYouHPpEw7byH7It7hKaq1
QJ5rG8UfmuhVdMj9x0lrM/mxBigr8mLFWHjkMHHlAAY7kecgicRmGb7Ji16/v3YRF487PXXPq+Di
dKSAJkuN/e5zMrTBbX8LZ3azq0jQ4n578kJn2ChkJcGoEmqdykxLXxM9A8tPbm/WIe4a96aoH8SK
Sl35odRzYY822GxFIqXqwKdluftC9xeNc5TNWu7NSnZaWcIdSUcOQbxaTQCk6Yptb3ry4LfEowzi
q6CFm4zwZbIXN+jbswHWpZLgGLLZwD6tlEJ013h2ky86fsiAfAy9yQqu9IjqA/v+mo+AsABMoio0
az+uzmV88JBN9Su5ubbzBAoOmFIiS8zYG22igmD165H9yLmnXu/Y/7izfRfCp9K0zbiRFCcjn1Pa
vQG6q9qDj/ZAFNIjZjxG75nOE9l87KwU0tdger/T6v65C8FNjybk3LwXGGSWJrPx9qdgs/bvlBH6
eBGDo4BMCgRhRtpRdZb+42zo3nXqsgffnYaHJ33NRh9j+X4uF6ysAGD5QWdtbUMGy5B5C9Hh2Qhf
7N6bbUXESOabky4puYsLxyqOkvjOpiHxvKIBt9oWOvPoS3BLUePoVXygL4OkxWw4rnpHycJqiZM/
uEBCki1ajhnpNs7qrHveLUxNdRHKIpiqOOFXvmq5PCi+6HQhpfLdtzyWtAyb7AW5/KpI/cO1VbOa
F5h5lklmn+iVLqUCNubsFGg+Mx2bUPnWTh8KjpAVc56+WCO0E6Ag/ldkHU/T1PbC2R9HbTvaqfTg
+yJ0hXNxJczbDfoK4ySLhWGAY4sqAkz7HG4l00XnwTBbS7qrli1izM3cve7Lu50Ue8UCd8lf3DPk
Yr/Awmj2Yn1d1pmG21gWXDwIxdcGRGH2kHPm5vsc2K3W3vXQdurufusOAjvMbIRumQej6oH8AoZy
OY5r8xL+ngUps/+h3aPBhy8UX1GEraoQneoc0HHgb9n1lrFv6/By/OccfwZJfxdGzkX7HMg6ljil
mPueL8RVeTvRo6zQUmHytEy7QzQJzuSVn9Vr3/tVcdntQrrTr3Meeo9pEMLIqxWjNsHlUZg/cYyC
ogpDfhJUs5ENVLOvUVU2g/O6fWa+gpGhRbCECWLIyqX3jznNq9S9HJF8hGiCpX6236uprhehYfW3
B0oU4z9qPwHl8abGZKTtrCx0Rb2Q2mbD8WL3Coz6zcnDWFluOGkKH0fijAMJSllXTZYlVj6MA9gi
Vjr8nsmGV+aS88aYvSiAJEugCBsvhRyZzJ5nhePlrcxgxOXYaP8H7GKlmF3a6XdCVhiYH42gvu0D
/SRFdIksqRZeShtMwbYBFnVkSOEaUoqH1ZIUVgNXIeG9K+f6rIkf2OCKmc1sECr17rIl11/xqjvc
MRvvGw4HfmhDxIAMCGKFaiWCtHxp9/x/3OCebHofJhjLK42b9mJCaPWf2+kjMZ4JxoxSBo2xZAhB
i2+ikFXOXCUoYnYyrHoSeFqClPWjCC732FZQEIswhtrVAA+RSbYeacHbaX2F2rtyB8vEy+aBVORm
ReRYtmZCrHl8vX8l3E+id+3N/kPDcxlZXZmuoPic/74VB+IWh+S7/d+83FGJ08vlOCL0sfDUw5co
FJOUpzSGjfJb7ksLjvArYlJPxyQu0hPD98A31433dhD+ibd70/Lo/oWHb3fmRpe00HGZ8LHBcAs2
FpFdwaww4h/9dkcqhCsA767pF5BmP8VYuqrbLTaph6IECfeTRMCV6W+HwPgftZUnxuKBLWwmKRSr
kDLKb/v06H+hMujxh6+9imZDqQDsWcdx00/9ACYPaCR70mIagyPjeIaBiE/XzFpA7uVqrEEca4eq
JO0zl7AJ8ucImY8uGqGlo8n8j70wPG7ilAVgo3AtPxqWsUZJ9m4yGc16Rd9ota5l1kIo9ROjR1AK
yzdHGyC/T2BDpQr/eQbRIMe0h/GOoREMRBKZ654zwXNTq5JQydCxWD+ehqYwspwzBALQDuDXhajY
95XmtXcz4rLzeFSBLoeZPiis3XYX3ob28xWqVy4IZHrgEWkTGTS8DCMoSdXik/ZyVphcx/JiqBZ8
4ydnSEfv7vKxMYXHIdEbYzvwk3Bktzo12mphuLvHm0vEEiLVifLGVo0WVZVtDy3hUodbFAxpJSA9
32fVT04K9ZnnmC3zZA3kM8sKMik2P1hTz7T5t01wru9ofDb+3bQbHI31jOWV9Gz3uhJLU9XLZCo5
YrIYhGHvlXQqaw2nrXNjy3LLkndpNqGO8WMXG+AcmF47As09LFiSETBt6OYhN84GTfTvTC67fd7F
9G7qfkY+NbDnRqhpd1tHlwwObk1tQ5U+wuZWgk0FoB2EhsCtCb0uWJJDth90qlGgYUCR4/RaEAGq
OoEQtGICl80LSjtBM/ggtk5Chl2cvOwsmHSPtPui4X4MYqgy21b4bYHBq+GcTuC1AJYZh4MszJZA
vk89fA7gdn88EVQnlcSnQEr+0nyv/0oo1z/csX+s86FBk7l3ypEscvwZr4Tff042AkoJN+wPHFyA
qlebb5OqfMvCOm6ScsTC5U9eBs6zDUnQo7zkoepM+TqbsYTs/WONBl+9uaFiU0TF6kB/Ii0Kq8f6
YCCVti7iu1IcLXHOWjNSloPGjWqPAsOOZYicse/l7e0wYz7GWF9ZmcJbVv9GdX2DXrrIt+gg8+fR
9c07FoytxWkUKb/B07AI6hhjmj5V+d1PgCu0EI61Wt0ZrcSqa3t5Uq8SZ3cjMdGMKJEjrQxIiQEk
lLkZ60b8R6ltGM2hNcY+xJDSKWEuL16jztn9GVetK4wk5+p6O69+eP9Nit0f1WyUsjB7wmgRz4jB
94OhDsLL/TZ8gns3J/7aIdRYTQvvtpn6DBcsAr0iAHVqFdoPISgvBcPYckVthgElXk/XxcPpkvaQ
dnDYnfzN+7Tlg9DRau+iSADGM9K9rx+mUqG6E9EqHOGYO1WQFeLW5UOJuLWJwi+JIPLBwebBXwDq
b+yWKG+W4ERIRMVXaRTC8mMsnUuotkXpULOAh/fWCfGZWVQMpWhc6ZvzPrXzJomvgA4qEoeELyqP
NTyLrGsy1TMYO+7v1nSxsdbFRb/0w5bsxo1MqWG4YFkzhYHN0u19Qp1wA3w6gA+43FGF/Z4mUhWb
MMDdnbvRHM1+hWvNhwHrfYVp6aUoyMZ+0rhbueDOxEaAR1F+giVddeJDFbC7gQUZgqGLaXOUYjSW
4obE5S4j3DxMG4dkQPr0rdyZBa1TRzWI2rjxGa3RsSA6XhI5IavQqp2D/xam53Et4qlatgbWaLm0
u8UpREuUGcJxvPft8OW8lkvcs1KaYrgTgtfnwTU6VK/kWTQkXuNiVwBbCMrAf91yo/Sp6u0OYNNG
IgbqIS/JN+LDPPoBonTAN2DvAVeZI76AxrflxwlkMB/On9fWiPuOLkLuj8+xjVj3sx/hznRHfXfi
o6JrK/i5GiUYLH12i05QQrRAQcMlGJ9L9zauA9JJ8urKD4YVTv0oEG9q/KOyA4BAhkhDEE8eSEEp
fWIZXFvkQwkZOIxk2DR52d4Xk7d4t5cX9A4+OALT2Jjd4AmTtdJ6iBrp6mruEeqL2ajXJ3NNVV1x
3mE3p0TkXndL7wMpW40mzwKuPe/gX6WKGc/L596hJRBhUCJDj6ptX+k6qXc8mTFThxgh62Mm1EhN
CXhrqDkDebLJ+TZikSft85BSRomGLT13qjvgkurccJTX1jR6+SDeC1flN4gJ/UuLaLME8lsoorJm
IvcuutWDxTl9su66i/5zb8YoX3C1IUZi8nY7gALeGAmxwvUZrgGAtWLR1mGbYgCMoHejGfgHd1J9
pHagUILAkWIlkg8lZ9kwO/Ecy6na5O9ly0SZg7Z8vU1dUU5y7OFOfTHHoaztn3peFJMvlgC+H4Y9
5y6Ui2UJ5VCxizq3UEr3uSExGTBnpnH5bc/KMtF0b/8a9ubGNDRqbWOqS+loE9izT24FQtoE9POZ
VJhoGdTJuhsS59v1M3AGeDfatChNJMWDn9CQ2AMTn9xX5TFEc6K09G1d+GBlEbOsw27wNFQqcAfU
IaBMY+ZnJQyJ59gps0k/I7Tb55GTLnIryFBNLOBMBq1KVk2BbqYLXV5QnycrQcO/GKheurMLW2Dt
XuYdLbMlgZdi1YEVXdr1att3QG4SSqk5NfLeDVBtdreICLfwuNVkAAHy70Ny3ScQQbVgnFh+IG4R
H3w1xY3oWCptNgKuAETgBCDA0lfRUkoaIHxpi8bk7Vt+HPQzkFXorrQX2brk9yPs23tJmlig50M2
6Y2K/P6hAx1SCmSlPhDgMMZPs+vpYXw72bWHeDSuCrdEZp9DVtg7cQvxjoIisCYruCIocvGLvkwi
mV95cTolcF06cFBIiqtzYtZbWGNFdvbOOoxBY6Xbb8VxuUi+1YvDzqZn8Ygq47VkXggJxZNbtcsP
Li/nkXoYV5sRd/EDeaVlCHet/1RB0B7epXJjM3SLfHB3z8Gy0JpfQBfi+xVybePLUt2oAOdZcA9U
/pxSPAZ0ATbEJVlnIPC30ec6tMk1je71n1KI1J+lAbalN8DbSOfx8o8e4RN1Ur3yPrns3GLd6dfl
YLuLNcOmFWk3U5JDXLPNQRgouzO54OoiqwMrJOWVeffkwcEeH38z30MPgYPjfLr3e2Jctb05HxbP
PFTvj03kUJKBjWLdvWP0EGf9jiKLxknuoNFxerJXIvGhg85kS2HSR20nphZjX4Jt48G8J3TKfVSa
ucjVCxWzgtD7zhzowkOY/dnvg0CPkhONNUBdan/uUjvhAFShI3bp9Kt7/uuWdfSrY+5LkgksTy6j
DmuVQ+UYniNE+nh0xSY5X90tAwJkzPjelTnSdE+pnmWfSc4XAaD0oc6/Bi2KEdFEGkP0+xRyGjMV
+gmITkY47xnCL2J1sFY34bj6gFvqRp2mvsUINq6+UVqXEHkjN3CYQc7NpHKW/BhTH94oOgmN5+AZ
UtnShIkYKae1xJcGFgtGgog3rejHmF4UUKsxECuv5+kUE3HqslxEZTNV2q26biQqmo2r7aVMsyZh
XVEP9iImBrTePsUMeT/cBUAhZsIoUjJy4zBDSgzu95rrubmA0VoNovVlTUknUfG4WY0ijD22d+bS
TgRHmkKAI6o6vnYTOBqHtJcMK9XB6wH3IHEzEqqrq8xeov2kHbtwNcXOp2zFMZg3YWGntAvB8a59
QIVtMrWnN/RzCjTrcbZIynKq/Uj1xyWCzakgPAaLudYys4zGQQHTzMzPMXN89It0rM0xmwH5A0Dh
Q5XfPfbi9xqhLAuw8GxN0avdRJPtuvej6PaxXLZuwGTC/LOPfdMLJnQnmGmuG4y52Ggql+/D61xn
uVJJlpa02jP37C6189zeFogV0vsbopH03VOQyGd7NkOn1YkFUOAwVE+yEeEtD4+F5+hAzcfXZwz6
PZjktFNSNybQZqvs6/wTQt1aOoBwyhntYaid+d0z23x+OU9Put/53tfJer3zb3cTcrpobVHmF2Yo
lJhuHywr9HkAeObaz5cEXJpwlRQqmW6R2JmT4gCedFM1t35KuTic69qYuRdnVDK3rnXF+OwCalTQ
kPeP3qhiIycPdozdcmgWC8EnvNnGo4466P6pFsJx81KvhovPJFVRyNP3bA7Yo2Sv/BVuTt4244xH
wi/3eU3YD+YDfdN41jM+Y9TBp4sfzB9IqSYL42BIP143cBL9aTNSkwNG09EhWHjT8NEsXjok0rPT
z/i7+yAQxerks/t3XWcNsGs4H9gEdRSVsFYgIHpbHhsdbq+M+RMZW/jLtl9U+Myl+mUezL9Lh3iy
ivxUyuBHdiUmPZWTnmbVnFoF/pgCw+yPTSlWY2HKLoXr9/9UPWskBRp/QVZfjyXwEDEjujkIREoO
eEwiOac4aWCGJCha1AlHj3Wi/5UmVNQ7duONX5DBg4T++jUswVPwykpMEPEfMIoYosNWtabQEVSP
2TM4lJxYVNUfH9x7XgTNxqRXf36WA7rubSHkb1QWR0gSZpGbBqUzevb2SnIUUcKNLRtB6wETqJZd
Wplytm2tc2ZN0K2dEyNeNtqiPw+GBQZ/fyfcJ6CEy4hYzIA4TD6t99+SAAwiosRnT44/qCQBbeCR
Xf+GABEj5wgZE6NxqGlBkU+RY1WH0SXkIA1Gs6Fhh4Nv6N15zgUMwmYbmCaRhVMoT8dQyFgVS3m2
04cFdrDy9HxVCs2CVi2MSMqvptq8aLchQGnlNVOPbycq8ElA9s5H4R46o6fWH5i2mT+BVaM0KbpA
cbhhKLW+vhJoKs6JjTHFYBYXf9nSmYO+0Xw7c/olBLsU8MOIaaAK/uVKMaEU2XkSU5mBQ0zRDKhC
j5nd5MDHnxVH8PKov6ErfxsiuIE6/CW6Uvc20KuSed9M1jHBIPFM7QMZIYq4GkpVI9UOyT9htJwt
ug4g/VUy0KkSiVCVskYMZQlrG13TZAOSVr/9Jr4PNHKXWcopRmcEnw705mhji4quQbSEZsJm/Uih
oiYGvpelpNicMkaryN2y6lG2QdRS2cFdUv8NznSYcYY8P3W4hh8BxvWtO4nhNbqAYdNDfS2LXS+S
TijqJ2qw98000q9X0cUBxci+G2I5SKLbJ6E1uQSabjXHWGfOUeKVPq0/OJ07F6EMXjzC/fNsxljh
Xil0zb3J3VUD7Dhs6+McgZ4mNxWgEmPhHWHFRHJ+p+mYFsmwvykk7kcJgQT8U/ynDnINSdmPjsrb
I6Hc4BpXch5Fuaq+kc484ikbVLVHftxP4e3qW4ktnOZLftj8jIMmBwgA5uQIQ9CIsXmUMEllwAm+
es1rh9Twuw/HsiRDeTAkpz8Y3ymFpQ1O1FUiENdXrIenzZspfb+/Qetm3Ibez620Ayd9+KqGYAbF
/OBiFZOcFWdY8k+9yUg95eAv4x3nUOeShtb21ASu1941hgvP3xS5LC9NJ2E5NvscMPKYl2JOm7Ht
HaN5k8xw5FWhL8Mx3c2vyWKjWpPgOCkV34GQM1TCeu6nbUUJ1F4EERfsNicqtMN4631W9OEb1RAk
fDeWfnPD5lZD0RiaQIH08GwsjzqD2d4mah6nSwiTR42qqbpZkqtPBT3KRjYEWNIanY03Ycnbl3i/
ZGMXp3fqj+0NDXjVMM/sW2U40T+MC5NJQNzI64QUbk/P4rCMYmVioYmUpgCp7hkaCmTb8EISPIsi
tOlW+fVFAEP+9Dp9njD4sPexLCV8FAdlnGhqxp3Ko66fX4j12b3W9oZoT4RTg7ncPj1agoBAIorx
WqyrIQiSmNvkE+wuH/hrMYKmsFqo4qkhu5McgSLAOkbDUOerncMH1yCHDBWGTLzgV7KAbfSIl4SL
zh0ZlNFOhDS1MU6PIL3EGDa1yL/B/voUoUdfCp4FmdAzN+Ri9df8aw0VrR/xeJVSf4eQU7DnKQAB
ucLHBl12QskISwt1bUbQ+PH0suGKsfmIEH2x4Y7OHY4uJNXhdq2YMf7hj92pMPav6aeLPX1PBdyO
ecQAhamp1MP+grfS3gGw3H6sGtGnt6uq2vMQpinojMnIchP6W3b3M9HF+5zRgA7z59sOB3S+5lUo
fto7E4ohmkZ7fISzjXM+KoY6mIEZNYyVMA4jKsh3QmljmmKLiKkVV/21SEbANifOKr4BlGYiUh39
laHlcdJWNjLsjsxxVM+1ACRxRTicpCBFcY0tMdRwr/7WXRAAvmiRP0YPZjFdI14UXATOVNXnV9lC
nJ+OBXe6QcTx5+wcD5NaRScGeZPAjQciteQE5xRXSaJiubF+pZuSTKN3HRcgrb4foRoGYzlxXuOx
1ul9OfkV72yjB1kN/BjEX7rL7FuC55+SfarWMmBPxWViOKufes+VF2PRsSmrzwdUq1pGrcdHaOno
yxtlxvHcUFyfaX9gaxL/kULyHDPtOVG/KGFztjYdh9JAZNrVqb5x4ifszf0m9+rIxuzFahXjzR0H
a7qpJoTmBmJ1ym0XwLqIcjbhRAAVOd7sB2qZe/+7fPmSDwL1uta++rVY4WMkpZqpVZK3xeuR9PuN
fIs2YRJehYQLd/Kg9gYNAANONH2MGkMiI3An657AYPIpWbXgCVMBnW79KIgYtqDKe3MPPmUMAKDh
/WgdZ7ZL0RWuhA+tcid89YAbo7jfUs5grbyzGE8LqrnjLXjK7O+++cj30win1m75aYQvtsqCefOm
+ZNw1lW6004jRCQIgVft+/yVpGSTQBMLrr6p1ZjwaA2O75tjv4F4LArEJCw7vqOe/qfxB/Rp54UF
Mw4OA6quAbQKZf7uQZdUxyaDmqIXw0oW4/yXSI4lwJfnDoE2EmEaDkVrEsOcRz/5aTHZjuAxUgKe
pz5fm0cNqkdBBk4hscTpKFuYtbuH/3ByDQztipVFEDLHOH5LmbEE+zOWM0lJB9Z739Y4SdxkXCDH
eTXrRThVSw3TQbw4RSvy0jka6lTH5UoEQRQoSi7Q9bLNBImhmqY1h3CrFSEACG554w7ULPovfLBR
mdPCCM4RvpLox7yafY1u3cMBkiscNpGNtyr7qErLbMbpAReUgi5sjPqjl3uk7xLx9EVg5ARKH6TE
7NQJSw2MilwsFYKv8N1rlwZ29TlkvNACTmRQtznEDzYmhzWBMq4f4NXDrWwEdXFDg3qeMibw6Qhk
f+jbDZkkzW3H9n1r7IZA9sizTqc3SAhLkhD8vyHRimcvZ1NTPcPrzQ5ZPpvtDKUAK8af4/1xEDfw
tV+p4NrRYPsl9j2Vf4BDzTgVz5sCNvyjiqp6B/oAYUgyAQkhNxzYqEhIT9DEwRQyRq3Ascj5lBEe
xSaK+4V+0HLh68Piigbybji0UVZHscgW3ZAcZCgLCRUlhYG/1PlsCM+fdUPIkvuxoTifOBL4wWXf
zSWXc+UCKop8y1K5KEjJ3NTpGT+ouZDcZ3Y9dGPIOS1hjUHL3VkFV/JXgwFMFI8L+woNIsHFRmMI
fiHXYE1IHzoMviJYRO0qCNMyZAFcNZKHgzJANliPOoab3KO06lDLcrTIAA8U4t/Z+4avVsRjFQre
Af0xit+9aeIuyKtYBOgeeA6SyfFfT2ss8PKdopcOdZcVjYY6fgJBZ35v3w9ZPLzfh5uRX+hygFxB
3ePcbEKEYaGBcf5LSgD0mKBbv/HE4Ae312a5VfcpL3vCJm5VSmyylkrs4jyN6zDx3DK2bOtc5m6c
4F76L4G9n8nNlPbWo0CWN85Oe1pRUPTNCqWXkY5zzzUvOO3sbw2N+woO2t2onwhTDfUceIQUJYBG
ALHfDIgEhT69QNEOE7YTo5z/59w1ZhC117A4Y9YU2ZFLLZzcNL7ekAF/t0WoFB/ygS5tLnySunKS
xTSDO5XRLqwgXLjB8BuLX89UOzjdwXqFSNgr0u7gVpvD9+5F6c73YL1Cx6/+Ve8YCgyZs0x+xZWF
+ZbSfl8k0Uc7n269nrck//fdo6WuUfv5941YHjACRHryP/gf315dMr24q+MMEiVI6/JQVZ18qdwC
Cj9FTOF0ELAnxkYjs8lNAEe4Jz3nLXsDPbwJq4nVehJE3YjlVA0iLBinB+dcdKdvTPuGTgr27Zls
1Bdf4hHDyDTpb6nwZrys24OV9f+Hz+ueMOrkjpIpYZS/xQGYy4lfkJO4TwrnWY73XRwp00cVMf0W
1hDDZB3eLLibQmlI3z0gsjQ0RbLWcB5mHeanXQO2AG+NTYAQtgZ6/2WPTxW0u/eILodGYSxj/xy+
IvK7lbKSIcHh8zWadxjwzXQymhP2uNgPIc28lE17sW/pqWSMExEuoFy+fS4X6G5o7RKx6oTuJAqk
F8M305tBxDL3twZ6yrbaDVbk3uERnCA6wRiL7U2wWA93hwVWZ6WAI5tcFYa+ubL63Tx+it2CUSnb
10Taeietcs7NGsWFbEzKbplC0o+IIMvmh3MiTA2HLn7spYJlEKcMftri6eE9wcCYz3f2LxqxtFy6
nh1IZnFIjFYU0lz8bfQIrBnh3eDY0gH9jXJ3zqkJkdVAAE0aQfI5ZF3VRc0QR8IhJ24MvpH+DqAI
Bs/Mht7hUAMMC9ablGR2SD8nOisAIEaeL2FAVsJ8+DzWMuo6GAGO+iXeBeJRSAvjVOqaHqCJFU5y
9CB+jVDxPEiXc8dschUoiPnb+jqSxuDk++qRWFhK92ztwUwMcUrnyKmtPYjj/YFSe8B/opJ9NS7H
JL+6Ml60SJeVnIiEzXFecFOHOQ5Sb8Lfggicgby5U9Be8njfKv7tDdqv8SXQZv2pETczQ51kXi7y
C702utQNR0J1CxnLJWACSVouNEZ9PjgHFlpordc04q1UFX03K3jZJb9j9jPW3YuHqx4D10MT2lV7
r31C/jSf/KZUdao6jSsa/thQLP2tM70yykQZAz+A85fcNZBl3sD6EwMdFelvqK5V+TKLQ4l3Cg5/
PEHB1BSuW9skrFKjD65DsDMYlUebM90Ld4F1dXGI5o91W+HIrNMfrPlz0pZ3MXEfl/c4abl/s5lU
NSxMZ2ewrLdF9UVLzVREWmHCeG9gvALJQnxicYQTOm9i+28Yt/yJlHE5dmjScrCuqCkw/gwS+hla
hryKQfYv8Wxm0Qmoc+9Garz54mv1YKt/j8GFuUi4ZPIjqNm1Z2/027FARzj6DRBXDeCLDhZGcAom
JtjmA6h0YuspkUB6LoBiecFc5kzKTehKF2UnsLlpWD/RfP1b6o7hqGcC3usbvyE4Day8TGxXsAST
Cumdcf2zrtJTW809spzN2O6IeitPqzjOYzaTZ6+Sc7gT05wQ6UFROOUCkTvmDosN65XMBiw2oK+Q
iddNjf6E+Qydo0Ze7fk8jygsKVm4JunI78yebOQrkjr2kVZ/CsLM8ARCIeUOLJlWi80OX3ZNwYfJ
Xlehocn+gx0bmKHC+3EFzXnxk/1At7cE9fbiuknWZj1chntDv+YZDB/BGJyd47yYnMdXpXBo2s3l
KwoQy2spKu1YLECuxdTW34AuwbW3b1OHAMYX3kWZ1SuCutRMtv72FkGcVm+BXmWbJ3P7Z6YfMMfE
xWyfnyLMbS3YySJGVVK5t+6xQzkZJbnXwrgBzHf9ZjShhSu7HkZvZisXr7YgNBiPBcRP361l8tBC
Q0b08HES0f52Ns+JOKNdqxWPIP0uTmwwYKFIfgziX4NtXHumjGqQong83v4t11KFHryqOzXwFgxq
cUDF1HtBT+Gvd/ltBVYBaotQXocK7mNpT1Yyu4dwPMOgHaRNRSP/+kB7H4iE0RVvGcgd+QxGQPns
VwDlwQAETLYuBEuQQxQbBOikAPQ5ak8riMii19VY/1sg2Ny6FnfKenPMhsJlI3/TuSZPyD2noJZe
YAnOwIKjMTLeRjt5ayyqr9/GZIwZpsNTqWbdDSH6POrePc++Tyh7dI4ba2YGUUxfDC+UjHmE34oR
T5mIgW0llpj4Qz1/SJVFUbU/pdGrs8T4EyMg1yEHzg9i85RYbniy99VC70ynL14EwGlm1LISEDXs
N6y93EBmwXBD3UfQIyQwBYa5QsAMb/p+Tx1RK9mUGpGh1V1N8tg8miRaYH/LMb+FLd7Wx1lgI+xd
Wps4FKBXs9Vr67urlAd96mM8YJvdrcwezVWZegMPhrZX3E1s4UOMhrmdzReLA1Eidf5Qxr79EKtF
2h7lW5CRnt5KGEr/u3MXKmyMliXgHdLpD2OpccdKWASxRXhmrTfJcWgkO5m9zgbwkk+eGP//0YE4
HsuX3vLeSxUp52VvmiYVXSdgsjNR1o8OQkUZ1x3Lcil6svJzh9AtBNNMTsgeoR84QBLCpp5dPD3Y
p3jlb+db+kn3rEuV8Gml0Nls8eLjTlrT7QwynsnNNhK2B3kL6P6AsGeyvOXPzah7xX/VsLWLmKro
2ujkMkSPrrS6S04e45x2iVWDz5z9YixSd1RJhBY//0PQzx5H3iKIPZPbsZ1quAgVQOHxfteYOtvA
h2Ao3J8FjJa7b5J8DGIQXLvQ+Je0hhlraLXkVpoRMlTZZj8P/vFCLykogROMdqwuPqhBDGr79IF8
BISBj4NKiEfDLItTwSwE8we+H+ELDu45gSwaqf39FL6ktZPlDW3hOYloB8H+gc4M8FUmoTGl8sZx
g5KGJrEd7j0+ceLMKFj7xEd/CMJY0hWWD2J7WEcJ7Ay+dlQTMfOn73M10AvYvDEtEKxX2+NE46/S
yAathDjKlpybxJNtXZDl173ePy21ektV4C4RmVTrHw1KQJA61nVTY35a+hkd5DmO7A/RS2SRaBNd
fU84QWnmxEupjhq7o0onhkHOmddJlpsSv2BloymSIK4WdQ036U73YB/kB/yGagPIrIGxrjdhZ3Dj
JEnIfCLv/xPd2teisGuHeVK+g+LB5fXe5bUETSdVZpUL6ARuni79kW6TWQ7BdYQEw1iA6q28cZzY
gT8n5xhjLkgHXXxMq9GUKD1ukzz3bMoOQBq5o8BybnjGOTNDGesbqd1AMaj2X19KG3BuXIpLqspe
pR3nV1l0DXwvi2DFUo7D5WwXlhVqbrKT0vsJA8qbv9ceKF+8xXDLNtpt9YHbKPehr3O6Fd1G+LSl
rXpj3fDdlFe9omV6U+7AcYptiXoGEGmsjdM1RlS7JgsQdF2AQRMFHrRsm9LdEJ8Uq5uj7CSwuUOx
m/SA7p2ZCNM1wAk5TaCZGqsC4X6ZLJTSFl+V1hRdq7gJIQQZLwrbgA3n0SPwtb8ZS/YIwA3BhXft
Z91AYWYV84Ua/RnS+wA/kv7/njPJcMpWPhxxYVI0bJkrtbamxx+UOr3cDUEULqHofYcC/t7do6MQ
wdtbQ98FH2yZbCWzDYBL+Ie0rfrW/S2iHxsyi/FqWwiGEo5q1GopSJ8TnhD0MHOw81kyOis3b7Ac
Ck/VsEzSPAaL5C38bNAMXsoRVO0HQG0XO0GYGuC6Hax7/P4kunueehG4JBnYUBlQGxRukvu37Ngx
OqhcoaknUPvz+ZQOmuJij6HbdahNfkKgCZ7mgxB9GajF1IbWdWuaIeUIPot8hSrlA1iEeTx+MlcN
XRYCs7pWg9FXCGjf0pz5Zjq0XCEOCBRWwsLUZVEJY0bEYE8vziR0TVa+jXCBFukSQcwaBOB5K6FL
LAgfOtz16xQqE229QGaH0Fvys7T+VIb0yxMnu7gLYXxE86fs+y3TqEg7H8yEb3U0xHIJ4bA9hbWi
KzMH0E1DuTwQMxkNFmKfEVifYLz43/Fl2jVKqfx/Nhmd25oX9MOZ4xgt1ziGuHqZVmvnmMAA3+wi
lAwG2Ps2k3a+ooD/rZmQr0MZzmAsoC7Y4WKHn6xK8joT/e+B22BjpxV+qFWxcyedF4c1PVIm/UYo
fwQcQUWrO4PC2adyyv0tRyr1Yzmr9qjHspSKgKXmBbh5bSoRYNTe3fdR1oJ7Q7M/pEw4er1eEH40
abqA1NtLsqRviKGQnNPbz/OTiFroRtuIUA6AVTIl4lg8ipVjwaj0CHokp5AnSNni6FHsrAl59S52
pg6l5Xwq0Nmcr6xKXl3BXcFhtDeZCA/twClYVhOIQIRQJ33LzDoPpqCyUVV6ESx0SaE2heA+CV4Q
0JukfkV7VCCNTcLCCnO0LpexzK8C2Y+obGZYp0vGRlLCC6Vatq0A0w9akMvMaELWxKFZK58RdFXf
YlES1RdNP04IQ/Yh1Ftm7pvpgKQmofLPn8sWLO78qNhQvALO2nMKngo2NuR42KfHhE6TI2uNhJAC
dwLudfng/8FG6PXSS+scnXxDEJZpVJum1ifpLnrT2Qn0eaXK0VYz7yjMn2edkFSTUdkbGBlDtUY2
U/8aoQXTtsLkHyY12IXCROYH8QSzoCk6fuoT80lE799QoxwC84QqBu7u44FuIseeYcD6Lry2a2IS
HlpPKXwcnuEWLOMFZ5UCJrZrFwYiY8H5Yz+pRZS1rlcfIKI+Np/sQ2hbJkv+/s0QHPEcsCL3ocNd
LaqfwZlyD8Pqh8ZIBzSEaRMkD6T8jZZuqjYzC7JLEB4vthJv3lOUVLyBuoZx7a0bhbZjyFTQkDoo
JeaapR0RRoVT7HDAjbtoDuPmHOOdCsqDpirZ8uQ9p8Nk+sTwzp6W1JXiiQ99EXd1cfiDPs851zcT
P7sePHcOZF25SRHyLZH31l1iC16qmG0qC/BGqL1NVuhxmOWmxbhogxq05axAN5xfQy10lgtSTfhm
1PlpkEP5MKo4ibVFY1TFxJR5tkCfywiUSbu/inL4O5aUiVBBuVKBGGyt8YFeFESfP/QaFdYbuttY
f6E8FyL5HsmBhHI2/Kn81LQuxId0rv+gcxW+cdEAWCO6CQgHbtJ/zHQ4liDiQNwL4M6aS0bWKGn4
9HsOWP9hK6UR6g9xr6bNQlDrblxi9JqYbo1qrY00IQvu4c9drlDkFkbQX2KcsJRN3Y1JoA+3n4CM
EI8ld6N4blULQCFTD8pkS7c9SAwt88R4ORizCK0epkknUtTnccy0n7FjQGIlVcZHdiY32YXJX/c7
MPb1pJ+D8vFBg2pwAurz+3SL6FyPGzqpDx5R3qbU+H2P2O3g8lI9GSmVBDEMbZFUGUQAFxUdizcX
ls4TBv7Fuq2Ws5N+dT67YUBhjxgIcKpZgabkYOyBr5kHZQeQVnRUXueMXqbUFK5viUr4o7pUWBlh
NIwVG3CCNwg0hUKA7OOXA//QLIIrSeBzy7nkLNXM+D82YC3oYi5prWZq2ljmjxWNGHKST0dFMy/0
kcJSjXsbInzE3+n0lzE+32jwTDtt8wkX7AFL4OpzzfVyI6xMVh9s6O2pLfTVogH08rVhGVkKfK3L
TzoARRwJmc+Yt62uIrCX5Ec5gbkJCTeCidmAavoZ9DT4+dF2tnXp8V76yMtV6NfsKkun+N1biECY
XWkOPk+M1PvDJ7wYFuttfYYk5NP0YsiaeJEvL/ceoToHjYu29iQd3CSrVXFCcamqqQ0eut8COqAU
4pIVOI5BwAnx1mE23GQAnV+3kqf+QHUS2ftwCjm4yyfWKqPCvNDU5gFfMLv7lWNuXdMh9zsppv8q
ghfurkd5WWxarECWr4uXxSyv9s0MEbHbAkkulK5vxeFRM2Fgbwly8kSZAydSh/yugmIoJ5zCNu/X
SRzoeDWPuC+kZP4pgXfP0KoGoQV+rw4ZR6pJsCv0TIfBCSxRPoD8Gzh03FZANDsIX4bNVRDODRJN
SGMuh1U6Re2a5e63EGCLD8OixzihO/sSb610RRRY9nxD6hISdReMKWadslVRYeyyWIPopnNAvgeL
G8UKQtcouDOSaChdSZKhJq3ryxSiwbPVh8d6hf66MUu42VK57ztuDB+EGDVMYt6wJEyUXJ0vajdv
PoUMNxYafwv0iyWNPRJYFRZ1RCPSaKLXhTdiW6UG+JK2jLKNmsOKLUDZcD7PWvPZkpSgriuBoCfr
SA3CxaEiiewpaqknqlyW4UdlKWO7A0pou7+z+gjMN4NYiv9dDneV9Lq6zTkKolDRbsl6nIQ2cYhI
Z574nRwYbrBlqoZgV1mDlp5snTZ2h3X8vVzx3UQvCC37KpMDFpf7xem/5bx73oQDwkuSR8He1feG
+gWPo7vUtagENeRldwrpjg3YQnwhr/z1A89Z3m3VYMektBRCao0GrtRRAPOYEMAhpMNBFIVe/xDH
KFsCK/PA8wilPeKJg+ElT1ZSy4r9Dj0LhB/MhN5/b7kuh5BXd218l9vxwYFCGcDDB+xsQK/1UK62
eQtwVnp4Mzw1oL24ojLTxlAE4FcThN6VYV+tAeMRPMPPGukFt6BZBtoMNj/w9qNw4BsheaXW/Vbn
ay6sipCRJwAcOshtEsARAlNpyqQLUmTxBXo0DMDbCN/n3EfwU4Kobh7nEXmvhRw5N1oYfcMzVIWp
XwT7X4TAUAEl5UiLkqFX7LQ/JHEpLl+OJToeRW4EvdRtoogaSUPPB8o6RFHWByFO/H8jC6/2SJlI
hzfb9M084+B7JN1SbGVNFm5hc3meD105AZzBmBCKtxhcDH14A5plXZGGoWXwMeuo8dsdDBEIFZnQ
7MNt+clk07YfVgT4FYZFuau+awY1AbqIejHAHJyu3wuPGrm0QNYVuz1/9rklcMvZBc/atrsLzpPo
sO2BpXNehQkkToBg4fC8L4aSy0wyoYyFkz3CuVRqPNcve70LiKx16Z9eF8vPenOkHqza9GeBvO4Y
M5iGUUaN/IbqWGuQ10AaXvJRqpyqegtfJ1YR/HiI7Xd2AJDpj1p/byr3TjMCWfxPnqe6o3Qg/MEK
Gns1qHfppZAcp2O2m8FyvLvXd/hzTFtg3RysjY0XJf8adFYCT57D9wIdat2vltwtOnBD4ImdhLuF
cEeRvtamaLaSL8WyuFLdm54xrsn/kAEHboSUCijbsfF2c/ZpQwhfwBixqLHSQNsSbMuAenr2DAc4
Kn0gQQO0M/8AXUrC05dAw6n8bd9wGjaZVmfiW0DPSQOxton/Cbj4HCx/QcJb/uekwIJhYEteKFND
7RjRUJZkbclAKipqrvuj2op0K6U6vViQQhAckwWxASk43cdlTX3LJ4uVxDZYb6PQasuvN7vJ9Coo
K2U7ZpGfZWMJTvWvHDDoh3B618VNjDdMTXaBBg+gxjUGC1qJolzievTGD9lvL7Jx9HaEEFBui3x+
dochgw4z5ujcT9fe7NxpI1k3H5c8xkMSPYEt5l2wu8XilNq0mPjzqj2ERBZq1mdIhncbyW84fiKV
Kpar44UEJRClfpp4+SbQ18HGgYyqGvpJw6G9vOTTqu5oy4wbvgtifNaZnWG7I/jRLoEM2/GcxIwe
k2JyFK2MuSpMwupdaYiyMh7+hp7u3UGlHMWNxWXLhYlx3KTGO0IiXSDz+TngKggj/HBQdP7DUYkM
Z+VaW2bL6vYgmkVsAdRujxPdgZO2NJ8bjrdna6SL2WGrs9tA9DhEsIObK7i2iQDSMnafkg+iJzB7
HD+efPRL8Gb9/OH8kPSnKEUf7XDkolKHXW9olO3ZWMOiD287ZtA7ic6zvhBhA64616TxCi7FmSbH
UFDfsHNirQFCo3uVnSWqsfyPe+43CoGvgGpEgCdcgVSOptYNtPkBOLMz4NPH97wUiIq0nJktoWwL
Q5mGKMqG+6FyF6/WyyqgxGvBT36MMSj9vIVaxtC+jDcC5a4NqGDOAVAdZVhhzYI76aYjbztXANlQ
ZZZh36GaIwWRfWshI4IfZWaYWM+ysjE0gC9EZQUPxgKKxYa7SbY8byvA9NioYn20P/1VlJCT+pT5
CPdAxoGgzLl/+G+wF9GmJ/xJEAISseKtD/9oyAbfE9hJG90z0OBhTQwB18NJ/ffyRQRuMEmhyLe4
O2mX9OMSo5x0vMx9B4ye3jsFiyJuIH8I02yOROqO6U4/r5A/AmLem7SbE9xSI2VaLk4NBFosM6Lv
mMXGSVnBR0EkwZtUtIL5QxKM1W5yduCD4sitvPNj2TXfr4iCaoSEzLFWeKpFpppIbvFuqtfwPHIa
S6i6YJ1Wk6W9CDUczh30p+JmW3qIpI/jV/woltr0SAl3WhQ4oRJ9NdecGAlaI3E77h+b4p5DdpK3
WRPfjOp8bDue9dzw6KCP3gYBCyns3QxjYHuuuSLjV+XonobON/T1ESd/IjGPlC9i9FqiuoSrECWX
9KZ7gtoO8yAV+I0QfQk8cdHCJ1OIjB/UIjT5pF6DXBpHLWOuL7T8fv6gC7sd6l0CxYUXHk7OHEV+
1mERShrKywC5QL5gGc0t8m5EDTpkYGKPhNwGskqla8THoHRUxeDli67rVtxgTKw/0H+Qn4HpMtDg
k/4P/TH7zQ0Qlybuf5NvgjUuNdFbsYa/S1epfYvlGzQezL8VhJf2THRpM1ugxiPkNWWu/P01/KKe
w5AHlABsOSFXGJaIEXwSJZ5mxWtzLWRBfU3xmCHTw9fg+K9FP4AxOtc/TCHDM30LGwkaUKLwgrDQ
otgkJmIgcFOyhZWCJynWFZl3BowjRAIkyNDZwe9rUpDcFSL2HMNhjvzTVYfcV87chhgOnypgqEIi
QJf6TtFNiN1JESV28ix/UJL7XBsH64F9JlUhaGkS9VuoBUi+gPQihQL1HkhZF2S+4Jtb+giGqPDF
8ESrHaiVEyUgNAH2iyi3TF6Gi7ozJvwlY9HPwSPM2uwDwl1ZTy82E+k6xrRH6vYhbQk+mNxMru8K
Q/UADvZgWvbqwkXjo/E3edtX3CgqSWeimuvQeUzsfSnRsCLATgJKwoAZbBz8sFjLajGNosR8uBAv
hOO1Mree9lVfLZNYvmtzorkPZocc45PWQ295o+3aCXIZjUV/q2K9mxC8C4CXxP7Q1jNjteRg8XSw
ROQVZDJfmMbhjWm6KqKJImj6iU2pa4sa3ssp+F1OovWF1vmPMkeTeIwCnML+jBDB4mQY/niHlVfA
Ov8v5DPKKVXbmZTVC6tZszLuxH46X2rnVRDvixlxGBDLIr0MvB8jznIMqupC7ku/RMufAJCv7Pq9
JXcS+hqGIb+L//cQ1EpgSUTT1Rgp+vinA1EFLfDgqyj8
`protect end_protected
