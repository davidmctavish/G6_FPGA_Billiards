`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ezlmHfThO2Un8MjJdXv4rT7MuQQcRdPWXb4trZUl5JO8dcJwSW55Zd7q8zUGGxsmm5KKn1EYwB1G
UrGONGvBKw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A1B+SR+o6IaBGUrz9igY9CNB0bWJFyCns/53ctROhMnOLoBxAM6Jfprm6SmK8OobXfVqp/RHQ7Ox
q6BRZ1iF6/yDLUWGK3odtfWFIpdEvccUOO3pJTN4+zz3MI3eFuIL/gPIpMDiGoYLiEjArg9ldgj1
eT8eK2aJ3isZTcbQkSU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
paSE/LL9LVyhT8P6gPCPVngrSZgpqLCD6j7n9uMAlaphzmiFQsqhvewMk6eTDeMbA6mFWWk1buoK
2Ow5CCszLZb2h3bnU+O1e76p0BmrDFzGt4FtS3blA2dcpT1MjEW2qMQv54d6JwHOOkKXMPcMxxty
WUQ8sHPqaTodiTGvxSrTbYOwZ/WjeGXYsYXm5S7FKYrMqsXthAoT4ZhEIbgsBfGmyhNq9tZa1DZI
TUQjxrjpsrc810gYJL9h9YAWx8dzrF6lTSKZEbhYuv7HOy4qtu0vgtKG9QFDhG+GHBSnHxm4d/QO
PLwTs9yjQNvfsvZ9V/yibeVJcm5amYk1vr9Ehg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y3mnedL1R+8DFRPX65B2EkmGLolKDP5A6/vOdR2weHwn3zktFHF9ghcwQEeXczb8URNzZrAEuv4N
d26o3znf2CQ11s4hi6TDbe/yLHHWah1tuVpDwlLXfzZXN0pqO78mxbmZtSnE21hX+NqUNnlVXiy+
rL8HASsZ875Z2w5FlFM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XbSu6jzyJWr0HQHPrzjx/CKtqiLkA4E5f3RkoiMATCyDadQRsdO6pYt8p/xMwcHP5FsRtLEY8VdI
LYsMDp3+8mlrsdKxKzFFiNB350NGihVuYYbFz+FYkhjB9Itil66du4H1PUFECaZ5tipGuOrR2wAn
cyR89cs7uv8FU7Xb8mWvXJA4XxvHID1TTd6qtz7xXY2Qj0CGnV6w/qrnhonTcr6GQawctOZzSq/G
nLbwZRh/oSnxOtqd5NzGtcAygiABKGmXhXfxfTqlXzuW4fMhm/hd7Ddgc2kRIQB9b+6d5o5lU6WJ
fhYimNtbhVHf+qLseh47PCrDdPxdB90yMWKE8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8656)
`protect data_block
HrWCnN/ttl44DJHrHMFqrAC1en/UB+J/ELgxCwDzsSsCDt6aKKzOgOU0t5V5ejxlUb5f0/jXHryp
Ld0HLlBNoWHBhruMP5aijL4tvhusRtORXZBA4NZ698OvuiOfRm/cyz5b72923mGxPJj5qc6tZ61l
BF+M3uc0Rkj6bbmOXRcZgTLl7Ppt54YHOzxJ19x5/Fty54JA1JLSM+4RqOxoG/3PAoFTYWS53eJq
ULXd2boAT/JL0iMUB1UAmRbbyu/ShY43ialoZzVzzCYCLrogDwhyubSNNil36LaJdq/MILDbdHiP
9BRfyWwxZn8blpzd5Rd5AcXRazYpI2z3Pq1ywRE5ss27wP0sstdQpICDGindE1aCqrt/BjyDlY9a
0iiP3BimI4ziECbqVWwUCmA3ARZ7yoGhMcwtdfjRNhMhLDl5WNjfamvpspvdxEWMNyzXj6AxshfN
eU8J2bRLcEFPPZyszTwpi5iZZofKaehOwMEQEJwgTuUgTA0Fh+fZ9BCbg87+78XpOIxRRXDX1PPG
clsLDCPu0x8WEIGtvWSS1OceN2qgM2Bbb5eLG3oh+I5vcjUrc34ZDlVIKGiSFxj9oBoXSWLuZ63c
Z23gnWaahfZM+UhRzxCI8FXkGmFLrnUB+W6Ysu0SSslWLGU8HrywnueshqB/rBlDLiEwSrtl2kMO
4Zvuu5AefIZKRbq0cWPbLTSMoh8EeMDXRF0jg8kPj6x294yTijvWVcqkC0xEs2C6j7X48JfLpeIm
LDnOJzygl8LxpZjNzrOcBvEaEaaHT8P/WD7ZbpKg9ht5ccc+tm7VaaCWL1QysMvB8lfjYx03AwdW
+ai+u239t1BNMAQbQoIDjuffko/2ivTS1XVZo4uVjHHmowPLimgDBvG56NCkoInkewqY6NpF2tGf
xDeekBX4nnRtBNvqkun9CpiidCzY1Ipny3jfMcNc5pETuJKwq2pnaEN6JIYQoQIrUXGbxyj8av1B
pmhKxBwS4/GID58YywfQv7ndEnud910EgCGwd3+qzB0TacVDAMDCVrkkb2r8Zi2wei/rOtklfzap
u05Eb17EqTofxmvvi+iO8uFCFaq2Jjbqin8S1AN9CchrakIHMbxxi6NS+/jbEQ/S2COV6lwiqQaB
0504mGMAVGhyYAsvPWnbD92Sz6M56y6OcsRZOLuFtepFMWOZqp0kx1LpBqjGUMNLkNxDtYat+vjZ
osJ+XFI+LWPBPOIDbmXAxDsHH1amBtW4G5GVh7p0M80Hkct5PSbggs2EopR8gtilt6b3CSEEaz4W
EcGPloVi3wcnBW/2ZOk42Lp34fUOXe+55H1inGqQP0J7otmLA8BCpsYm8eLoG7BwoMqpf7WhMvSe
jHaNi9PTuyqidlJl/JYFbmDXP8nbhNkqnFB9KjF88/ik/jTOm5kzz0gguDtg5cYVNludxWY0JUa7
cOyPW2O+Y0fFToyYOftn/SIPr0wyrSrQZuijIiSG7ssUtiNeZwdPffYb2b5jfH1vYkNkrl84xxdD
GTOPCsyZmFoJ8I8mL+rpyfV1N/zrZfDpu0QoPPsKuVEYXJHQov2EcKvyiItm7OBUw154PdX86uRc
oamfvKEdTqC6zvTmbPf3YKQQwswNSOqcLkimcF7/bYrr6d1KoVYLIecYukkplMIw9vLPtN5MKiRk
ulEs8SDEo2Iv0qoQX2sU1oYOOzv1XTFTsrHD+rMxdOZraQlSUtQ71IRQewAsQK/U73Bc7OEVaQwf
uzGpNwhY6Byjf+FSZgFGkhWjjie1VYDYvm5RQm+/BVs28ecK/fKJb6YPDlmpL3r6mqLbry8xJkgL
AjMu66wyaeByaveq9H3EqfcT63f8rnFB35CJVFnZVtrdofQoyYO/OFVbIeMBwOlprk5RvFGr5TUI
gufpzXPmjmUZJVBLAMEBDKqvbfKKukhbzh/35NSppl/6Y2PM3z3runDFLWMMA5s/gV9nKJJbAEPy
ucaPAlJhCRifl9GyBebYvpWi+M/chOJKw2NgVnLG0jfG8g6tW4Sngw7XM6n6UUGzKqj0aVeTMuZ0
cZV9sFJTXW6eLQ5Tn6vUyBMYCMoo2tdfuZj8QI3p0GEDH8dnAmWmScvC/+WgSm98/a2UMLfYKZSJ
PrEbPIV1wR73Jq+eqUAfaElxKqA1hZD80m0KPClFnYRbISrZEYnkfFsi0Rbporl+Zbm/YYSYSlpQ
rPuek/TCg5SwdftC1WNs8aZBWl7H280+h/yyboPk5BlMmWdnQ+ZwHQiSTm+hspnTw4iNHezCn3f6
IZSAboQ+wst+ojzxrG9MRebpx8kzPiapb6L+mciw79fnGjLXQAPtMkDFLWqMXbzNxD02Kg3iKc8+
X15xyhteMK4du0IVUKr5j3yyM8S5C/DKYanh3ntpvipSCHQ8/CZCvd3tXKP0+6WqsLTPeefF1wsY
0AaHcc6tDYaiWRQD6pJeqhEiLYT60jVbVFTbgadsFM7Ce8cNitQgfHaMZSBZDvudn9pSoqlChL2d
0xtoKgJJT9XeXAvpMNziwDKUZ2JGpeLhPCwwLO2bMNxNwNn/ZCh+2sBCOTmzqByGDNZpbHQKkJlH
FvHxMJ5K9Nfrbb21elrFP8dxn/cLh8pJCucnQCiC3btbi/WCCelRYYu6/8drvS0OHA6VvYARdSbf
LUhpxcwyjK84l7nSEri/0sD12rd/exBhTUMyvy5UqFCfCWEHQWwukYi0h5VGMFhw4Gz+WE3glLf9
wIzT11taDHDIe+roGQNsCohmzF+YdFOfif8nV6j2i19entD549iCRYLn4M8aQom5ryKh00qNGBG0
QHB+f+egn7TTFyEIZICnOpOz9Que+wPZ9Hzgq+Xo7AtfTRd6M/2RXOmmsQIhzQ90LPNVXD52d0Um
KQjWgZb6S22GkJBM9M7sRuRqHkSFtAoa1NBdWH0u/ptSrQOoOhXOUuVx0kKg9SPX3Q4/BLCEAgED
9Q0hLpBO8Xy4008COljwSdMXmj51kJCNvt3Ldo1wTC5uv46A/9raEZWNi8IxLWe9e1aqZNUtGQDU
QBbFdcz0zstlhOtlD6NPP/HJ1XHLddXoixYhCufpZ+AOSc69ldXwNKq5xUj2Qs1HQ3VLJ/4uFlh8
ijhS3yvC7ytgUDYZDfs7Kn2T3Y2i7kA74fsXlUptcDM4jMQKIPMR25Xy92ZUum/cgfsZgiLlKB6h
se8UoydcQ2DWOFoo56DQdidb0rap66zwNOlVTqlDAI5xEB4sfgCYnLu6eh+7FX9+Qji6H8emdait
mFlBFjDQfK2a+nGsJS4PfOBrydIvXqI5zi46dicRWwiI/FMZZ85F5i0X8eVQIjeZszn+C0Uwl+of
s1EIdU4j+8R6pfffH2UW97L+Azpl+fNlHLXPn8+Cn8xG4qat7zkHfL8GnSBt/AW4qi1yHJ2qc2BF
h5pEUCUmOXKBXxcSIM0/WSxFYpUi321c7P62otZGIR2cm1m+iNKEUEDm1NLFnhGxAaiR/g2+wzXo
+wMzRuGOCuDF9UEmrhfY7FCQKsYcf0kVrYENQKULlb1jLvR0HkgA/s+uFaseXZSi/tKjOOdnHnAZ
1vnG50jEqI8nITWQjL2dY4VTgMge9ge/M/3mK0qVu6cG3HLOntYIBf7COoVstP60DUfjI+gkCNf7
iLJ6MqLTOEKn2LAf//3K8gtGSxcEhsUvspwfU6q1mTCoHp6wGnRjZSgJOEx82Gbqm/5jogZy2Bct
+JjVQXVIGHu9YyR2VhClP3is5sTzd/Cow/uHNCk0s1OXiTwY+BazAvRoXBZDOBwOD5cn64OOjqkE
Jh4x26olFmWqVjY5odAR942pZqMyaVYTbIydzLnBLC+cnr/Pm+wdG3D+Rba2a4DzSIDIUCe/n+HS
R/WkAKvMVPRyi0eVZYlSR0XVJ87viprMiY1zU4EzSsa4BGoYEtkERpVHo6AOpJRciodrjPgEGaD5
iqNlUCUR34wKRbae7TljuJT+1uFye4VMFfhn0RyUEjlUfs9b6Vz0zQz1hY9vHHFF/PBDORd2uWbk
zn9gyc78s77mF8jgfxYI3SHDQWn8dmG9JyN7ch+hkBNK4oHrtWlK8CteM/qjNiff3J4/vZ34A1qk
T8K/ib/hLdfwYY4CTP7tuFwaZZS8ZNJw0Ak4wEFlJOiFgzuN9qJy8sC3a47RB81mdYE5bWUe2tnj
Fmq96KZymUHWWNYlMNP13bD5ztnAkYZ6cKdhWJR3vuVNM3sfq6ZfTHjcuetkJ+JH7nPthDQjFn79
0tNoA3R6pwy8QE4n33AxzgGGRQWLt/F3gmHCuqL5z07O7O9iVkfGgAs7D1b/ZuvchuPitUCh/Dgf
CPb3vciDp3SnawWnb/iR1HOKb1GtH7jEBfb25ibb4cyIJBY/siPwed7E22ojHNLuta/qdn7Sa0gG
XD8/8zJEOOvprkVTJtlXp7eq3RU54cw1UyTD+5YWaTqfDcRvbbNf5KsxxBqjiercaLaj3mZCsGh1
pF3OrAw9POHbr+z2xKGSC7ZHyJ4b3IWwb+ek/ddBZQ74BFl5WK0obt2udRLHlI76zCaFQCSqZ7vq
hCX5dfFIe1Obp3M7i7W3K6KYY0pP/SFA1JzbuT8n8gjpzk4ra7qp7yBHLDymftYUck9GDHvuI2nl
K8IamZ7Nn+Pp7Ra509OotaaritYT+NBESqRFUaDtw3O71qiYopbuZElX3RbTqOrWeOr7va3Er3Cn
ASOBUeG1FO8/HvxYfWECByv+i44+fSgwkXM6B6kUoDGjAsRB1cv4RXQylYlTq8vc4+S6XpvZVHpD
RKDJUUwhHQlaMzx1CUpYK37JCHFePdOHZwxc5aHhH05pbnfLOkMtJKVl6UN4ZH+jFxdvl7dWaBZ/
qxqxcOQkzMUiaywJmZlAwNJXOcYCFnM0SrhWwWPbiKgBkXBPNHJ0E5wR/ihMO1/gDXxuAHuHDvsC
y/A02CmnHdzvTgtzy/Mkm+E6rR8gH4GIdr/Z0rVvy3ooTcStugrdQkGOYFMOBVdyEa4QoU8prsdD
U2EBcZSB1Q9kVml1ohOzu1TIG7BcNb8kpsDESvZevuAjBBBKSlF7oUlggMOQw1Bx9Jgfi3/7gtAh
giVmJKnlrn4W02ftKw+hiEn7RDSg1lQ9EodECXeHfL0QaC2yrVpmYOk5hM0VmPa3RvXNkROOIPpW
2kXHnGyPmJmUBKRvcANzaCzVDUlmtBhrhBnRi363o+hA9JuelcI50NVsQofdd0k8COgC+bMohUF6
cowmfdpBNL93+/nt+s67mh6sxHjcCJazvUc+svJZdNKRdxQJUp3iw7YyDEIrrI/eIet1k1GkPpwY
A2/+MWqK1mDiXibTw/cyZoAr2x37OxFKrSzt3klKzKRnVsUrb7I4jSpKMivGzovhAzSGw/9s/ulq
PdfZ+qCy2ClhG0rm6SM6HEywZd4/XMriO/nIqX2AIOXToZXizTE4aaOXad5iJOHAfSCkM+cKBcQH
IiZDTRI/ccnoiD2eFm7e+KLBNk3scXL9eF2toApTqhXvMIUERt1zDwpmd5yTSLYXiqa5mg9VsQfQ
c6292v3ssK0Nbt0SdxIPIfVpPAhbKZmwSZhKsVpY6ukzJJ9ULNRDwv828gV502Fy/kWAJFbiToLa
w+oIIjMPlJtijus0DnWSrgjJzEELehiEei65+jYjc20HVTss+Ge+a0MYkSwrFVobm+HxvsrqM/rN
Lo96QLOwkN7pekXs3goMXSDOlmCqTJRwNQfuRDkc4S4gPcPKdTfPpjNeOy/6FI5Rd+sURzIh3Cxq
qcgS7p0XB63jyZfT2zArIC870YEvQUzxclR46hBH0UsbRvlDD6bsUv8lqS0iVZfD9qinK8DuP8b8
LnrI7o4RTg6nc4mk6TLEPUBT1oCk1mPA+sGd4cPKOiDRz1fPiuSM2qe/ZNR3xBBdQ9UVzI5R0GlZ
1qBRkfuinYNEGCF1ObsmwQEbUwQs0OwI6hc+HX2/fVfpEpJmG8W24c7fb8XXe0fWM4HaOkPRxZZ2
GhLZsbaCR5YOBSwQuAWSmrwlExplarJLGxQwtma3ZW7dYk8xOFACNSWQyuYkELqhp3ph58qcbMW4
bwypbhwkzisqPdwLqnNHQPa1EuQq98e71Cq7Wv0KTEzbC26/I1Vo4mR9wBWmcIm07pWeYswn+zUR
zF9eD5csIsLB+cRoetYemoX4N20bMWNdUV/vGsbiZn4KOWVWfytnhG1Z85pYbKvDut8O34Tbzc2L
L2AwGY40BAY+xa+Vv1d4gF81jmaGBtIrxPy/o3cWK5IWV5A3Qi0n87zKuSgbHO1b03rxnmkJQw9l
Ys8WyEBSu3s7SZGQqw2FdR4gK2yb+mavgUsaBuHxSZdMi9Xg98zxpYEmeBvLfUwYkT4YRG9ONYTt
qQ5LgtVU0Dpoi6QqXzBsyKSrD9A43FKtw36pBenntjdSiInSlU57B7+kKgxIQjalLX6F/zXRSsKz
HKb+crycIVtBt62vbF+i4rQ7DpOanx7YvpVlqp60ozSTlAgg5zXzF/OIdKut80oYB8ZHMHwC1aD0
P3From6w7RmhBArKrwMHu+YKBezNFI5U8s5OFsu2o5TyJowbFRCgko5F7mpd0iIyKdGWCc0E/Nlb
dt4AglroR076xZ3kN1uvv8S5o80JpVp5XztpiX9r3ZSBMxv/tl353seEj0xpYfZf9wTSPcAjNm22
6nKyEwQW4+DKoaO2yzCjPWRyOr75QKbpaSbxDehrmvaI9WVbSZGLKdMAcuIjn8QosQg+38QmSM5u
fw38c40/QsuYQz685Jq6AzTAGC+JIqwUKj2kS3s3TGXttXtHJNXdQe0oQVhj6vu9UzLPGZzxve66
rwPO3mbFwE/jzyJC8CYyw7cnULpHA6Nlz2qqwC9efUyvW5c5hoG7eyU0ffXZY3zxGytucnqRuFZu
PENaMX0nJIZ8lH/lvLb4HyGz4fDn4+NzWi96lXZjmGCE5u7mvfmuhIkXs6FTp47PI8CZnGZ1OslS
8DHg8jPITrWtw/CJ8IzVgRk6V1iT22NVvhj64CGdIUdVk7KXC5Gkeen0JC3CGMgSY64glYpfq87j
948lrowwAoQ/f/T8u/L7m+ehiv+DFSkh2gQayIuVLL0wot1ZsYkVaGw4qoDSpt+pJV6o8P3PA3Gj
i3Svxcsovh/9AISp0pAssXK1RCQlXwsvY5fHzTb6Xboo3/QtLP9/id+j8+q7Y/8PYi0iK1Uzl2jq
V5q2nDbPQc1J7EsaiK2g4NJxTNcrf7ja+9ZQ/5GMxS5lkOOAlCYeXnKSsmUFC5EJweCKXLKbQho+
qWKbPiWc/ruGVy02TU29kqKG11Fi1FYXdxNqaGFKff67lU8yw1vp16H1IUbmg9t4sqWtRv6rbL4n
xsmvKzoTvx+Q3i/VVNOv1umbyGc4+jRDkQZeTkQvJldFtPCNVy4fFjqhvGqpTimizOgEIGKMXUFX
xWlKK2K6ZYqFY27/F0+wtwJPCtiImWhcq91ObfAkB1oLwkS/BBTGw3v4FjxNYl+I07K/kcW+udx6
kqbUlv9VsXhtlixjywBuLm9Rur9QFQYgmSi01R81Sxx0Q0CAimnhh5nDwgiaqJQ7LnyrLF2jJy2r
3OzQrUvqBCHlxWr83lb21sxslmB7RW6p41lKVAuMZqx+BnYJagVW8g6AM3RiYrmow7XfrDYsYbl/
GDGOJ4sPr82IJK7/Z+LLgXrjQfePCXCmDZSQJ9vePptQ8/HQWbqlWug/SE6eKfQSWjNPOUwWD288
9IVrr2YRmEs0lFwyb54Cvr+FFHMLyCbZ1eofF1UY+AKk9Wr6uvM8D0WelziROnvPdaDLBWNuPUZP
Hxc95bt6pNuoOWlw+kJFnLqVHjcNBF/SfRFNnT+A4JnmzktY8WYQeqvPZ4/0+6PHK/iz1KE1U/0J
5Ytq8y4cM7OsTrU7qCcF0m08Gg+CnB8xrV7SdyW7zdpKiiRR3EXC0h7530NO4gTkxTnnhQgQPSQu
XKwuOyAtcJshpKWu1RSK1ExQoj0dE0zgkeXTK87+UZxyjA8z1KDuVKe+p1aSdm/zWADvLGAS33dy
ftpB+008SF5a02GK6EFyp+mXKGCYzaivxOR++avBo3Kh3cnfQVihEIZ2mM7/OvPSshIpvcBAFB6r
ndoOFmH+FNXQGsAQSGfWZjEeqV8fqz8Oj3bgUEpa/8BlDGcVSzVKk96BTWQXKuFT8pUE3y3i/gVn
6rD1nRzb1p+AeDpt2O1tjlFVSd1RehwQruIbvKRP0afUX9sPhsv40h9OyxfFfLxImbSLgRnJyKmR
7+K+oD1yJQSGjxPo8yfYIKno9ark4Ua2m2OyBCqSEgygXCYi70TpfNQK7mv8T0AMd/v46tM6Cgdr
OVc3v09B4srhl/2SClbImXLbfXHEvxq2qjFKXUaewek4BofjK7tdD2BBXRxJOd5pGgBys1Z8J7cH
Xa/e98r3DSwVR1g6yZOHCWUKOUTOv1J9e0V+0u5EKG1LGGisvoU1XA4o7alxqRxj6ehIU7K5+Mta
DrRV+RssGrMYme1nsX6djwynLmyqj71Etutszoj6yC4O10Bt9ZRcvRSLlTbG2628LO13zjMdneWq
b3RJIDrZnx4ImhBSgFhD05DcmGn2cOex5TztJr+3jlH33IIHTDd3ZWPvbi4uICrdLmWOJo7xTCHU
n7j6N1rMe+4F1RKiGPaTDA2vepooRUmMHoOCXwCKIDb+4gNwLy1pEFpZ8CfNLq9POk1C53wLlVgL
1b+eAlU4GnXFNl9sjMAet72b7orgwMplVu1STo0ywObVSMwIY6IXu+2RW6ESF+3KcHXuqVCDfzhZ
g7X4sezB9MI1W0uxE52SJThoSxlpZFqCUD+l+HR+AvWpFnB/OlTheVlh0DHMacKeGo5akGwOsEjX
iuD2TBz+XbGyfb+xagtQhNPYY74CkWtPUqmT+4iC7NuKhYb46k7SGECfcFn4TcXTuQMTSCt67yPG
vEuyn9nWLQVzliyh/eMPHpe9ULWbtHFw4NuaMU+QccMCOsZPmKsrzEj0hC3VGDbR0aUjGrq/YJtR
iCX/1eEeOUMklqOOU1kfxuviv7n/a1LqQ/RR5NhpnSSblyng4KXA23Xi4oc0muUw+8ySelZUiwSp
ls2N3OtLnsgK4dXtPteXPz2FTvnBGcNzGwGrbT7CFsutRxkFBZ4J5x4dRIvwTkTpcvuV+fPZLQTM
OaCNvcoiwjBYNW8MmpQcBT+9byCfdbfXFyvZzQkdoT6/YsOV0w3kkO0hVlrHLQ8B9k2hv5fJIe++
DqgdvXYpua6ldJVSCMkd4+RvNk+mOy94sGokY7rw97gndE+IM7mC05e11N0C0mjy8bFocxp+s8n4
0EcO6Y5wppQOOBwPoCprqFf7tkuhV+ZxW25Xt/2yiX8lYrFDEAJ6wMtAn/wYauPlO5hIO7uDI5Go
N4yL3b9k0RNea97c5NukXD8f/zkfLTjZXTujZSEqnIBFd3UMqyiJpgQfOx35bwiJWMqodlYiD1Aj
1nHQedXGBYUPYynxIfmjmIWctDDXVsl7tmmPD8dmP62gLARot9B8xYLBo/YVH21f++Llb6P/7iXi
7SwuCxYle1mIvc1p87uaGGXOKnFmwlUfXFGT74llpBJibEbsDqXmHVTw1oPQ0HRMEDaiFpDlcIv2
jVBPaVEjcaCIwUx6Bp9ca7rlXbT/yroKr4126NytfDsaPHAznY/X0i5vvS8/MN3yWTMKkD65aUDa
35T1teyDRRW4YSMgJawLElWy8sNGLflLC3rLsb3//PYjE0L+/pzS5cBuZll8nnp9j9ps7noZBxdx
Hl2LRx+vCCYW8B25VhjdocYLHbZgveGmuJO2TUInoYGVHRAZfnK1qiRYeRzK+HjbYoU2QUTUwe6f
LntTu1z4HI+aKb3TOaNVPuibgccvK/7u/fxYlzDSlrsQ98c1/67pCbAsDuaDcBTKFj7/NdkY1adJ
jqsmZ8tQB//PMjmOrMH46Y8k4a1CocCTPyPKXcdopQYyUHD+G2jnYQkkah76+qNSUxegBPx6j4i5
ZAMCLz4Z7wLq7l8WvxgZdxjniCZzN9BcjDacDTzwiNBiVVGTcF4ffPXFrQd0haxQQjrM05u9rcs4
4aEAWBZsOLf9OS/GAw3tjHwaEN6lWm7dTiC8ZAooo0WY2KrEaoasp/57D+Nt0Erj9eH/GbNxvUDA
BIEykq3zy5eUjOcNmN2s3o5f3vy8AByTfDwRIydUVTm69MiSBA2KwGjBnP1bZGpIIDgBFRRJQXgT
z79bVRZw19cemBuSBBaCOvk7EquEeLSMWhJw6sfDguJrspsjIeyH0fUpp+wDUy7Bqt4fI3dI9SVn
AYwth+QK2wjqey9aIrI1RS96wpDzvzQ0W7FUEV1YkBqAfqm5W1de2t3PQDs7XO5A9sj0ZbXuJaBg
LThfmA7kWrQfYVbHiLTBBYjSK0TFaBZL1rZ2Zes3PNoDisBwGyM+QU3ygvBf8NDobVMiM7AsQs0Z
uwURtrhoNcrNpb9AgFZ5N3CANbUlVPWHZmkD7XOld4GAXKe+PyOR0a2dpbS3ZTpJNwA5nb8rB4jZ
LukoQmotedJwdxigciVkKI27IlV7qj0NWEVv8hdq4cbRqUFXp4MwEOV4N77Qkr13k26cEQA+gJ4n
37ahFgmlgFoF63vF8botKhKU8Nk00FVu1/QSm4AhoQUSHTxDMdCkc0itP4/Fr9JFLgaGCCyjDt+5
qveTdvE4qlQBjWEBGS37MVjVqi0bEDBtlvlNpAtzLN6eogFqEfYKWsSd7HKvd4GBU3twiri3anui
6OdvoewfpO6F1eXMnu9lWgm5gNoqg2WG8EHMSlHaopdhVOtvEWFuMIJmTcl7BCdnNQmBCRBEDaxk
dHF4LXQq6Z8HdWpQ7ULFlx3gazL8mWyXxNFtweReWR4QTCCdDWkAbzsbO2auz06m9Sk3h6I98E2G
2goe3NJ+oQYf1d5NhGxryoA+YXLLTZ7d6QGEy3MCWtgr4b9I2uzPV48OY8cpM7ler/czuh+aYLQr
cGi4p+muuJSozPgbiOHGwSXTB2VEIGDg2rQqAcDPdrBs7TvwoINf74glENwmRjxFSIZDTouxvGQU
mR0AHLhyU70rCwGec3YhssrfqPmbC1kCtrInB38E2hKEPwYtx/4UK9l8hDvrISH5ubNZqoUEM0nm
DX631aDJuVm4wWHN0SyN4ro+3kPZvQGOMlKuotb6veWeEPEFZJ6rHeb/8lLTktSMN8GlHsMkiZOa
fn/ThRsguJaN03ZLPkvuLObWVrThbnoSa1dkka3CWorNCYMWMgt97D54mKTjDSI4WdsJAtrdbx+8
hu+VXtDFH2K0VqfsA2ahc6W5ry3UyEWy1I0NEIBd9S/Y+Ynaw6/fSxr79YnqIzETLELYoolYIOFu
fsAFD5iKKG/pnOVfjRa4/7VWBCLBzKjCNHgaJ7psA0zV88iGpcFcKMMuGSAVF9ncXbepYmhhcnre
RFV6+0tIrw4/hAUfQ6+zTX7iJRt3RRtn/H7W6U11f4aIM+TtfxAVxUw9VJNTxbx/Jw==
`protect end_protected
