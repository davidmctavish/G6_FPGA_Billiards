`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FfK7r4S9JgKwOuf861Uqk5cJ7S7TlOsWjthLLN7V2B/Hii0PW/Ek+ysmCxHmFWBU2eafqNgAtu1N
zEsiqUZNfA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bn0GtkGnGL0LNUKBmV8EA4PY/EEdWQ5AqeDEl7pvsNd9xM0SCnf/nyzUWvKLfAU5sX3YRS0oXvGM
gKskq7urT/q2r8tr07hlRRGKzfKC6YCV3uT3U/nUAsr6jXdSMNe0AaR0h/qqd6yhSXd3tO+bVX/U
XDg3BsdMPp3Sf8hsJ5s=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CQcKj0Rf0OT8NXdcknnkQXLzsUfEiep3kTQjhot49PWpPzweNsKRcOel/QHmmFYRYk0po9rhI4n9
1FEXzDb1/O4ShCVyP253wUajy016G9IyAuUmseQeU/qF3+5HqIPzl8v5Np2l2M6iOyJ16L0+gWyy
tNVYxLMf4LWOdkG7NODmvctZ+83LPZ1mzV2TJkET1F+K2LIJmxJXVdZgC4r/kE/j9Hrd/9/u1V4v
EzleJ0/iZqAwh8qT6TfLscWIf9c2tijK68vIyxxMYRytf+GmVmmitso4aaDV2NrSr3YL/3IBwdKi
WgyH33d0M0S04LSCIGpKlEhI10ktGjc8ZO+FxA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JTljA+bs1EOEpjVKt3PQVqytndphLEJQw5fgfJ/XIog8SmQt5sb0AbowtKBsZ+UxHtpeJyYtAFZb
PZ/tajIX/J+BwOum9MtYUo1FhPmYDHmhY6pFxs6hGKcHiUevTqrsicsq62TxUih4yZ1GA3gZI2aP
3xgmlVx97PlyfJKiUZs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/WMNqakGI+2+f4oo9l+u6i6TjdVGaxvZLaQEJ7xpucEy5ToB9g2ytYOGlUo6TrMtbiWwoCsM3fO
QthOHk01giN7ZezXPn3suLeYxx4BomWYIN8HzznN1giRpKmtJQGX7JwoaXXZYJxVfvoUuJptDkFD
LyDtOorZk4kkbMSxtsIkNuGChMcOQUm04elkaeYrnMS+HM+iORruBvQOS6oFsyTuFeQ2vmOW0zhw
aaVevjip9AN+Af2auzug1nXoyFGFnEyPF1LacuBoeDFJO66SCDnyCcGDlFegTwPsiqZbNCtqQU7S
kpmfq/fKd8f5n4uBHTZdFBHMjsruOdD4t2l1bQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62832)
`protect data_block
AAQRq8b7M0FxlgL1rDaskPffrZCyy9XBS/jX34yAUwwOD86xW1n/QrYy2PtSck7dQ6rRbaA2NaP8
D/wZCz2XaQBTf9accWL+/HZ1h54dDNw4gBvfV3ESvFe06Z5hVMfYy0BHcSsarH0Gex+8VdGD+7iX
iWqJP7dVgnl/IvfG/yWGOnX92ID3kUmGpwKohUdgkRIIy8nqIZkI7U1QexIP7q6tD9lUvDieYcUq
aKydDhr7KcYeGL6W4ij1zZWJ2fdROBk/WthKxLJmpw1CUFqfHXKTisDAoN/XY6Es9qO5RGjPwd1p
j4Y1JE8MONMq9hKWckF3nJ/LNvNHdZTQ83pjymdrsjjL06I4Uv+w75pkjUJmxL3MMR40aDAp2N0I
4/xlSv3ka2o0ouv4jG2ncgZKPW5fyJF8KTQAVr/PkWSUHe/tr5neeilufDDdpBINxFt4nosh9qcy
My73QhtjWBFYzlXOSz6NxkAofyOPpKYRL46UnFLP7LYCvAD8BguVLrwfhB60IaNouYq2q4s7XHud
kklxS2iaWFLoDixGxLPeFuak3Z6z1v6S/LMZyCTTEecBkil+vChtYo4xRG9Go11R1/Gut8YwQ62o
zReR+/WJTMB+Qqh0P6/t37hN1Y9ih8AJlcj4IgKX9N/6+luEtROgJHuDMQ1gXNze0pvKrMUd08+L
7T1uyoyS00roQ8JAdvtFAXJeR5ESqDZF32ks2oWtYlpXDp6Du9iBlgI/gXXXQOhSg4AD6fwD6pop
jWDEsWggcxFPis9ITLmpnflzJwOFo1i4KOOuekvDZMCKnig2yhONzxXK1hI/uwQqo00OaJvVdVS2
qY/NqhZKXIIZAjqJSmkearsi3RSiymujnjz7RXbN68yeZ9tg5vPBdOpIZBojIlRu5JuDtFEJlPFd
/uycxPPJtqHMdn+BJ6iOKXIT7ypy+F+cXMuAc1LnmkcaNegPVyW1wmTXtzy2NDkhFstj4dPMo8rs
Ml+WiAof03jYMQWvOAJOlIICFbWGU8wsC1HCdMRtdvDMUnnoI2a0gvowCId/Qkl9USbncxIooq1G
cNXChXRTBxdq0uy+mvs8T2PjYodDl3NzTvzPjYm97w1fU5v25ytHRUTLD7BFkE4Cj6Tej+JQyNwr
vyDZPSb/C9DsD37CjeifqbMsZZbNP3ZdDCL6TS5LnD0GV25t15jOsbt4mCN/vPECYAbiw107BPO6
jM7nBUeRxXT0saZ+xn9aqGxlrg344CkuXfbyo6VjTo3y5llnq1EqP5j3D9vBSud0/VdKGp07XBrE
pLYgVMRrbz75kV6uC4zN0RS/mFzHRQtaedWMpPPOqQA/+J1nLHHC0gSKp7EpkmUdiTkSnin/1qVH
GYb500yk1cawXsIb7WCAA4ClIY63SsHXGWxc9JxadWPyjSyzg8Hzuysadd474sqzpMmmcg/Rq6ur
0RHzwNl1etkfYaUddPLk9uWW/Dc4a5RE4OCRQ9TkDyj24RH/b9zlRT9VYD18Q6QI+yB+R1pGzSdO
ELNkb8TpaMTZKsjk+IQvb7TsNT2j1SNFcZzNzbNTIZYuRnJhSi/+ghyVGV4iHSNPs+OpdUFopNeC
amkxqV6mlU8vZ6huCuWc0ze7T6AqatVgvYwERUZLxoJm5+0sb7mkFqMCF/rL3GTuJBQlKTOy4/QR
DX6EYIddSfXxQUSlgozgknuisTDv8GfriXoKM8+vudDVAjwajqGMGihTrA2WEDEUGcqagiMfCE5q
+1GwgabYByAxtZsX6dqDUD5V6CwI7I15kulL9F4+g2yqxVHyVsUTqBZm9ZUcjChFIyiWdrHUhOrV
5NVcKfLcFgU5TqWqHOY9Pu+vNSq9mVv6dZ8Eo1zGEu3929m7qLFHxzuigHIJWauGuuu73C68AKKE
A0HYEzEA8BOZB6h8il/xwaSkPxTD/C+rO2B3pMqNd9+cYTGwUTEaOsqkccYjqjloHdW117JMKJH5
+u6BisMGfS3I2SZAf1wkFoDF75TWnPYkf7N56YPs5oTdIvZUkoSCVkTrMV0E6BTca7mk+l2ebpZp
RTuWOaeiJa86aIIHtNUaBmm+2TiV/sNYqpTTvHw95b90I7sHMdXUUmuJwTDHBDyBw3/DC6VnKDTh
dI7rGjuKOHX5b1vtZidFWXbKP/PV0KQ5Iz1njnJsAqv4JJZMNA5tBzRuJjPqguBRcrlvjBxXaIdu
jf+jQhZjCFAQ15B3qseF2tSp+Bwj4cbryL8Jwd6LvYeujd+t7IMH8RdPalZrfuqQOvp6T+V3WVvt
7zDBlBPX4jjrWkd0eoKlX2W6wvW4dMOPHxUzfeQXnDGODDOa+Fx/LUnVgXmeSQ4hprbcAIUaqcCL
991WTPPm2w+NyWOm8NHpejup7TkVp39E8FVQje7BUJX3V8BCocuzqPItApALbcj13gzJV4hTP43N
muT1jl310VIemegXa3IWr5lTp9Nvp3t1Wjslm7WPuQBZ8y638RzwyCtmg0ypynnaoUcvjUkHP92p
9m3t5uKrwMU8Icgb96q6IRG7WNP8AwTIdY2RJaWhytbSmQyZAsabAEMi1xrJsAyeGs3e1JSUehQT
7qSZAQA0r4fDCJwKEsNl67bPMdl2dzSFtLXUKoDUGzrS2LpVvfBXBNTHSudW7hOyaChJO/DXygo9
fwyLSGN+WUSXhDSb+So9n8IiSndfQT24HmreRO1OedSw8zcNCh01WCzaiFeCsCYbe687WpxhH7S1
huZjp77FD6FWNq7PjVjcKfKtJ1yzarAMkk0YVollZGltItkZSc71jyvnHoY8pAqV/SY7biUJxKTu
+0GRQ+JgcbKt51E+UucwX7RX368P/lmuMemvjHoDLlO8dvYX/918f7I9kDwbu16mUmIlZr8EdraU
18/PoY6VfkWkhZHP0HygTioerI7WWdDs9YTnp9elGb5y+hn01KQyLF4hXuluRqdlS+oFUE3x7liS
mzhHhNuIPFEs27hP4WlNRLpYbhRddr1AypXluHNqvQ0+MQ7TwKK30/lKAXnasdtYGdLYqIJTgT9R
UgDBWCcXRfRFBqKZgMmh25LzLMxg3udbyScFEh2NGMv6MTsZvY+6Rn2eR5z0MT6yRot9QH4lcuch
3dj4CaXmjm3gVhZBWfTHOOmKI+Yu2n4oqoCe5dU5u5ggl4Xhua2OeK5/jXAtUVPXJok71op11MT6
FrLOnlqGZhKTbx6Bw7ULHnHll/j+ulZAbhGxNWGxWP95JdAnK9I1EjENjRHUB/2258VBhtGIYO3Z
6A1Bazcs6oeMIv6/xbOunkS/Y+mLv2tElddGSXPIfIF9/epOGi2cI0h09GEpCzd8SqQ6ONxjHWBl
ju3bZe4VqRKa1LohuALuh+1U0LRg+T1xJiTbPE2WFdfHhXZb57FFyvSYykODoR7E0YRO2NebtDfo
hUoSe/PDirK7ymbfdGSu0ndPycsElBIktVgEcJ2+2gxvOGBfaLhGoS+wm3zjcnuas+CSGJIUvV5w
vlTmbQxW9+bbfi98QNRMGdbTCK9DAuG74+YHnWmJ/ZLWhibNIx85pe8roPXvi/mwgrrk8wMWsggv
mFO0HwEcTAgitO78h+jesVt5444m0SVJmMoD3afNvNphwuFRve0xBCTRWLWNMwq7GGoOpqtETwNg
Ac6zDv96qg9iRw6RX+NicpTWoYvae4ZHIfHgPDXa0zbgFaJszAsnCtqmqEd2AaXnwOE2A3DKZl8P
816zHyOxUi/aruFCgdaZTaHywJZzC3acvshd6K3/75wTOjAjaI/9Fu8mx6A7XRNrWXBr9YRNfHQs
3u83BPLicJOzWjhbhYOHXG6d9YxvUvhQyxVvsGh2KfE14YR2qjK4ZtIBptsqj9aDSl8htJtWgTHM
cpfmDZ5A+SLYar5WbyrEySf0GyE9/O51rBThdDHXqaYSxsu+Fcpfub1lA2Y4l9nMyEM5cEmf9eb9
hhPvxRNFkiuKorNxUy6XP42NHHjanKfXK2TWIoFlEcbzqdo+vwoceVqTaNEbUTkyLOTLc1JKz464
wuPYMPgjw0JEqAX25TUKofDIPMqthUQYqcERVbVXsYNnihu6qHZlvuOLXTy3aaO00ttmQgjTVerr
HE9pz2FLVvckKsfrL0eLpAPAzLPiKkBWS9Xlul1A54geYi+8PcbNrwF1s62bnhgsEgeGR+dGIeNa
3sa0jzzcWnfRB099J41f/Rdd4DWhWo3tN8o82Ov4MprLxns2EALmZRsvppUmyzxgRPuwsP8A57xK
O/Ra97aQWhFDLtjFXJ1UldNurYSNRKneGzwJPL8G0WBmPQIigBfRjki5lTN3naLkTprAbH89oNmu
CEAkXx5R3c8EfsOenoibSJ7O4luQ1Mf+D5VkwBzUqan/I9st/YuStvkiX1qNGoGXdJpl1HZrM26K
kZLaJPN5F08QYL90Smo3FccuL8rS3rmTllaheGRVm+pXdnqCm1K5oUtAOOwEEcKyuVSL6oPcsC30
8i+l5In7rbilzd3hKlMHCVAxTpZCVdWVfFRgFoCHfqHJyJUOaMfuyWBQLkvSwTmBiDNsdtrxT+zt
id9Z0/qRkRaqXanEbHzo5fA39yEjlldqhUBJJGIXlag8LS3J3HGd3CVqMHxU2FIIQfxGDKKVD+55
rS4IYS7tmNLF+S7bsqpACqCFziq1Hqp4uPelL4yblDzzU/0yX7c1bq6h3/citYzgcxnazugbt2sb
oLdXU48g/X2z7xGjLnVl/I9ABuwcQMjps5f1jk3RiAnfmVvb/VvplvyMaxorfMHUjDtQqDOhZK5m
BDx0pi8fRex9Ypu5NNONS662qH8DL+dmDqo7122FNO8VDYO6TwbBFul/FrirAhcH2HioQn/ZKBXX
G1gyqwiA+KC3SMlEhVP+JbBtXae+djZxPerEboThLJNqEZLFoa5YT5/ll2WX5M+7xT7BDsnlLa3b
wnL13m9V+MEhMGA9hJVDztITwpIV3fKa3G56v5EMMw46kfwsjfkml+WQOHPx83fzXU06fGiS3+u5
5o006G00JgpBGN1YPAd2uCv1uIiB0F47XrCIf2qyYX234XjfD0aUmFPJ1wITBHYCbVY2DtyuJcpy
r+kL4zI28HqFKvGiVHSDz82qlgiQvvVpP7RISIMR/1o0QMPwMI9Bx9Tpg3W+23lyyIhFQLy1GK5/
MnuQBeX4soKavil48ZmCwWOUsqXy9jdaxjxw5dXgAY19+nXBYVHYj/l+w41lqYO3lGI/pu8SyNoy
BgiGjs9vc4rAx5QFxI+lVxoFvehfgbZKnOlBa9egeoK+mdS4k0Pv5lnmdr2yAWnyxGQ0hI8wRFj4
SVmAsa+yvjCZgykUvD4cQbLWmyZwR+OnEV8gbVdmOnOUiPRhdtC7NgBydSAnF3WqAnblYPGgt96U
yqgQ3/T8KPP8lPGgBR8mGQv89Ho9yCW9zrWOnQeK6J7gvw05O4hzmZebs6+GslES5ZRBJbYPnzxG
/VxGmGrebDFHRKnCYXhXHf1zZkomUjHDz2F6OI84xZwD+uslb3QKRqFep8EauqvpwkdYAbF3toeO
48GuHVHtBtukdtjFjSeollLZ0/E9jFFgr4E9N1ikUH5Y3mm9hWJlt3jHgZ2ds+///vICnjgwP8b4
MZkcGqK/1ZibjNOeAmTZJi4Pyi0BejinbUsubyx0hW7ttD0727A0S3shYdDKvt9IGWU1IFvi3nOx
N9gxoQdovcxjqmd+RtlL9zxtk90AL8bF64cfm/no8Cr9eGWlktnpZmxAzgf34dF3k8bZGUHN6+wS
b54id1/I9n92YFPDmAXjYSI8DCSvEG0iSvCPGwNarMhlREYM8WCl2HXIIc8oaLlKFSbTOh7idBbB
1vpdfx7rKEKohJWYNf+V2scSC90sfnVHYat2imW5rpA/RNRB6nYlmcYy8gAoCsIytP7vcPw0HyIe
3RQSuWN4U1v/+n1xh1C6vd8qPqZXpIR0X/z8LlP3uprl6yQYZnx8TIm5whCk3OO7OWQIwUJImGnC
0LLv4xxSNRE3aYZvo5689COdZqOjeGw82Aou2JC6rScGOq+TvpsLPBwnqvekGhzc0IPKMAL27xA0
pmnQOk6vPoy6BHOtkfbhsysogyzs24LZHbHC/IxcQPv3JIWZyiZwNCgDwTH/U4kK2zITQPCOoTDw
9TnksNE+jJXpCK36u0iHushrW6ulfoHCZjmyOATmQaOzXekVDPSQah+Mo6HeKVMstC98oIzxmf0G
+1eY1U1z6fo/IavCpAPoBEtejhQnCGUAPDPpfAq5oN/n2JMD0y0QoMujStdmsqTLtuExpX6DKNaZ
d9XsYZxFqeO64NThBEG/RxEWJr+lIG8rIYChEwLnZLac0VMxHjH5WBWtLXThc+RYrDfINoLHd/MB
9ubeGWYPNM/XH1TttlW8hXcj6sM/nuhy1UtkbpxNQMsWqaPQJuF1fAHfv7k5AVJYBjOTv5FavUCB
nnenZ92RELVAj3VWsGVLc4pLDEXho+U0bYSFd/WwKIgegNDdhfAJVB2g41KDOJuncjacOIPGAGOj
uRDIrAGm4G4QUkFwLjTaMfOP/Jma70Q72TM2hLYzyaMzglVfbenIepxi8nJKWD1FAONdCQfS5Y/x
5UR0WCnL0XrTJGay+UFmaCH57+s0DXoFI0UBu0uhi0+HF6bP5qbRH+x1cXjEd1VTC/46vxSr66nj
LL7V46XygmRc2gL3T6HG19ArDNFc5y0eSuwmA6T1ewiUC9qsHWyuB1xNLvlx7/wTuyX1MLH8V6yw
OBQuudeTCQSZxfnwfYiWv+W8+ZGTKgj4WQe7Qv7dsWrGT1yJ13A3GuSxBQnYGMPvTZ1j0AsHqBDY
B769E+3dF7niugW46DuiHJvHHWrQLGjbmumNoIStIHEuhr9xiXDQk9lii6sxiUG1gERd8hijmmH6
ibzuG/YKxdZs13eiIaRjH1UONKq/zQVlDn4im8OHcSUxhHNiCw60t1Vg0xv7b1nxO/qGcXSOxNHD
fZo2gv1Y9yOOpHHrZbJ1R1d7dnl4abMI066kMi0UYHyapttwFiZtjNexUtyaHeXWwQditxJ0dJkp
VfYRUZhfzb7zxbv+9HYKJkjQdAFiKpSzxkRnbkpDMLY4G0x1v89crW7cozbDB0xzg/O17fse3AsQ
u3er0zh5atPXoiqrN5Pv7QeFQmtG+ivEJMg9xXH9m7SFqqiOypQmBbwhnD3Zaumqm7trM2zUhiXG
PM6ogCUsbJmoBsLj+4X+OQqhy/5WBEhanMdc2aLzOJRe5wWggRzEc3iQ3zlc8/T/NbtrMmQBAsSN
9Opz6oLdsePMFRvMC8zdVesk6c9LFo6UuBOKK5L0/SmQCim6qAIDXQzAW5VGAKnQle2R5tY6DzHV
9iAUuohwz15XmY09VXdInNkBSsnEC2KXfjzsp7F9LqyO0pR4ZVQY3gVxDN+YN0cZ9i7QOSiIJHNy
I6em25J+OO+yIxGox0Og/CnUrmLkuxbpLoTGFq1Z8AWldSDKVy/SQqI2zF13BKjcZvvrmOuRDvO6
ipOayu1wk4L3ES7zK7qg9Hvu2LtzDgVJha6XsL8RiXd78YDi3BBiTAtjnSjX/UEqtzvV/Ka3pVWY
AJwOH//dl9wrl2LyMpOTEPQOJq+iwfju6Mn1tusKfpTX4Gp4FOGyvuirG3MvsdeivdTxJ+sYOV7U
woTnls+0mvcsWQzQY3cTcScONG/AK8AzMnaKrGLdX+zTc+NZMZjo1TbmEvim9QmjzGf1i36NtjX9
sGnxln+rWVWS6p4cFRo31QQuAxyWfq+QaU4OsH9j+uK7TgXvBoCQ0cc+ECHGCne7F7kouPAx70AT
m+mkZ+wKOOzm/kKY9JPf6d36Dha7CoFJkCQLsjbNeekslS/bjssCB/Lpa6IFaV8TAjnDGxHtYW83
HkQOicE5sKMk35emHsMPiXeGRuoQMdmwgVFE0xOwL0ERmO5RVLygtpWhbn0iuRw8sKodoBU9027L
/PvQZFi2Yl6MfK90OfTPO4vYDpXpctmD7e8PscueYwXidqliFT3/ISwBHpqWAL24H3I5499meBPn
/yXl7iT9PGVuTuQZRVC5gu5BJBzKiwiQf3p/A4HQLCaXlyhb3RPVOeFQlVX4UMf317ZQav15wM0O
/jbjdU+5NfYSVpiV3q8VRMT+m9I/S3NX12M0X6PrcUzAAkyjdurx3uVBqe+z6gkBpbHvawyDadao
5VZUFUA/22FC5xy6a0TEdUijKjYJGOGpJ7XZDG/Ry2Od/z51gbLodBVlfKrajSZhbqA6/rHbHuA2
dhO/sEvUGRkobZmZGBOG+BQdJdzZfFKGAct/vRcPnRoUpb4fj347CbyqUYe2b/ydxmkKitcKCZ0U
QDtYU28S3fS/eav8A510J1WceuVGw2P1ZKVpxSWatOSlaXNSW30F1H63QjS8FPaxD3knUgZVtQeE
uUwnzB6eam1/s+9IDQBlYZ9cpoRI1qLOEPj3bBj+sdlPv4MsNWrqQL7tBFnwz3yYCIZ7cP9RNsjV
ObNXJGUUbI5DeishA68QG5GKlxpDU+zvb0rg3XgxSs4eEoiYfZ0I3+fKSnqH46TaUUrtI1gIvwHE
ypUT9bdUCehj0EuhZU3h37JIbn+mGb7J4N8O44TxIPPt7r7dOxHWGZC7LGybx7h2lN30k0/TNQTZ
ipxsVCZWaD6xaCCAX/tgby9oKaRFEL62yHEidjAimTEJleVVT0oBnG6m9hN9jWCTihesF5p+ebzb
5tamj7jVt3ok7MkKs4dPtgqH33ERrT0Q2Mwu0jQM8FcC0mfYu53KifnXkRpYaNKtEK0QN9ixYFe5
fWWDIqjuWhFuaL01roPT3swW09iqbGoMxrmTO/NjK6YFrQcgmTkZbDIZSQMVEENZHASlRV1xAdfa
SMh7MZlmwea+Dhm4Gh634nIQPxqRfpj11chWCV5dbFwWEa+R407f9FPTLgpoyU/GUZ6hVjbpni/x
z5oJLY8j3Q/QGdtzXTVF8zG1hdqOsKH+JS3eGG66qxXljvN66VW0zK8YGk2n6Tf6eNeGJnkhYCJG
sdtlpYGVk7YOsrbq+SvNDhG0FeUQUZwFEwLUaqlu3f3FF29oMvuC6pPBWd0ElF0aK64As2RAMhS8
CgR5uGBHfiS2pd/cvjQeEppsomMr8Z0DAxeUtfJroF7gav6PnIHJId8hdeXpqttiRfsO8njlet5e
D7OfW3uP+nvzhNuQt4poqvKzGvu1ulrFznnWYwwqMf4rbuvdfy1aEqObsp8/KlRIuZRzA7RQnbTW
T+aW+veqJgCmPVIKmL6Uq6Ss6fP+d8O5puB1glb6kdE8gqYPQPe60Y5sfjZNBS3OCtyp1EHOoSxf
4wNH5Ce0ozpwFhZMFYlH/mP5ZPM/3rq3QYZwu0a33vDiRoSTglhGwiptrRcWBvoxMuYfhO8BbCBJ
n2YQE1wQ4XLu3HNHd7SR5wykHULS1J8eqa8kALeN03+p7jD1mTXJvZzd5E4nUbLoCIw5VUcKMpGf
tJHZjGRUd4ha9pwcG5AQIec91dgWBx9H8xLINoc1OfNVI9WkhcOn7QWaMUXVlO56xHzseReDtjKP
npz3nWOVxylalci88fCqoraXP/DXYOA8ALHIJayrDX3ciP0Fxm+DMg+B7PndTiPzheaMxA4Zatla
GSaMbqg0hMUzK6QtTAQtj/44H3mmQ7RfXDRXAq7VUEkUwWzvrldApyBEGHP84k5lj4eR7F8CHCKp
34yoo3h2XRnBzgd0+bLsmRLhxoXfRNpazznLK3L13yW4rRuWGkb3HUyh4YDO+Nc8sTjXQXnB02UC
SfXc0fkExuD8/6/Is1NSjVAPBkbxdG0f1BQm8lFmEMIlWhQs+64I+xkhX3UeCy+RpFSydWQc1jxK
FG7tT1yyZoKdvuWx3hUG8jQQyOcet8vmpusBGo/A2sM4gOH6InXSojoUPl5ZDGL2GlHKUjhzNSqz
OEPncUgmKEg10Fjm98wmMh3W+h8xdUL5g3s64ckpdzyngLBJbVyDPLfVWRE00DnLUQm4ufsmv2gN
eJ/2lAERm+fJTkKDd0s1ulA6U0pekulbC42MxUaOsJJMR3yUdcjAKNFWqK5sq1mJB2O2Zxrbo+j0
wfNDbp0Mjdz845maGnjTcMneHSYwxvHmxQAy1rlu1fjMznYm0AZCO8vtEnyPq3dJ+fvMU+BcyNHJ
NQ/cCOsuwubTVtyJx71wOpR3EBtSRAV8vnAqvSlT4HNlye/Jl/HHevXXNJcImhO1HeRqL+lJUh9Z
L0RNgAuakpk3RWKmIPcNBEUcSJ6Yj/VL1rScX8x2QIFVgA142sOpBo22xMpXlVnMg6eW6q6wQcWy
QgIIl1D3yxJx48+9NVastSlGEd6OW62bM2elIQ29RFfUH3jzQ8Lv/KteIMjPDlXvsSmBLrgvdIV6
KnafXSKjH/r5jFZ5hf5TzH3vraSkVpmzf1Yd+8jmuqtZMYp/FuybjTPugiD2cj/KJ6wDvxG4g8qg
c3WpjD1Zy/uY0YlzHSpOCrTbZQAln46w00zKghrtfsiTd0eyoQTZAr4tPr742jJc7JrhbOYGpNhA
nJiUuqkiwBU97njoaKGuBDY5PbKuYGUFW55Nlz0BkLZ7iHbzvz4hVxbag5xtpY/dmWTtswUJGCpQ
DPMpVbHEe/0tiVO4dHkishOS9HT9wpiQLnBBlVnePZTKakOLoz9JLJWNz+8UWHQBPZp1z7qQGybK
xk3WW/wKEORqMEU6Cj1FdqjNLBDDs5sKxdV3KhnNudUIb5FmrfxiIhqmJLuSIf94xqY5RO9/m7JU
xAnJgPt7eyKjn5slLXmWil3THggbQ8wx+eoLgXmNBogzB3C4+oRI4TRX7vMzYdtf70JYetR4Sd3y
JgTUz6ZW40Yd4E/0AX0Vok7uI9yi754chqjYDNH9xEtOYe8XWx0swjUHy0SJ5bqo1azui2SEPo56
ekeWsA/F3m0TsbhijuM6mwy+N2GJbLTPgoAlcheU7m95eGkRSO/qcrJHy0YslpmrZRudRNoUznsG
rISGErSjMO/4I0lQgJexXAVDYi5H9AAt1DnW8hOrzQ1MNIMQ+27WEC5Sa86QrEuMWqNs9J/HRvqX
mhLN8PK1zNZAndKXeefnlmLpj+7kVkgxERtUbAvHRdz1fVYlOWBgksXBvqCSYgQqnL+nNZwCBIEb
D/LL7knpE5vqxs0AteX/QNtJLnGbX5E6adXJg/IfWWiM/VWSnw97YPjqG+hF0DwTFQcfJR5jKuka
m5Uwm+psKuth69lC34xBhipuBtMkcDgEReSP83xVyS4jt147w3YO/uxBpAzt67rmD8ofVldgGdtt
xw/UFq/Z0365E/AsHZvqJu3R6S+jcdmcCXpssYWCjO/pmxtrrTrg3O7MBQB5/EtyEMdCjM31uY7H
woB5KLAmfFkKlNskdHWpnG5dVODu8RKWLci2MRePLYusuxaEmWxKDD0XQty28z/Ul/XG+Y/oQieR
Ul2TnMXv9Svc/CiCXE8Hcop1LSU6afaBNxdQiLsJ2fjfB8sj88B34RlVj/wP/Ub5Q5ctH6VLyO3V
RWWXmYNk8HyNgA72MOgejDj+L7YRCSKbC4al1aHgfcR1dc/GEPJYU0yey+R9OVWSzaSSPsBFY5bk
NhEjy7aXM44iQ5JBjI+i8vTjRs6c1avv4qQWZk56OBdPZpvI+gGgXcOHSjzJpRsuSvJTEliRu4+k
pwlxI/WvTi9raYlDJQKSFAxDV+sS5L7QlAsidPXr5gWFQ80XANkHHc3dIzARKjdyVt55AnUQHM1i
LPSB6Hw/e6oEu1dlnFVp5B41BgBMh70J1/LIp2+RJWxecwhG28MfoJiNHCHHtKZOzzCuqUgiX8DX
As+biig4B91r0nmnUoJDeS9jmH0GEvGiHVGuWwaonwVm8ekkxB6bocUf/OYiQGrruso3I3jNfBin
XTZ4LcDR6PRp072RQWY6BSxRV4c7+A8Jg3JK7Yn5OPYgHX1s9K4gvZoWi9wtaTtJF61VfprLN1XL
/poo7dZlSI/k29fRSior4R9z/ZLKrHDNF+DXJIKfgo8fRZ9L+nOBIIK2EhRYDXy49H4k9O/+S1we
mDdLNFR2kaYVHdnie0/wO4Zfuu8t8Xg4wcUsJL7HxWb2UC2VA0bZ0pHr0hXcnSt07ofNzrhSze22
JPLfHzMNpcFK12JTCYbeTjcHDn/27pXwDAtrKXlqrSC7I1KsulSJiOn7899MYiSVNlRecoXqzG+/
1gr6ZH+xXcdvW7k1sbE9Sf/S/fOUhSnCNvXs94SZLjNx6JWdhvJxJbaYs4+WvYGRndMo6bp39f3C
V0T3M9sHuZJ8gPjh7h3wK1Vqk56luD7oMDzFdtJZyh9OUWuoXFoyqmMig482wQZN4Mo8q/PXUw/p
CvWnW6ku5TqMIi9NSPXkDIZz0xmBkQwb/nZLWKNzNH5pNInvICkKPasgH8cgRrTQntEF+dCAO9IX
F8I23IzVmYf+SiKUCC3BD8dXERUTXSP1JvPwfeZAjnSWlASJ8n8Drx1qRNfHUEJosagxn+Lsvv6O
rgARE7+EclsYor4JCPCfsjnOMawxLItBqSZqBaSBL+GgY3af4L5UlxubAg48bW0fsGayrMKNfZ1h
f3lpuC9wOgHJo6yKr8f0Tv8c/PRQSnmnyKMLxU+jXdV9s8WBJSCgPp6E3sGflCyQ3s/WbqImmR6C
36wG4uoIflbmUZ6B7rRtublhAMoPFEEmsfmYAiRmFgAu1HD+KaiMhAXfH8jZfExNIfMeWU0AXYYJ
3zZ1hcKxQsxXuJRFBD+9Fl+lmU5lj+Db3F4ana+x5Fb0zKA01Q9CfHF3c+QNNOZuEwFKB8RPkgMD
1VyObTFJ5rtUCUuDIPrdd9+LoDbKffg1V8zz6XBYlcl3kX+wZe/V2xu84bJIevUnzzupGo8FFS6g
YFybRf+Vs+R8NRrkPReIneN1QpE2coZcyf7tPwdax9KzLX8rxVTqsmWjCq+Wn4z+PNMMGYJVLOjM
kaszv29HvtKTZmTpxRunDtWLT3pYYzFj/vqT7kk4UFTVB5zvXRPIultxE1yJM+6CkaEWpbT9B7MO
eZsfLnDr53uM6vvA8HmdFm7VLt8toMcRMZtXdAfqM/Hgu5jurAk6/bJCMbrIeJ6niH/l9LuIkENy
MDapRx9HuU6OYTyjA3hmJg0oVZlyOEEQ9oziyIytyk5h3K3C6lOmEbeqDNCDta3DBgV3FdxzCBJ9
2IV83h1aMRZyrdAVOecbRad66dLatZbQcwXA9030CLYT1hZ4wrVqFKIgBDKS+mI4jS8TEjFTV1CG
U5jGWvL9Ivs42R1nesaZmOkKEmKqkyAT6QIsyihdXMcoh7jirsKhpN5lpXNV5JSZmSlTbefXd/Gb
+cVdcYIcToxPluxqRF5HemzAL0mduHHokPVa7vfbeEKsXJVpkklWZBzR+/GroxhDIuCz6besZH2M
0P0hyxrwbL0fYXUw+HSMgRkiZ5M17AdSzu6gWuo6N9XWylTyHfH2L8QsjkapUuzCXAPYxZh2sWWE
0L/vc2cXrafym0IXcWJeDjFhdkUzhu8oomYpu+xiTtdFbqm1aw9mvIkDXe21TCPt/37rMoU0j+/w
6D8k2/Z2jybqLOqzD+BUQmoaUomH9/i9bg3Jb+mqg8xmBBPsJq1BdSfHdMSIbSdARebwOpWTBy12
pTa5CaOOCFJGVuj2qLW9uOeQjIEVsYWxRqOslHuKG7XnP8xfXDlb8orHX3hxaZsYggj0ffxZu+wF
lqmfp0rf7OZTAxRB9UDXfMmCjEEn2SSPf4YB5hd5tDnai7WEb12ManuuuaL5wBjmVQtG7NhdKlWv
/m2KlMUMke/Srdi9NV5owmnftEjrKCYTDhdHbhqVk0hy1+eCH97rx0B1viXVPYpIfosqlIAKyuC1
4F4M0K1rl0PAi/DHNMeEhdOpiA1Jzn3VefOj3zrsE/wTnePQz+tvny7+EojgUQ0C93ycXC/ex3xj
yeGK0KPx/ZRRnYhi0WmjgzmDd3nfZarTsgMWEpjs3tKGnmuzgVIqqtp67suKYp194S/syxHm0z1b
L755VWhQISAQOdYpzHbf6YUKN030nhY98Hlsz7GTuEEc+5IJlclQGE062P3T26XAvcoC4EpiGkBy
KtfIM3egvEHcjk+ld1p2GXwF4tXNU/Dib5WX+I01/EJmjEY5gTqlR+wqLq90y+aV5WZW5mB9duvx
A4lS8LlOwieQHsMCmQqMHInIRqcUb79i2Vhb3Bq0+5EQoo9FQ23tT8YYdqpNxCdfN4lZkr4rGLx1
j0MgPPXd5D7to2clkVs5XxumT7gMibfMMwE/1F5sydR/NlzCtp6Kje3J5LYGO+0TpSOJWVMHXiyX
FDeT6bq4ASoJY1FCsehS4I9fUNvG5YH5jNa+OuxgTxhu5879P1Zbg+hN4WekQLY+fXiAOTZ1LCZ0
eYqjBmwp/+rtiHkHrsBpNY73NXtv+CloO9DdFReE6U2hyXewKpmA1VfsUUvx+XOb3gCHHGgEsy1s
1hhVYPxMS/zWnI2x3r0kG5Frpp6+bQ5db87i9zUsU0dGYaL/IZOV3vFkgpSqVGn/xv3ck5XVS8RC
q1bYzROPRPWoGmHbx6hbRy1AbXh5Clk842iPO1OmPeTC8im7V6O7pB/M/00uS7s8gFGBPd1yXOYH
puKMSyWBa0FCiyaHNarkmMyQ1TWpubO3WNWoXCZGPRwU2zqgwcAoNC6mSiqiqMbvXsYFpo6FPKD5
tJHkmxeWyEU0gpRgVNLzBWumHTx08rOHpWTVr5fOFRmPFjf+LIiBUGYLcoXniAdJCM1oq0Yi1WD6
xcOunyhJJqFPBjt2/dfMMExbS/SVXWeOGtzyvUfvh00WChuSUJ9w/NlZSTAzVH1qoraPDi9BuXsT
eD7nksPAmrxNHPeUs5DCHfh5yz2Izi4uNZJWN6QLzOH6h2n1h1pq4yLxYpNEpAUKZL7mcX3uBvit
78GwJC18CaaO3GgyfNfUd32oLy+7hzrW5sAhvteoKar0cdqUctLPYgYXt20ICsHpg7P20YgSV0XV
5QCkct1uHDpp1sSwzJ2rEHez20k0FvLXEdlgUlPypdgqLSOFQB+iHjrXciSjTAj6mR0sE5dk1Jes
JksyOP/THEu6laRKP6VVVKeBIo4FDL1WXDUUFAwO4LYVokHs8Rujin2yNuIesSRxG1JvnA9QITQs
sdhAX+WG0C9FDLbsYbPrWNXWknQrqMNwy+PcYH0IZ5BVp63jXoMBOAqBNT6ZDNLfYC6A9NLr3RGN
/krwwhvq+ZraMklbCgbm/lot7TC/nD0SefeStwgLjO5fexxUfgB5tSinN4kVSs4b41rBxmc9/0Qt
UJHYTgwJdX0f+JLorV6a2SizVBKyp+lg4XZ3fZz+RE1BQ/bt0mjA/UbRzryzRtKNIVQSjVRq1FBS
qfA1mLosmSMs5POyhsDkHj7XZje68dtUWt+zC2puB6JNx4Sue9xVVC2O/1kEVvTPUGxq31KteTFV
Kv7BrLOmJ9Km/iHpi3X2xIXJIAd6xBC8cXNYUDXjvBIxr/NcaGdStfIaYwno8BrYN9726O/dVG5K
8/4GQZhubrQHWHAv6Kf8A2EBzjbCHvGWB0+FVwIfGks7f34RVUW0Wd1XBSDBTGptfr3O2g7zi97W
w01WkFNUaBJzZ/E3NtOgxZEBbYRU38iay8GZmC4a8qsvOVsmjTz6YwTwhcF87TjpJYqzQ7Ql4G9v
7XsUEdHncHysQIq2MxSzIOZ6D/ECyH0wRx0INmMY7xm4uYEY02ZWqM4XkpV7HH3oAAsaaHOA4v2y
AMBzLcJEN56LIRaQhXpHsf0CRWTrOViAK1Yug1gBbvzxXkg1cWLAJDPTgqEGUh6bz0DucAIFH7Kc
MM1W+XSNyYO+WIP6Kr90md+i9vu0t6I/l7Sbv55lJe0ivEmDmRPzM8K5caHwy5n7WAOUyGnrxnov
GqmFw/MLqALu7tPYGvtAoBrJH/xgZP7dWO5BUhYq+tWJD7Bv4IGUkJEotwBEuY0BkqK+zGmBv5xp
E0k9csHwA48mWjYZc8beNjSjrs4txCzHUWxnBTVSkTeaymMC5MvZcsn9Ldt9UAPniubfox6cJtP2
QoJmth1Fd54/tIhBumvWD10coaY2mfS6mHU+G70AGDJZR1+WY1KZZT9RuuFL0NPBPMK18my7k+yz
mpMYoJbbVvSn0nE9id7akyjO+u7Ntbp5LXYZcfD6NmNr5jtwi/1x2A9U3/C4+gY6Cy0fr42g517U
cwQ7+2y3p1BmnT379fZmNV+5bZ1hCkNchusAVVu1ZFl/mgXtvao0F8g+5EzijS2SKHchT0nwH9Zd
lHP6Wgkbdsl2+sD7I5/4SLoO8RvJi8aB/cVYSfOI5TBAEZ/vA6x0JNof7EHYTbCCnpmfBfq0XLLi
bPUz3r2AzVkrzA2aCQk648V/LS2FfCheVl5lNW7e6iIcH9B3uxZwfrKNFjZ/RrnHE4PVVjndJiJm
GoIKekH1FA4UIoMZ5w9m3xSO28jbCQRR6Y6z9qUXlq5uMiVV8wpzd0IXYtrB9koUo9yv2A5uO2/s
OMSJYaS8pgxF5RIBhI7+CLBTSaXmCmAXQV9m66l6WpRnsAYdQCQPMAmS7JoduJHc2D9qz644f61n
1uLCftsTMHd1LKbVIkv9gksfPooSWcB0H5QMRPEZ3hy2vzP+SZGl+Xhx7xsUSuYi60XyNTVfvYsp
4BHzeqDhSxyitqUFi+J+BxadJyPGcW30PULbwze3BGZghcU5vwWgpJxw5KxY/3+cvJqMC0GWkLlO
4UREnf1aO3jEm+oNJxTdyT8Y5rS1EUYfA1DuGsG6tvIZE62C13TeS8NrKohlGFk/MA1K55EFJACZ
jypciNigGK9u4nCTzXolZxoPTm9mQBd8cSmE9CwduH0sac9HlV/fAVoyhsLMhznO7ty9CPQ2YCbs
2BL19V7GAVKz1BL2KEqw9uWtzHjQ3+JPKpEuTd+o+EZmMVIx7xjcaEqbXEZd3rAw2aPthBbt1eEC
WdQsi+ze5lqCZ+P/QFbBaJyKGfhTWAVi1GQ55LxEk2oX0X6DDsh8++I71WkHTzazqbPim6UChyxi
hGGTrSCtslvVHP2UvaAWhsSvNk/IwHfe5GOW8nurennUZDvj+xvWEvouVAIZ6h6+7SQRfxALLgM4
lHr/Te0/Z8gVDQCalVcj3vAmjqFEWsU829t61rLt8E4JdyRTsyzBgAIf3IAP2j5QqdgZfr+LZI4+
2ZLZE84thp7mrespr/V2euAfjTY80i9RIC03NYHtnqALp4n5Ia2DyNvAkOsz9abL6IpGd7OVz35W
kFfxRot3A40EH4T+wx6nPK+GBqFv56eIg5RaA9hfdf6+6AGDPSDJAoroMfaKEi8heL2ux9ZPSUrP
AQLizpogJZgmZT8W/X3RjvFMTLyO79jUYkUU0ZZD/pW6/70mvMkEk2gRzMiqUQKc1SrL5i4egMKY
3kQxgnCTfJCRxDGSwVJIFqMxHmsAr3eMk4xID5TiK6KvH0pbFj0Ttx8eblPulj+2iZqUp5GUOyhL
fteyBC6AFmcE6YpRemA/00Vq1f5eZ7Hgri6TfzxPlmz6FnfdcyRpQxoVcJdlstnNqrkNisaG8Nh3
TOiybIHWJwuKMTMQoF52OYFQTuA31DnMG9LE7Mx4Gqunf0ZaXi6uM+OtzQdyclKvi90pkJak6z3w
PzwDzKrLlWM3cLn4ngQxzQb+erGwvsfscs/kjAxwzYxk9+p6FfiLzm1APTC1DcoKSa2JolbsUEtm
EtAn1+BWPHX7FsZmp45U8jZRuc/CMdIGIY/LHHJRa28VyV4d3x1Vuy7hoV5tfI55Y7UtTlwJUIub
e7PABBSBdzI4HJCFmqSzuE58gvJuN5VbrGhIxRkiw7cd9xqp31khhYP3N1xzmT7amv2bNKCtzABN
c7cbLOLoO+y060wptpq7G17BXpXS340GWvJM21g0k+EQL6tMOkf3UiTgAg0gdkvaajGGPM4Jp3sB
4bWw37b3szZwDZcXHF633zQ5dcKa1tUHzgycr9z7UsUzP5ZmjjVCR2gRpxmUkv+gVaRqo/2DN46f
SgxP4X7offosuiz3/eTKj5DvJXazJIBapzfYj3FhQEo8eOt0gihdLJ999Q8xuMzPaVGOyRB9QcjE
9c2/Vw6AN4Uxo661PKfoK9EcUpIquDzB7FvngQCHkTDjyNSWUH3B6sWZBU2WEFlcvU6WqrwDj/yE
i8iWUJ3ca6je4nTrjnUVNOJkZDax3xOiRmKRP7JFgHCOq4lXnYUGMmb3tUZqvu91iTykgx7s7ng1
5LL7zQON08ki4LD6Q3D4IS7t/pzH0oBRS/csoUBr6tKCk6FPmDF7JP/m++kkV2rijNhGia6nOkjy
JfkMXX7IZjf9l0a13qCRKYyDY2lSKsP6YNET33CkHCZFSi4xE4jgjD26E9nFcmctjuo391iTX6vJ
bK66xRkbJeDshHncGRT3sGhZTDoRmWGZlcoNjSXKyTzBUwpwzgG66u07vN8h6iVqkZx4BEwV0TZ8
0kPQIPdPRdaKU3I+Wth0wLvNJ5+V6vC2Jbg9bzFcxOCM5lhD68FXEuCdBIMldIvT8iIAHFgAazRW
rxeHzN28G2lpkGAnoQu+JW1/mQ/Nj2PGrvQP2XisrBiqGrzG1K0ZnerQY5+GXRVZZ1B+ldCkrYtk
IpVK0zOA2KBfGsvpvJEzsuMT/tYMcr7OP0oEFUxFUrglFInjsCyHBQhx3URAPBUXgCHQh+MQ6UVo
V+CQz1e0RAk6VRB9j/F32ti17r8YxNze4pU/bqXwSk0satN6S07s21oUWcp9sVM3gJZ7bI6EPmt4
wlGzoMzCzGS7tCVgaiD8lBQBcVK7PdnD1YvchyCL10dRkqsKa/sJxa45udj7WlYj1t3tiTCbZm3H
q7lfPCfUNPymENN1JFZjZc5BIbIRTFSkyCgb/q8UvQPeJS1+VORaoHAzjhxM72G3QJeQ1F+tifYY
/vGqZhaW03wLdBkmVqi3EYSttvgWZKFvMElbRu1E6XLQmI1Je/Kyoaz9Ms1udWv1vPslhkNtIHwa
eDMY+CfTFW8yvXKK8a4I0L4XXsE+EzLUmuqWnMU1oOvUGN3iTOFVSuKpN+f8THk8+ps2VNclGJj7
1dupdDTNKIZSiVyRIdgAJorCjdd0mFHXh4sKJbNh1A28xGiNvBJ1fIu8C0/rY64gqg+7hh2XOfnq
E4Ru+RF7TX8YQHZcTGID5krzm0AuWYwh7sHW8k9q+6KPrqKc8jVebP70/Hcn25bpbujgRytNzfQv
XphGsgD9m2JcO4hKtJf2eSsjNQ1q+M/4NegcScEyoCt6AfUUYW+8KWFmwVE0kmRZ9Zcdf6vY7gZV
rYgyAzAS/50p2VpVHujN2hiOCoB9WJ0wxCn9wNz21ImSEn5oAFY49aNCKDgxYMhcrLuYIT62Cqef
nk6VgaZTOKpJSdRrzbbgDr47s5JHMMN1WLP42XXBPi2CxhZTcBpbYozDGEHmhR3Z/MWJ4nxdEB9h
QvIkNCn6uPT10d+YfJgS9sxZ0v5d8hQckRwfJTeNJp/qA4erkhL2Z/2skD5mYCPfflQraBdNKofA
R7t7GigEAXiaxOWkwd6t9FI3ZsygCutNqTy86nHMNPOWrvgJl1S5dByQcIHbbloVdE1GZG9cr4nS
JW9euIWrthzWkkFhLptxMjxXK/KvZ0HOz/b9Tdt1MMK5AJw4UGXgn3KjgANAVImOUOr60vT+7dNn
CmIm1nsb8D/ANM2rm1oAG9nmzgnG1+/Q5MZGpN9bkE7c0JbPR2z6HbRxaiYncAziWNiK3fiRuudz
QuqK0nN1jdtV9QWvbt1kE0RV5EqmreoRjKmAuwMtQwLxQgevXCpaWpiAdgZTNYjep8bzb2cdf3vS
Oz6WXNa9+lBLpOofwrr9h6drGOI6BOukl01ZE6wL/QajfK4TGgQaSTsaDqNoegw+R0KtGkQV+L/K
uowCvuvd9c4018gN4ql0eP51icb8XErKEWdPsdaA/ejOoOVV5q2yPW6OFROtPBfwR+SBjPXEJP5H
S5PlJGq5STkYL0rClcB1sHBBT5C7QuYmB+2+rE028Y/rNv4u1VSZf24xoUJBBB7mvwFGiV3DnPci
7e+ctlBipx4gVdDzcTvRpuddfqQOLUaCwVERsXBmj69jzofSHTbahzV7VK7uIK0nyBR/PZX3J1fX
5PZuvy7FT3jGeMRqjeHqFRUNanaujMjbBGfbC871HXahCUcKgd+poMYSkqF/vjTxqShN3es+HR5g
B52x/zeCCQQ+yBQRSt2oqapbUfxYaYqRblUzC/laojs+nqu6psjkzgUwj7FxQ9ByaJ7rnBnY0Oje
pKQfG44rH0MjsnikXcm34PyUWZ2YXOwhFle3rDDksEDwxOhPMJ+4ABeVBUBiqEJ2ZUFdEEWz+jHN
eu2mALjnD2lR9ml8BtK++opVlM/UsTNoghhtcDk3XJqlpLnpCifIv3FSP9E2K8VQ6W/lUHY0KkGv
GaBpI086UVQLcoYt6X3+mTIP796WI+FnClTPiilvViGhsnYsN4O2LjgwsZVxFTb/b6XEmN9cEjEL
U7VI/nEt5514BeLAqKEv2XeK0DN+lrrxCkwXef7AKVOd8qZnvnv5iaFjvPLaH7+YtteZJFf+OLMi
+OEpYOEnUcALe1BgT3GTOHsavZ/9LtT5XjJTQKdQYwXTGJ17bZDl365sMPm62ePTVL8taJB7xzYq
id3HXn2f7sTxgNC6/+Q9fUzaaeLsweK/MY9xtBgABshKvJmMpIP77FQIyUN0pZD6OtpbcicQAMfs
1kGdc44FdZYpkDLEtI1AF+YxnPGdXxFBuPNruedCd/bU9NmlSs4kdb09QP7gHszrPqlkkmy9mI7l
jOWzeb5jqOwgVSMnaLej2o3iTya2qKOaRFFW85bNMp2On0MfNKsFe4XfSoU5NEJEEp9NrdrR8L/2
YnungdISXYTELZdjHkjagmtmXd+j+DvOEjP+ZWAZjyZTG47Oy2qZQ8lBf7mTThobrweR0dtmO82V
Zz6vnKYx9GuY4GaH5CBPQIVMxbn24vjJ8QKi9DhB0uxXKEIqE9IzY4dxvU4qc7YT4+IGSJKkvNNK
gGWbF36h8UTX312igkMYC/c+85CkFt5Q+KB06H+7HQbJ2cA9T5Uvj0ZLpv02eiOkUiHILhQO1bZq
4fNzXm34Lj2BGlm0DTiXPsAO+PPViqS0WMJvqgrvdfbbzKJWyoLWkeo7TS+OC39vt+RSlKah84tY
vkzd6OKhDL7uh7at86sslrL+P7fyvDZcoED3eNMrsgljSThjzql6DcGZl6MfvFERnSMosf12y3lo
7uMe+iNe2SWUqz7LdgLHhFhTiiqHCtkodRVzkl5OfU24Y/WsvBv9UCUXAz/xcvMo3Xw1Lxdv0GBB
cJz2MUI+7yAHhivpfp+PMpzb8rf3O1/LKe/M0C4xQ2FaSepuLE141LbGF8uhLzr524q//WUN9pI8
yfniI5VcfIqHFUq9fSBs6M4rgKFtKMAPFXekjLnuu4rx+PcdvApJA5ovOgGTzPdLesZc6fIdCKXt
TxZ17soFIMU5eC3yxRF37Cay80OCAT6lxXtCw2Ch62+dzK2EGsfvMi5rieBI5dR41tkEnF6G9ErJ
/bSpFKXVZA7iT1OPH+CelbQac4CIC2w3RGxVfEw2SvPuOjTiei1V1IbjcH9+syiBqY0Rm9YnlQTL
CP+0VmdfWnHdzz6xtUU0+0cnmFAlcfPT8X9nW6uitPQ+GSkngGl6D1m3+sAZ8T9GgZUUp/JfI8ls
7mZlGV2A2XeYY0LnvFKUvA+agnxhxwnpYC4hFRGpbiFazVf7EAKWS6PQxON8DgUupP43CFTDMxa2
T3MW32BAS1weuXOqj9i5AKw78tAkLjXF9YX5VKrVyg59Wjnmqp4wmvOOMWkNnI8BWHvV6nPqxece
WdqYizANewM/9C5hx+SXiDnAA277Tr1s9fNSGox+yQ8JY9lbsIz6/fKhk8LGdDF4K6hNgQA+50rX
grjR23JinzJPfPnkRtzooItcNsDfnOZhfZ6QDILPpy/RKYZ3vSy6MqP834nbnyBXfSzCLqnIWbBk
IcB5fiDNb1gWHqXp6zRDGjkYevarh9oPMxUk+bf3rw3BOnTO6ECMGxnCm5f3AexGcSanu11uwV5C
YRckUhFnMOKOt95Se3K3hPf+ZUBJ/KewWqAIMHKy4756NEAWwutySrgYf+ZLz+AMVUeqi8Efe0Xx
Xid3w8yIsOJ33Q7MsRZ4hklOxxA0Na2mNMR6dyAEcIro+Oae8aX7Ut1+RDmdVRWiCGFGFHjbinAA
yYNHqWGYi2Zeu2SQib2q5NXzxanWR1EDxNOqY1GQPhrsYIEdxd1Nzflala24zguALoAUCSR8T5Cn
rIUxfXMscUftPLOPMzr3DbrCZNlrjTWLbQX+1mjBZq0EBtWGQW9/XYCCOp6+Wcb2hBzE72qucard
kSVEzdG/mfFhdle85ELu8fq40HNLbr0O5tTJPDz+GtNtBeLk9nsU1XMLBu3opd4cNPv/gUnhv7W8
mQDPpd7lbLpInAhJZGcnvXUWLLY2O5Ov3Net9fLdX/cbIAJrj1qp+LAuuqAZgcnlEQQ0i6fO+7i0
AembqbrcBvmjZiYgLlDQN8PlyMFDOAGhStBqYOzBRq9cw6er6P4l/0ifrVfe91Lght9+/FFWuvDY
Ur5FIFNWV1aSWetLPR47pSgSuzPWKO+Q7iH5myBZWHffhQCo9SILjbqtgQj3KgcsDMzvpmtyWnlf
CooaKNkCXKmM/Bp4mT/onVt4FBJtElrX3dxZzDF4K8ShQ6E15umKiHcXdxzy2bqqhGQVPEs1uV5i
itkRXLQ6wBpDNDkD2m6/TEH7inixlXROoclXxAEi/YGRl3Kxewg6edulHmB+NnMgPoNuRCc1hlku
VYy+lTnPxAQZj/Xi8211xd5zhddNzHE++74wfRc/zBqziOEq33pkcEdXc9IFzhjN8ebIPW+N/dae
9c23NEyUItUliU5Ohr6xm7QmklCOoTAKGP/OM3to6+Mcfk8TllWBxL9Mso2pA2ECyoGVOZ1abdGQ
+PAQJEFneRGH9PEsvLNJ8pwhvK6XIKQlXgXfXJ2OYeY+qWrcoCE3w5cBDMvcBcLpnsjv5e/s3wuq
JxJWwyStnXUuXGVzVW41U/ELmrkGGJxEAgffs3vNLGiS2yH+sitOd8rY54Sv+Hx64rfcznMD35a/
FA5qrjPviikzvyqs0JiTt5XY40tIESPoE5VxmTbBdsACgeMGmpJZjhxMSePpGtdZ3W0i8KwORX8N
tyDebIfoOM7pZqHckj0BECtoTw3ioVSLIKqASCTpdGNAuVc72RazSOfvkocl4QgU+6/tv0TmpG7N
+C/JWtKjXmS4mzaUOetnHcAx/vumkp80nyZLh1rnsniqB5dKJ5+AXRdKKh7cre9rxACfvUEtUiNx
HKAvGRL299rmBzTpE7j2pMvzsE+/ZY3cDX1A9U6rtc4RqK3MGsGc721hAN7yopSt3llwaBxv6uuf
iiK6TcTe/C8kykgVvtS0xe0Bq1C73yH/fd+bJXbWvkTXTQUCJAT/lfFtCVUVQk81ZuuFLmLT+ow6
ygY4Yb64XyH2Ea0t8lrliXm7oi54GRpixJZ9lyZy0I851T7eQzZIm0nKbLEHqN8u5eT95CHb2SwO
tI1Ti0mn8UwabXHpP8FUw1zniIu3N7toxiYEcM9rq9MCUor6+pdOIWuvnCwlrWclqXFXX2DUBwan
BJwUWKsaOuZRAkygL5BY3h5uUJMe1ta1D6GV5bUibianutpzx0heIfLx31b3bMoPs1BhbStBqvJP
dpMz5g20+YqUDJufNAxaPMq48F+EjuX6zQ1z2tQ+/d/2WKy7IpbM8ziYHTd73R1I6BVCIj/b4CtG
LtOXeRpPX+5BJGIi4nmme8szy5wPD+J5ip0VJmmV023Zdduf9rxIKFJ0LLnr5TC9vbPOKm4SbQ/l
WVmd0I6Yaghm90jE/nJ+mytxowEsPYIRzHU+lXzAdCcUAstPv0VqXTO7lPXDg/FMwMg4C9TfCu8w
8ZzhxGd4/ywM+cKqfMQwq7r9+WDC/su7n0jNWDRESebIcdFt31SBo3lQYMvfbE8UtsK5mFUSYeMi
+RvnzfuvA8TNafVrvTyzdtn1pVDL5J5dNJ+Ts3D5C7vliNxnK8Ld640KqZfqKgQv1FZUGU4nYi7f
jKFC5FvjIPM2k5TPhhQ8Ht8RN+CDUwdU9xcSCiw1xm/3TgkaJPKpo4stIQeoq2ogwyU65w1M6djO
H6HfhvJkhuIFHIbCYdrdzlk5E+EyGWbxXeAmo9Ego5etXGZdt2R+azb2ETSwjZIn8K1k78+IrA3j
KpitUDQq01j45kWSnGmeQz1IAMPeSLENTLUJYECp7R/G1M64f899dFJ++XEnTCTvtBCqvup7owdC
rZzcJvFxTsPJWoYAvdlfeVX4CmgK2frUs4ipYzEONI0FO9c6TiyV7rbXeLIKsX+Hau49YCHdoCao
tvwQF+Nf4FiUcPoANV7jZZEOdBKgFpGQJvOaytWqUbtJPijCNsnSPy0d6zSxk2UDoMceRyG7RLWY
NjAXdReHLujU9CewmJcdTu568eW+21nNAB78H2zRUI43HXxa7VcrHbrusAR5Y17GTMYp1/X8aosT
GiJugfDj09H50jGZLo9NcPvFqyvnNuNOY1TGr4vro4JIBhqRXApmR6kayh8D6bfMU9GjV3gTzLyV
vVHUyltvi8ExBpTKjztusDuL72zANUHiKqZZB3SsPoMqzw7A0drL3s+jxIEUJ2yt1RPbHlDE/jBX
Q4ZL3g/xkQfqVRp4HlHSHKmVtQmF26Wd0/WzyvEh+HKscNP9W0JHzA1yOmTZS2uu28dT+nQbeEjW
zT8MXUIqZQuwZwnlxvYeFGtQSQ/6G//SGILBiCCpodIcSK+UKsm3fGzQiA62SO30kFHVuonnH0P+
X+iXlpEvPTcNQnqDVSIMIh+LRXP/yp4a6WVR5+DfFacG4mEYVeSCSMzLPqtq4805C2Ue5B5DbqlC
Yd3HyShpA7CiLd/gi6omd88GXIJTsOeT5FyND4NWUMVBko2uC/Y5ooxhNL2YBPbYoj0EeuzkMadi
E1YuLO7hbvWwdvZjgWwLnwJ6o2pm2/ou2AfWJSG42yLjQ4mwi5VEaEctPQHCfh58xGKUHh9GuktP
6NLLuKmWtBWY1b7XLLhuEwGmARkkVDZGdsdYf9xXpDPzEOp57zSqRG6gM3WgMaeI5k3gfl8kJ45E
H92p6G8tAk1ctxD3vuXdeqnOzuDCQRuiSPTebz4UQqOz6ADF229uNJNVl9exxDyzKaDrTW3BECjH
B0K182z3CwQrbLCdfR60SPC9GIkuqpAL/OYDBy3XlSRxXl8mbGjrwXxgnD9eo92Wgy11vC91UL1s
L2Kl2WjQy4xwVXIT716+51qlHXIk3ICk9G9v3D6LOcRGJu3w6N0OBMIeITEimxiPQDZ0l14G/V4D
u0QxMSZZsSSyzJbfMu+LOl89Jqir6G4MmGtqZq+JR4pf2M47Q6qItztfZBiiv6eyKNnvMLSjyQjy
p8SswX2l34I8qVtO97H5660VWxZmTBYo4fnsxBjNyVOyn7sSJGb6VD+SUuEaE7KYMw53b0qzZxGC
u//n68sOQ7SNzWiIODbge7IUF75ZKDJa+/3EeHcyz309C6mEnX8XNDgSgbGX+CgKNazTJ6naMsyU
cRDemzRgJ7uk+7QCwK7o0Pvyy5DPqlirDoscoGkvSqMbmDghrRMeewuRdck0hkyXzFjJL3kVsnu5
tScfq5RiuwdZigG7fx2cZ5GMzqJC+pOF2I6EUK8zGAYFFGTXCN2hU/qGAUvG3/EiGECtR+AUa9rB
1016Bsisu22nKjIh9KdmAxFoip5ExH8kBfbfHXAAcpsI5yGJnc7Gi273PGop2rg675Pmf+TrkEzK
ydfk0qNH/LLBCZBS8YieTuKyWBUDqXBoWaug5ME8TdGbskbw0SfBQW98xGHL13k2LhlfXL8gu5Lb
jdoNFQnD3UQHJYoPMU1G2hVYXRs77jByOiJqQlPX4Ghw8JooXMW+VGG4Iusb7warHU+wGdEo4zF7
C3l9pgocfghEOsGKbl4sGDdCo2cNQNVE2fYqV3B0D8lYEi5bFh+E1H7nA9YxqEKFKwdlOOPFM2Zx
d0yCBA6QhVuXiQPzO3Q5SQ6AYC9yTkX6+v0aStqQlwyDRL0CRj/W42A34BHm7vnVSmSH5PH/oqxL
rrVOHRQ6YHNu4ApEAcKhSlLtc16HFnuun8Zf5FmaZrg6L4/47hb/tYlHMTjnWI/1H59SQ6faf5aU
U4pvyvFAaE+9glVmlXKJekdD1WEqOSLZvtYvUNyC22XWBhE66jkyVWlTesHAfo6rIDcyXOF4V214
j9p4FoNk8aHUrQYamnVXiWM9GfYuSzzNe2tlI4vquI1oa50ByciFotIEbKzQhpqg8+Q3zFYMvpYO
yryfburoLq3hBtq3HnmmA5AfNWkrP+vclm1Z8Ru6XNoQaL18z5oL3CDlaRWPkvVXHNqR4DZhhl4/
bpG866J2qch4F82CeYwLnqK/vumfvyItOxUMV/sgkdVC2KyTLnKi07PqSDS1Du4TbZ366EblrG52
m/lMrFxHWQGn5Kjycn/q6pt3+sB+q3noly58gZFCNc+c6Rscr3YBV710MiJemwO6xOAtAd//gLVj
CzOR7E+o7FeWco0oxkLbregXAC7bB2fxHowd+2GNfab1tkRwAuO1+BPR2gh6sFGZNXr2Fan5JS7D
pQMGnBRTEeKyaDVjz/gXkpJH1QEpEMTmkHR8Z3IoTGahkqj3kWP1eqSBEnZw9wJg76sLkROM0SpW
5LgqMMY0WO6GqkKskIuFCk+4PXs8B7aLVD6EMLGYl5Ls7HRfswvhNMshBOintX4LRfzbg9qVRt2V
SSSfPnQUk3loS1sCR+gJd/60AqAc/GnEiEmc0Cp3hSx8n6BID/6QU+t1Ql7Hw2AlvWin/HKRCQBu
KMe6KAfcgflqJ+veRqMmCleb6jBRwu3tFKyqEyEABlO3fFQbOUyb7Gt38sx4/WCIl2+qo5WhzmWD
90ruIoEG2Mvb4fGgssspoSj4ho6GkMZIL24wQl7CjcTVgnbO+xPXHhkcvuqfq87rwvgnS1CzkyqV
gRAy1n15b2yFF39UDvmds6obN/V72OC44xSfI5w+uVJQyhXIe3a5dypsiSQy6qeNY2jdcrYYViQr
PQZhQ+p6HYbxqW5aq1Cz93ix8JDd9wbSzEJza0dA8bLQFqpSlKSBky/vpa4ENqaC+nNkB1B2rGmR
KaolfSp+he+xl4bQBQox7qDhBEgG0GTip6nv/YGRBpeG/QjfrZ1W+E9iBGvcj4UrED+WK+TA84BU
WvZfMb90de7CmrYabXEpcpoHOcz4VGRdR+3Jkc86UASdpRK8abqxoj1U7vzcWknNbOlLSFv9E+tN
WEgybgS+zuLvFrEQc+IBjz0XbRJwX4oRSBCsjsT4uwah4UZDhZBm3JmUKm6Xxl7TDafUkpq4CBat
FJlu5JCtgjanR9pPSbNTP3uhKLAtgythFwv08BnFUlN3pRGHDcTC6jhblkWUsGqwn8WQo96Gfh5y
r/Q6OJ/oiL77x4frWYBmxX3tp2rD9p/x7GBRwyDpCoPLuplwORfAYMgW3aYhhwSNgmR2WTIbYU0M
7GeMrbNosVa/cs16GaDd5qLmGSqCUxB85fDgyD/y4bsFrpUiJXLn2Yh+AWr1gcONFLUH08cq7FTY
Ki1IpwCs+yoSYd62/CAl5snhK7BJhI1VUrcvJmxtiedjUM4uwib3u+Uf19+UpXfanA1qVseebTqQ
MsjXD2U+gpKF/bMt2KiAzsZkqUY2z0x2F2w5ZQNe2rZltgKtqwQHNt/UoJh3i1XIBIKi1swfIaZ+
gk1hHpGKGtHBlx2gNxnNJewnbKZezyHm/QWCfkM3Du/xi7lpsZovAF31+hgPncO3GyZgUYYVYxAB
aDC1bBxIDhqGADCkuf07uFM4slwwYlvtNNhAE3lH/mObIQLbZNTqg4lVdkEL7OADbUC8lx4mP4eC
EdXwC1h6rGFosWSpPRYopHWk6mt9SavwQYMACeAYHxjKlxqCuy884RnrrQ9FNJc8K+INe5z7hwvB
zLW0Eg76eLS2nmlvcLazHQBkf88luSOLchkIHsK0hIkv+rBHWNJtq4Oy89nIK4e1x+8HsarSKMth
QorKkhvFHi8R8A0tgK4T6zwbdf9T/FOuuqo09uluwjrLA85OID4QOQvjo6P5L2SpCeYEEvN58F4i
Kl8oTzpZBKRKixuhynSelri6N+ef5QAxNu7YAU/xYD/2N/Ltmc7Lq/nXjATM73sB9kId1ZtHL+fZ
32gycHc4aY0fENgZwq5z5VT8Ep7HmMalA4rpPQZwtrMY/Erhv0h0Ysofmg45CbgwimvJ6wM0z2Mw
s7hNNq4giY8okjWtJ2UhVQoRRHlzJIyFhnK0qUuGyjPuTGPTcp/IygYlFb6Q4xS9huv2tFovJlwe
3gOl10mfdVCDCdAzBnGERTRoqHlXQE2lexjXSipb7pSYLPBUdedz0p5xxE2JDlnD6IRP1V+A2Obp
NrDdq29fW7xpRGb5Pd6hhufmwwc04Kmno9FBk9g8HoSNWTnOtdpiLmAjyt6v6Kio1dPbf3J75XyA
2EQbd60yqbEvDOroavQ+CRSNfMSgqARaHm4II1sjoSuO60hEayUkiORIQLFqusPu8EOg26bXUQGi
c+emwxgpEK9MYcLrnqAyIynU5Nqrly68q5d+H6tWE9y3oKDfVEzecIwlc/uOHAOdQxk/U3tmlNmt
OFr0wEHbIJrzgWNQ+dGc2aAaWmGvn0SGLMfGlz5RDCSjot2TYVUUAvjlMXUbyMiHp2XdDcNKyjAM
sjc4bBQ6woKCaFy5TjuDke6lhEVc/LU/rPNiZPygxVlGXCOr4A5q1wvWTAgzRgcKctA7zhN4pRd9
7QnJa/X872PrBczJdCLbd88LHc63qA9ju/7PljPzseaZmrn6Mme8/iOxSucFmvRzeLfQ/eGOL7rg
micEmTJrxPbwOOp3oulQJx9UzAm0fLDkCeoY+1B5YYLiKPYXLmBPrAKU4U29fCWdBJCfO6KjNFpC
+qsDzQ4Xjy9Ck/tsruS2FqlW2MIZGgJ10c2fOlk8WG/IOR2BlpGUh1iCE7Nq6Z680yd6cTdZjlii
Y+AyPBZ9NmEQppB1vs7oImghDWctlAcVdtNtC4NYRObr8tUsvgunxfGIb0T0ZMLzsOuBTyAdGaBD
U4iSLejUCfkSCynf1PNr1v4dq6RrlcJrqpQv3FKQFGE481GhBSGzip3fL25w4sTKfGilmJ4o1KmD
4gy4atrzlfBzVmAlTsn1DbqqANP/+7ehyU3rjaC2kp5O2VMp+w9kSAEwKEbDb/1hnQQo21iHO8ZO
XoO+XKZ4Any609GVnpNGL2+OYG5ajn/NNb2AHxW4sv0WxCeaGN0xEhtnD0HTrmk/2ZP3F5FpmWYS
aSNnzY8IpKpDbe6BEgwGIPkKMoMu76uOOfPImyS89SosbT5zdE3l4afso4dapNlAsVbRh+vAJztn
FQMpnGkKiFAA75EGyq5DSvrCO9MHCnGqxvaeLo/Go9usAa3Wjl9RBd1f5JuAePogRbaD9rF2Ij5U
vMVyKEBgXBaKjVx0cElDQ3RkbW3eKQ2E/DxAJUusTafyEb8rZOLBLmLflLR/dNwHRP08O39+mVQL
q2dBzulJuMmfgdeMoXeggS8AU7cllquZJps5ALTHfmAykVp5iU9hS0hp/DvSVYJZJXpxpZZUNDZj
DS/ki3LCEPWoVyub3kMC74Ulx5epXPm160k5NDsCs9ncHsZCxXVblgVHbY5vRLEePCvUa4J/f5Pt
tUemi9vwhv5RFba2EssiBK3T/Gki8pj+jZ4BcZpcqxft/5+sKZ65GHztwVBhos9mwkEXlWBb8bZ1
jlyT8NR4QqoCp80FDSHHp+QlMMbOq4q4rzdN4fVzb33Vt+5TfUo5JtEov72MEy9c3yMZcfRzhF0t
ne/1cw9S13AEUI5oYw3GeMUD1SrqdQl07cB8CLjsYbtYl8HP2hGzSkxXz/i4SPmgc2KTLsgnFO39
iBP55d7WXRSblstPLPYjtwfphV27D84YLOCBeXEYruz40DAucFPZjvGWUp9/BdzH1CLEtcSvf5xk
GUaFmclG7+QKbuqF3IaRRtBCJ0NEBysFfjK6IEQhP6oizY17uwVlFoshxIHR0OjsF9R2Cuj7Jqg+
FMlUBA7QGXe1D/DVVHOYcNVC8OjRDGPhRdDVcJAgcLNECnZI83dKYdhUQ58FeZ+yCFKJIvJmoPdA
6UltXCY8ePDESvx9FVxQ4xvNyqdY8/unfBchKSJyC+IJo0vskugCrA7qX2qfnOZATk64rLSDnKce
cZcL1u+vrqyZz+zs2ihTgfL2vyWQilyCfzge7gs8fm1dPYe7kqedt63pTFmrj6VAgSFUybGYvi0U
r4ejffzXmUVRoKVtWyieQuhRiI5NJMlfOvRXD0NFjZhcMSIL/Wj8QNinbwzU6crVB9vndudnK6bl
GajXZLgWax/FEjpj9Be6YgKQXVlwlW2xt2VzNdvrwYKXUutpSy2Z/c1xxep052vaiRNbNVjNM+3m
474wevHzxUc7k7hnsKflLJmZML5Fs37ra111TkTu7rAIV+v4OC0bYaw3dIHcA+xk25ek0d06s9ix
IDIAAF4PiDOv3k+hYrnuDhTHNW0JZHCiEzwnPXQ9ZwBvS5rtZJJdsKiNhWpFbvsxlHFpkMZnbzih
Oz1GsTq90ub4GR6jCr2MmxfhXtWU5Oyp60mtHVHVXw1Iltt9tKf5Oe9KSKIFkFqUrkVr1kM23e/W
GijFLmvJ9ZyP9yPDw1uJVa53h7cJ63ZMgQwmWCcHxJ3P5Yq+UojLewMK24DjF9Qk2OhW+6N21IlH
qr/lVfZpdCa1OSXcgepEOfTG+bzvIM2xPvSkms7pmrwyEEE5KE20uaTIywchguT9tAEl05RPYWp7
B8CjBNrTIFZUNWiAdK59Q/VwVAV44QaUqdEU4kiH8/8kNOjcIYUhjXtEBwEkF4I1EE+DLSowQyid
XIuM1jmH18WKtUUtpFAK5ecarBJ8/O+BxkU0r9ZXwRDaAmV0/GCwxQ/P7JHuM2OkImWUhNAv11C1
7Cn4NhEF84w8kVqxbHxM+CplL7KM4Nh203t/ot5SKpiAnkUeAsHbkyQSljPFhGzIFmTiJibL0FKJ
MAXuqepvxZj9EvJnWo1Cdp6cl0tmrraGPKWoKLjPsqs6PXrbbb9t3rFnfu5ZDqyr2XFYgW/7GCfR
ZSEtV4vqCDVJi+ffXA6Dl8T7juNzLwu3GDTdXBhUHlG9Hkn92J4IK+VSExLIegAUmRD6tkO/ZXWw
sgsuWtuaUgU4q3XjmYtHIOh329tqnoONAhXSsRrOUuhSt40Arm4eZmgYTWkaPjojMxMqlKBte2XO
jtzIL3jTzQkeOi4q9/EmBKsHvyhbqcrVTjf97ku7MCShTQNo+jNXnwFX0Z26q4v8ffwP1Qe/Jvkx
QLWkuN65gz9TSsBdQRzOM+95zlcuEsnC1ASvZf2kVljgQ6LrXuqcKTkoRPAFFW407FkCDo6d+yz5
+0kwBldAzjuQJRQAsy+Ftslc2yduTxAfOFAh/+s1oa59f9yFF8WM4UEsT/hilba08+tp8rUbX9L0
xBPUKuAUVcASTYJE03+MUmCwFzGCY487IVmqpt4ACDw4TbLwctCIoHvjN5Qcd4Yz+LOAk2wyJUwK
MJ7Nf3yXkfkmjVmFbnyimWYoa8XLkS9huF6vTxNfYISEngikzRKQ/VF+bhjgHcm6fTtwj8ZqbY3N
/Ahu8FDVISUs0jAzHhcve4cElstTqUFG2UR4BxioGMVobCOL6izybon0SpiQG/hoh0gZ1Z1INOfl
y2LB1eQYM0eVfTIynjwAaKkbTLY5dB1Sfj/PDuNaFYKeuiQAr7W/JsqbWUD5LXBk39itSJAZWov/
9D4kwtiz2iQTb2uDRTE5Up0XIGIEPWFaR3RTMp3zDUqL7cBK5wda9tsxEchoy4rT4GsowgZzIuqK
c51GI7yvwn5oWvjVvlKk4qDqr3WeFh4SqnoAvhBdsmNCtVPX/7ikQG89L7Ot+y3cYNqo16jBloCT
pZZcNNEUxF736feqPZ4t5AYc5ji91N2hbOJaMN2FQaldXqnjOXrmYkuO58kameHX2vKIAK/mwyOm
7B8CXbJRbVqwWVs0SmBZCOknykL6tgdWnS2eNOGrSji44D5T15tUtXunP1G/pBqqk1u3MJ1QAgBl
ECECA7kNfqv5tRx02D8l+W4cPoswCeVPsK9Em09dOGAleT94E4wPlfe1cB9cXF2LiECBFDJs933M
LZ8RSIe4IpJVPeBYgDrHtUPbS1rqTgfXr9ZvTumBK7dnbMI05xtC3GS+PyYgAFGo1v7K6ycmKlfX
p6+LAGahYHKOXX5MgFxVjojscnVuyvS/mgnD/xxPHM+1vwBHvHvDAlxRuYcqx/KD3VPtDAk/g8LK
3e/lcBG+q4i/dTJtulzX4MEWehDy5nhNf5THYx0VcPbNectavSQF6gNtC1odoGue8JUmJcLLYFVT
Nw+hpvgJAxghZpaljh2jK0hom0CuUFOiwnityNbnS6FIH5kd8jF0ti6iSI9MdDZbF5gTt+une/KZ
N/ra1usjPnLKijteKqD/luA8tzQ0yoKTuAT7qyJP4102lwY7y+D5wA6UXTgp/JsSN4CjTjciHhgk
zmE3PR3/wzp26KDopg6oAWBQ7WUzVWbicp/+xW4c5YzoZRqtNmudHJJFuTi6If6gWf9Jk2YaUqhT
ROLkNtw07CVfEpudo4IqHG22J5Zk+kLw85uziRix4c1qQ8A4YhTy1UfxMhnWbv5uofwFNvevVynE
/RQnaA8C/ra9r+LAn8R3knQhMd06lYQOfjIvLcRrM6hj5VsJUleOYZYKaj7S2ZQE2fE2uo/g44iR
VLiAJG4IGoWOfdmIpFFlIZNqJmy4J8frrshQRSRDOwVHBItghVExhiCSMZf3IpSNDVUli8YZucNO
C4WIAR7Zdvs0boZSYZRze5R/g4zvNdeW62bJ8jssDuRt97CTCNqL6hwgee11uN0zUUHvi8Tid+g0
SDL03Xd6jW1nBdDTDZQzUpnmp15RRUTCklSo+k33m4bRbs3kjdZo5dQVAvdQR3vX6WMCqTi7Y2l6
9Zf4NnACt0DIMstZV4RMPIK0XOQkQkNHMmqo16gb7ynPxvnmEAVWKCuZX3J1arT2KMEPDGj+jhzs
bDmD1W5XHkWM9lSTC6/WFbTyHDnGxZ/x2BudAAqGTEPpKfetHOvLU9EjadSSyy6AmqRjoT2iDGj7
towACsnKMj9/tHX0y4SwBcN5sOKf0cuDGgdoOd0Yu8SHY8F0XKzLHgY5mfPqUxGoGbu0YPYwNFOo
DyvwylRH0X0wB0tokCQTOknWOXFlqzpRgqtxjV1g8LWPySXyOIas3YXufGUl19rLX8SQ9NoFeLzV
4+9VA78jMm9pJhpBwV/UC/tNWVsQTpAWAE4NZ8LyfS/18kRtZp79v44PJnXVdnn6qQp/wvqFTpFI
+K2zl4I6ranvihL5fvkGrwKoAEJmYHvLI2ffvFNEEwVMOpPOs5OdpDYDWqfjMS34Fb7no/NY3Xzm
FoGCc1pUSqU05oRlbiq3oN6qQfO3D0/PwwRyEomx93iIvG1kC0JXKPPZuDW0WFoHruAJ3+3Jp9r/
Fr4pOlpBDMLClhWnXQBaGY3Csitmdoz/UlY9EBFbU5rNVanoFyHJG8icb20oZ8AiN+zaNV9m+Txb
TlNyj/KNMoqSkcjLXtY+P1rP/jpG73mAgh/HCI6qK4L92HAskAQGEdZ0oJhX7cyvH8bar97EfZxA
qUFZqIiPwH+b/4fdj+Ahcq9gpMXAzyzR0mQFnYUBTtMYPEshnjckdJimRbtlylz5pOhAp0k4G2rC
tl1G1peXEFscsik4qGHQN0dAD86CHMw1hGlH1ZhVJ1drmtZUb4pajNagnyfRsUf07FraRPly+UIR
bHoxIDomSVesmJnv3ZW0smHEZvAbXe2M+vSME5+RlZLBN3utSfarsC/g2hBWH8FihMCQ0+yjP44F
kmEvIoOBPc+O5hM2y+7Obz8R3i4shIButDKKsO/CpeO1fKa2s9ffDkDSWJV52HIbUcyFRKMWk4mX
pXcG2BbLhcAvXqi8LQJDfZj4Hgzt8PICjf2lhx2Ts9aHJuELAfMsljEKDPy5Sdex7Nes9eVmjbKD
GnuMJ4Kr2SarHcRRnORuzAOhJV4uRTQjhWp0vjPMuhLWlAH08jtwCH/0EoOJCkC5Vp7acGh//tLO
JN/+fNdIftnTSlP+1lSRHpZofcvSdJ9NS6DT7YOlwR5yv7ZucDDkNT9nLEAh/W4PW+5gssZPbGKi
4QrI49nIl5wkQ/XNYvkjmaG+MdnQJ347nBG+uI4ZQZ8nesoC72NyUMhlIjPgPcXslZve/Kx1yBPB
SoJAUIrmOETlOuAcMFZ7SVwiMgj913u5PEgv7I4OGprNZOyZDziq+FO6dh8jDtejWGqt0qxh/OZU
gQZpTrmiVff/n0N3K8mZRynv6c4YxuVD3I/Cyxqw1Pdvmo6HHOJLmnCw3TZesXKEDVKf9IuEgzDH
PJAG0T0tErOS9JjcybTbt3KZ1C0Nj+hsYHNuK6Nbg+4LXMNYvAS8GLGMwaDQZa3I7xZpWf2iBZOB
EobSqKFxpdHv525GOPryzIJOBos6EonQJ2gExJTcNEfNGhJ6PXK6B9QE6IcdlZoPCnWhS300hOWl
MboTG81PxqN13TypEpcIioqVL6AhAw7/+4zxx0FkfuJebZSRBYxv/B7l2SJnojIaRQtEsngl5vzF
WKd0Z+0cnUrFMTy6+2LDObU/BmyiR5BAClxaJgh/b9fWDmNHUsAs+GImIyZJ0EmmTuTb6c8msOxG
tVKr9hnkMAGJfA4zxL3WPwYlWcyaBDaaojm+JFedcXeQzEYAZEuwO3FzVG+7qk3CAjHo3wZdLiLw
IF/ss2lvca+lS4B5b7wir0Zzzr9r/uvHk09t8y+QxtO4sqcj170ttV3uUFvXzCTh1fSMUbLauP/6
wxwmQ9yw5HGrJja5qO5BI9X4DVcJ1wpSLTVVYa5XL3c71do/c5nk4sT4Tl6wO3eXW3BdmAE1ntpS
/9kQFdKXZTMJQWyqy2jHUN0oJaxQ0EHQt3PNJWW44A3I4Fpu0rf6iQdGmZx3wBgzOHmWdPoYrim/
alB8ktS2NUmupdGsfykMSABzD3TtuEZ6HT4fg9RjMb8lClIy20uV2KIuSUdufBo3TuXE7PPjIFGe
WF5eVDTNITFLsnVyDYMXkk/V7I7iXl5Omxh6ujhPhRqZuCGQNnNZaf+mP+XOR3DQBRKosPQs61fE
f520Swhq8A/Y7Q349T6l4fNhPAiuPUTTB1pN6+Sr/PpkGXmtYDZ+I9lztouSIXv5BZ8or/Cq3fnS
DHmElBJRMUqGqZHd91LST/CrHMoNh2U4DIpMpzX0feoLDRqddxODKwuUvdy9d5Uii68csvcOe6a8
wzCcTMrF+mw9mOlm0IUGxRsqyqFX2fsFz2hfz0YTngE1KWdhTI1AIYyLhpBG3X08E09NpZYGXb4U
xIhH7Acaog0WDmYbn47wMg5ZUz6Q4/Op+vT8uk9gRx7XhgxrkzVkPyhAOOj4/B7klzKSWSeogqC6
mYigcwnlhAj54Adimt+4M+K+vzr6LUWiz0yv6CbbyF/q4W5nFjsM8mnDnO1oDlIKWXz7TnPwzAv5
+4YE/wpVOOaRw9F8HIWDLwaxO55P30zHdVivANIo6ny6/dEetB7P+cg1uhVEBhE19Cm2RnHg889a
Cl6ZuaSbFrvXVBjpbx7IPDgeIDi76DJjFaAfpUWVGajfXqlsiMztE/lEcUET7e86rvfg0e78304Z
lpI8NyAZpBb2dRjlJqir8dzoNZYH1te+E4Ge5VJ2nI/ryfK7ioFgHaqieqPF2QkrdQFd5sZqBq+1
guQuQQaldutWwxCF19890GqFuqDpU34IAJT5W/4h9EAzlQzvYiQkF78qkkVvlqRvR97sWS0jm7/Z
fDKQnxDKFKT4OxeEUbbxeOif5JXDEz/SjMUO1yLiy8sUgdNEAo7c6mpBfwn3YlGokFEnH3xGxCdv
SkduOMPbyUVhwFoA5GG6TgdWTdDw3jB2rnuSNhrZkmZNtxvXaWdof1by5xgCugs4WB/pIWZXpxJn
Z1pulXz0jrW/BTXpwXF2UBf1oTnGbLOb8hF+5fQKAFB/R+s967J+4avdYP032iBVBFEO7g7idvPt
9jv0cFQ6+CEITTuHbl22fsV33GxQ9fdPXh5FPs+F/v1X7WSmsA35/iCyC35V9/p5jgWJp0pkJ5Xm
Ut8OzLQ4sbpqbKUqjr64V0gXTKMMCRVqFRjF5eBqg9rMxqf8sIGi1YnEVR/R/9WniVPnvEPkK6r4
+C2h0O9+VSEXN7WH8IhVmvSUWUv2r3R0kBEydb8BX3PkB7oref5+l50cOzl/elRlze0cPmppYvpW
irKPQA9hUFGJsJQLsRMutezyFGrLE4v54Y+oegFVCmUdM3lTg88GwKbLFR63rpiZRFaCRPT5/xeN
Y2kbfzLd0HSLaMtk7nAHlUQfTYn8xSXbrc8AekIzQpsBNNJrYPdGVCP8rb0k3WuaU6L6ukvY3txV
Tqy9nVdvvix2pigEyzASH0eyzmWvQX/Z/24Z3rLgyNbPXI2NE/f9xNYIjZw/b+38k3Bif4b14bd4
osk0TPqjHXw0QNunKTJgOZW/r6znEaBk8igJruR5M5FLvtC/iZ3+AsTpyQNjbFpdYcNee5V5PO4p
vdXNI0rTRoHmA+KVVyj+VncLP7cVpspKO1AZO8mvRQWQ3oRxXX7+mTGtp8+Sa1jKxkOEHHdf9d1R
0bHKOAWxC8RzzpjMjD8mnfqUbXyYi1Ud6dn6taoXwAwUooTdiWQ7eW2KlQtQxJ8EaPCQKWkAQMr2
/SH+AEwcTdILdyWA06ONb4scnv+AMla9zvvk3pPhVuavqC+kCHHkmPKuvhoyysfr+Lp2dqW9XFel
cgBxJhsIDcrXfbEr6c8EOJ5Ta+ELg9jyqdhhhiir7+a44t7kXDazTzpa8pivusJNg+FzjqR0QWlv
N3JD8J5dvKZZasJzyuJVECuhPUh8cHVzAOZSNVVMWIBfK7/dZkWLyiSgrUxz5yQ4HQyOink7ZNsX
Pi4EY2m/1DBhRE8MmGfEbWH+CqE08IpFRQwsS0eflXazG8ePKBjH5JrXy1lYK2n8cj1m24HH79WX
oIK4TeXoDdiNUML69a7Lbbez3zRgQ97lgVSK/hqNjaYTukY8q2u7t13w1Wh60G/tY3H4WlkTDxjl
/nvTa6jh9nyFgFwHdI2iDp4fe9W4hb+2bQcBAfgU2obSR0BC/jKCl7kURUkz2Kni1DgLdPoTVJSY
uKF2nUWl7M92wS4O54hlKHjjKzcTdtFRk9OS+zDjaLasJjbKJye9JQhaFNbhs9RH7rYw2K5HwonL
TEC6ivYLQY4XivBkSF2XIzmsc7BvI1TYCVx/w3E1ngVooDyXUzcbbUEoQa5NkqIyhoEkGqviZv5i
cU16vgmqQWQWPB/sZaw1pNw34q4BHwGhiXzEUv0T78Sed17S/zx3a6njEegVVtaC7ADfgY64yJX7
YI2tlvwUhQxm4qiDiI37TyVXh3uj2IlnY547fALxiP1KmUgdaeeUMo7mCNrkk79t+N7pHd0AH9oJ
+SAyD1ZAFWNMhiqdEcJYGwSCzIo6/BvrC93sEjlZnfcfp5EmhftbQXex97ssbYrpbaMC5rQWPUYA
eGNFob3xayZ24a0vEyLs1mhSdatAaGUI0H+APNDN9C6qwib3D0gHsv6k/pR6fjB9bZZ4pz7psBr1
CdN8uZ8Rj3G9kJESC82UTJkchgIMsII3Y/bfWDPFp4frlCp6eNH4PK3/FST6zXPJsFsdGPCukwjJ
l/OrY5PK4JRRQD+hn8l5Fs6tGTjtOockga6FFU1WRQRDL8mnRQpgT7A+QwOqqZ0GTw6poXHlfCWK
6dwQHgxahJs0NepS9c83Ltg+myyKKNuHtKRJU4KMLNi3Guk3jqkdskKF4lv6RZ4M8CUG/N5yqZzs
k60SmziWxi8ftJ7V/p/yhblj8Pww8l60mpkb4ygQhrjPeUyVPu38rrnGOk/iDKuqZzCvEcuk1SNI
dFK4/PRU1jfZo5uljCMBeU47H36gJjEZVryuCq16EMwGPC2JNdIuI3X7HvVO0p48En1j8lSpdC7R
NcGF9IQUjCnt4ZHl04LnNoYHHTH3hNU398prjGDeYvNukAsHPoLZEGb2CYpOVFAPCoBDNDCdraKR
AFGm/GIpjcO6gsz6RM4dX3vYdHAmRNA8uu8h2tzBFp3O4fxO+qDeZShoIJ4daETRzUjQYNhVxd/n
bxehAzoqaWCX2RilE5uKCBdY2FvK+dO4cVTEyXzOKLzF+wGylcaQ2WCD1h6ObZfVMfEBv+2K11Ze
THIbG/1TJKvg3j3TaVWx+D/CWMDC6kjnzy1K12QNjdODLp2Tmf/JNb/4ELrdn0O/JL8ftIhDy9SE
k+3XIcPhmZ++i/WgPg+0+cyBRyctFNTYHntJv63uv7BOg3s530IGMZ4cbiqNAR46uYNx7Fhzc27N
+DACHp59k83cY8J3tUzxfSLkFDiR6UCA9bEtygCLFVSEZJ65jxPzs6oCd6pW+4f2pbzKrYn0DBkj
NuFlA4ea+fkzhJWfU1PsYNBoaztocn602EiiXpmHEfxH7ID3AjRkFROH+GLHeoc3YISEFvqQ5NM9
F1zwkh9tPVaXXMBJQ26y4WHSoHmjTYuFjT2PKw06PnFsJYnn8SINtPM8BJXPtXqECxPXwY/8t4G+
L+L3alp3985JWQqgPXPep4Kn2YudgIvB2BpEqjOfRFIB41eqkpqJErfEfD43OvdUSYxYEAw8RJRp
GdROy2MsYuIKCN4SbSPmGXnrlz1N8fGjg/jraMkhDW4Xtw7ni6sSUBYDXy1O4TsPd+4fcj19S7ZZ
bwSivdSpReo5q0WA3nOfzj/EyVuUyT4WR5h7CW/4kCIYLuWXjRz7ixSILtnG1YwMNDbjleOMILES
ewMzzOJ63mPGdZkZtrsIJTK3PyeJCUvrzyRRde5nRfwAfANx1A1ywYZxqzLLHPtKGwXWpogk2JIB
sy1Kiwq5RqBvxoSAop6Hqdrr+Y9843czfbE8A+yboPt4lR3Gfsgc3TDvtKiAmjQBiWz+LuA4j3dx
iYXIZQ4/NRuB/Xy+eSt34gjxAC2ti29XycQ3cyJ6JcA5zU+S/Fl4kuaDWLVBP8fbJ2Po72uvrkhX
uNf7a45ZPucuaLisVy4+40NU5VAhWIacYINB9vpBiCweXB1O6BRsoOrsKWpcScIvEWs+sknM66A+
Xsg1sA9I98kDY/pRQtywaquthoYefnh3wSGr1xJlF/gX2/75T34onzyMmLHPGf6ewaonAgM2IHfR
113XI7uvelGbt3vc5TWsTK42h5rMeRV1NjucbOhAHsi+w5IBg02MhJhrWTahGy/RMQx8pQAVjtW/
lTBFh/fIRH13gNNaChMOfpr4eQIY6de1a9FfqaqcLjzEMPzXJ9ijcLcqrpVPSte0uIEkpmCm0MXD
vdJ5IT6U5oWwl3TUWA292sN24miRl5Yy3JizklAfaBpL5ft4PVmAOcNaKIaq5tdHh1BKTv7m9CN1
Bu9Klb3kiQd2zt/Sno5co0OogwY470R6NgzW/xgFfXgCzM3tUgQ+uf4n0NfKEkHKxgWIIkFJtlVF
ewJ0eqy5f8/DKFKBbFhDjLNKkBVQvxnsjq8E7ea9jjZkRJp+J2E7DD8cZVy/ceFQxhVx5ZZANA/0
IHJsZKUWAg+p2t13j0jZd8MWyBg6VgpVJPJTr5SHMqi1Ya3auwh/gXt/LEQVCyK7Faetl0ByzuEF
vYMg9vw11aCbDSseiHwwUmyJQSWPsdTnGbZAbELgvcDGhQB8t+3CDJjnXBXhNEakh2QsmHIw9G8h
G+OnGIQH7R6CxWJzmrEJZld8TGQ4liXunrTQoWvKIHikRGnGJzY0TxSMjSr6gFjPnvwRP1dZYCW3
M6BNP+i3k0mCPc38Bh3Q8NFeqOCKOysryxSfb+SYwLFsz5ugkgNFMgUg1oex8Z3B4XKF+ORRueRk
VgOHKyC7w2uEFMdO7SWi0o+/Xvu0SwKaLmsvdUAFrnS5v4Pdy3XEytiULb8Z7PxeltTDQ9VvMFof
zgQ08PpHL2zQERVV0L4OXstfSJJB/0V5aaM5UI9XdUHBrBx8aeWiPn1ZqqIlqUcimoyMmu5y/OHc
wAkObqCcsHkaHfYto/cUlfm8vNqVW4PCV/WL5idOM4k8QmZueE01BLjXjVZZdbz8T1Ulu7qKHkfQ
laY2DPYmmfUkGv15bwTzqpU/z6wT1bdkBOnHSSiSzIVP+CltT96RjOjDQYy13E5NnrxO3ayDuSmZ
6B5iNpEXxqnoRMM3K4L9MYFK3Pq0mJtEFqo3ZKj9S3KHjQ3q3ePAqnTpe1nd31kCnjGxlgQw9uTN
bRdevogg4dCu9TjIqZyDwPmpkmcZCfOghGhd5I5ieMmHnhwAE9Sua3TRoB6c6l1Jj/Zl/3pIozmm
emcN/vU0vAVU8muOyU5LNgGwi6MqBQyXWImf9HDw/5xGIjqdwEgJYnspem97TC1A3OXlbBNb86YR
xbQ0VELrnzSeqPPylOo+TWED719wwQY1QAywQ33K/PmbEPDgLDT2UcTKLRTvXAATgSl6B6eK6ucX
7PKMjvSrx90aX4fAK3a26XsPGuRRH63QWeCmPvWlDzxQXQHQFzOoQtSwlbw871YcnTpGopaYxbik
eSyQKpMTAdcts7gskqF0+xzp9K0GXsCrn3ez4naAhcOKaz2rGPKgitrTq0ev6XANS8Xk92qUKJet
D0OeYePmF8/Us0qiYoTWKH3/+lDOa0AUllrJqP426xDIQHOkKPJEyt+aYpJoAWJhUs1Hxni74TM2
nRpL6VUKhO0TIO+AyrksE6YEdyP/OzFGyLgGyooSEpYa3pxOORd+ohy/VTnNI/uOwH5bYKnPlEB+
8woJC5xw8p5zLRN88mi2Dt3ir4UkO5OLqZoh/QnvV/RbH+A3vKIVSgcswEym5j798QZR0dbamUGu
+WK0Sy3Bm61t5dwns4aksZdSAXRxuJf1GFveZxy/98m5aJkM6JiZhZN/gXQmgMRouNm2dapX5MU3
jzgrVo1qNn35RVqKm3Hslphb8bLBmExWDsQ8UWk+BiwSwY5Rs54dUavIQcoLwzeky39saRz8KQto
Ip9QeB6h0wCVPe06QzYahcGfF0HtWuq8jZPY3uRGxPclnnD+fv3YzKx5hH7w3wL9KGYY91lQAojO
CM2Jfb8KxOFC9bpSy8IJAmn8rk9nAfih44RkiRGWkIcsHcYDcg6FV96HThO3o4sksiDIXDjoN3pa
X4fka0G+5tAeMYlPrmbavvlL+uQPGElXp4MaZ+or/IEAvSy892fdweu4USvZxYS5NuyhbQ9dpIFh
3Z8Hsuwh/5/CULXTL7rUQFF5UC0pgWiNqKtULCO/60pSiZAJtX/DMYlQV/FWvsbHI+Mwi0ZYR88C
0yEpC33Pc8Intxn8g5YwktHuQ5jtkhGEOiDjNmM3JnLbYhZt8OdULT+O6wB0tqVImtU2jhk6DDxu
yMfFgixYi6CApCqEW7Txx6O5g0xFreaMG1Q/BaiucswH69+vvpaCHRrh2StCzHv13wo1r01dtWqb
Vu/JBggUjHKgONoCyh1jGVrR78hlua7umSGO6eLbRsWUJMV9ETZVf0UgvSaihk/4FuwENKkBUgzJ
GUMgzNQFGxV2V8p9VFChntVhMd0gmfGh52cpuX8Lna1+2M3ZmRiyvMexcRDd7gqyeRgG8Fx7QxD2
66tmsCoVawGZFCxc/MeSFFype9ISNpLd0r4eV/nnRTDN1UUVRhWYfSp7ZoSC/rf0oo6iEsckuDuq
eLMiQ1sQUe7PvoaLPLb3JllsloogyMyJTLRICnocZ6d3FNrQb67DvpxXIZ2N3ZYjwDX4jKmsXyND
ikqcg6HW2W6IM0aieF/n2CUdqn+wts14ILnCGwX8aAJD2MW0xSsy4lIKFZDXgkN9FtvAVq+IKevX
FM4Y5D0cuIODsK73al6YAZfyq92JDIBOzBX1sSpukUjqekzP/jfc8d/EWfhTHPMdY1RLh1Qp1DUA
Fme8W1MoHZkdNB3QLBRkYpfk9JfiaKJkTyEj3dO7SbrVGinlF0AVTscwsox1b+1942JYkD1iUb3/
U5Hcmr3H2agC0pq3oUS2WBr7BC7FQo3mmBwhVdT/D9z79Qg02JLmeLrGCLfS4hiyFTMrALknz6Xx
TzL65ma95OQkCv5hujEPOQo7vlJFHSKe+D633IFvRPdFHU4Ctd89p6F7199BAQczxKzCX7kDyvrU
YmJRvQAP1NkFtOhCJ7xtiDGw5QQ3o6E1YbOy3gkveZdsC8hOYrFgfKM9a7aiMireYYBJ1z3P4Vng
lJWIYfrrLpKgvq91GdHVZn/neginPcwGAJ8i3lkXihcTE+k8VB8WPRaFQMW99M5i/FlfwLxWYjRr
vv7F9GMBLowdJuRXj/FSHptNQgvPs6T4J8Kt6koyQ6KCEgQZHiOpSQsJ9klImWfmkE9so0U3mWLj
TvC1zY+j7NLmsBWkvHApWXUYJCzLfoXPNf+vFypEaLhiOPvJAvPa/o6s9vN+4MmLc86fhogFs0Fn
rUBQJhfTVpYuZvBRjKzK/Nce7FKhUcamME9bkHeOSyPR/xWQPJRYslTBRBSQIaXJvScwscDScWHe
jnuDgGPxxvvyzk9183N+0wVgSvNmconO9EtHPH2Kur74vuzCXaNiCQbRr/X9dIdY+g50ekLe5gNW
aFBY9RcgJD3SU9sLP0w4f9yWTtAjXP2tYLNnbVhsiZEv493nHNTmUJhkS1JoCzeRsrWrxnUzrA1w
BFnAOh8d4gGIq//cjK31swpBehw9XKVlLzvX8zFvPoiYPPXt0umheG0kgZKshsrd8vXxFHB+C/P5
M7Mga2kfO+USgHd1RObWbGpEn3x3KDvoaPcXNrZoXjaMwDaHwFFIw+30080gkmWD9KCYDLHW+n2K
U2NcUCK1NK4Q/UvoC3C2Pyrac1WpUT85QxAbwsuLvmYrhMB7RByYhL6memE6tLPsQn58e9+JAdVs
J6zEIL6KZpfx7L1noPb6iyC51iZCBsIUTC1/nPre0mBPAMOekXqxhC3BbXK4Bxzv2FABFjG+u5IU
1xi0r9aMB8Q5IKMeMNWzdOpY+jiRorvLWZGn4lV1kQ10eYmqCWLUZTucYPSvNYWzFqUjdAz1/dV/
FzVRL5Cx4YVOJHMXRC0aRzqt8PvFs1rF/9xRXWicNJCqw1w3SKpuy7QYdnVHwg/9TkY+DTvHULVe
evrJ95Z9z/iR7UxJCEfsp4RBYaIDoyGpmYLvpXKDc5GRq6VXjbT/6LiXFZU2hM5RjdZ1aKzV+tWZ
jpjwt5p7O5ppxlc8Wb5BLQXlb+ogspdZb5Ftiv5jd5apW9pMUX9k02Drla8Mbo1upnNY2lG/gZ+n
MstaUZRj1M2hE3XFue7VsxZra5/ihI8JtKyHA6WtHtmo5b4VyuM92/twsBbA5eXb/LoFU6IMqmWK
ePLvuixoMw6uRt0DEiDuxcXbfpZETxu+b1+3jINvey0nqGBrj16mnYEwxiRpdEM4kCzOxkFiNcqx
xMTRKKotxiqrfjs7OlKHNnXZ6L0F9jUVbm7qfR6YuW5Hh5+wyxD+IgOQkEoBisAx5C/9FVKQk3oy
OzYCDO1lVWpOFsirNBV1fJTjZZKy7wmYc2Sfdm1lfWND1Y/Hi6jzDRInLZEvXfGYrMbcp3pexh2e
G6WjokAnb1gBaIVc0x9QS0J783lc0riyC1+9tVMO5aWqDVzuj6pD9HLDN7hrda8lksk804hNiJFV
7IBzl42dFkpYMOT8mDvewFyyFgmj0bgRaXjpD1Fxd9cHuX5cmbsMGzQ0U9QGsSP/x+ps3uJ/5B90
e34MQDEa+7qmALNxfQbdPM1Jra2vTCwBylz3tCmNT54Vh7hMFHqDWMRby6k6JugPxuNd5cjtk8GT
7hJCeYKQIY4t4RnFFezpTYyo0vwM3hOaFHPSr6x4o62sO0l61dFWSom8gOVGaFzEEV3oasx/RU7U
+Y3jl+w/afZdfqAcyurXAGkj/FT8orCugCGp2sOPkT2cvy1cn8Co+TnHGCsgo7NAViW0eVZF2NEp
Ni3y2x/FMru+au29yds2tx+YqGzmj2QS1CY5vZ8lB0Sl+z36qIAtWkV9L/DhjNrtxzQK9hP5PX3A
RP/I5BWmwBO0A/fHnhu0cduq1ytjHNsJ5Pb5xuYX/8WnOJY3BG3NqOtdJw+Mx0wamcWMrQIp/uiZ
xK6rJ2rurlI6l89M3fZYxaM1lufBvo177sPRDOr0t1UdOXwK+Aciq+WGWY3ls8R+ZyENY7tm7ZLQ
CpPsmqWhlDz8PAQLjXBvMtv4lWx5gE9MZXDeRUmlp94z8gpHN/yqHZm09divHocmIRIWFy3lIUof
qCr0zHqdmoLrTEGOIBvEZnz+kCXbL3b//4XsOQ00ipS5kNTDkyp3VGR0Pn5kMpJnkotUZU9uv6fi
+3E9Z4mXxje2bNhQ8wfszYKxNjjwCx00pnKe+At4Fe1IjSx23CAmDIGniePW2qX5D96g4NNssyBl
/5qFomtM2Ct0YfK+cDPZu0EcJLB0zY+PqjKzq7ZgQ4aZtveu0PBrPfIX83u3JM1Lg4L2QH4APOaf
wNWHeoPvbtSE0jRTOIo9+nYIvZeBf4T9F8rqTdwMGhtSvCoUS5iRTISKgf/gtT2mS3LyGwaTRycD
tmuSDjpYXri2yz+VzwXYlq12MqwnOBsjW5VFuEoE9PzZMdCk2qdYP9774nRGmWWAkM40PmZBdfg6
rOOexRDe3t2XIVDcexuxHuYibZ0BAmn7ZOhergF8oQtAC5uRMI3kDOyssnW32qo1A62NPnu5sjYu
TRfharq3BfoGvrYtBjZKr/9wrJQz3f8+uZNqnFVDT3GdID7nctLKOm9S3eIAFvoVjRIkuIwRm9wt
/JR5QlMw6ubgoMYQxfDdNWZrHKR4y2yX/D4rj+D4B16UnkWVUHnzQuSa9W+nckZMtSXsHWOcJ9nK
5OIRYcoVCUP1bGDDI7rvzzg7mYLaNHq8LA5O4Pudf2jHXzLbSgxuf3Ojf9OgzScYSI0yh8FDjVP6
XeFZp6Kr9nIeNokj3fg9OZJxZDMQCTzXFc+J2IPuUKiAeNdwnkmqhSeoFA5httHPmWPe04vWy65p
PAh+N4vW9BiqrorZrVK2eUkyBkzjQ2ARRLB1/h+GdkSdmBHJqycATy6/MstlfBzamAglOnsUjZam
nMj4O/lw+7iC4+DW/sXwSO5zVRdpTe+it0rJ2Z26IMCyFNmKsX18dYsYByBMchh2rrpFhUTnltQi
g/g0n9Nl7nAIOFxPNKUxpjspfH526Pp1WjUCVXNxbNu04+DV71TU6jZJmJUsTUvakzSdbMMyWp//
x3UHei7BvIPtE9Fu0hnhS9pIZaBlDPT6pOXSj9i+RmhiUHnL3Id4NvE4tOWN75eSawJutCVw8t6z
U4CMKq7B9Pu31H2fvwS7nHEELa7fzPMb1XI7gHOgLPTiYVgVFtk4GZtvzcG5gMj7s9EM4/13a8p8
fo3VY8GVH2Wm5j/V/M6whEQAcodd7MParzIhPaN++0s0DYKiKqqA7fSctvm3nio8BLjwpw/TiyNG
h2NO308LqoUazwG25fGfvWy4FrXAvxywfWR4IZ7dFWzwW41QeJFUAMLaBIsa2MRDVYL9DvXI6nFu
8FupmRdWEg66p4/bPdSTqg4LevNMhksK5/MtuVo1nNUQBj20WgyUfxuJ+QWgQ92USpc5QAgHvcou
lzM8kkqIFn1CVgZrTooVeZA9pSwVGf5s6D8vDDUtiaaOSv/L5qbGaCikVIMhu0CKZtw/DNiw4BPc
7OiAd1M0sykJUL9mKI5H4JhiGWJN4Ld49vD+quayTiMeYQk1vzBgLmQVYZDHYDUCuAN5ag1FsyK1
aiM4U3zhrJu+XxLxHgcjDPTPCqmVZggfhmRQXPrkbbxYqiebzMn7GblkheGTCH8cT5x0SP+6Z7bd
7BTidOmfNAmLP3CIAB/K5PPABbWm0HpRQyShCmkX92gPiZ5wMmEz93bk6TLdkfD40nvoUAxfjh++
qpowjnit9MpuDUwC0+T5D6kvcXtk5X9dNH/0QiReafsobQPpPBpAbdpUzEjSBVydQv/8BMnJf1wa
dbpV+M1Y6TJc9Qw9wdlCYvwK5OTakM0VD4kY00COiDsrRPt/Qfzw4fpK3UgAsWmvshiBGN+DUL2W
N+3g9oskTYYWonE0d21aH8Ird4Gp5Q044CJkBrxAQuvQddGXg2dzN61UGTGRR/MBPvdfzv83CzEA
UL/NXzEAHRU/5vbNjSPdmHvTm8t2TCDzEoSaQTGO/1xa0HFddU4mG3oMvriQdcBafhVKIcg/evvZ
14yymRZDcEYuWTobxT+4Av7DmtSC2leDwoybbaq5ZkuEO2glRNne3eg9JoE2K2CqgLDOhlw2yIeZ
TAyzh6J4WvfqIV0yMDjGYmRXQk//u07oljtCFetwAMg+WODiRDlp1vlXFl0TpHgv6m2YIBog+ZdC
pdmusuohzXdSMcIKSVZKVDaS/vZM5Qsp5xK3ushS7h7m1fxn4QsJUPoUIuxPp2hEQ0t/DKi38RRU
WCSx5MKze/hQudL1f4hjurEBvwX4Ro3juk4fXQ0Q7p/4g3aRm8bDvZFZwsUeKOBbWSDTv0ByJhcf
bNDfqIc/V8vJjh9DOM1Qn4IzeV7frHOsMBt/r0/NEV6xHq6yARBQFNqKUk6DIL9gb3JOPK/Uk61x
ywDKk1H1IaPzoZOJKdHZXhkPI6GZFip6Kckh0P4KW5qh6eZ0F33gF1seQfy8ZmjbtfUhLDcTydtN
5R+KV25F654ReF1kCl5Zlp7v9m828646nQYg/JJ78XpJNWIk+vlZnBDpFcMDJp2URt5Ag3WCapIR
h+7icLJVHF+Oiva0BGILstJW0zdh4SNOlvhzXxijkArcrA5hp72Ych7kjOcYd+hytZMCkxK9lsbV
ol522VwAUePZgrfQwu62Lm+VXdB2xsgFay15SJwipbUmCw/ggpo1nPtVRBRbD9+Pd4XURBoLF/8+
p1TMYsyo624dh1h4xFgZ6ABL+ShQN7G5JHdeB1rcViEk2y28+Sm0BJAaVCtc+9eS8WuNkSnMeco/
SRO+G0shzSkCI355UX8VUbq7oPF+zFn1kvthxed3G6C3wD+26IV0YHKtEE5FsWHO0f/u5WETpgBI
yAUe71SYQQscPQgW7hCZT0ZAPU2AGDOEANa4hBsd0dYyIncptnoi71h9kndhl8WPJVPDTqsi6xvo
qJVQ8e6/573s3XDV2TSWX2pZyJwnQc0ZeLi7cDbHQf1pLn6vrGeN6AY7jvlyO4uUnnNmL3YMGbja
NpeKjWBW7/+Epvaffi5SLG+sCViOLz6XnmD2tODC3BzdXmEzW88L6nMpE8ZL4ICcCBjT2mE6foD0
s4VggzaFssXiwKxVz8YkwsmHLZ63GlT03SX1iZQFsXNdpOW1PTWVWFacKthuzB2KsZTHUOWUO1bl
jPifppMay5+a61Vncp6us6eHPGNxIFUWyI5TTT+8RoqJedp+3XznvHL/k5Lz0/FxA5CYtKrnSqJl
Kq4HCFfZBk6RDw6yonrA2fHanMBVDy4S/irwjaFDYOsXdqFSIkFU2UEnzds8kGqyP7XhoLEr9YQf
XR2U+k3ljMwdOXBCOemgMt8YksVtrXYKdDlbVoYFRwED7zga47LE3H6QRZiEbS1hFsuYGJV2jDdQ
x287/aha6v/gpPlFbX3gEInWMDNl7MU9UqheQ+csWOJFQDBIYAUKXy8lE4sszlOUUSmke610iSwd
6uZU9s8y2pcRAV6CBv1SjKtOz7oPgdqBUGmBWjd1tpTgHru0jneNUOPyfeeULCz6JC7Hjmlu7znB
17hBjqHCLvrpTFaSQ/CrQ1RY766yWZt70FTy+HOEuZhhLUtFzNr55RqF8wMRlXb8h6m7hrkLSEsc
bShnn/jZoP8wi3nQ7ZZci1wNz/X2odRA0yZQJxbo9unExxl3Vuku4G6gn5hMfm1de1Vrzt9cSECq
RDICsZRZ9VR/r1Igw1foDlRhqPZdTmURkQXF3sA7PmRiW9OmYyAXmycwGBO8b94M1h0BbJH88NMc
c9wJKve3JZoNiYwAmx0Ub/k1jAnFdGUDveGEVvKUdvZNLpfzdKiq5gVTO2u8x7qSfbo+LdwOBOf9
tjPZC4Oly2es6kHGVKPFTOCHA3Apr5sYDVsb9GP7aodLmIVCIllWFEUAxGvvQ+43O4HN/TzVJJ3/
veh4mD6EAihbCoUUYgQQQPLyVbTMhpjDoJcvPPo5grVPZg3g2Y6sC4x3Yeu3Vk1Bn12JAofpzX4l
YQtjCzrUnM9F/YenaU3QNsX9z6hlqYm50LGZJyGQ7EG3xfnIq6jNfFdA5ev3w0DAn3LckOFykSEP
lv0NuNT2ADB9D+m2sgJW3y/zwH23KCKS4vRzfff5B44PzufU/xNpHOCteMvcwjJtgbRDGUuORf/Q
eKTFzT9zmkOd9bmM4cx9utnvgCOcTpgB3knndNlDnuvlqrZjESL15pOT4IUjM3KJi7codbqx4poR
LKu9SX84nHzwylRSLo1sSfgbke657Hk9ZYiX2mNFWYzTlfevZ/USHKw99AciYL8OKxmEF51ToEei
0hvOOd/mWFHWAseD7pFvCXicy+ot5Fegfbop+uvCpfq4yjdADxli74c//Rp6Ck/6s6vA0R9FR4Kc
gBwyw+/fUsCB3bjgx8I+fxEwXkJXkmAOTelbtxx+ONGhQct48naiSz6U3jwboxB31iuoj+DpDgqP
qdQn6lW5hLtaSj+D4Ci8t03s7XKRxEo4rZGXKbVys6Efr/l9ruQ7y9W57OKl973Iop6WdFTH5Vay
Z8LqqPDGPNcelE808QFeBMPN7lJId4Eh1abQr+ysuFHJTC9/vzyUIin5YvB70C0QzEFqIyA7MGlm
3Tp0xV4Q1nQtHS0COVjvua6Gi0IirTeLDvZF6jkSTQfVIN/TPhwwuXnQBB3nt31kGH6VXgG6zZGx
Hx+n2EjpajGpeTPaNCbz6NIgobQJy9EjNN+CylfvnwZp9C/bGDFuF55YTBiGfbse9OJwWBTN6ipP
X7kIZbK+IWGvDwNipcsnAywe+KO0eTm2ZKBJiy0x4Ne+JHAac17cKi8HJ6KgRbCJd8M/U1RL6J9P
/JTlFM2b1Xc6em0SY9IUXthZhKKXtUuTZpRufBJYF7WzLmtY7W+kgWVq0jLfF5HWTPzjtntNcMf0
jGxfXVYb0xuuKF74otajfs3oX5GrrR6+wITvfB4w2xhNxjl8oyG4uyxwmxExT49WbCsV6s1q8j01
yKJkeQON31lhsDBMR4Nn9Os+H90jFscH8EWl9e6w17SPINYMvZwE89eTVL51jt94Di6utLBi9OXE
YvhgH8S9FyuMR8QeMObR9cLR8piAHEMm66k4RnEyaaxgLdbstBW9FLwCQX2mwlAPKeg94CO+mMUt
TX6LKEK5fnz05f6EJ09HBTNhmcD3Gwr9QLi3pygHZdzPTYGcd6aJ/1zcjGQliVg6NpaImKxaRQwQ
n/dFz5kto3tlGwT1ywuhX3Z4zo9sKtbBAH9T78YSW8dLRPhSAkfcoLhzk0s5gXMx2Dtnzcz2SdYH
5xxtWquZPZjXWh8ahmezhTWqcCb3VGnsi9zS/kmpXC+yJV46OaX4nFKYp+f6ewNN9nnxoAQ0Bp0Y
vvPM/rPSyYuVQGY1eJdCtfo8K4RNNIB3dkrv5Z4FbU9oD68MCo0SK287n1rm3RXJzGq+SKXdWlTG
e8Y9AeErcP/e/59CVTHfxr4F9jujeL9r9npZXEeyLMZ/JGfCYY45uFnsRskrckDbBX0UQH72jt6r
M8gYRrraw7BWDOQ85hw5ilL/CNmiyuqjLr6XYfyqG+deM/Pm9BK7y3k0moldYyUdl3OzmXcylwHG
iuA1c74VpaL6joaTEAirfUITuL9B2q8Q686CecYTSvrwhLffvj9trpYCR2JvvGfECIlq9vX3Aj7y
VmLbie5mvOwO2eu0aYUO97vbEnDtW0T318PGbDCjarJ3hWsxyAKxgI6VCwrkoD+6zNlEijnpzKtW
GEKrUMwGYLmm+jrjCMpy1sxFFiW2S2Qxf2Lgx/uplTJ8gZSV2L6CaITG2H+YHJiHPtMSrsDtF3Ml
fVuRCayvCKvtkI4rqpTd3f1RX6uhNYWlfYpwio3iKowPT+Ma2IqmNs5/MC7ympV5hun+S80ZGOx0
nqumK6yfbvTKITMYPcAeUdA0T5votybZ0TsqAVr5QaNQPTAp7dX1NCpO8b1hgJZOYv21G8qWYwSc
pyUbyl44CA+GffJPgTFzGmnW+8lTT6n3gS81+CHxkOl6Q6y/FWEJPS/LcbM5hQ7H+zIgiZjqjSt9
zpvJ1RW1+by/vEbd2jQUHOT4rLF0CEeZSjpaT6D3sT2FVsI13xwmdt3tHhp/gt9GAZEWCA1w0T5o
k5TXFD3SMApa4yH1QIJtx5T8h/rwb9SXxkzjR53rz6mAHkhdSAC/yPSpSg95xBUEOK42HYAm09B6
FBlRf6mfe+5BvrxoUtHJLSuIKQZIOiRlmLTKhSAbdYop5LibYqOfB5iF2xidoc6pWbxowrH3hjnz
h3SP/eUyr6TCIHlABP4o8sq54HQ26CC2ivpoU1yBC4o30UozcYOgBcRgnIgSwo1Yq/iwMd7cQzad
AA7+ZgxHP2K3nRprJ5FhNQSIoXsT43kz3VKB4duaRPentaSNgmlXHJdUoebD51F2Mvwjzk7Cdfn/
AHe3bOpixv97K5/GZ7loUTmsWomcBM2vlOBwUDWnURKXLQWSFb6nYvfVgaaHV8jOtM3KdyInWeXG
OkCg/bJ8yaiPLy7Kmpthn+YK9RZC9zCN3Maulf3jG3kHBrGz4K3JsDDJ7RrefivQBT7uOGcz2HXN
4t7JrNvlmzUF2+9g5jbijU+PnHo84yvrpot89Phnyy6SgoCfS61Xd+tgEJpijJkQz4nmLXPGkssv
jTDHqhRRu8NLN5HLjnxOv/TDJpfNITwl71cABb2PVbfSJomCILLkzavACYkbOewcHYHELuhRiApD
INCn+NdzXbi8ossYN04bSqNRh/6M7kUmjgSaYurax+eoor2guiE20EkEn6aCl7OSJsO964b46lNO
kS/j5cgJ/6WpJk52LI1sBC7zYB10j/SwnOmAS4tF2wAO/sd7rKaEjugdKO6AHMPHj5vYnt3Z2jme
ckOgTLuNzuokIgrwN9xm3txwfg5oFQgmsE8orhbvaHYFiQ6a9MYqZBiVARGXWRl5oRVesgEcs9xv
WGmKt/tYQKU+Lt2mnkSYc1tM4DbJrJxo1G+u8e2bjNgrtDfeJDvLpaZEAdxmuaB8JhPwQBKfXyf2
TEMvYJU/bnxnRLkgnqdSTbkcKrdWnlnCULUAnUTfAjIqSxN26WU8YKBbgCu3XpdH0qc67QSAEitJ
ooa0aHqC4C77kSqvMVC5ArcRsYG8o5oTNAKn/715H+5NJUQnvRUmHIb+HOLrX/B1xEKN/cMb3Hu5
euwDDmQxsPTuMVUmkJUqhjCZpbFrhhGgwQ95qk6qjLT2hg49x4lXvibi/98AYPGEMtk8PxmtrVMA
PiUT41w7/5q9r/4ZvwKcULMzkyX/BW+BtEACPq0TiFGiEN5XT6U4uFbBmywP9Or6spv3+A8+uBwS
Qurhm7VmXHW42T8W1kod+loLeqc50zCSz+5qwtjxmY7fAXnG04GmBibWbSa+wv8W6W7yA2cg74BI
FyPsArtz8JT7lT6HrgwpLRNfcnmxBD1R+pJQrLezyEnUAt9cLOd3cEsp/+K1udtX2bfqyDtXm7W9
+/biTIA6i8l+eeYet18ZBI6u4Fh6qIGft0Iqh78xj4OqRMWMHNC3uW1V+0zpDKTP+0I+8wqkOfn8
fmxLjpz4KkqDoGe3ShhxN6Tf4DyG9jRCnqXb1gFI4C5LclfrH90Ro+WehRaiibQl3fxmhDI91y4G
ZGN/OomXI9weGrsP67qn2PhCZ+ebZZkXOtCm6Iwqat23iDvNVOSm57evZbt7fFIf6szUdla/vDBe
tTifQ8oLgtohLgmGIe/YoFxfkbG8Jvjhk7cRLns/A30YOIrgatocd+9DWer627I3LDA7Y9ozsB4a
SFE9LXv8MGXZLaMo3akKlLRi2h+5XDrptNegxE4vGbBy1agFTb75+HL7hHqBgfKqU9HynlDVyBLC
rsJ+1TDzI4ilwuy+9bnOjp28irOaYBwHLiW4jbWLw4Xr4Y0YOo3WE4khkzoUZhq2nWbx8+lo/cim
275gxtlL48QDiWGNukGMFkbQDF8UDhzxcLUvYudFM8A/+sAV8UbWGut6MBIWKYAipvM5fd6beEvB
s1ha7cSuvkKkYamoHmeXM+nvX9HVHUbjw8oyaIZOovylikYPK5rGtZOFtmXaNLCs1Nr61BpOvGxJ
RE3gsNx7ccOwUza8e5eErreWkeVAMTJ3Hko7RvGSuOwC4LmLxGygRfrHcNXtRaYcG8r68k88Z3Zb
+GBG0TmGSFV5FvzqexFI9zXLt9VaARa9jjHIatFYrdygCsVB2aF9P9MKsUzlr8QPXCelLsrXRj4/
uOaQQTqNwros1euHTJs5Q7FfbNWKO16MkUBywRZLhBn7OJ+KxiMS2JOwRF1W14IkUrgLEWi5z87x
BNtYY5P/v0ulDg6DvotAez6b1NYe9Dk4/PLO9NUPnk32LHTGazZgrXmU+r+VrtHkst6C1mTsRkza
GGpYEDvRG5eErFvH/ToZvKVKdFNn6t6y71wpnLhZiRgF3LfFrxJ5ucV3yV92/YxiRRJN+/pw9Dvo
Lw5qW41eQrBuXgY2EeScpPj7CO2PM+tYPHUym8qwn9XSQ97O6MPSfZWfq8PBa3k7HJaxhpjMRJ3+
jsYvhEcjQi9xbf7D9c4WsvklIkk5p/eJ1pvENUIcNOV3dI6HWqAVYbS9XIHOIqrLuYEVe3zaZ8cD
JAdzveVOwxGIWyqPXDPo9/Y3GbS+oWMpuujYgyKrojczCNiWQEV30gsUItQWicWR2M8/G2p5HDQv
gki6OQe6mBSUk7RdPFayf6gwvgOmS4jDpoOwPoqs41qwoHTtLKBHFEXwoYVSAK1uzpjq6JZfBH+r
A4KBLzi5NYwJIXQGqEG54EUWmkMRac2EJNnj93JWqJWn1sMuqOm3H1hgNakU9Xhoad6fnDFejqMs
bLpwnqXwN58Tgpo0QMOYnzy7P554jVQdhKAG2/l3K6I2pfCW6BLfFTcphZpxWmEWVyTTJIMz+5C+
3z67R3uIEc8mRLJ/MJ3njIc5NMb7dc684h+PUfxcKoQSwXtPwglA6IIImid/8q9BU9dq68ykF9+J
Qv0nTuB8jQ89NHUQrnJ9CcGTG0aFIFpCf/uX4lzeaxgYVvB4JOMYsGV9loQh68DusMmWIXWkCyia
pn3JgnWmouWS3kJ9U8nXUrCSrLqZSeHEqMhqJcmFO2xY6xJn83yFm6BXUuzy6F0a6Eg/ZVJQGPMC
AcYJUAcAr6B24TNLCsJDvwBIK2Yp/nUOit+dpjTozXcH286B6L+kC5NuncKocuaGYM5gb7SIw71Z
aexUzXsYET6D/NXLBzFTVY0eutbxEN9vWS4Ufncjhe2A6FMYHiJ+HaMb3IebBbzgTZOeTbBLMeMm
QzfP+SFkKnKTeqdFjtIPGmbq1SPmk8a9Mj/yEXn8tqPlLQiv5hF1RgN2d3Tj04SCtcgRRzwCWAb5
jyCW/vrP65k85IXOuASrbrntSukupNaPomYvaju0Y+rmu3j9K+/QS2uw7NbrldxRSK1zNTFM8UDg
1LqEJtJx47tST3Awr48oISz+SBasilF2mGR21lY7ZXzGx2b2TsRZD2uaEdlUrM0MMle832L/rq0c
tgNIAwhfnIK1iZJPozAlA+OBPM+0BgFXhOngYckqfvBu/wXeAarMKuPYq/paHzW7lPTPMvov8wwb
SIgv74151nbWViH9jjbZiJ4Yf91HhoEyJDeoTu/p6RYvHte3h2Lwhx3PMKFS9Rp7hEhp/+68AqUj
bqqgKVAi+K6QyBuZkynFyyChx1aLyCHIJeg73+axNwxSK52KfNmiQ/JGy4YxFHk+ClsVOJIkZ0ak
O6HVNLQjukia8cKCw7PFlmlCO4Yg30e8hPJCPoRIKWkIICy/8EiPhj68A+96hH0Hm0tDfbN2qx63
g5cBgS7PjZKIgvwAxBTAhUYegHbJpbbFWCLGpJfVYESu8leBwsB1U10Z0Ylqv5PTs/6kj9SkUM31
JVFu5JMAqOJFOuuJ4gtXqUS3FO78aXUyeGHYHPKLvuP7BatLCsUqHBdGd2I+tvyFtXkBaHRZeIAS
pueNDOLY+P/U3T4RcZkknur3e5ADOYRKlL3lIKomwZiJFSzq5Qlb6AO1lA5zkcAhAoCCnJE5FrYH
boIyqichhJNjn79aOBlxmW6uIOK27cq5NJQy6+8W3KT0w3Ee1B9jeU4H4soax1M2JOsZlRkUapJu
HifGjc/DlFBJgFI5cMsk1/3wnq3ej4qZXjjukwhIGRb9jTe3wtvBAoHtfolHWf2Jc/FaFTL5QGXX
8JHJWlIXgw4QmIB+PFHVmEVZba2K2DFOPAEtDcuhsPlbmk1Orv+vdGPokSt0/GTi5hNIUgUa2FsO
bFTZBpNdQgqhOZkxZMnDoF3dMm8Evhjt6O4XHFhypxwoeP/+oGafRHIVYyUcesw3auDaODLf0ahr
Ssk9vw5RkwcvMhYnn2hyEG7JzUQ1pSQlJVNXfUrjvw68/ohJJxndR0zSdFygcvIGVLZ4UVaw6Gy0
F1ZlS7/uKjXxNjBKhEwsHWE/3QQHZtJfSWdGByG4Aq9Wb0/e524VTjhjmXvcoFzvb3KqocdrzKUr
vTzlwMdBk64YVvkHL+ixac3bfTMqT+VbS4r465Nzw5CSSyOY2R4iUwF994I5qU+fhARjrdvXC4dw
Qw4d4ZBoiDHqrvwstb+K5I2OksGSV2LPbc1g9kjBSWT1CK7//lKk950XbQQAukgKG89KfzybchC2
vwyRBkmsi+h8jXx72NhVcY7VIl0YiOg5jXA80MBNW+XrWpJB/sC6dnnPoUinklJVNmTZ3jSTzmOB
DZa1upEYNGX7IEGDNuM1Y/88kpL+WlD1m2uTCjWleCNpvfL62X7KHNPxo5i7BnjKmjN85UNKySBr
JzeUZNY6ArrnywqS3tCTmeUEwr7UInMeQqPPdQ+6CmbF9l1/j1XLfgAd4Pjcwl1uv2jScjaVQ2VI
BggMPpz4wKSw5FWj7ZgkXTNLI5c7RPzwuZzjdt9huhRFfbp+qJ4MPlXryTSBKzUkWYq+fEfEoYa5
ZOkP0qwfGECjvE3+oEAge6C1SpQif9ksT7i0TzEwgWXowDX3xwC8oIk11x74rAIBqUsVvBpCRpqP
Ni+//eHYEuVRUhoihB+jQuNkMPkX5Cv51xS32rMS3McNdV/tqwxXW6wTLZkk+qVF3KchMZriGBVa
rl+5Zk/FlgERWm/UehcaOvWikZ1i3lXMHIC0/SARYhb+cgPmDCFdhbmMFaMeBjKnw9AUowX7KqP2
fXnvbQ2NFCAGauAA6b3FRflGdm3JZoGBU053VqJwoav+Mr+lr86wKQAO4KgFWs2zGO5yn8AF4y8g
z3RFcvlBBsmXCtnozExY+bapWKh1f6aTOIEhfqwMbYFUyQ6ibrhqKyHYltS8p5kbNQCiMs2F5M3c
Ludd43DCZlQARC1QtlltSCtz+jNB9EyqC2VA3CKyPrN053O1PKucTk8vBU7DPuVosKnUjNAoFo9I
OEItmyCK+yZuIGEl5V90Mt+W+ZOYmf/7UVvnY9T4muF0xPhfr/s2/UKjJZO0DgpjVo6kTQabnLWp
1WhFwMiCHAQy9yy2but9rO4ZihHvhrAUtdBK7wtplrAMRoF55Sqjjni83cG5ccXmO3hvkO1qTBY/
lTByBTTWLb0yc6qHcD7YV+nRi+xdOQ1EMoRSw1usM+cGe4SqOeiQDcmibXjSn0vug8G0l2aFe7dM
navsns7s+WD59Wes42JLiOS+2kZD/rBznF0xO6cduxbvxugiq0bAbtG+Ehg+MwEmRg5nDX/6IKVi
2bT1qDGE+KM0YLIPo7tQ2ECXAa/6wTMJrAKm4ci6Or4Co9gZcPJ9Pcy6QpJusg6dMzoI7Gcm0qxa
TGyIAU+BFAeZyS9eFpK0odOiSo5l5ZehxxAx5Ya+td8LuLX40qD5FY2W7Y7ZTI6AHm8PFSnuD0IJ
wYROi+hYj2agPH2gXoJRUhsx7Oaicb7ttpyuBLb4XUePghkVirayMB5fxn+oUvhqMxiW7wW4mHMk
EoYIdstxorIRUEqCKrJ9tC299UZ4h52cgOlbrbYIU5LSBE4XAX9W/gUfOEyWOVBKN7iDCnMFIPZ1
lOXmj1qWNlGUBPJ6u4Dlng43pr4I2WQBzsahoz2c2euSfTixWxZ3pxvQA8+ZuOw0sA+wAYjdr702
Oh1bKF5tRW4CT9eSDzoybx4Gry7RqjWIihsbtNQkEki7bR+LafookFdAnNAWxWKZl2Y1G3TfqWEp
Uu5YggskrPpr6LL16GNw4YnEI4w1Pte12ntDMpvF2WFgsAFxcN4GBr4sOsL/4IPWNV2/5euyXpTh
qwFeLffR6pMOnFNPNKI3tSRvSGBAfL5M9I7KiYq+9lwEgKH0VYF/6yU2gSmfXqmBME11mV9JlPVk
Ev668CZSYBvX8AM/G2k1kXOu1muOoO5oEkVcff+rL1XfvgLd1Bjt4LzjIIsp2BRwaHwrfWyvegBB
X0cEvLUIcwFXT9ZU0VE5PK3eU8fF3QOJJ6T0ryBJVfa/VXbURcdmcqeqrthcW5GzvBRnkdYVZ8/w
sDkWg3scP/z/GrK3D36J5TIDzhJCaxt6NZGeIMlw4bdJjbx+PnCV9ajmDdFVHNA8pLU8/Huo4kGo
SuaDnVAQxP2q9Y2fWzmonJQgBwUPVrzhIeHOeQsU0duHs2an0btwDYj1649LZlBOpN3CyGSliwWH
anbQ6ltYjwEa7t0yQoDxPilvDzEViXO4FsHipEu/5dryiOftZc2IATFyxthRmFm8+4ho2j5APpNl
Befudv++hJuR4z5e9oersJ6xNnjREPSCJSg4HfOjSttiaYEbPAb4GOKZpDni/4q/TQC8KMhP1Cq6
yGlZMG0RAwszpg7NV1JBTBFD3Sxh3/zWBdebr7QJkV25iH6AENnKQIUpUkdYg5aMpDPW+3hGIKe7
pk+GnSfOMXB9jUUkIjoC99KEjJd2uKvwcEPk1gEBL/7bnoQcSJuDYd4UmTZRK5vfdoQ4CN9Wgx5w
0WMklobrVrULIWacxD6F8hflg79sF76QuzEdzqGNdVpx+zOKfZ6qzELZFK0n9vdX26/G0eQ3dDFM
IyswgJdGODwzA8KiqWUtI9A9Hmzi06khx87ILGBBUisCKRWLssRQHy2GvARlGUeypyv7fE9GaeRy
1hXxIS/yXrzSo8t0CAr8n/y7CEoNRGCpfsrvg6JFpS/eY4Kn7tBh+NhB+9+taItlw7/avgKg8gTN
6O+YDKJfndcJEFPwoTHNadTWZuFHPJbwsE3BNeqFqT6ogyQiljqZa3LBjlaq/vofaim34kAYeY8Q
kdT1qXkLoVTCt96aaiZcFmeuEhJx8l2v68Dy+HiaX28eU+hZ8VqJs9K1oKCq1Em5cRGvV0en2MSV
1sm/PNfRHe/HOOzidfXH3H6IYfsjUwgwIVsh14brQJk4QC4GHjO0FJ/W9fOKl9gU1AsYYzqmPw5P
Fed8Rkn0b60OpQEEVZzywe7UwwSqkIFBhS2wSQ/tCNjW9egXaMhnKlfi+auwceN5CrkUTna2qSDX
8RxDLcVBio9jOrNODLlDLoicviJV7oSUMfNG0wi4pu1WGMtTj8ljMok4CnVqMAKiTOupxEgznRPK
qyazV3zfpf4quMxSvMGU4Kohikth2eZ1gCxln17/YG1ox4C6dN2OmGOY71sk+7Fp9G8mci8OLKO/
PU7ktop/5f2DKltyPxPlyvGBe/Ml4lmxKMQ02c5DG3CiyrJRe61fIJPPrxFg5RCurCs7pDZEwiyk
RDVvmFPl+rGVt+3swruC6EBcdzajfi1mw1UbpPXFtkx/sgjIHDMIgeiqJhg0MRQZMkVJk6bRcaTF
c2Bh+iM8d183G0N7KUSawSxEJykGAwcSJQc7c1GY/EH+oZv6r6laR2iOMfgbQu0jOOhaqGIYIdMm
wPSUEtV9OAdpCR7RMLYcRRguBJTc5s2euwq0qsocp2HRwcsp0VftvDdiRzRMQT6GemkahNhX2ON3
YrL4thcesNmx2sFxCJthJcloLymAM3j6LyDCBrciBwFNvfQY/XyBfABky2z+EBrXIM74LpuOCuGf
f73YKJoWRDXyi3pQJ8YHH9WJCNnIjJNsDRp3TiDpc9MEd4VVa253VmUkjD6IbN7HOoPJTNQ658hh
azbb0x0WGS4EmCF8b1fj4kAqITeOUXYoFlfi6/EvxZInrn0x12qxtzulOwbAYrJUZNUCUfxDzyl8
Xj8cG/RP+kN6ZJEy6nXBot1RgvVZVgaI1Q6hJjeWTGoFbPbrNNKmQStG+Jrq+fMGHw3a4lC6nLUo
0j4TuB8gpGvW/gJ0BRGPOhERZ5WRVjuUgbR+ceJQCtazPn8HYOprGcSDG1DeGIVM+MKR+GpZ34NE
R7be14GRQa7vJfQRaJVkEs46Gz/DAMhWI763yRhNlWCLhkOyEWjzx7zre1M9HBeEwhSFxNU0oP6x
e8OkJhUlRBd8q2GEyQsQLstNbRNtoYW7hfcLe/M0PPR6TfpvE7qn4ZfYCHaRkbzBqTs/adjElPx4
QQhfEQ6Qaeh/i88AsnWW+VSCcpPYVh2mjuP3XiUkQmm0+lyE0ExXrUpRdrkduhqNSsZnIpOJ93ip
ewnvP3MJGTLbuVZl1X4RufzjWduQrolDkl5q6X+2PHS4Gkg14sQ8u/yO9lb9ifaaxeMI+wkQG8U1
cS9upAiLQ+ipUgWyMnxLedcxWvYgZDg3lxSB2iD7yvNI3kr1sQQ+Xvuoqm7qEBPF6rE0PtEdNbsr
A0TB/xEN5t0ePVdgxrbTusEon3aZoazy0D/XEcnMfe+dBVAYcIX77Sgy9dFDhD3AHFMlOljiLC5Z
mC6nF/4FC9YafDID3EriYPZHGxhOFyfpot8HNbK5eUZ5owOSf5hMHkdI2VhbkNHFIYA5iR4R0mfr
YEh3mZ4ihE5gJ0NicsUQ8lHh438vPBUiH9FW2pRSL//lPhZzJVbpCg5dFMDNzeBdow1/PScO8T5U
lMvqK0JPCwQpRZT94iKrXpxjE7MHb00soYYEVjp+TjEPuC8nLIawG23M7IjTPptQGufGG3ESljlS
6nT038XXrEFE/QBqyw3mA84wJ1xpnJkwo0eIVGA1tHJpeVF8scN8eh0VHQ2Th6bAfLm+q9uHeBQh
GvcmMinBQI6MCef8+sWXGZ2MF71MpJOYcFh7mk8dKoEI90/DY91eP4KwfUHg2hsGKgoy150QDafT
CZgO33CbKQUmIt6Nko3mq5HYa/HQ/YKX54i0UtdIbIG/ftF4uvogH7aEuUM8vVP0iKehqO3xwfFB
MNx+rUpKxLIfllW8y7QzmtYfC5XaSf5gDf9rudjL2mORrr7rrkKrERh+uLvXBk8fAkquiSzcLm53
nDcNfZjuKC2LosLOJBCA9lHPQhrEcbfveb5eygztp80jF92deZvwOp1uDN8CB65FkVK+xviv5L8K
pkTsnXFOEwX9EP6Eb+BwmrSWsJ2H0oTN9ckWNpC2dzpEY7MNC5Epb+QTcLCynjzJVdcPWcf1Hp8I
gzBGQxtWWhF56gFIU3aAN1fDQA3Rpx2b2B2rNDhqjQr+2poQXhBxNfQ+MfpqpEClYIZpg0MSKHjr
n9hUskzY7jM37GDvA30UWVq9FfNmfYk0htxncdOFvjtFv15Q2IH2q+6ycO4h8rRWN//GKFpxY7Sq
r8cVOM2RohKGbIQZKRa1lOqUdUZVTaAbQTLm/J7nBddzUCYUJMAXWl6yGHgZf9m9/YguGZpf/6VZ
pq7Izq5sVw8SBmj0U6GiUptCDLiXPb095M6VX5LPNHDN6TWTrA4vNJ07FKVVBTmUtPOARxLC2KGh
aWCpRQ3lwcLf9liYXOLic8/NsR4nFGMCdnneYbayDwPAWqKFVBEOFhk5xGA3bhh6pj32pMqE4PsG
i4LEjRMhUdjXo+HqvCekcNFwe2uCghEzhAEfZD84dL1Xsws5qYAp53eO3+U4U2sVPf+LQ+yNOUrj
+w9ExwWrcC7YcikWIawtIUkpC9bHRWdt4GcW2cc8RM9po2P27JNkvwGNdVc8OF6PhtSuoZV3fXQ3
zPBBXP+geC9B2Kkgjvs1O8HFcKXe96YLeaoZ+M1qTm5ynYfCBFwhPV/IAM94twftoupxuuM50nf8
8S1/slIPsFsfbskJyv8PffmwhujyyFKt0qsQzOtLMNiwovtggZgFnJ58uyF3g2sLekaHQcmrKVN4
MQFT0eLuUdm9lxeMJd39xeOwpQlGvvIc031REXS4V5Y5f81R8CUaplDkgteQYR/zUp3ZMGoafz0W
5OF8MJbtVnjQPbd2ZKDCc0Xd4sZFuHXGlhSZRa//Y9/2irjAUh1zNvjW+aA/rY0oIErifOdCSqIO
t9hjA2Lcm9zvsN0CM5eLLIsZKjPCHPJJdQ0R7xjyoneAtH843C++F7gSRwwlq2sBE5xgixkwbbEg
lWPCnTUiX2+X4OQ0nO8eZNlFAWfNFKVozvWViO+EEfbXCdUkV1TAYhEesG1nmzCrjBX3mSbloCAx
ZET6Q2xH001PiwIPDxGuq33ByE73IAp4yJMcv5RwgKyLtLd+0x2aaSbTPfC7w+Nyht5nHz3nZmHQ
w1YUpXJDzljrFwrY5j9iLv76OQpUm0iMICUDfvEQh7q4OqugXpxgUMUJrtixjpw/XpL/i7F1hkIQ
63kBZsPqjcO/YjDTStNVGoHiYvgUZWVgr/4WMFfteULathDbkbDoDQzdB4qZXCDYCrR1Rh2O7LGe
ri17FWLeAIRPBuZy6bl9WgYp6AzirYzOmFGx4ibcabEMRwXlL69xa3C4JHwcm+w0Ytpjq2QXfow0
15WCwmtyj5NTg1Ptjj8F2RFuoBu8BBVV0nLlbyik/xwpfJqF9Ybbq4S2WeU1ZPRdZ4fpZjWwZslk
6+ZVCyOZXb5+0ShU5d0asnmMSg+YbuxcsnH/ULz4g8ipRg0wLZjIO+oZTjXC6REzjC5cl1l3HIHw
hn11OHyDhD0xLAL7TduhjFF2wzKxk5xmMmWBDvsy+ph1I1/qtUDPsoLH7/zVDMHT2y/JwvgxJAVQ
YogYCEvLMa60lKA/OwIEnssBx/EMZsK+fjsyBFBkn7xPl3Td6/6wI0C9YXCmJtDR1m1twcSSd/OJ
KoShG6++Uh/NK3chygxv8qphMkBV3q0lK6yUJpGDsihg17yP/xrkIlO9/yhPu+kkF0X6nEJaB/Ip
FJOUCtBnLYA1n9QvDftlwkWYS6UV+Kng6zkHBXnu+aOcuq94ywU9Ko8KCDd5VSiJQBa+9tuZqapi
aFTyBn99s4OCB/Yh9m3/K8CjH2LZz0EDD8PMRMeB44Ga8opUZem7IgXWmjPwudz0S3rZfoqU+Jb4
E0CU/BOI9PkJKPVX741HR8FthmI+id6t09ohgMYaDZSWjfbtxw6aJragdKStRim9u9QeTGg+o+lW
SGo9c5kmofH0vafwEfKzMHG4Qb3pnry9lTeSufGI5ZS8QCuvFxF/tj+bemJaHUNV3Xm9DCwID6dC
qxve6JWhxoGSt9vTBxXFt38ohTXjmtSnfzf2UBuBXJG8uWThCX9iRLEJAhOYOd20ltNptL3rHrYp
v0RKJ8uw4k7e7nnk+zTMlr68wPBNUqDGnQsquEImJXJV5Iz35Jt2Ghqz1x9NQD+fKqYDB85a6Uif
vq8kIFpgfGCNZ9PxbQQcQnAelQXFx2qDFI6oACw+r9l64qTSyKJrdJJJq4GEsp+VNi/0DmobmnXm
MCAA0j3/uPfXKP0506K/mGsAwE7S5Vpcw+5SfB00aBaRApwk1FkkaUW+OwZPUkWCkBmV/VDLLbn2
MNkr75mURTQnE33aivg9FWLtDg5HhLU5fL3yWqM1Qg1C8PvINfq/7snoEE/RmZaEGQbhgYzJMBCh
DD9ZADBipGZVf5YOdNyt2KOBBeDhcB3Vsid1FMChK/cmyHkSbgC9skaTVSHsGOOD8H+dUpZxnK0i
Q0acMGFLMR0vd24etIR7d7+WZFgwpNZikZfY/pbak/mJa3lImL1OpBp9DG4s018CSaw+QWvijrBA
/JbmPK2oEN/+XV3C1aL+BBMbyJYCQy/2znAfrQxUYXAl/vTZECECCxIuZhNF12xckHKqmGVOzIYc
0oBNtrlGrOegqGi+bAwwKTQvkjo2CZ8WP9mS/8KW69wgTo5fMso1Qnv2NyCH3M8k+V/7RFnvEJBw
mYO7tdmF3Xa1BFoL6/qVxFdV2RSqAfX5Y83wtqyLX+6/rGMrKx28wl+s9ILduQ0F1EcuCI2hiueU
VXRADjaUTDzCOdEyAVNmW5o4xAxHTtVy4ypZtPQ4XtEIgR/Kg/kK/smn2eotEZZty0KeAts4P65Q
9qL2CA4rtV1S6jLeHZcySEDMyqbYJH3fMAV+7B/7rROwhWehXVPor91R0qLvepLT5cgWCn7KJWua
KGEupZdXJzXZKVpMKQE8HvXd9KDFQ47e/MVzxBKKFxHh4NL8NWBhhyjOswIM7UmkHugDxBKmvYXF
7P7bI3uitGhISDJajadwP//0gz3PH3JrDcvFZ/nC9YjYbaWlls1im1Sjzf2TfBd+wnyCnYrnuSd7
vFnJeW4UcpgH9uBHcy6rhKm2yheC7XDsr1Kk90wSTSiO9xB3yGNO5Wd7/Rvo7RwlhC7RkDrFnqmS
Upok3GZKzGnWXajx6gdQ3kulyCo8/FG9JKQzQoLJXQak6A+xoIBh892GCRcORYKtwD+gPYt5QYkI
feF1CtnBiHCL//MDMAGON+TGElZIQqvv5RHRyvsMARkBqjNE4wc8P4t+VyksjDOVS782sD6lJWZL
gOYnaWGxdlNC8wuC1nrba6Tlz+277nV9EBoahBPeuTYm6NkkBnJOTRI0mi3h0KbU+auEDEj+l/ju
dk+XEfiPEz0FzcUP83pAk6wiV71rs69S/ltN1fz8IDbAObiz4Ai3vamFB9eH3B7WsV7ZzbzGBPlt
Iw39lU+SiIOEb4yzty0f21e8jS+DmJaNOaRlrX7iOgDd17VUg8JpKMoS5x8mqJ5vbWdrXWzTYWcG
IOVDv/+aB9jm4Um6e57Q+qDOqWQrn1BJtk20MSHVFi2Na4HG/w54WIzEc4NOx4+8ZS9oeptUeC8Y
jhpct5vLmBF5cnpXIiVi+atctJ8CkVoPq1Ys2mcSElBRJIzcQDHD55rFiYT+AHl1BPVkGIPiKcf0
UrKdlDJc0thZUkE0WEAAkPtlouchZyMOwwK6odkqdfHP//+jJDoik5hmyLKXNhNS072NlWLxuQLv
uNf3dNeCunwO0CvMFE1UXcHveotG2ZRTBdHkQl361yIWjC9j5ZwwucRKSy1ACpd13Jle8dVKT8At
jwaJoT/3LWnwyJ1+/n2Ni2FF3ziEL7WgAyHAQvKPkU4WyP6RT/pa+9k0yPzyO3Q3FsyrZ/y3CR8d
xwiF47JfAqfX+T8cQft2lnbtyRQwK3XuX8FuKghJvyvAK9y52SJnstCVxBf6GaFFSAA/Myf4MTCt
Xay5nlw1MJscFRfqmxQYw2kxgmcfNiOZ12mOm3qzB8j5IHfyfecRw/K/m74Y0b+fOZh1n7TH5GQs
9AwSQTbLET5cOLMkpj8pVEKMb3IorZaV0myxu0HOolB7UfPHTF4Xs4ppQkrtiTH47Yr3kUZ5Ui39
yNxMZgRDi+32Tu4Pr6ud3oL1+rXRSwOLJUbjtuZUpllitHpLswb0Cgj0htwCEovAa2YlUfmugpZJ
6ZEcAqL5J4EG8JWbU5a5/fHmGeFKy8HmJNsP/GNMZ+GLNJZj3nIiCbtYWEGZUj7G3bgi1pG71r9U
m+tLbvdAYXWvxKeVB+pavF63E+yA7Jj41lxPddtcvMNA0psJXC5zPdj+zxHvCiijYcBfBNeMAL1Y
1dHAoR/hUcllqXxQLtstY9990s/4z8ZaR3z7jVk0kdJYto+3aXP3zc8UQ7yLTMP8ByrNCI91UoUV
ytUfD9yHvFxDqu4l1rysncujrMX06mRfiaY9p+l5efNsxp3XYAVjkU1jRKIbkDG61JJSkV0dZq+o
Zpd3xQyjfYMZgljBBPDqUnVOkJqXLxynHUMkZ7rklJGcXUlHcm1QlUB4lz9Ss6NqWGm7mPm1edEG
LBsdRJzEurPR/oDp+YIY3qMQ+JCXJKNiE/MTGu8KFmm9cJsX42WOaOTNgRnvgtUqC19k06pv7DML
+JvGunlnXJhqhqMWBzK6wcFZ6rFNU+qAnuQ88a9g4YyjOMeZQIwk2sYHXpQpF8F3s/rTjkywN0/r
cy7hKGqzf3uzBkvyXhbCTEElaWHu6M924uwIZuTyBOwoSy2G/x0S6sLPWD1aeFViAK2bTgUob5+y
PkBgUrhbDy2M7TJmaBW9QGBQdleMP4jHBHM0IPbBxYv0wCnziIe+LY27QGG/1qLzbZtxTPXV50rA
DT2jS47b0gDtTTqJY9aHBlaUN3tptIG2cb3BH6YLYz+fDWuTQfL6l8yGzil4p2FnTNyrykREJ1CY
wr5UUyjpRj2p6BjKJiTCVq7v4evTpT1LdLlNkWCQFGByRs+sjO6POqhAl2zLh/R8JA9lAz/h1aA7
dC+Jd4IwsYaWUfSi5/R97hwGSJclRxpH0dvmosInb2BFC0niFSpKT/Q5t2Pt8p8jjDl999HV4TDr
4Z/oo4C1UNXdR5bYMqp9/p1W1kte5wJGi2XJLm2l4Rve5cYLv3LJQgoxfnVSDoJTi58Slz91KNuM
jJKJuTdF97g1KULdg4nAx5QtTh1HApEYwEqA8kmzRj3HaHmrSQunabLBHenecUhFmKXXe78wb3P5
0jQWcAEL3Mj7Kng+l/HoNtypU0vXL+c1NXTFahDGNBmBGVmFoqJ1VnjcswtMKaoXh1D+ZfiyCMBA
1zY1qRbnx7YCsswj5sN9jIQJYK2NNxykNej9dj1Rz2OIA7JOric8bvpn+wK8fks8iR8SsIcYurft
sYnxUGcu8fg558tpNowOz3NAFORiXz6D4CXEgFPjuKj+6OcBfAo40nPvhuTL+ScK+23fOgR5K+9h
OzlB2dBQXlw0YPi4rBSRZJcqVzviK9zlqZdwiz4pBUA9vrPyWMzGgFa2U2Cx8OsJDu+ed9pOqfzI
+AyxWvZpuFH0f0aljV5nunK2Bcf3FLNLYyQgPmHgPj4pnHXhOiv02qiL/ySVh5ZdQxFIeYv3dWxk
2DLN9bjld56/p8PJcK1Ef2b+oSL51OIDNqUMX25vDsTGzgCHGChrO61NF3g1xRhuaOnykLAdlSjZ
jVh6C0LEVYZQMGcXWZnKStaHHaeTFov4nAxdrtFa/B6RqkOHOrHbJizq7wLKuW1Vbw+xHMGOYbOo
kqH2RSQ+xdxYz5b2yeLSUlxcoES7cRBuIMOTc8/86anrZr+9KnuDStesccB4UR8aGUX7JPSQNwLK
u9TMVgt+hf9Xzy9VpOfL+oqEysJsBP9ikAF8t+VRLDTJn4fPk/Arj+ZfOsWWxqrV2a66MwLFE8CZ
IyiyOw4UwzUTYGojaMjmkpbsxg86hl5YLZgXjW6kdqRDBLZrCbmrO0ANpet8Cd707T1flcQxOQDQ
kN4Xn+vB2kbwbvw8Vt7eLuxVTo5GlXJ0sWwZYHvxgYAfgxrXDF2awV76bRrCgGSaEvun0RVF4WTO
Z9fhgRctaJZAUfZnzRQvYV1XovG3ujNsvUcxU1Os4Kg1GrX79sps8L6M+Xqra42jGexwjqj1i/kP
1vwDNfXHgGoqfntMsxU2YmCGqV72uKBshwXsX5+vOnosckcbOXtsFG+Re+MGaQIyQsV0SJRKtGSq
qp2do7jhc8XpuxrFq2I/pzzeicdrs2Z9pbyVdsCggfM1m17db5/BNOTQFVjThuYE1cbYTYvW/HmW
FbpNZuwB55MAx6t8LXiOrDCugTIHfzrOsNBI+5C2UoM/b/EF2v+X0J+Tr7QG/rDyWrerD6htlICd
EQC7nu4FghIIt2r/OXr6XBOkq2Eu5rH+/9YkcUTchxAyF1IOdlPtDcUlCF+A3RvjMe4oZLK8n9iT
MzYfE9qSCZmstRv8+FgE/cf47San533+3QTQIM9QxxlG/vBXIcGkuPJeLTsQ/bhjab8QE19B59oH
hycgt/J8XiiU9YFADt3ZUu7mgRzedrwRVWUbRd4q1b4W7WCP+svMiVkd3l0JFuKI2yZELP/uuAc+
UrKhpSlg5e3wB9LI9uAvEV6LHocFz+3fNYvXyHqZxcCbXCs1O5P4p3tQPwvsl2ehZ3dMO/tbA8cm
YRdzBhCyJVqFWp78MRjdjoqA16NiWy+lTNcBJUly9MTiyi34xONZcUS9G3RtnrqUCuM5K64LotwZ
fR3OfTNy5dI2H0C+jPSVBy1FYjE8hZ5L4GTCqCKUFtl3Dac/Uh6X2A6sraZ5k0MhRmQX1/4HZQE4
jylafwVpv4sl5UMCTmA890Cn6QOlP9Y64PEPuYO8kMoZAOrGR7vj+tmVFPRUKpJNzqGGrxPgg7nE
gxWSewBWxm0i5c88tFx/6lzb27NrRoz4YaeX7TqMrNdhv5CtQzrzNO6RH/In84+ybSW3F6vqDQGA
1X9zf5/IxLpz7C0HN8ZpwSIgBsxmyqz05NcR6CHqkkMDiT0PSs8XLMBb7plAKYRj2BZOWiGIbGQk
HRzD3cE3QxjO9cZFSZ8ZXFoqU7l9Sg6ShF1kKGosqfPWTbi6pa2H4keeulSX52gdksQBazRUa0v3
UZol31Y2/V1KEHRwym5ncxnHN7MQd/PYhgucdsC007IItIESWuW4j0zVFzkCnV4nWB4xKfXu3N0d
dbAJ9zzNUptJnZcc1yB5RSROyKmuHD1mVWHrUivYo0sdjvXVF7JwqlwhG+PeC21Tw3sjA02pgWn3
Rbrgz1jfMaliRHzX2i99e9wsKYRDcGCVuPj9MOnm8jI1A9TgJkeNKuHQgiZX5syFwrMViskQKCfy
/hFEbr/UTF5K2fkY5Bc0mxbVddSof13KvtdLOa+Bp5l1DupL8O5d27Q/FnkoRAXGD/UUg75p3JJh
orqnwSH6hQgLRNEi3pDpeJsrD8QfwTTRb0LSNLUa2QP28Kw2k/lslj80zIJAJ4UwYSdc9qb5OTPK
u062xafGIOdQzd0SkTHbhTWrM7ccMrJeCJQ/W4ZYI3Kub/Jrhd5MH1effhz/KQsAy1GeUN7Rei7O
UBS78eQq01mLgcVtbw3bLMQClhZeu3P5xRcEx1Qn0G7P7c0/1LVa4H/dF6abJxg4DlRATdTknaFZ
VdloFD8M5ug07XNq4zTGPwuSSt+YjHN97Jyf1VBwlcnU8GmmtMRdmc3hlo+jo8WjqZjmJhQ1RDvj
9wBuBUvS/jJ8hjc4b19gB/QaAGD+UTsvyaJQLDP+GZVcaqNBFlnwbgvfw7xaVWKOAJ5ITVJoLXQ8
CYy724EUpdnNwYLqXCRv6C3g8nmLYlLKoivOmTwbN4xXoDtPROL2CLPoUSmHQvebmvLXR1Feyhm7
h0IlQGzXF4O2NA/LEmrgQ96YEwP4++tTcEnk7pobL78iByM+JHMtiYer7T9M6zb5oxD4Ez7O9v37
LcqeQPCM/557ixcMvnSsKCHnp3yiTvf49Mo9kqMoih3Rrex73bW50JfZvG9PueafXOkmY6nQ4jZO
SqFnAhJAg+Hfe9GCN6bbadXDwnjtoVmMdIUXw68/TBsuYiUmUVPXmNz6QZZNqQTEDK4CGfWVpT3s
TxI0Y6KO6sPproZt7hf7o/VDBM3JbP70ldebu8HwTNRiUowgag/9eqekyL8AzDoRk1ohb/GAwcqj
NuTRj1LE3uVH8AbVxbLkIguuQk084NpwXIheFc2N5K1kgSKC49y6XSIof7rGOZIqZqRGP2gyoOVg
gNbziZz2EJoy1F/vpNLqrRRuo6Sv8lUPBXo9z7uLz8IlcPhrfvMcQhitE6cg8wRvvP1QKtg4xcda
of7StpTYCEyarcfFv9OeYqe7NqN50fqHNRMI+sw1Yr9cjtbA+MZXpJjUVRi8yk/c3/HxH94zs2Nx
NVpu5hNb/t5CTvv9cwSHIodbUJwwWwao6u6PaKCJP8drUyWAGIf9P6b6p77gcLXmmPo9EYy+nu7o
MfWVwVs1VWUT3/ng38x52bCnzSlt4BWRLARV+vRJDN/AIQnZIb6p0ik6OfT8Oxx/EGB8Mq22N3Qq
DV4ImEaDW/FhRJy6CetHdjiJ8A6YHQxlRSyZ3YftUF/1qXPxY4JZWvpweLIeKq99itubXC8bJup9
7smQrLoLa6RWCuVwragARrgAE/1MrUzfAIR9ETxZxYU5o5Fz/xGkAkHqZRVai9mWSsHxSgi3dNq6
HdPC1GYczCM0HNGkdV79ocIeznm+ZNL+rBUw/apdcI1UOAHhMUg1w8+nUz6B4bhtBGXT4TGU91W/
k95nd4KdQKbCwcDWG0L5Kwg3D/xqA2QPdxB2O34m/kWoMR6HUdck7k4thi2JBOq3Dek2L7PLdrph
gk8HEoOFZmFvQnrkzyurzU8kb0f9xJHzXe8HzZw904acAPCY2g83St4zCBr7/chi9LlrkCdLiTYU
JSmyJ+DBfmKMWSwmpXu8ACxVMgkPIhvhzlESkgsLl6gejwrOBIW4U5NuJSoq2qZ3YbCVsPpjB3u4
qBPRQBwhcKZD7xR1qPgVhmYuP77e0Xa6lPgBKJEsZhdjqcVHD965fdRtHJPOqfyVndeNEaAppAsw
fFyxgDFmQCs/FFD+iefJQN1nj85qrU9mJ/vOQDGUjrb5p/KA8/NhvOMeQbi8978PJCC6Cm1E0gVS
sgB5ucnpfEybHjfdARdftTK2hOzb9QKAq9F+4FKgXZW0/Zb4LSaxRxus1MVAtG5FWxRjl5V4tZcH
UCDKWqwVL53L8e4wWlouUoJJKvJCNlrCrjTwn3VCt6mmtsR3Dwwb6Ebj5NbN7WYwoxKDnWRun/Ak
ErpVMMADEvxN4EXsa0ujK8VPWLP2XDHzdmFavzxFIUt3Df/WCwml5PmBzrmWWaGNyIJQNRpOEJ3f
62rn/6N4j2JI4DoBFRXKlymzPs3GM6/tkVCKHOCoXsk1XjBInvHwzq1fbhVXem0fN30oiyRUcoeF
mFFasNJUsgCCUlpP1PNI+WXiuSvlLl+IEDa/w+/DYA50w1bY9LrXR3CXE2kVHXCg7/kKYGCxQQ7L
kmOYHQOnK14mq7kn6otp+euAERO/hC0SMkg+Pg3Db4B7ZpIodOnJogYdlhXYr+6Q4NtifciDUD3d
ZIV2m9ptKQ5j+GMt5f9ss1oEnboReymO+Wxwg4TOLGaAfmTkOL+Chpj+z0cNu2RkIxRUIfoibrOV
7BeYrepcRCxWhzvKPAuiDdW3TnB1zML7YO1xOYQqPObwqu+DqMiwDRF99Uz2ACgq551X05a8PzDW
AcMwp6UZjKXN9oOl2jzK1xQEL+Im+da4I0Tl1FgsM0oNLI9UHEd1+KAQidDbc/lWFgqbCfw/mHRT
eldDHDzpnAJfcYd8eztK4xnTY5+0kY/U88cIKPEUj2RKOnc448rVC5d6NXau/c22ShpBk2o7m5kh
LodJmsVY2u0sMCzR23Gf8nEl2rlT4T/+K35QqIUnDuNhqq2GNlg+5Teslmf/1LS7OuTMZZF3UVVV
JrH0rK2kd3O0sulpe8azchjyFadfqa2BushuiFAHrnXN0Hn8ALn+VQ3Qy1GRT/471qXjPiM7kjvz
HlR7cqsrOg4ltHICG1CQBxwY8WsFOOJtAD24ZbftQskkCYbmNByVhW/NRSxt2AwulLgMcMib9qQL
fO7/X96B0wUXNdBJiI5lpS6N7cPpdLymfmnQUMni0xHOjDaG1hafNBPrLMWkMCNvBV6saZhrC4Ob
OZnIRkF64nk0EevLJ4qfXeJRsTw1+T3awS9jkOq+6ek8oqpukVA+V1etb04hgPExgxVMb4BE2SrS
1d6TIHgspikmBHvu8S+XRN0s0fZez1A92xSMSyhXKVDngx4DNx9O3eTOM474bbZRZ2n2/HNNhCZF
dLxe1NA1KtaoFFznaOtmO+iEAwQKV3G4D+Fb4sBk5JSV8w0QppFzKnlR1o0ye01gcsx5fgrgZHxI
rJX0MuUiA3aI57QBoj1qbRUkbee/p0KBlb8cCMohVJLRZO4IxG0wGsZIncSGV+Jlm+PlGOSqswnB
+0+q/Eu9fDVjDIU7n9W2KwfZQfJthhsr346QA+np4FFwdd0K3TXSVuJWCxqtdTbkQaQAvwMX0sWZ
5K4z245tR42heQTXszcRw7Vld1cNFtlErRBzJVeY2q3OQ5p13Oy8tgp1XptldvEpi0aPwlEgJR9k
/z/pzQsJWxDs8UNNO/d7oIuS0KomDduXn3Dx/D4MAMEXDcbzEqahNAO+FgUJ+MJ4ipGu6+39u0op
UMS+b9AOoc2+c743Q8n+eemYi/TWntx/cgUX/GYENteBtAOEOSbuIsnWfqjMSoT4VZe3R1BOfwDL
LNsY9N+X7c9nA9HlJ2b11BWt0gKWWo6JcyfO1MecyZJ7zdkJ+J5rW2myW1qQBS/82lpzmidNm4YT
8EkLmuYwqW/WhLaUoaYLB0SjWWuQrGsSL/5Mk0wS655hnIshJmQ78SxGZdIZR5NCwtn/lPs6mSqf
cziHuLzjM64L0DO6SPeRbT7h4rGjepdmni2T1KNChNgZKqIZiq0Pqeai42da7UPKEmE+CfJjqbIK
2MpSgcB7VlaFsQnpx12lGylJ2w+SAe3D8Qm7dPmsNZHsReCM78uamlQEe2t+ADnGGq0lE5kCJtIL
2oBWLOJH6kW7ctnGsY4xwAoj/0tBJwYDYK122TNQz5ZmpIl1JQwoJEvOCOKRQinetnoBnuqqLHpW
pvhSmVLmpuobAu0ereYc06i7gmTSrINJAI1XbfBGnDooKOqveB3qDgWM67bDqY3vRqKmAaVt8vih
mTjbSxZ6UX4aZjbNmlcFsE8wD7UNhZ//2w4dlACMwUfssfLr+8AjxN9B9fNbaQPXkdKVyVOdBB4c
R3FOg3A5HU2AjXf178HBC7k3E/vVzo4OPE06m8iTtoSiD3x6M9jtB7n7iprJdLnLUljdLGNXKiSK
hM4Zu0P68xIGdP6GIlb5e60brg9ztbLVXT/+MQDsszhc9ARc3GIPprZIEDEqURIJR/pgCEMAkyVB
k9x5vo5Wk/x+cHVEyHJjeuhln6btZhiKokmoJog6nej+aSevHxwMRPTrKoXpAoAkdEmomXX/7gd3
CEwTaRmtPDzPjfNNFTC+oA4iviqOtH0cgDRhiF6rluPMExIqkmHkVmSw3/+ftKMsL0HlCYbRmlK9
eX5Odw1A4Qn50/Y5T86sqFKYfWm9r1K1pkWEpkAlnZws6pP0dACJEOozzxuqCPg6Q4x1yf/yCr/D
nA3GahJwuupvyJiDBLok90WpZS1YmrG/WVFJVURfLoUCinz/c3Xn1ossxvkyIA/tPgD8x7JjMWPx
NioJntuOox9ZgV1Pu1Kv5v5Ch335mwpLLnKxmvSqFreUAAuqYUUxntxlUz5xjG4K3Ano1THFbgrL
hdiCnRcJQxSnb9Lxro5LzX36uJqYkOs/frrNMBfVRWuano1ER1cRxY/y196hNgCWMp7RyFSMwmgl
YnZkYqx6R4QYDdd/kdFq0zRxhzf/7WB+RzKgbVQQufIOlyi0AQRvmbA/i2f+bAPmuU/suoQxFHMM
/CUAaKAB/zf1d9N+ounbtbltTL42m16zF6wuvpQbS75wgc4aa068+4Vooiy9M10KvJlppHlB4CLm
UK/YDS4gx0yFaPwljQRFOSbVA6r+B1cRt3tTpaRTrhzw7asU6586VI9a2HZJ95xRkv43/WHtdFnU
7a+AFDya5ALgr2K3AzgOEDXdVoXP4222g0Dlo0YuFd5wYJvU4UTFtMHHWWx3GbeIJQkYLb+sajYH
sFbqazlaubI8ChqDB4Z1H82TGHKiC4Ygw6Ajpd/BsDgWe7d2UdgLlpH6EBU7H9PXr/gSUKEQQazC
8mHw6aDbTC1aA9l4wqSrLncxjslzt7x/5+1I2qSVYsKPd/V4yQwTna+svt0ilsVVZAOajYiABrgj
pH8WaPW0tq/Nmq9VoZ85Ebn9ZnZ6T30EA9i6UR33dT7IS0LyEiJkHxnyiUX0eCeiH1olezq+57Bf
4U1+oYSopPQm63KqO75vDZSF+hTwbfRX2ElXHTxfQ3pvn4B7PeDM3WKFdzlLTe1pICJJNxh1YG65
khyrooQOplM3UTkw4egY0uLbfFdXWt4Qebq9KLSzqbDvehDEOa82xtTw+UOXnFuhjx0UX+57pSvd
kDgbjmtROgsprHynhPIgvjKMWGR8Y8DkB7blLyHQIXlVfW76BvVAEjtQxHkW5HecCuCxiyy6NVPn
T4qk0m479OK2PnbU5UWAYhVvgQShPYF8kLUuBf83bNCOc3WnHojUMuWdQvOYwo4/xuQ9PQnlRKiH
uWqs2BRotfsLXsOC7funtT18hOFVspXxGw4bME1GxA3G4S7xMbrIE841cuLrK2JqhTTIzDkndsjd
aZNTV70EBP0KxNoa4ob7oo4cq6hJE9lOteYxCiHxiXwHroM4qXuXrQ++liqYa3kONks8KCc04TMW
XY0IBbz52HtAATSqnPkoEwn8w2weveH4nfOX5COHPtFzdgMMGZJw9OaAqA3wj4fbzRIQ9duPniPC
AT8qj1oeN8OPpqyvbkuY6HoHUWxg3JUzCFz78tKVuUuzK4jvZuH1O8EB/kVzEnkfhlYBbVrhzLG1
bLnAwrVMvxf/s2/f4t+/RvMI9U6IYt0du0iAEsegDRAoy7IA0hk2Phz56hOcH29j6Hb8JZKmLi+j
d0U9dQJH7dptN/7epsHBu4V4Z/tGwfoY02f7VnIfCqk88tne0bHjD1pxp359v4diAwMkz+dVFXSW
YIvlXmZ8/yYoy6g82KrorsswwQZhMXoKMgptoL/8+WW6h9gPdqkEfax1EjMLpBsrMQ1y+y25aNbY
mK5LTjFyvuuWo8zlotmzWYpL5N2D6wDBiII7RbiAVHSfRyAtDONHQL6y8Sv+YyfrRlOkK2okkmBM
Bw+ohXQmqqMDAazTx8HpO+2xb0CFVzLafTLWqN2Q2idNsGnxjdD1Gckf3eK0aqtpx4M9ItqvWZpu
/ddD4wT+ZQIpDfSmo3W2XLCsBWbBobUITSfhLe5prgytFnG9P1vbRP6FtF/nvoJVqa/hf3gkiZSY
tpdq+NAtNCFoO3iWLQAfwfjq5hmbpdPM221Yeu/4hDHVOJiewpVBz6uzeZJjwDaOKjXkth+WT8qj
qQCjjyEVOE+fKWAB5LKyBb2EBCzl8IEf3qjJ2gIeMy3UHWymEJV+Gv6dJebjla2aTd7lpw92mXzP
t5EjrS1FosN57L19qByZ97rITLuFRSe46EnX/7GIUlcTQErukxfJiuLVZ/CaMGoLnxc+4uLJeGfl
Q7QGj4xVUj61zKl10CafMiBc0MFfp4dtS9S3jzX6XdsPesoHQOPR4IUgwm5xCJA3Bm4XD0qBKVZE
BrRyIWysUSKIDtKj0QX5R3cowFuV2zffjPk1J19UieAVOt91PIAIQDd5J4DirczulBB2idTkgQOo
BrbvrwIRFQxx5sAfGSyKRT8yS4SZ2HkY5pqSPqkT6qhgeNU9xtf2jO+9NYjedu4kkDIvqaDdWxpF
f9N3cEgWAItKFDprS+VTxvwyETMf1eu/aXPBucah+54qJeJPRl/UME6NSZ3S0u/tvcV7qKjRshKU
FHYvyG0n7f4PHpJADFPPDak+DtAx3WT7OtllMrJZlak2XCq7HxCioay3vBDd++a2sanNKl83ICVt
n00L5gkHVM4bbCG0iyPSFX0TfWOjeVQDSyEDOEXv7Yy+kflIij6OTnT75V95UV2mGyNNGGDeyFTf
YULanv8+4h5NRw6mug07jixYOGGqKS35yuf1lCdDpk88KTXd6Y4jztG8FPfuU4EeO3xNm36cBzj7
mVjHR72rWlN9VfZfO8uwPHM0se7bpdiyI+CWNOkVaec1OxQFEzf7SRtmbsMegk5lcWKyO5VFUMyF
BFGCQrapl2v29iA3TsGP2rW8JLSJt3lng2J2f46ksfNoapjvH/jz/+UcSJL8fGD/iXSfRc85Gnl1
pvDO9vgJEnGWPTasUffWOTiAMsQkA2obUbErijcMPR2DrqiKKStTYOU4iDa26Dpm+NgcdahWNFi6
G318Mv8CkkCQeSsvx0Im41gQXYJWkpGA6EKlCq1kTutnWHNM+Jf4v+K9PUbPaHXcc10rX6Dv/vZI
wXLNyF8XA2dSHZPIWZ3LqjD0oEHI+6TkZTvxvBDbbHLOgVK+6yCePXFxx3gNBa7sXPR/LlIlUdEK
nQphX1MOtLedAjs/Rmj159fFVUmjBjwrj8Ophy2w13BK8YCA+xfujk5wUMSikYlQuqVPjXgjAj/0
+kINYxAvIIWknLLWiBhI1U6gzzdJp1cBZi7R8E8oPKQn6RCQJtMw1VKSc/KWvSsPqgtZNHoK7eU4
gH6DVPB8p4jTD7bA7JuDsDHkSXJKXlEjkW4dQwZNDOm9KrNxdYA95TzrW8pBL44ChlsyNm64kL/Q
udICukIYqa4UQUP+yVj0JA5Ciw01GTUthReR2ysv0vgZssgqb6eedqolmGwb/vGNZkHtCmAJ5ozH
zutxSclueMN+0VajQxivJ1lEKB6Yd6WusfovruPflceKa0vK4bA0WxMEl62x8Ef44cDl+g1i6j+g
2ZG0e1hnbPsmsbY4+3X0wVi2eY6yCSZx2bwzv6m3Xx0SqgiiKQw/rnVGw4+4pHnbsmcJ26DzOE0R
EJ0VqK68HRnX6Nzpv+4W+9YXoHIWJpw+Fh19F7yYR+h9vogiSQT/g4wnbTxjGz+NxiQQWXvYO/oK
2ulKI3fNmWXTCETJ8XovzDxkfBybKaZgTvpQt28eiDagKxMRnm2/mo+cFjhZ9jWfiGgxftVB6Dnx
2F4QE0mtptzyZVJHFWLvRGS+7qu7cmPa1zYIb4PznuijBQLBCO0Br8nSZFNEK1evTuWlLoeALhkV
jSY+JkWMwn7bJTBsqL7iT0e8H3ksKHKChv65DPb+j83igWbG2u3XTgXb64UePNU+lVaGNqJtcLzI
h9LT/b5l0zQ9AIuXtOYzXe3idLmtMeD6mIfhHtBROthTVVBaeZdN2VXIiEg3Y4TC42K177eXn00E
HRVIyaz3gpiJjoC42oy0Xnjh+cE7OLed9DkPZh0Qq9ckZn+EnDXjX9p5xcNi85LFcnuJYQmlJLNC
sv6U075PlB5rchpfu1+f7+Svxhb5Ct5/X0vpxBBg6pv49WZidvts0drOZwgmVUh1S9w1qLqI500f
+5NG9vXyVKNLJGGxJ+Np6Lvp98aLBS8PKnkZDvCKW0PobN7okL840U4YjrrwsgXaX8krJj+Khoba
s99du36Zzu3odEfDU/s8PXb/yS7fHdrZGLdgyHx7pjhq7HdZ8hAmwSzENE3PF2Q5Aq13KH2Z48MK
0rE5Y0/m4uRmP8+hAYXVNf0sJO7YF17fV3tz8s/9ggWBn24biVERSz7oIcFUp+G4AusJDGv+uN3m
bxV6lA/MyUWQafv+Ejr1SzZBb3tutT/gDtRQipJXwfzMBwFHvuvIGZq+s/K/dPJlcXJHVQU9f1Bk
vBcOYxdtOP/5GC0l2VezhsDdiLhaSi42a3odgNJAsDIi+qLimaF3qdSQIsKjYZhflffKhbxFh7mG
LXsuzLHJDbWIObZZIOquSlsgbVnXPQzQmM2gLvFMObB4crjsOXmwI74wTZQXL41aW2K8xb336qv0
0/lQo3WZaEuwXLzyLaAU4VHiFED2N9eQWDi1gA9D8rVK47GYwt4s1IK/bLUpk2GesfZWSnznVg6C
WxBBIUuLKszgSiCgK2jaYTvMTCqJJ5Gx4lRRsSC2gUV405tBrvioEWnDEFmhlKuXkMOrfQoQb9pV
wBcefTp9WYE1jogWw3syX9pc2SkDZe7paZxEB1i4RvzEZ+Qy0QQ794xPfdQ5OqwsmMcho7WgB9ho
Qz79ISnRys28h0qtrrrqRp5EpY7NEfvvYwRHLAme0OABwkkYyi4IgcA7VFn6Ff7ERRSJvqR4RZh+
s3SQW8O1F1ii8koi13V6OV/DzjYTLjQNUtQT7VVswrtCJ0U9mx6L5NJYcpLp4XGcJKNhVrvhb7Ho
i+D4/PzJTIKMhcj69WjOSjwUejCPwrF61c8jWOnVtKkXU6X/kSZYx6iLknuMfAOrTgJHwY7hFwB8
MaNViAKfPOsJ/feKMpl62gFtKIvDOiALFvrtoW5EgAjG2JYEBeJ4AjDNOz1ulOgQ9GIt3pCPxgfI
Ouy0jLZAaRh/vhie7CjBuzM/NPAkC4PAdicmUTDDTXTXroaEq3pHS6/rlW+i/ZbMChWFtIakkrkq
rQuknkbORtb7i86AP6inTkjouq5M5GsnEbdoajLZDRXtEe7if4OaJ72/QvgK7bvLGS+yDCgsrXJv
WCB5k985TJdrfAeeeGYuTArwsF5z6f3yMGurYZqTSqGrtu0/I69GVgCGhaUuLyl5/iuL0pPJwK4e
C9FxEDij8HOhrx64xADJ+Zkyo+aqzhIWBo/Md9mTueeoHBjZBODbcxrNIGV5ITxM/iZWQBpOdxbh
qbkfCCLUXAG26ttmBhUwFrQYn2p9+lU7OtH09lFkKKjJTHdlbc2glDxISSwSG0td1WcoNN/VzfrL
j6SDaLG+88G9Pi4DXXfx+MEXDtQ03y7zLm1uEMMa+Duf4G4gqdyyS1OfeQBcPw5PjKYINSebIDj8
ccG8Cab1Y92qCTiwckqRso7RZfDg0ICFgurXg+YdBQ1wn4t5briVlmyEJbYduwbSjYo0W+mgmkQA
Z9Ap+Rs8jVq/SJA10hI7wcVyqOztD2oqdOeC32Odlh9vJZkbo4YrQCDlZ/FGVOmMs5BBA+2/molv
MLvW6e7+Y+q6wie+8ZonKEDGdpfwTfZM0WC9t6lP4L0qMXrF8/pqbj7z2ZLaCKCocG8oWGhUY1Am
3Q52/6/HVP31UBfvIY9O8yEh5YK95g9YGviXLCRgve9J0h/xWcRorw7Voki8X0O3ukrGCjjEpRgd
abE3aQquWHpsb4LNwpXXMmQi1hQ5uMVULFfbPmTuroyrwWPF8o6XhwU8tWFatCg/wBFeZPZuHzSo
y9VJuqagfOwwWzC0vvwIXCKskMAU0QFNjTVim/GEu0wlshRuHxbax0MsLTRvM5CUXbVrHG16BYFn
N9Q4+5BX3vB0rsdDgNcm22jak/ZvmVFLHshiYiOfVDKX4iVIdkYjPJSpq4Z5w14cbRylw6qdfeJC
VXdyzFr79Zzc+DQHafszDJBb8vAaOmm5DvujwVk7hwHssCBKzfSxCbhxprf6IRy53UjpcXrGpLIR
ZWdEFUdgJWvDzUD2Mxs2RNBxxvwx//4ZdO2J+Tbkg7t5g1dZIaAVzMwEBFEBh11JXzfZUyZb0uJ8
eyfyAoS9xZ+uginpoC0AwgHpizZUGg4c0oHxb9SuaDMIt1k4gbS4nDLXQB5MB1QdCzuVhIuaXfyl
Vg6EsIrIF1Lfo+U/HxvlMe6XCK9vVYUp6djL0ek50BSl1DIo/aOix/f8ExGbNoQ6Epj4phnW5Vst
RKdysk7Tz8ToFNWD5cNTGldZ96fVvhvawP6TT7+lKod6TLjH3/hprvvfAexmRRZp7h/ASpNpiGKO
EfEZIutr9YFlfLy/iTxBnm7KSLHgKZD32MUxl5ZGDE4u8EgNjm1Vbn+GepOnt8alarsvOJb7ogPF
X/mlVnZoSE54hNx3isOYFk7IbfLeaUQnBBd7JjLy8DyPp/KUV9MYXNkLJHdwEswglYcGKcMizCx4
FugeY5SoVkSusAtwyTxXjQ5BEJYMNA3ylqqwqYbVx5vxsFCGZxcrCN06aOi8B07G0amIymBoU6dy
9QqrJKfyz4/XJ3cANEW+kMpbV7P3GvK1hYmHBWgryIfcy74Kx9P6ABQ04i1VVVuAe0+me1lZyVq7
nxjCNxXl99KOK6Ee+ssAVV14xYLRJQCe2bH5Cwd+ZnEGAMzgWFtGr0utC16JOv05tmJbmzkcnbES
r61beGmTn7pTKiIWQBhGsG4+jPlKscTDqrSqgbxKUDBoBkRYnz1zTVcnkxxDMdRI4h7bx7uXYhGU
HN+A+7ZjpWi9+U/wXAbq5vqwPo18GQdFfQc5igtrHRSvtixeInX/lY2f0WGNle5vuUbUwZspzbMG
c4NJGk+LZQNWVaiYzMcE+QtLXIsdfCJCa0Q7k2C3hutsff3HBFCNbEjGrbgwKc5NZKrpCFTIVL9s
5inZ+PJhitZezLfYXUr+pBppubsuvqVo19czwcqYM6L4rR1CWvjfD4Y7RGPkikpUvkiCCIkLyMWR
RjfFscDRIcyDjC5fzFrDyj1cy5rK0iDrBujRcM1P1jkcfzKPQty+jxuIR0A2jnlifxm3z4zBQHPg
1gL7q0w19HIefn2OIEJP5fX5SVvzEFoh+z2M2aPWsUWDtHy62Swh5ByNy67zCkOMVUldw6Q+pa0U
HVN1Lwzzs69CqWp5AMQl3mARxL8XcmFTkIgH6F7HCThlemWzJkO8F+s1AxJZUwFe//WPEec3g93B
fSkVvurQyEKYNjeN/ZQXUCJbkxeZA584RG6r2ugxvzFJus4gzJolW0cxJMetxSW5JKDJO3Y/BoiB
l3OutfTSmVTk3xGFSOq5T33+QpSZfUtRhz0DFgbIAbbEmDlBOZPYfqVBniCRrioygvrleH72BUT9
5nydyewbJPad6xkPYaaf8+UagA8ggfxy/PLSol3AnE1qgFUEnqSYLSypLgYKzQoqjsJQKzPAZG7G
8F99lt7BsZDeMi4XeYh7ngKCL2jwlrCSqlKngqgILRB1sbs8miq268o9FpMfqpmLWU04/Kqrb+f5
JQjpFhAjv8USDTIsVH6vOc1PnVcaJpYLe/NO7vz/4UNUxFeG7lNJ/z1lfZuZwMu6jjIxFExvca9H
t1i/3iIvL8G0omo7FROmQNzUNfw1ctEuhXml09FleKhGQgbUeyh90PKIKNbPqhsTZclXRXF949vN
Ifmg/nRYqrOWc25y1ZY72pSGjarDGF35VPh3uG8QUePsM1c6AMND+M/zOdRqtaLATgByup3MchGb
1kk+C8xyEP4E9pfgLOto4rt421AbFkH/RwLr4yiDc1SPDVgGq6+vRSoXssVCnHuo+5Ap+xGgsK3L
ckWWaCYERED4NMsQUHskSChwWK/1AssvrItHTaZ+E3K+wZdiC7VYqMTMT2hCy+49tpV1yrW/XJ0b
uQNEphS+t96vRBAqTgR21/2cpJFc+dODMm4J6AF2DojH2l6oXix1YNRCBGpvo5vJwQXUatDddGRr
pTvRXEDqZKNFIMn4LT7OY+ZnR63mHP/iu5z1gqXh5FD0dquVvOMa1VBLrgMbikKv9uBQGOpuD4a8
SwyuWfYUJqXiq2clfcU+m/HKZBKFJvIOgMN46V+v1c7xiwpkrJISG1wrGtOsSbdIbJXiAbKoT0Sw
EqVC/BotGqzR5mK/Wfc4o1fDzKCCfPZbPsKRaTc2ElXPLtgeXSf8Xs0bVtoMndCzEBmJWdRuPVWs
/8jClnpYBtg7VeilQ7q4UfvlfUMsKckbH1qrAlYZgXqrEMQLJJHb0aMDJfYFgZpcM9wGIfqiJT1x
Iq8IdsfW5tp9NaFQ7aD6MnvmVnw8o6kbDqNPxyzcBdci/A9TKGsVN6pdqwNBKlyHkoeY+WW07T+F
yDQSsmVlsdCHuOPzAyZ8uTExEGEQU+hAi+ymD6SCIJFKD0iEXMguw4W1eO/7Lmsb/xRp3z2eFkZS
a0niegz+Zj3Lpcl23EdGP/Rmf0q7T5ShM5B84E5Umj67jsiudBTObvPxgRfDR/rkiDctJyotaNh3
eZHdn+kv2CBH5vajew3xLmRR92WbR63apDtNGs50wfRd7Ou4WqhHkW/UhOfkPhve5QBtL/ULmfrD
+sNMU/4TI6NuW5D67z1rgDQhyj1RT6JNQk3FW0l/hqA8/Hz5sWCXCfp7g/MRGqXmzQQmEhctjHdZ
r0fywNvZqogYJIJDn69w3O/Lg/m5Op+lH+vAQjerOsDyq2slY1+vPBYbCI4jCPyyXgzZBNSNYuhU
KmtdwkrgcfSu9SyrX5cz72cOlMm3KbGqD3sgjBZU1NZCdulwUSvxOqix4ak8Q+v9rNwN4isK3a+U
SUELQyiTLLonXPt1k8wHIo0hlTNFrnNlTHiVZbL5iIulsSfj37Py4ONFSfY8NqcFFWDtFzYtvXTN
NSPCeQrbQshk4/bqrrYCGfV/2YnYjp1JQ0WRLWnpXbWehShDDkEqwC9DTh8IHIzQtHi+AOM+iny1
AdqdDNYhPuUW943KOUcZ8SUBN5SEoivSZaPMGlXFtNwemc+fH+FL4ZOV9oXU1NQTWDXmH6QhtMOD
pWKllFP8XorNwUSw8PlJ3DiweAxNQtPh9hw/83+eO6AEiZSw/JT4+o31VNO0FpTYGINZyzEn4Fzq
KFaqw6IhdCtaheBeDFaKVQ4lpW3vmIlr03mq+UQOugwCQmL86wFxfaoRMEgjC5jlZ7aZKxgoAG0s
YVVJ9fje8jtgCwWfQv/lpEshyn9DYzeISXNaRjP23T2RwQ+fdX2uOatN4XpIaLehRei/9ficD5Rx
XYhu17o2yEijkbUjTCyRQexGn0vb3Rnhnf/2FEKM88HKD9G04hLn8kL/wAvhDTeKINkKzUS6SGd/
UC+BQRy/mqJTfPPR5u1p4/b0BZyZAwXgQ7Nr78PknXZfc7Jf100LEeHtWZLz+77ZhZKAojuqpgli
aWNcbi5N4opoyAxTsXpvkWlbHQn8yT56Ucg3G0bsFqMrlz6UyErtnFBTdYFw9L276hvBwUMhNaqe
NsFwdpsjk45y7Gxu7wgTffIi73y/WF3Fv+xNLNqJuPN4ctzGzVq1KBKyMSjv5KRL/mKX1qwJugtK
YTby8X+MPv20QC0S5zhMhOYpgj3Hrzf1NkX6DqVPKt5IrKJ7xs8aITLW2wRQgLd/9OyeWm0/2MK2
yZO9pKtLc96PtxYDJsVAPCK9RKjhkTLSWhbM16m04TjWsEBPN9M3jGk5lL08nr8pTTcBTf4SDRSq
a0IOt8HwwJkPNXTfNvqKLUZqtfSuGNkDT30WS/Cl701ip4IAWJ4F7TXLc/ym+soTsfheTUt37+1u
bmQtxlTmM2264R4OhJ/waqYy107UQwvX32W/LdCaPGWnV/xLk6372+M5aiO7K7JeI4Hl5xoQsS+F
+Jnej/3qZYTL+pad1Coa26Bn/Mxc0yPLnV74E4D+9MGvQVJdEMnznooUC8hF1914FzdHQ4fkwmJ7
LQ6WLPxN4jZAC1eq0WpW6KAAIa+A0FOCnkWmamFYNsxV++SnCvoWarmcheFVrTC5ZGVZlEQxFrCI
RU9tkVvlVEUKuT/dNs/H2bWHtoajJ/G7LmDxjkGpWpjK1eRiZICDrEjzoDnvVX2jWPJVP0qAwX9I
TwCxWpOqMUn23oh/8Z0e7jTnOvCuA2KUurwLAWQtoq3wRt/sVB6dAIVNyRoVJoM69CD4jNnhfvcS
jqwZhiWhRW9q3vWmPme33AD3ll4xIn7I0R51Mz1VU7awJm6GzLmaQHU1fPJJfybLIbMIXx+Xung4
4f9Jb5pMZT2Y4Gt0CV93OJy1nEfiS+Z6xYe1IW9I3qrxdLxV2ez7lOcmF8xfhR04E7pB8q3rbdJf
/9hzRUdPLXKPUfYRAUKYrdw9tOEkc91UwqwR2fUVWBscjfkVei+jaumK+k4aKxd7Vd/pwI3DczPQ
D2EfB67hDRNvFjfd2ICPVJnTvhub5O/C8AFp3AXubf/ZxGVNJ6ks9QnumdWBjb9yxwlzl0i2IAc9
bpDsXRrfKKTY8TBl1iGftd2EUCxL5FZ24uyVQzI95OcaMgPDK68EDQTttQPxrqbY+VDiedke4I5C
3njbclG1Ye3SlfqCP/XRrxaZbnO3829E13BiX3Zgj3QqO6QyBFX6nE47oaEhzt33bi5wrGYknw1N
TsXm9WgFh0shQVBtxrC3seFEoPGbzzNaxvc2073XeijscSfAoJgYDXa3GkqcgDLx/UmDIxfglLyp
c/2KqGRGgHe3vvDBZ5Eehg5FpmYoAayeZ3XfPNN0vzvcXbQU6eS3BjuS+sfWxD5V2YgE3QqMFaBx
I8XVzDS5q3DGzL3+Wj23/F0qXZ2yMUzTzs5dRyuWJ/9DVl5hnoNykHZl/geVw/K+BQGJ7WMiUPQ1
3Ay7u9vjpyD8qfRxud0KlIe8OjDr3rD1lauI3LxRuc9ei4PplsGUgEqeL/12TniseZY8rPo6xKk2
G9vhNs0n7REP0qw2jKWTlH+FDA38A4Qel1b2hsRK8GKUZDzqfNSZDhPN6lhV8OufSrLiauqKiVYZ
r15KyYqUtXsgZvvg5HFmhmFG7vahsn932GiL7rX/cxoEeKzBELI5EfMLpkIL30lIaOHQVvx6upy7
8E3zKnu7ZpNMVs1shGjURzImDTH7MZaehlpGUGyuZgbGnd3FWkcJEHAwirMxziG/LgnREPFwZu2I
Qx4IxMNAzggAOUs0SyAPNI7Ss5uUz8Pi6bKUF2C6IV4IhWDzgd4TRMcZtGIw8Mkb6suDbIMehe8Y
XUmplkdxnKnoEMzNQZzoigrN6UV3uod1/GXYM6Nn8vg6UpXyAXaK+t7adTGXHn3OaTH2nLy83U6k
oEPFzARi17eVV9AHzD0n89il/T8tUkr8Wr/7EH59klzF1K8SqlI95EfUMgpLDwDyrOkdH4IYw3fR
P7Utdypc1V/grUluRZvEEtN2VK/iV7Jg/nIQyCbgqDHPEMgt5wXpNg7FN5FQcvFBsjVrEP9tSmRJ
509SQurfU15Ie90o+5gI5QgP3UezowIlBLx1QkgLDhST2DQqoH5CNy+5XTfst6ElsCvEAzTj+CI3
hHPoSGgYcuwiDG10n55N2pmPWXZqbznXNKV0aSDwJO3jXT5xFBSQeW+yT+VqHKz2q+KiXkQam3JS
SuonsvsD/MBUTq3kJHJCi/QAFQefFmNvo2mu0sEJvKG48u60kwu0LwGE9tkNEpSeC0sHlCo38H1p
zSz2GdrMd2ZhV5mmckvi1DBIrbkjd+ZBvP1VpsKLr2rD8iZYPdTw14hgaJEPtCrb+FOeglmp1C15
ic+Buuqa6z2RW9+JzkIVGIXSiBssIrPL/qIAhl3yJPc7PTkEbdkp7GdCZWwjn2463xYmDpQhWY5Y
AoTUM798nWCh5oWkPJXZp9f+
`protect end_protected
