`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RdHTLNptwuCrJ2ZVArWQQpbEow/3o3R4migBrOwX9qQ21gPdDLYDmmabPxFHVoJ5ghd3pe+3OcJC
VOGpWgIQMg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CMihs0YJEa5oTzyWspOz4PCc/pS5yHo/qgJTdyD9xvpuRonRww4bWZPADpUxGNMe/x7oybI7X3sX
2J2wc8WKpBDJsxs2jp1DB3pFCKVN9V+slitIYPXp0O2Ov6zZWgNA8Si4ayBovoItGw/qz39+go15
mHzaZ2lMsPezP4FyFPU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J7cWW/FR0QlbaLGnBcJbUIB7dDp92u4ieFHNfKwmV3RgkxvuDhY+BHVuoFTVvFeSO1lcCowEMTy0
LpHisTUjR1PcTNLygWvoZ+AVTKzQEH2nGlEQKhb10oNTdPZcK8EwgdBfgKjpdGVQEzKbZxp9rvsW
mXDYTlKCFnqjeegsvskasG8yKkPXMkrMHlURvQ5a/ORXIKWSWyFl/UOWrm/mOanPLkvII4Zq22cv
MIW0+WyIIinOS5oOsOB9cLgcIPdxempM1+vgMUgmtF1joJZf2P54PKZhYVBrzlxC3E+mGdKGHU28
NohsjowDI33l0GH8iHkAwCKpmOb1Ir9OX7ZTGg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fya4SyDzn1pFlwwWWtWi7gYOmYohVRReX3xPePEFR9Ft8RybjmUUPFpBEvyNhthGtq8ywX4WZYjg
oeHZUPonCWBLOC0dognGHO1Pejdy96CX7mSlUrahE5/NwlLi7Fo3W8vlszu0KNywlBjLDwra+m4w
jTs5sc7iTwjAbK0K/94=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b0qRoBptqX5HK4Ug8CpMH8HmcaeAFtqEwIeB60jDKRDjkuwNi6scRl2HvZ2aIUHVu9/aCfo826hp
8DiZbq2n7m8+gxDFyv2QGLrkkZ2mVZJ/8aIBbb9qk5FbVFYkBGvPRLzWbGvum6G6wIUZZxQgAzNc
/iU6dkhtwKdbwq34R4HUGOBUJfpry7ZQcS967DF2eej8R0BF72DoTZi08PAxK2pVFZdOnSb54ii/
4CJus93DzxiiDKI0A3GHqoGFBAxfDNE47fbpRFsiRUgUj60Y4zZAnojN4RSxCtTp9+M994vWTKRO
B7JA9o9SGYrxaCe6eGxBj9K8YjNDJHutFplUPw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12080)
`protect data_block
WL4qRE6DlkmEuXocW83Yewit/66QY6hmQVHjkGztdczn8ncwQ51o+HOTumQ6kI4KBEAIxiznKFLo
wx9up2Itk+No4iSr8PeMJlF61+BBke3COWkuSI5xSbKfSZqOSOh7l59Qlla4q8C6zOCFpiTlxkQN
DpN6c1gHvel1C+jaOPZpiVO75IUw2lTavv+Ss5H44gYvLluWrkK6BJ9muFmXtikN+1Sh0Oiii8yr
GDNhR6y6U8s6T/2+vZcvXNI29xcupv6b/bdnsYwLXiM8QosWOIZKfReyTaO0ScLu8ArP3eGtMlc1
jgWPEhBs/TzBwmP0Ipz1dwkSfF3y34axOlewbFEbH7I4ZwwqEvXSmoPvGwZewHAd3ypan8Tnk3ib
QcSCUfNvU1GLN0Jr7vhm0ooJZpz3rk6Yxtju0WZQivuv0CnayNw7Otyd0rg62IgGsLbZCTUxqoXT
pjndw3ngjmfovxn80hv6/MJqjfdopNAMs2+gXrd7+52mRRoQYD9+KKDOdxC0qp4csWhmjbVW4563
Tx++82DwZmvVzq4H/wjj1GEsD7srd/VGLnctsL6zSTjH+/Ad6vsHQ2B/TI0ub+23ixZZznZPCDFP
q4QkbnMbrzPsuYeY67aeGeKt4wCadgvg/q0qKd7xYrtzprVh+7rUYw5f0H4AOuc6Wy0haacDI7GF
9HhlD7fI1aGLExtQaBgLeEztnDVVGDibARC3iKl3eLsfalVVKSMbscsJQLpzZaw07j4wrdBYBhPF
BN/BV0sW56hZJuZtle0Xlqizr3IZGdeW50dmpOVBIyWJKkcVfBIjbvB/5mS9ETR7EkrDqofOgsXH
j60j+3UMrzXB+eUmLmkjXgwVHmAAQjUx9McOhHAn+sqmihdQhB497p70qC1xEZPpvNsCkKBCaScd
cDMonst05inKFVm4yB6L0TnsfUOUkJMQSj/2d9cG1muDaHQPpazLmkYbgpRGPeGbceoW4x9nkXcD
dyeQWf5yTNXwgO8ZabB4C8dKgIx+nohVy1wNMz+MVtNPVUfIxfUJg1VUwcCuTKGt/SKyaCEkvemo
y+lLY39xVac5VcM2X8AfllFSKnusnvHaoz1RTjq6bzILLVFkxnzfcqJuGmyTykVHCzEhajSdBWdP
6lUE+HbVWqH/F5NqwBrZOCWhPY5VxnOprnX/6McYM7y/vV7FbE7RIHQO0Ltg1y7E42iZiDevZp5n
EFcqjfcCo+hMFQlN6ICkEk5dJFHBUUaFkeKBb6lXahEssqa+CA3Md4ot+VQJL778k0TvBvAlZXUQ
RthGf2uzknkfBvpZN+RSvjssB46f8ysZnwM48Rp3EPhEHnoClwyXmVrYg9MLBAikDNTaIh+Q+IWw
Sbw08FuMJFuIYZ+9D5hy3a3slcBwnNg/j6IEBIaRwEXBUHYjs2o0ENK9x939DAEp6VR0510BBcwv
4lcv0+DrmOInSwOeW6b7wvfPuhhnHE/8fmb8F4dVvYB+5dLRSe7kS+fW98q1kPLl70aMVpQt0TED
ErW9H3URAEzefx8gxBLFCvE7x2Wh4TWIdTxg8SRxa/xy9LvHW51//QBH5E6VyTqOD2NsmPTxFybV
gnubGs/ch+V33j0i4i3lF/shTA98xAUpZvntndJOwpmx2YqrzPuhXxT/l3S4JQzBqeWb3s0g4xmX
kLYIJwHNSRLyoJKxCGkx9g3mF1KoL4hB1VUuXqHdbJ+3Wey0uYBPzZsH3qfd9N6glC6Cto59d9L1
1SZNMOVLsm9bGMXo2EMrH0juoRv5aGocNE92W8MpxNxOkl/1ZAf8phfnz8WkUDObWUynq2llcXw2
IHLTE87jb3d9NG5He350vWgziHd6Sz5L7XbiPdT3465Px/3q/+T1i7mLSak6qOoTlE/kp+6EOVxo
Bh5gyXTVA0HebhKZfPyelS2S5bRd7oFaWnLcWrbaUJOpJ74elKhQLNLk9Lf5ZhpUhdJupqbwdr87
FkkG4JjMjoWiYhh90MKLJzs5FwBDEr11TpAtHwB6o4G4Ln/se7vHqaxofkQEax6P8rFBNKLMFwhb
dP07wr9hu4ViGTyZ1yg9DDMmG+c1PdyYkpABeGxdsyNSbuX6Lp0+TPmb1MBGty3UYAAnoiTzUdy6
XffClT612P5nkI1M1hMB8K6DKpLwLtr7UsNxY2dOxRzcowdGGWTTErc4h/eX9K8s8ZCHSIBMYysw
JXc/qkLE5m4c807yDwDEtNaSWsENNcWlbEU0f4XBGUun8QbA4YG6wm8drk8JN9/cIwKHFRX4J4gx
kgzXByW3GEKNTBjj52+zWk/RQd/4tr3YIi6ssLXKwqPDX+VtTq55OVnImbj04nP2W0xWJj23lDLU
ayzmfWCF3fRqMk2biQASlx6xpd0VMrliZE8c/S2dOylhrjTnf4vvs+J9DuE1swSFfk4o4nepkfhy
f8e1zXQV16g5yJH3MpKmWKfXj8Ie6RBF7JO8kIyJdCKRhCihdLWZr1U+xtymoSu6MMbbsTbOn+2Q
d2M8KfQnzM2h8XPrmr/CtleNKv3OS2Y4liv92aSLqsKA9vMqS5jZl4Lum1uBQHNjea650v8R0m3I
YL939qsqCswpgD6zYrlpn6CuCoDxmlvrVFZz2Q3G3dVYxB7+TM9Rz6AbKo6/toawdLq2yggsTlvQ
TlhpMwVRO+XqvvfGa+nngay9YdxRRWV16J1DkyfoMWlPOq6ffstnp+wRDRfkuUOuuMae8YnH5aeg
4kaarJo2FlmEMgXfOkh8QiKyUcJvzSgNyLykJ0aGaJGU0UtmB0RI8luZEefj0Mi3pK6FhTHMWCaL
A7ZFnZs8OTIiW41Qrhzdbypriqk51eJuu79ttazPZV77ipGHzVhFgqCfCTZtXlP1VvVrq/FEKXpy
jG2qBGr7us7a/yinLmiorP1PyjR7O+WHhID1exwl6NLJmuAP0+0cDDQnQFxiWdv+Z5wL3PfxYjXQ
k88DqJXJdBPbXH5gQ6vpe36OdYzuRmUEz+iQ6MmBJMnOzZ8WAvEixeOyx00GiBmVIBLiVuaVPyXG
oL0+OseiexORQ/R3oNlJdqctPhvU5TBs2mL6/rsvFZPItgVlbpYuD55Uhy3fkmg4DIgoDSgKEsPF
659tD1dHKqEzNMP26873bYbS9nDkviFk53S+XCTCK3NfKCk5Y9Jj9MNQLemyr4WlL/2BYlc9ituH
fDJTgCfiGLSi+IIu955si4qeO1HlnCYL4UoRP/xiR8hLfmwTy29g+6N4mnk8+Np9bN1pPlQ7hMu4
fY8baKeWwAJxSlQh7UQJ/cYsEoF64VnI7gimNvQQPuBRBTGIHlCgxsn7pwzJrnlGR/rTPfjz+wAi
2Mb4Hk6TWlhQ6Nrqh+q7Hb23aujub8/Sr+EGCorCJbOPUY8lH1Ng6vzk4ex9ngwooPMB+bHK6tg7
v91bmpghq2oZYOAFNJQ+uavOSY4A8NeDunjLg4ke37qXwbJrLJXaW3dJyXTl57JYAiqLv3lm36n+
+J3nplFswbuV20t3tjN2znk+OpFg1Tt3xcpm7kx70CJMyEx1Hhqt8YSVRs2i0/f7x1w5z98sYMa6
1jaSravECRMisELW3+yjw4Z4RXOudOQASvpUyBMo5Rx0gjCmKQK4OogOr6D9SDeVI0EcMKILr2tB
P3/gPTk62gqQoEexcLBUGnWcGw22WfMb1/m7p2/LHD8UUwdPaBOePszDtgkHaEpq59lfObmIsxpZ
5hBB1J6sQjDnHUvkaOrKAoCcuuCIb/U7tSRKqDDG/dQ5REO1Drq5n3oFD4DrKjpcbP8DY+PsJLXv
IYFWYllP3i6EwVFyzuLvu6ap0i5bO3SphtXCnTS8WN7lq0kQUhaddwmJ7ZlrMAyPulyKl6wutnRG
rlpFtTfpG6FashaqGUsfy7VbwnRm4bn9AX1WjzCBpkGsTA+pmkvhdKImkpMyZOUiMEmUqX81wxKZ
0OoImqpNA5fTZAGOXBb4VYxb/lMVmehek0J8qdqQFfsvh6lrRH539iWP24wNnrH26Ec6YlApHntD
5OVwsvRB+1XRJ3IxhpzfFKhNjM2tw7iwryDvGsDS/zwwBm6bwCS3NmjD7wLB+gXPXvr8krRYSX8x
35RunYxyPtlpDxtgpFDW9GsuQ39G18oy4ltkrkkY9x3MZunzYA+gzJ8QV/7W5y5ZfdBUvxKwKqTv
ZAilg8bF+O2kt3bK0yoVO3i4izbe6kggP9LDvJ2LgC5hWPZOCsYSFeL4AAMfN54MvzP7us1EdFIK
Je7HSUSyMkdNAAUcjoldcuFgdPiKcGq774w4izR/hiHudXnUG3F7BB8EqfJQm8V/V7D58C5cL2fM
xTgUvBGoNkrO4FO85pWAKN2Sn3e6CMTLkv/rkNIFqcsZBgOJqT11BjjUFHBm2sAWC76cDWWLb0lp
7EZyqYfqf/32UvWrZ3rRcLRHTog3ZxgYsnlfXb4A9Jihr7d8nKTIkEh9i7pdyGIlt3yODJcVW6pa
0GcIRi2lFF+1fH8Nyl8N/O9or9rO9It34zmYlruZvI7WB4lnoxd4j0Z9oGuyU3vdC1KK67ql5nSq
UcO4r/0B9LLBZTZufT+7PA/w0X2/YxMfQx8pCsVygbJqUsomzSMKo0YPaJ4pPHnlJB7Y/7RkIRgx
9J9zkO5Rppz6SZ2Z4k4UY3N/M1jUnZf0h2sguZb2dvBl9uoXlI3PRX4sGq75XNyZtru/uXA/T9PR
nkqGFY3mZ+b32eFJMCn+YcpoZ6PseylYgxxln7sJrIiWVDhh7Hdw1p/hlqMXl9g1Zm0+PfwEy1uq
cn/LArHBjIHzfnLSgl6ptNXIH+dF0XUz6CvcQfzdtsquf0dqb9o62cxlXQwCY5w+BkZ2O5gBRKod
hIv2tSwow3+AE9u82Hxo/0ay5bzm008XF+rco9IZbgDJpeeWahPEruSnscdxf9p82bKTYD3GVePx
Ul43LNfTv3rFbJqsEpIZk/TKdzeTrMxIw6sr5OZuByWW88ffOJoqlYcRPmsUICvg2ExDYv3y5KA6
xif9OpmKYMCApKL4ngdsfGG7WDLklejJB0A0ZRuyoi/Wbl81eefrUGU2N/H7ix0gL1/8KpQE595Z
BlfWFopk2a0dGWtBNp0OXTewoxYtmlW15A99t7byIbU0yrlwoS0+QnvF0ZsViH8L7FuZjEOWVdbO
YAj+x8fOWccJ6XbRBboAn7yhyAEAt6Z7KNRGdAG4238aRjhpA5ZpX7tRIQZBoyU2y6j3fKyslpZZ
4zU+jCitTxcrkKlNQCLQiS8PoOM4Vmor+VJPd+lm0r7jjY9Lt6R5IQvTedswQHarxvwMW/xnX19i
S0RMkSAsv2M0yPSNGetd43StiD5HHl+IOfZ3c/5DD26BZAiTSNlX5oRUCNbRV0LhHMwUkAiYCNkD
AMWjl0jV5Q1E8YukTodMh/YyYE/FT6ixB+ULjuEDOHCp0P/4YAasqtI6DqzSwn7VPWkqQDv3h5y+
bkbQYq7cKdihm3zFqhSy8HcjaPPyPS4w9jbsMM/BecSj6bAJ1tEqLk4MBT7F0Kczlnif7pb6h7Ze
HTbHLFwdNFX039tPaplVFxitfuE2HsFlQtWnUK9J6WOA7PIfn8giFXTSQuZqKX4+gOaAlPUxs2bY
BgAjqg6hk4w0wgKp0q9/sh5ROvS3M3qLmLzR2MWTJtS8XmnnFfjqvl94NUjdOe+Uh1K0YlN5QdHl
XPWV6B9iyIBmYCDy3H+sFBxrRRwUrAt9wwDo90Y0dAISnLNKmiYSOaBlQHyj91xISIlaMRHPKc8f
eZeGWMd+YSLWG+GLGKGx7SQFXzNDU1+WIQ1mdV7evUDcA/1aES/idZS1JwFuKJLYJhgymUhM6aiu
lZ9fjLMM+oK9U9eborBJIsN6Uvntn7otdF/S8Wyf6H6W/ucHCAg07Q03aVliNBGAFDm85RST/vB8
iRDRKKLjBCx5aMRtkPwTtz8b9Faz6GRRWV3bgFUDG5a/YQG+y1m8UVixrsNsEOa2j8P6ZOb6cI0I
ztuatLSrWRU3r1kiqXcPF3P4OXnDb9zU/pB2BuRxYq1NO0PzbYdFkyIWJySRfE8wk3Xqi1/skqT9
/1ClXM/X/Pwzh/ik86AzQBmv7059lIj75kFZwFVUjp8aEDZTpIj+uGOeYuKMXfPjC/VSfpX4JLRO
lSpJTePYsY8ebIPvIbtnIf1RZDs+I8uvxXmkgJAD7Z0LuLyqAkQTrrcy2cLWG+ywI1Iik1tSo81u
fkuq9Ryznu2qXbki/ej4gB6SB7I3Luv7IuABDj61QfUBibnbp+M1C4GOOa5D0A4+0vpgR+9KJvF6
4nVS/hN4aN1KOmv+WycXHatc5dV50aOzIfPbL0EuRCoqP/yFlmGJoFM21SM8KB8X9JlyHhjF6MuJ
UTNfvgkmR/KvsJkE5EGBYafyOZKcpt+Lgo6i1gg0jaEbmNlt7TA5nJWKjY4SlKSBWwDR9UWDKHab
Pcoe36+JxttY0Q6vWTawHy/KzA2Ru9pm5Vv+PHO3WiHY2IvlWL0rocsJZC/NgM4q3+Yj/WRA8bYB
RJJ8FKyokN7PN0UbsxUiPLyepXaDXoXgLp8cBsmBDmglABXiWkWIrQ9MkDUmrh1qtr1Pce8r0DlE
mrZEGijUZD3RLF3V4zGVIxTdZ6xCeKGUfnFrp/RNa8qp7l/+Go+ExN5uhfjlDr4S+VJZxRycV65g
Zak3/KJln7CB6PU97jKmPClbzUzrM5sqC6Xwh1F3VV5zwO80SasnB9t/ahFXKvDfMFEfA8hO7/1J
YQf+S6RhAbiUKBKsFilYT2kpq5bBJ4zmMWbf4EZI9owaEV9TPsebvh/dG5nZ0nPP0J0J//a+5iCI
yz19PtjUnRL2Jt/NHDdWS4t4JEIcSvbPCO1Ih5q28lmwMNY6swSb6/b6QR02XcEAMH7yKJdUz93G
rCgVtu+GasYh1sZVrNWbur33NCy7pT/qL/16kmlAWtarHMdzEqmQSlOI68TQCw8xA1juHy1BWfI+
Y/75XV1H+5r352mMdYj+eBqH/bKKj2+xIBNgLMECq5Ys21VPqZA18SDlOZ48cZ0tHPkeeRwX6wTk
VEp+sVoQTO9M43WgrqXvIDvqguUetPDIGh6iF76mox+6LLmtOg+4jCs96IClZjQ2qWdrhbSWwtiN
YNN2zCuy5cSyAMixkzlGoNNXHtOvESyznnP9QrLSur1WJ4vWZkHv6NWgLmxKDqji1PPNj1RAktUw
n/x5CvfxjDW1bjkwGkha0+mBJdjBSkiwtsw+hyFXrHkNGYutAuXUUFiaC3eyD/sw4uBZ/b7L7XMb
fwsfo7FffkXoZxJV0IAbl3G4nKvt2a+PocbXSGbG/pl+S+og+0hZGSGUinpPcHKjEFc9idRL/gM6
hr5KzxcWYqs9TzL/jkwLmzYniyWAu3Goy1bw26IN1giD2Atwo+tIsKmYckBhTQv9gzJ8xrNnTslm
SMjNMsupQCM/bSUCiNQSfkVSX7p24XXysTQ5mZQzufzF+pm0VMOjfeVmjRKXjAiLZ9+v3bqx5P4M
vGZJGn6LgkXkQWrumL3e2zAJOI/VCO/myHG3c4IJMwIMReBx3KCZ8Fvg0x9BEm3s+C4cfoBWx24/
t96xlxShiv2rN0EO5LFbjhSnY3kh2RVAGUmfml26GRf9wreX8qyKxMowHcKkZrDu9oJ1JwOOtk/K
oRwa5cA6fYYX0EMpFqIMKOdpolPRlthWpzw0/oH7v8ShuyDuC/w4keBZZ3LE2v10KagtSNZbpZZ6
wALsHbBiEJczCbRkxJUsrj44mSP2XsC4Z2PXjaq6VUn5f3bUYL7wr4wNswCg5247VOeW+YZiSWx3
2DmCf7h7XHmiznyVTEPNsMJ9bnwM948l1Ot0TY58HD7BoqZxf7Y9H1H9gpf3UN8vOg6MGKlTETUw
c452U6mpCANaDA6ZXXtc/0LWB0vJEcUU5M95k3oIBh4RdzbM2MDqodVkl7rU2F0VlijJxeiXta1f
bBseWI4KkX34q66q6Esl56dlPC3hCjEZv+GKrhX1jyDV7eVQtbhqK8hyQKkhteDTsy85T7BG/y3a
KwwpA0vMAc0GhuNnVl6tBjXRqsQLa+FsuxCoGlYkTBw+fcp37PqizJ7Z9+mYmxp7ckar+NrtQptm
NOEXuKZFBbnn9vTXqEIzUxUkDtB0RYFbLjrm3Ms9GmScMp1dpsMWi4lRrkT5QduSFTl4x7IlE97z
ZjCOP4rfzRFf9jVaody4XEx50qiJcscJds2TBTyfCHYeDdtNQl5Osy8WODeUZgHdVa2Ytr+RgPsl
mIKjc8uGehHu6UnCOQEVQ/ltjbSyMQBJimdl4sBtnuaF+uncqX/f0GFv9nr9EDilnkon3y6MCQg7
tsVP3cAaud5f8eJdRcCMAGRI+POhzaac/+6HzJ+BMscaLTFKUeCjwvSkGDWKPZNhQ1HgHobOornq
Wd1mX6ODwES0EnPmzPzQxjZ6/tyWcrpbpS53fVALRgewKRJXzwc/6O8z66nADrAUUdRiCvSR35Wn
ddPgpD0rtam+zJ2UOlubFT+iM2pie5fbDaoGb3+HdzH3Ek+6oCONX4587n1/gjouys75yEj38iDN
NiEcouGyNAjZ4N3qjcgm3yIJXCaYaOwPo9qx8Ya64OlS8+16lRrT9bDgFdT2tyY1LpoM8DrBsNFE
tISlFCj1kyP/sp/d+d7du98B3BPo3wSJyxrrNJqYpWc+A/DhQ/Ifw7J5UGIMK+BwyO/xr/BYOQVr
7CC2aWu2LjmK/4XxcBQVF+6fj9A/8R4asdGEbr9oxK5lYPWA4ljHg97XdznfJyHYbjkbokld+ND9
/i/r+s/2KJgyMt6HUCkuDxdZYSMtw0i5cLIrgOEahDGqEY+E9Q+TvkqyGMKewRBaakJXTW96HasB
CnO6YpuctV84A1AWyyWPw+t+3NDuM03XeZoAU+Y9AvMMVllvUo+ucCBu6vdJlVnvb2rOdN5NlA3e
asfVH3zkBDELzdlSQg7oUS2U+e4mTl019aZB5mOYfNEP0+HAOH58daAOFCJIQW4BZuyt9RTBMEeE
0KjNXhfjNoRv88jUy1F6HWjrvll0wpi2Gt8/uE5mwiF7hoD9rVO4pLPcxhRA24UeEsqIO9hVOE8p
7QfIEeG/WzYHCg75o/vAsQ0r3U8Giks/M7zq5IK8qQrxHWCOPwGJM/b3gqv42GUvDZ/IpuEbPQGj
0KWMrfThj02CKzPa10T5TNY0u1qEypANR/iNtd1fpZQFur747dMhslL3s6FdFMR5JqvFB5A/WYB4
TWH7jJbJE81ize1ieNgDEB6gX93ZbwZMCcN7wSkLiwpl2NWFqy3j21jJ+oLjDSMvpwgLJcxQ5XKH
EWWSY/I4rKmwWMrlGyAYgGBeLkHIN7yCO3p5PLQGJheWccLzXUKUdXVktX7ezlHhhInZyYhCMqPC
7/SbTkz8ak0G+K1K/MtcVGazRsreRIKKePR6Yu9737Po38uv1EZXs3Ia2AhZySrfrRR0Rwn3jP0t
3WjqmcRCxsUEJ3QIzkPTlCQ2RkjYW+6tGbSaqlFuof49ZfGXcmfY6liOsb8a8My3x8Vlxe//47hJ
mLdirjsAV/vF1Zoc9cu0JS5Rb7HzxiSlWYg6Duf67/ci02a9bZhk+kmUOl/06AtYc0t2MaZvSIQT
sS1EsD56OD4RTFPLjnzcIeY7QpXtfXR5oTmrN5GhsCL2SRaRGOGkxfDVMH9eJMGcDaq+zEiTetI0
MOMTnan8Vz9EvlBu3cubIVVzkDo/UQpChW7mQ1zMhouQWz58aTtzfeCDc/37jQ4/DfqsnweZrmNF
j+Yy6uERp8N42Upo4hxEEh4LHxWCYcSG47zoywLZJouUFbBJbOnZSBKfSkuZDDC1Vyp0DHo6NRHQ
NnC5fIAX4qFiMB9qPLvSYJYSfeEHmMm88vx6RWKDeioz15nma0EDWudmlim8T1VD1eOGGyhkrFBb
yfR1SLalAfEpnyDAePDwyy5bcKCVzjq5hPIQfm/9PW43GhN0hffAh/MCWQ1pI1TX6cZbhDXur55L
i39EHTtIqvWwAww0HnR0+wrHKnJ1lGXbHvlLXRrRwUNlKlzqCZrhty5cFXRt4SLV3cqknjFKL5bE
Tt7UQ51SDYj8t8vN1pQDxdEv1y9ScXfishuurK3foWn3/WxN2f74XjYbjNbCQHjdz9TofirAuTf0
EI1Tq+m8SFeJt4VEF9tNrsrmYW++nnS+R5KTlOExWXlaEFuIuo1mL2M6X9Ptxn1DIP65TevOTSlw
8KIceRqVg7vjjn8NYKd6mWzorJWuRgPc3himgnxPTnVK3tHMTDGqSqJBlDfUU2xsE7+BOVHCeWdL
XtKUN8bxhyFhLLDLrGAjQxrf0l8B16B25d8MzhcCRKMBaGyNe98lp53zOyFIYnIJexopjAMPblK4
3X3ODIowcxggP9OWFGukEPryzA0+mdzkhENMD8P1Q80upi0kdjUw0/FZpLpbHBtTQf527mVo+n9h
y5dt00pB6JR5CP4VTufWe0RadxJi0Yd0vEAmnPnz5Grkm+fTQq4DSZ2n0VFK6JZ27QlQvDl6b0r3
KIJcUgJ7pvjMrjfMaCFG0mON2X/n8uoPE0cE5p7mXcudnC463CY1CUianWcl6nxObXNt/8HwYGk/
w2kXlHC1mFAIfljaE7gbn284mwGiRxBMYPpk0eTEwaYfNa6wdDt7F8WzQthu2flZy6fCyEkfgdtA
43Ovdx2jv7go8kKg/p27bi9yEZb/wI9FpRqhwWSQ9QQDBcEafH5nYuCrQCgT07PUxzfkbWL2KiA0
0uOfN7oXzjnkG5jqnoyTm4uTCtK2mXF7/SAi0Wt2GB9oMqUZ2OJPv4oZPOR5w0b497wRCwm+CwQd
pH71qOUazyWUipHrpGDQqW/AcTHTM5AXoXfXzJqxx3IKbjNVMGEFkn/CCE7EIrMcYYgyGpuNrPa5
BaNbp/R3jgbpcr1Oscb6g5k9UrNy2xgDT7rqtzTmLBFJUs7lnanQ1+wulbBp5F/MPYkE/H8aKFhC
ie7Tg0d0wzzNw/JkuJ3zjisH2ErVz2WGobs4wFQedLz09wvxx3IB2xvbVobs+f2zdgxdtRh5vJep
oGvYRkJlux9r1wdhPpm4d6s8+02pkRQReS0v2prDALUbiS824gFlBAPpCFg+ZU2NGtOg48NEclN/
Xw9WtVD3GkIw9kN8E+aQZE6nBe7Os3iCdDzXKCI4sVvZBL1c/6IRQW8DgHweRYyELQNyPZx9lw3Y
/Lc1Zj5t2jw/7aF1SjHf6uKaa/xZVa70lNRwAu+M2GMdLdLEjcISyolBG4T21hV9c6n/rvkIdhRm
pimvoysFN/Cb5YvOiPUeKlTVE1Z311QbK9YYydAz0hBA8u4cSIesd4+aHxk/o9Mxm3Bwj0DQkjOF
VR1fSeYop722PkXuBALepgWR7VNaEDUoikcoW/b0l/b93VWWJXP/5Cc6uI+ywFbwAUSLsj0ggtUJ
LvbmqTXfHjjFIbJvuHnTexBWh/uHg80uECZywrg86eqQHChOWj4Oqi5srS7vNUqsinSPWC9zZO9F
nhixsEnqZEvb/UOJEE7gZ68rFFSSc6A6P25C89rthqxy9DsKaMTuwMZWCupRNo842hRNdcpqo2Js
coBozwq6qSILY0GvU+h9T/uR75JTZQJwf0zduEg084MJvC/QY3kQOwoXYKIiWVXvqD2fCA3D2vbm
9j3R1Tg+deZRUliQOFEvD+J6Tq+sXucbDeMSTXmUjUgKLbu/Dhj60OrYpyTreG9AEFCqg9/za3jA
ubs4xUsxJeMULCSoQMpSVARYXcNtB78CtW3yTzG2QtHTV60kz5vaQymMk1t3ArgTN2UlFT2xsvhK
NIApjo1NcWd6eFlgTdcLKwq4cCMo35GNSvjsdx1rCsnOEnbiE1wd/SAaPiRngwr+4gR5+aoC3KS7
GR+3Gda4nGGraw6Vf7/gv4mlGQNjVVbfolzXTWR5fmPKi+3UUr3mGKCh0p/TcVEjnhcG8iTW1cK3
h0levl/YUj7KlytR3VsQnlfoF/2r5CwxPkOglP6xFq6/pmEXBH4WgBZF8jXgkBK1eNudKOeE0uTn
sELQiGGGw5MB/9pfFloD6uFCAMzIhPy6GEm39veYxYU120kV/xfReFRmgXDU5IGzmPIw3GR5dt8H
bMkMwGwm4hbGfZjCKigC8QmaA1gW91AfzcGE5Fh2hNL5eBAQjCFrICRjyxjgp51Fhceki5ailKWa
9eat1YTaaNqzVAj/REcU85sDpec4BVEP5aHQDruiaqNR28/lHup9dTSQAk/Mk6pY409dYbIw/ua6
YZp/25BbVvDNoqj0C2QhXlpR94wn3hvxUrXCAlh5a3xur9KhHTxnmkpwN8ats793GGXgan1fbcSR
3laifSA7tu65gP8qdHvhP1cxbDe/cFMAOb5gWbOr46GOcLiVmg7x61AwN2Jy9N8TsT/V73lPcwSs
bmUmBBMzmMKwcSk/wK8OzO1u0OwkYPsN7Y08l/jl43KEvG1b7l1COLOQTYNuO/5GXS+jXzD3IN4y
/Gn6LJwrwM2zA6wyNR/Bv2+R+Jet2fzCXN8g9l/67hKUNsvRHYYqpGuy/C1oIZscORobOcOv6JHJ
0rKI0F8nXSOA1q4Jx2pkaGGIh/TOL3A3P7zcFrd2TFiCBjlbinm1h48OVU6ZWU5+I9H/k4heelLM
FdKGZZ9emfL7as77ToJT7JfNQwJZk31ksAitKGOAe+3ucUDdWLLvaeHNKanavPW/knFzaGFiIQyk
ta36Dvbqx7zvsK/KS7BJTVSLh2Ssp2G69ANqV8k9A0lGK2DFFYNF/wPJ0BMR/zqRgf66wfFQsneo
TyHucCIXe/uFYi4Z1gnRHJ4ohHVo4ycTZkbKC5VTWnvOKKuT7JGAOfGXc2nRDhynzjXkpjJcSakL
5Za6IEfwFOZ2mm1DUlBUsYoJO2tPVTJuy8Zq7YMIc8+HWnmESANleHxPpjQuTMDgmBaMw1HU4woJ
Ba0Jq1ulE1zEmDyWVwkGR6d2jgd6aVv+Dv5jHqtNGeJ3AXWFoqAOVF8HQQxFSZFxcwu0VVlXArZR
fTDq1fsbzqT80MOFSVUi2wZifHQMa6PsIhRqLv7ab0XjIlUIcwgJKOd6Odzt6siDAFiexRkD2oGN
Sg1aAiN3BzfWwNrzYmEpK3wVeWgA+iplU3pQp76jkFQewqON+r6/wj1PR2qyr0MGKsOLlxD7SKLP
1ReeW50X5YOPXJxrCKpyoS8IKNcJcAlHGXbxk19+qnR9Qq0oEqqbRjOgFlRMLsZOjThx8BpgJx6y
vOxrYJJeWtzDnzqdlx5Wvphr0+K3/+WtxwPrnvvv5VsE11P6B1j6ndjvZ7jiVxjxTrn0+brRGTfA
pPwRQ4CLltbgJDRxRyMT/akLEamfJGe88llRh3xvyw9eydSYXadackDmE5zNy5NDhXETjD0SFLvn
HkFwlKgt6gtUcwA9PvlvUGyl17KiqOiPiciPZgwsXaHlV3VwOlQ6I6F+dLAmNMFhseD0imr0KhBN
eBiurkhW/InC63FvZIuyb0kB5prf1TQ0TCq9FTEzUQQ5uEd0fbCWjjr5bZmTBz5GHigry4zpeXJO
3hmqPVWT8xBMQNxEHoi8UNdp68xmmifuyt/et2Ms/wnCSY4AXbRw2XNYdtJ13591RkGfSkO6+JdZ
oxNS5h4s+PnQnbJMXLSi7W+fHYOSAK6Zl2cH9SBhiAwGvmXflWoOnU9MI7R6AzrVZEjzINdP4paF
jhYwxEOxsU58tWOuf7Yv3P350C486hY0kGrshVa3HlmYFIFe+6C0kFndXszSOsMcrbGGuELaRLJP
vIv0Qg7Hssu2i4jYs2GYFWh+hSHvFi0X1rl1wEkPeQLtYc8rTDphcs9un1gWDEB8C/1heuUnm8IW
gI9+x3EBOdFhaysTYCyvAUMFNPFJRge0Cwpm+g4WrSq8vx1M7EJcRqCgt2Ow1CP6mNhCe8rVKBSV
zCtiay21BXCqLlXmF1/8uxmvrnphWObFzvK9XqWdmkGzfHny9txTnYRCesDs5DTIkUV5yRQW+se0
aUdHh8YUK/JKcnDk2w0l0Eme91TjTYSE3IyvTCUuLX76rOsCii90B5L1r9WSLwcGjuAlDYmAxBiH
mqcmdyzGD2nPa93ZH19Ys+acgdwiSPNx7bBMVOzCs38p/JX59nshdRXw+nLqWuCxSK5YwxcOXdW9
YnbBofRap18DbVjjhYEXHZRsxYEXE2BQtBSNajEVgNQfhf57xx49sCQ8BMsV2758viCil1r0Hmkm
I/QR61J82FLhbTP/PZ/MU6CPPva0WdL1ZzuzomcvjjB7Thuwm86G0aTFncYjPJnTx6C86/Z1TTwP
AcKxqQVuqe66Zwus2dD9z/VfXl2hIgg1iG/smwdF/dvPyDhaWgmTCwiUrHqjsLeXsFFLdPI+q667
TusAFBtQj7Fulmdr1fKvuM/pDy+m/MVDnvMpncIrGXVLtH0TlsV2Uur2jinCs9OKwHa4FB5j2vsV
tluiLYm3yVgWBkgGVqAyzMmQdyrvgsGDiT8ct9W6ZpBSfgI0vcFTutNwRaxqMvnU966zW9Ihqb2j
EloXDFjibgZe27quaKJtzEK17Kw9fchrT1+EzbrQbJ3rDrxjCLIXyzp0Le/OvP+OFvHpfqm1vZGO
10BFrSDdhb7FvYVLF/oySKC1ijJy6IFQna48s0rM2yr5wwaMFuXsviVnNi4wGlkfnXCY6qshXPKh
L8f+70Bv5FgLk6fqKvnpoX9PWKUVirOjMwQGwYZ6mTrOU/f0TmbaakW357lE1L8K17czmn/GVVTI
mQVGKCkCkDJtoy938Znf09L5g0hdQrdIcAJ+y9Sv/3t601ptwxu6nwowpfKwkoqZMkBbM2Dkqev2
Z9Bog01Bgp7sbSYCNejpGvC1mzMmTuawblWqDfwX3U4YFIM/12eIFQMmQkJGVGpSGnt9ber56aBi
Pn11LTBvUyrMhKU6Om9vhbxBASMcTxeDrp92+YlU887tsD53nCh6EKyTN8/J10dq4P45enfbR43V
9HxKeb/aKX1G9492KcJ41jw8ZoHr58/vhmA+SWcRNnBdTujEqBT6Y4xBudlJZbRMdK7GBHYOivE6
Kh3qDpy2ndU9RQIsz3ydlHnc0Ku+gYJ8r3Q0tNyZSz7JBVYZI8vQT71A6aNNfajdO8kzgAsk0c8E
Ln/hs+a2cb8ohIcKoBaBVGpMp+x/FRBFeLfjhS+tyTJZoU/Hpi7ubJPRiALTlD1P65LPh7D+fux3
xHOliB0MFavSbMrMxLdrZw31CsJO375oLmvJOUB6bmVqOBH+2sQflv5zLWvm3AM38clP3mfAtRxn
z0GfSX39nY0aToTDCCUFL/QdGo+vdP08pd58u3Jiz5os1N4g7yB2CREQpIHiAWIVLewDqArZbXHu
tSNCTrtwycAnqZhP2BNyPwJ16JgeJJmSM9cP8B1xrp6oY7BQM5fMoF2kKldnxk55GEMCe3DwJLE5
M3anbIrZXtbbjNZFd1DQhCYNDFraWNk3ZrboJK6jueywqRVry8OdcDP0w1xbwr2bX9RNb3s8g0Qd
8soA2u5vf0LO+4cqMKycW/4bh70VBgv5AKwiMGuawW6XSZTU9/JaSlq2VcZ+ZMTLJRrnhyOh+K4Z
vW9NGS+ym6PTGG5oELaXSQXYXGeL6q9VAkfvjTq4E0/ImvZR8L15zHr95/U6TIwbXNSI36UNJHFW
Hnc8hWdRj7gapI9Bl9atViiqkVNWdst2o0QtwCcirynBJ+Q7hknKrVOowegHzDqukPK9+1qD5b/f
X24ItpM6YrPWCVRJnd+nGbelvK2sOzBQWrsKge4KIWms0CtHqoBzJqDCUbvh1xV9j+T21Au+YaO+
3Ygavf1qvWAl2eF/8QR+Qi2lwR+wimgX8f87b8zdu3eAOskfh3l/jrG2Gs9XZl6Ra14fuVUEWjQi
VFQPOG2p6AbjgeptsJt9jYOS6V/nGh21nFEIzLpOl7UJx2WM2c8NiOri/8BAGAgQJs5onPZ9uutB
WMcdNwp3UMc+KkxEE8FVHrg9FVwbe7nHRywKrAb2etYaqc2i6ZOQ89YhRcxUDX06VMU1sZc=
`protect end_protected
