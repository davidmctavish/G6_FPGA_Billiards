`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
c9vsW5JBCvThyxOUH2PprRXrwDWuKZW/Q7qPv429HnbShw4Uk66yycd+J5tES7AzUCyGeanqADbi
t/NXtBFOdg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
THl1Z3bcMS4H5t6D0G+kJ/FC2Y9oXN8UuO5gTyqyx046tFrVCFbF7b10tz4zI+nryigVgXDuQjpn
REJa68sEKDIsGl5JYzOYVe9IZ30LgoXUIOey68bvuu3Fnu8lEQh/WChcCnbyekJTFEdRaUW6S2O+
5xce7Ha8Gv7YClnhp04=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KL9gEW9UR9bJ2V+rRImGqHBVYgwBOrGPetNJZ9L5EOgu04h1LECL47Zq26De2Obbv4OkIEGfGFbZ
muWpwFGMSP/qDDeS04mLx/tWX4SnYgQRVyk8AGGlepDKbn1R0w9YaYChqwaqdh3fMk+xJZbtgoWp
4ejGlCOtRuSFxFcOTPGLnPLr5saG0n7SH0iOlkdKRcxP8k1FnXr8kYqxu6g0r1ZNWNYlDcRB7pBC
lrlL52/HTgYUGboGp0/wpS3BU8yKiMyKpm/Nc0Q701u3QL3zraihgQqtTSzkLZnBFXKNrCd6K2Zb
gw1krcKarckcDY4W+Jw/vlWaBMsrX/8GffFxsQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I9+ICDzIgzYMfdI9n5+7cSfa+M9K8Q9HlZVHvp38kWsb+jUXV67Oh07GXgNqpn7RlOPdQSyhyXf6
AZH+fL8ycTHV0MoCLtaJieiw5P4E1Pm7Fdq2uCENFjt8u7I2RH9/lcoRh4KurkxCVCe86Dtk1oWB
bacFgZX+QZ+FCZn+6nI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pyasIdA/E1o2abIoUkxhLYQwvp5B9zIwQEm/+EGPR3u06a5SPM2I1E62WIwSJ7iN/bqdRmd03/xZ
zjSCCiFFaRUwQmJJ5xZcUnw15IQqIRd/WQQ56gktCUx2rEJwJ4BBJrhOQsbLLnEDNgJUxpYVfXAy
ix6G1h7tonYt5pC9K8hh3YN8608V5TRujBAEsLi+3lAMFCMgjGqgS6cpljhaHIjuKULPnRb7+Rll
fIJqbRqDAQ0ubxbSrdH7w8ZIqWH5mG/hnLBefDFlIZJh/pHjOIOLGPh9RyUn99n5SKT8NF75l8Mj
ggHTuLkcPsoN2kGMWMDxZ752vU2X39SpzveZtA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
TxmWdQtoCa72lA+PjmaVWNzez4mZxpW7I8VWfPbcGicMeEL2MwwAS4LUnoxwA9Uhmm5ot+LUjCmv
eDB7SAvMi2HMKnvkVOM6GyDSV3gAIeNsWXHPVpwGySt8l+veQ87+wCB2U0M2AjDDPy5G0YrHv7SV
3hwskYbNG5I35qHpm3MFyP0vEDTw2Fa861T3JSQElQvkHyiJtc1mCK8c+3Xwu2sX2tdUav9HJ/w9
ZeB6TCc1chmVdFw//m3On54B7bmWN9Zebwnw5VQGvAYNMLyudEgVjYJwsgwTfKt7pZ93DMozPsEb
mZW50l08EWStM63eu5CZx2XBarUhqb053q94CYABjIYCo57BhlAgWgkKSS2f5WQW0T4Jc3rrfKN3
sLKdFCmMZrqfr5pgPkkX+nvfqUlvDaNXr1tYdehUiUwQuHo0YktKmaf9b7G08xq2O+KihhDW8bJL
JxvKd5VOwLu5iT8eD4v22BpAwoc1xjn98yzfCmkC27huSSupAOcJw+AP5OFOkoRBWp079P45WQOz
o/hkgLdSsXaQUNYZhi2sEsKzRYQK+hrxajBLt5oHEBJbf7wIUiygAcdixuv12Dd/r5+WcBPm4SJO
EmUMYhUA15hnaNALn0dGvrSkIP5NslL6zWERTi9G/OFbUb1a799ztM/HsHegshJwRbCxHi2xIz16
z35IEn7CVUoWVCtQlpFDFlgUxi9BshVVTf/6EayE6uFNg6KX4HhvSmuwujoT0wRmbQZ3Ia7MGLGS
uyxfc7BJHDjz5MQ3coKQd51qJqfHTeRGTAeQ9SzqASPY8ebTFMlp1vqFRPbOq6KsrHx7WT75pRyg
8foHSrwUrb/E8FbwnLnYe9umPzKEjGCTo6eXMWpVIyglksrRWrHIM0OOlju1rUPs5g8RID/+aWQl
krguToDL3/FbiBN/OpIpzzDFYSMSIhrq7W2k0D6X90tLdM86lV4BCaIna6MHSucetYvc6zrnoGID
ZdXRDktS64+FUnZpecuBvQtan+SwG5Rvqymh0vB5LWrSR34biGzmqqTBL6p0TkGzPJUxr3lqAthc
KMtK1x/EDuNMioKMJR1MutrwOckHFMTYiwMKhxvYePPfxHJAgRzDfDBKJ9KWfOFooBxhHPeirSD7
ApSD9kcvPzrCWtqheCAAtKvcZP69vAN+sPL4o8f8ZwS4u3neFS/PPgIEyPAjOT3Rx+hphXuRbR0C
xcg9NF/xUbIz1a0O81Hw+8USWdyB4CQVxN5TGWS0eU0Pzoempf3cbN/Umb4Z+G4nc6TVnd8Gzb/m
jLUUtvYTa++9REXif4S6B/jCByLNDOxPQ28fB9svsp0vyMkxtzExcTVuuXpp4sLmoIH0UguSwDrE
x5YlFE3mWIf1OcehV2K2ErmJpe/bx8/yRbJ+kETpRKlv8D6XTVRQt+Vea+z/vp51qlFOXkOir/4z
HbT597Zit9GKjTATbsheBAZFsu2OizevmfFZYM2WDfnnUnMamAUqxaKqV8sBjWCkxt7aOfu6RZRK
yRL7SOf4zEEAFHMuE+GPm0rxk/sCx2m26oOMj8DaX8AQ/3s2oNdxQ2ddf9myEgQlGerb+eAV5o1a
5LqAFtKIk9Wa2pAmhmbxUpfE38EhmUl+234E/YoxdQLzujssw+CNBvGu8kay1h0rWYV33KjltIfQ
e7KSp27ixG50GEf69G4xAL3n1v6tR1ouThly320lFyJ3Wssf2xL8OdqYZSoLvRF/z5Km2UbN8C+7
b8ffHHM55SASUZgCBIzBG1crH+eNXgiO9efb0rlBQrssgT/gml39YobX1TcOcgos3QpPzFpHw6m7
nZtdH/d+GpWJzbnPCAuEPyDwb4nftuTZZeEacP2zZPvGGROsylXzm+/InIrEx2Ja3Pe03gKZ7kZI
MEAhq8wwkZ0DVk2WDBZxVi/MP0Bbu1xA2CYb9Q2ylABgnzj8gdvoi/JbROGOoF0aSyDWizHV76E4
w1W5PxM9E8680QSTHrxcNxNz0ZO0XGkV3wokatX/5drWMmp+l8vRqoY0zc5+XDjdNgmbt4Aet9cU
9c6Gu3Dz7tgMbXBJsu4EmdbZSNKQLto9ZAd1zOPonSwPo6bwiU+LqjOV94wy+eH4/jYjYrwJiHDM
HyNwJuLi+ht2lBMKmwj6gZG9yecfGBvmcchYOpnyXKAHrE4iJyQuqiqRgL8TOGuMS/BWEZoUV1xT
i+vQiLWtToNOm5bAPioM2s+TcGjzptmZQsmk/bK0sVLLcyXBBxlTMsYnpOl8TnUXNiBNSlg7yoDO
UFvNugB1iR9yTD4Qy+bX5OT2j0OaP1aSMr9OK3fYCxIfl9oUrqQAz1fRc7UOniKSxDClSdhrt/g3
2w+S2xLd1sPkJLh1Z042bk/BdmJgWwfvjpSdD9cA2H0bd9l6f1JmA+XOCcVm8aiqBP+AncvFZkNi
zTCIrFbLsPiUkIMQ8aGtWpFmxbJ/TFaR5RavOE77XkqCyfjvAS1CkGEmQPu45C3KNLMljHvoTGoM
K0WpaO6nYpRhoTp3pB/GFYZH7IyrzaWSCWGVDfmwl8kwuw077+RrBKytLdEvirocgA0XXTckkOP2
YlEVy4zWwy4ozYDcU3sZItQzhUk+XUAtuRyMYQaD+kMmv3R18LAiwcGKLZW5sHBT11dPSGdWpJPQ
JUoI6scMIZZkhWcAd6RdfSUidOpWtiNkDD3wRwbkGsFBwFVW3fXckKO7AQMpCwqeAZq7xzyIDvYO
wNsir/tIa51q0hqSvHP2aaht0TF52ZHQAl11hXQfGtlSMcfrCP3EXGW7Dyrjtk0bPO+U5jyHiztH
b6HKhOdFZarKHPuzQpOYGb4fVlcRAYz4ujhTcfBZOB50NCcympkfCerHKuQkjR7CtJCU/FuOJWqA
LJhIn6vd5ZBZsZKQZfz/Vfi4D8HtvIAg7efEMwCF4sZoWND5Q8XUITLBQ1vm38m7jGV5WooUzmA/
YYHZ5gNMKTNI2rjx6dOapKVN2kwpUgmnqIEw6NLjCZDHmJuvFzqFI6E12fndcObS1LF/VMSrKmhD
F0RLzCARmlpQ8YQaGv3aF/i+jmYcVLvf353fL9w1QVKn+8/5CDSVzjE423D4nIBfbngJneJS3+2z
duSI7FHGEzdj93raYGcZe43fEhZ1dIF9H50A84Rix/gVFWv3NhB/Tcjk2f8AmFp/M47dxGIRkmOX
EQj3EEWq0HXDR1iUyf6YMizK70jMfZ1r6iOGMZYy4g93/e3FBklX7CleETlXaDWS7BC243ka5P7M
jhlhSxTflKC6x9toDQDhWVTQOhN24qUSYugdEru8c0ju8NYZvhRSYvCgnPo5M6tq9hAZ+zBFGOgR
wA3czXQUG4Liq0Gt+Npgd9LUYwhQFo8ahyVu35826rbZybwbX3HGwBadXf5m+yGOmAKPzhu7h96x
FoFUeJKhCU6hlBeCj9IPG9Q+DiRvBBrlgGi/SsjEP5HYTGXP3XLdza4E5gaOqj1PBR/8S6e+NLA7
rQx4Omz8BVG+qVbNVkQpCN+ozDK4WK49yuLCyMWLl6SbOC05dZziMPbSP4IULW9bK/o/Sac8rZtn
QbhQojrvXv7qj6bzy9mUuWQHF8m0ZR9T2hqwAx0vVEpoWU2qRpp30md7+/4WU6ddq0mn3zNwdAa6
nhI/Qrga2D7peVuYaFKYg+iC9soZccRmUDVi5AepG8+oGRAEmvIadnS2Orz7J9PcDEaP7/wHqnkT
E4+0+OKo50zH7D9FmjY0+zhOkinkAmoxLI3koQz1AFVoYB3Oc4FJQ1mAjBn5RDxciAall4tcHmph
AHjIjF6/npOI9rqg9Kv3SYDhY8CgNSqexhQSyxe8FRwDncSGYRq9pdL/EepWjjkbvyAfAN296S3M
KggAEB+SdNHvqqstJFzRBc1LY8WkE8ouoHbxa97vRXY+hopaCl37NXjHDseFr9iZruDOXtGtPs5l
//oZT0Gd8qEzmegeShrQFplZCdGwtEHjMVaZOFcaoEri1SYCzZS8vFWuZ31NrfAzbR8yi/zay0qG
DgZ2iLXuVJWE0DwQ5GnozJl06xnXQiEnUhF3Av/XcnvLLupy3IwVDjcpAXsPQNpYgaNm8ZHiukYt
TjNlQxroJDKZKrBQTC7aTDeyTNAdBJfWQ1NWqryxz/tVKNHdHKNjdT5ubWF+moI/KkSkIv0mRI+f
4KJEL5pr3wdRXTuAhP+2qqEHmYoYNjfFikVfcZjHOeFwunZuIlbYHqaAR1zrI6D60OK/DHl6GzRO
7lhOolznbM00mA8FGOjesVn4WR79qgO7a6W78gkt4OJ5ukjp+CiX8uTm/NA//4Ep7QF6JdB9q0aS
7uYdsBb0qpSMfUiT/Ukq/OEbLHBCcTRq+9KqtZA10v0RytoU1K/qdfOhsgSwj89iQAYCmYHreNnH
Pk7yD1F+7ZAhRvP8GMu/DGcDO6d/+k2eACv9mZT5yr4xzskXlgzrdBCD36hL5KdZSP7IKNIHcHNl
DSW+wenxH1cxlfl5OMfZDkirH/RR1FQnuVJnngBYHPlv3JHuQUqE0ZF70K4hSKYYi3B6t/ldaCNh
WVGOdbM1SO4fwlxXL9M1AmCMX7zOaQi6EkXzzWvmaHmRtYeuvi1xX/byx+rII7a6qdzETqMkvlln
n/2UCz1AFSzQjVka0eJ3b9VVDJDQ4RQhQ15cM9IeCsvqxd2WlQCLXt08AUGfHZWCjHdzmmgkrlG3
e6pKulOVGc5VwSWWbnkxeqXfpzvVQN7XZeOboQn2IuyNvWkdNmqgn0tQhFNeIanvT/GiJ0HmBuMZ
9/65RLl7uMHcKe2Wr12VGmVDyDTNZfN5V4YZwESdWABbU6vztTH7VyNenpCD/ZFUbglx2Dc+7hyo
ljr3KnNPsq0hV/9wB5WoXClZxy1KSu2ofTRwfSQi7+G6AddDAeGKRl+oVQOvWevsUzoKJBpz2q8r
7aJoFF3U0JYvZVVFRRSw3SEVeG3hpUBcAQzJFFqLweGy2vP/FFryOcmCOC89TEVYMm5at/r4uGOY
gxSUhg6RaSAuxyQR+nKXbKjwJ0rA/P9lhNgMIQ8/lqKrWEINcwADetLUHzzwcq5cgnzq9SoKcKkg
PuSoKNIM7Zt2niydQCACx14PEB8696I+r77o8mWc1zwcMxHSk2C0WnQPAJo1iEIS/0WEJfUg+gGh
QXAe8iirvQme7pLOHHOuphtSfEqf6rXqQsFPj1zB16xcixO3lOJAdW6tjrN0/V8vrSlu3M1intJI
lX4cOJxn7cTy3UrPhSRsOxpQHhbofPKNNaQRPOfzImO8p4ldoWiNK9M2S0yUsln/61pJi7aigg1g
hM5OqMT4KwvBucdfSZDGJ8RpHmpHyBniIvzbbKyiumThPmNvL4H/0NbcQwjl4q1lZfeSoiuiW1YN
k2F+vHcbg+Lrmd14d3249JQ6wdOT2DsvRDDPFwhH9jn5K3DdeEVjJAeHoHnV7wAkZ4QvYIlzU8cC
s8wqUyhmDnKdF4nz3/HafVAoKzRxa8vJV9JaNzIpQa6R4PpMfK2xK23PY+dZbtXshrkNfEap5322
O5W+MaLd/jqts9orI2TZOiRAgYw4YYLoXN4GTjhx51xmj+7R7jHGCQqn6LrEVQyhWxPo+0ztK2QB
vEG3/ieXSJZbijN6TpTMQBH0CuL0uQqNBpgJJXPFWzGK87oQo7gkVY/iEfP+j2vhyl7WaagNDc+J
pZByqjDUoxq3/5pG2G4HFj/+wyIaJtre2+kfm7li5yy6yZC9H+q+85Q3ggS+owE4nuyURPbM/J8D
1Mkfer2p67WoF+l+njAuRp6nIde5H50jf+TlnFJ7dj7hXKPDUOIXEQc2KQ23bJNYbzs6/bpCUZLS
/KDNykC3mrPAuwkxnedbELLh5X9PhG+IQo4KBiLAYBLvpkwryx/+c6iWP0MdYwwWdQNlzjUb6zFZ
xtfyu5jynJuSOtUWBYgxnDL8gssrC7aKybNiwVC0iRGgFUtchhb4vCvFcdR63Coqvmn+IpGC1UDj
iDtZYnh/W6U3ZnueY16l0SbsW8B9iEzO6M/jhFmVOkG4tmmaS4IhIJoSJCu7LKYi/JKrnVUTgCS2
iRj9hq57hJie8ty8PgaUYvMtILC9g65OF0+m41kFH4V35QzagJIhWb/BQPSAezL4CPqcVfPjMifT
p6V2xXY3uUPVVAMbyUQTXe2hPWeem0gAVxx0A8OoTMz3oTY9Eg4y+KbM7rccywEmWVGqJU1/BA+5
hvkrvh9NOuCa+pc9W7WgIP4U4cUEgsKPae2Dz8D/izCVCT1Ffv+jwqjnK5wg4N6gEQmqvl9n7ME1
8IVw3qaE2GLoiA0EsN8SqeGDmQ5eOY0unGvarzyaJ9+DqjqMbZYO3bpr7sdB+ZwGKzBfxULPLKWh
qi4XbcaEpsyBC4uVVC4650BIUJ3LtsWoJ6WdHaDGRaiYCAaeTf5cs4tkZlZI7ND6XIT738HnO53P
raCskxAjLHW3pCT+na42X+Nc2zZCJktIjPV9vUvxlKup2OZxbVON8b5ddg20kSM3GCZcOlUjDWD4
hluKs6pY7/hpxVCoIZy1u1UqYeAknkKqlNrT+p7rjw9HfQS19efLUbcDODM4GZwtP1qijVXxVMzj
0dbD3fc/7lyRhY1gV4W/YP+y816lRKLfckhCtFB2ceq375fIds+HRqMQQp+3xGKPt1pgEX15V1ZO
4A409Mdqgn4D3cOSfo1SmgqHcTTT4qgIMT5rVACDk3DaHu8NYTJFWkM0uAm/W6CZyfty1/zirW5S
EBGBWTTk8QpMXaqtIT+SEVYj7PpGt4gCp0+Y1FjhP+JN6FgMKtM3aAjfK8+jn3lrCU9YB7WyFJ8O
pVupNv+2vuMSrmRx7tTcvD0NxtzU7UxQHWOTSRDA6cGh5Va3hdeDLiy9NQsdrF+C3XVnmMZveXak
hJXury9lmwuCsfX2YJcT4WxCshnMnptMoktyMixUIP6KKEn0S74GqhRvlWIbCOrsuR44vaGP9HfD
ylaPsFHGfzIMD30kRu981jBtX1v8bRK1Of9DoL9W4exb8ViaA37nsevcLAcBKeM5LnGAtmdUHkzg
8T7GEblSbuCRxdUxNWNj1LagRugvJ/ELYptjU3NcMVrfeWbsgEop7/6glwofBO5n3BlXe83qe6Uu
zLCt1RHh2XnO7lEF+K80CcufmJfgEgkFvwNIcJpkRHzrSucwXhoWWCseUMZ6pvwVpxpfpj7GLWRN
SO0Ai1D8D0AfWQxzQgoRty5Tx1TttNtufuTxV/TfXuKUWa+rbei7JuBL4gESmEOecV3+ngw0hNE0
2E8SQdT8JJnToRzCf3GQIBXLGmAQiTmhYhHRM7aZmCGe0mVYL/0b7cpQ5PQEObYKxSW0RdMQ3fXE
MGh3IJWIOVl3ANBxsPU+E3U7fVYc28LvTwNCzYeiW4cl4bp53f++fuNiRL+SSrRx5ysAFvor0ats
yma3/Fe4kaTOncKlcpI6vKXrW9MWrdTeJ1H2x0jYO84oIYtnO+hUpaf1HrmMAus03++llgiG+yIJ
3cpG4E+xFDgFs+MWKOL7+khzfpTmhw8x2LSoMnrq3Qjr8FcUKRTt+yJBELuPx/T/h18EK+gQScfT
cxrYLqP0ejDEemLcIjlxWn9DO/WeWw9Nu38d1ndQ44AJ2JcQ2LqbFPkejr8GkpeXaMnu8gZPoTL8
fx4lGaf27SCsX/h170tmL2QmMdVIwL8cfa75dINrKeThC9W5C4kDyrpKkisXL6hRQ9nUDYdILYk0
suWBz4K13fHx1xSQHIr2UslOri8bd06kcq48G7y+nLf+clQfBC0zwIx2dtUBn5aCm5jwlgpV0kRN
scCeSrGEa0QHnFgJLZUu1Y6j5XFP4j1/uAkLoJOmObyfWdTUL0yaBxM4mXcwbbzTPXLJX/AAExc1
WBEsjXGg0WY+usAtXZYXLtpJVzr7COG/ljnHPKTUB6WVgzL3yBR0JN+Y4TSaQHWH6IkMV8YLcg74
sw9b8HdOcw3ZViii0DP/
`protect end_protected
