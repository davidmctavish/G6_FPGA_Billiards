`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PMDKLwXfL5PreXX3bLgGi6wl3myxePQZFaEMNd9G+WJDv1G06nQbGhr0aLyJ/dyGCbhAHq1sGSYx
+jD3o4Sb9Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hk8O5bfJUWWOpQymMnsc2rWJn3efiJHVwmxZE4st8SH1Xe4M/+7q8fRoWNMIACvndDknQyJTV4Na
qGAUcPG52ybLXwkaLb5OwZnFG6TcIbvQzOiE8ZpTCLx2CE94ng3JBK29Xx+eEn5XHIhNrOZYfy2w
qLCs40NzbR3avMJcT1s=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VK7rvSvi0kvoh0mpXUux9Vy2p/GkumPw8wML97QWFS4dU3sbTSF5CX7qgxUtuC6rdF7zVLlhsLWG
C6Vd1CfFWx2HImmEPIPYX8UNTuq6aYcHBZIv/GQENOklvlNJBBOgzRaxJNmV5eD8q1DwgwztOMZl
h5zRUURC/CoJvxv6fAiYv3ljXmuu8dtKukIHbeC0nueVtDKpVO/5jGCcS2a7kqzY4kE3dqS7syQE
SQqy5WWNykZPGJjl/paidxgfpEqvMUnylTsG3d766pzfR9EIsNgo5UeacLbW2f0L80eSab+Hfv+O
AOUcfKD18EOL7As1gL92Xk6JyVjwaC+WEdbz3g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M8/U11oSYY7anTsIvxoyRQHNwtz0qmvOukg/ypI7NgYdgbeVg6EEUxFaZ5vI1y2ZrhcVI4Kgou9X
Af+IjAJpOSJbbePjHAdVhlGnHhU4tnjWVMWKelchvj56n0dnQNIMz2OhZ34ImDfDjtSSAAj3c9nB
S+nF8XBe5j7J3onVnYQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mmB3Z5FAcSNp6wz4dGOGL2oSWbP1SdGQzfXl+LeR5KXao3ENPpGGxUAfkTkG/1e5+Sty/iYKi4dG
lk9nr1rvvb/sDG0ErC+uInNffX7yXMXTrg31wCphzx+C9bjfXEmWxMiFWaKgLXhPoNHaGRq8KnN+
XHoFnOz/tSMfQVM//hShf4eRapNaxpJXtk0oir9AE55jSu5+7OYc7JsuQWD+L5yGtonVF+j7bHxL
v5H1Hwhe+or+EHQ/Fdf7l8eXl59zyfh9si6cL7MO/h3whUzVu2Xh4s0Me4aDR6f3dtn0bEufEMYM
sQVfDiLMZFWqyIsCt0MrSPlHmhMxFSYV4q6cSg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9424)
`protect data_block
pxZKinn53C8zLle21m7VRT4iAWeJwdOfDqSBeKpoxWUoW4B7ZKtty8Gmu0HmPbaQCqHNWziCxYoa
cRCompG+TVq274rGH264oHyKRUrRXu1AbZkNVRcTEvQ2RLQf17PQRuv/X/p9LVgvN1WFVKxxqsF8
Sb6bpRgm7LecnUyIEhMQ+/IhHUd0dXV+SCZ9m7qtELkG0paJ7xcU8SK4H2tBymWg/s6plbcyNaFM
iAZEuv2l7f8O7oxCIgEpYklL8r2/itU+b/5Vbkds+pqCc1TWD66qyBBE5poerapAJB3rTtwLwhVc
uX1JRX5dWjxVNgq72DHiwJQ1F5C9b8GaDhvIuF4HvWJCWfLQylKtiZ/0wi7yRu8QUB6d2iuu9sjc
SV50Dg05Mm18+CGxnsVpwshA4vR7hkbic1HsM3bXCa8pXbtPFMR76ELcFFIqM79xQJn7deL5XxEE
Ph3OXp3wUFXId/jUSZ3cjZGA8hTiouJMiunwnAWOqUa/+4PRAws8rOgodBhuKBePRhZa6ia2NgdA
5TbvPAfhU3hf/a28khg+rhxJZpgbgvNgXttjHkOdZ+AadPS4fKvCOToQ0kEYYX143qf5Opux7kfF
163ZbYSYqqgiMM87d5fyQfu/tEMDs47qVtbScOWbS1TB5lBwsY1KPd+PvKO1/2P74t2TR7nTS8ob
27n7lfBIa9fNnSX9eOuKY+VTxVkf/qmFZVbQuIbrRVN9lJAtvIQN/boSCinXufRSoN7T0OUhHy3X
R0797BtXUftngfJTlSrIza1Exc5KHa2NLrwZZXLofoKrm60n5zncXabtWm+O+qKy0RJD34TG9iR1
P+MZsHgagUTtMjAW3Yagcjx/c8pgMMTBBxKSi+AS1Wuhjapu4S8n0Ip67pxKjymncBrH+rXSzD7L
wlkYHrzWnaqVFExLaGRkRK5sS7A9YHNIX2h+7JEgy0NJJFBb2feCTxCOkCffFzckc3JJ8Fs5+vgb
yy4JTnXIF5QBs9HGdGY/axjn0c6LxkZlANIaaYI4ObP7dKcTT1stGL7Ol9sI7NyO0seJGZP+4NjV
CBB+rKO5Iq99tyeJ6/5vlyMcA8xvipwtfrOqWzx+EcV5WEKGmitc+uQnqBVY5MHKa/KGCqTw2BM9
QhdvjFhPb11qcC7hi6Z4se06xE2/8dD/RVca+LhcfQFAFfFimIViTKavDH3fHoFbcQrrAwPhi+od
TXtBq5ExxIZ+tT08nKZhReJJk6C6BZ5dUrzQaHd7Bdw04ROyqZuxhpoRIVnxsiSbHv+iCHBu1tAG
mrSw2WSvp+JJPFIrt6Y+49+a/uW7BOY7aINev0RZbCi3hpCH2kDJPtStk5nuVIutcZ3ZsB/Zxd2z
XJcHimpkoC4qAVT3jqdq82snq/ZymZb/8I+HMe6MsFPk2XltT9IX3uq6ivIc5gQ+izVYyeXFz3JR
rzGt3MPPnsjqRlWBi2KB0S6+31aCRHNUqhLo25+6BSn0ZaqBkXK8UEB9Q9Jkt/8JxnN2eT4FZjt7
4BMNd5MXhVtF5vyWCDac62IyGEdXQt1H/8xMtGdjUsoWAvKdUHRZxTZMolokA859PoZPz63y01vw
GWrKyTr3ZJtf2GvUYL08uzMhrWZfG+tZNRsptIDkARM13SPm+AmeSI5JkQqFfTz8FaDKtNlBgBnd
UmLmcdaiPMvPlebms6qMdYcDCFQvw2hLM+ksMHqZOGX0sg0yf9OureXuV6dCL4tX6L9V4+jX06Lx
HMDtTK0U98iZF/dmDF+oHxMxKOIGojNPlNfiHZn0+/p1ZpFjEM6LzlO8dL/fpjvsjXJ/Zdmv/k+d
GYjNLjWLARUq3kidSZcBFcGJYQ0YP5Ama2MSK1TK+Ms9S8M3VgwvVCGVOSrAUlSWOuJaQ+fIoQcI
RkCzlLAxmAtMzmvSdKZkqiUtOmTzR/atKFDz0XxzE3hRM5a1rN27DF7EMhGKnETQJQxJUQrvkQLS
EKyZFBIzyx/iEO4NR2rmTovdR8fHRrtuYHxn3zNgaQqQp4Z3jq/mtWmPS+iWNWkKk5bMyr+4Vewy
uy4D+nIYlsrAB1y1SA19AV3zuJQMcM2KWcULlE5PCkchhMWBFvGGurelXrBXrtE0Rf6sa926X3Ss
s0UMGZRxeCVpaH18Qy8Q+SwPM9pCZ/wx+bDUD0lVjv+ZjTuhdDjW7fbUzuka0kVVa2Qd3mROMenU
gCppC5LBGRUiUyUbbRSe99hAHb6lCWS0fHNxGZ3OZZ9CNVP+KDBlsTNNr+hvlNvsjX0HXbbqEb00
E4KwQNOn/q2PBewaDk+AaOBEle7bv0BsRlikjAdJXT9Lm7K9XTkalNDyO5aLhxFiKLqeHt10SNy/
+GSPfeKyIuxVnl270jMhn+Ou3gsJO0SOivHrcz2c8359NJbd3MGMlFAa0x12JiLRZ6ZFykBpvqwF
ZM8ImJd/Ojgu07MRzCshoDWu0GSu7W8eWLBlCEDkg8xwyx65vA1ecUD3WhgRJgLrH0Ijs4H8JR6D
mI+eSchXJ/phOzSnu79tY/EKi4WNfXgMA10p3sjg0Y5G4hQpvThqIp+PR4QAZO5EnZUtpqaxAwaC
6fgo4e7jS9VtVME4wiscBwxcw2uza8vT9qQyYpkvDYQ/LU5aq4fcBAulLXi/cQaogiyvT2y47hm3
LVZDvGshF3R7/XQtKnP67c8UqBgmsQSGEXegMOUMKKQHm+K+fMw3cuqbVPgheN1EXcs7pWxNna9a
T/jeza8Qfk7ydE0rmNbwCYKGKqj+EqpMQYW9l+uObjmNEL3mshdCw8plgK7kvyk3360IIyUcYHar
SxOBBD1Bp3KyXhbj6FymUBk603LuNRUsvxCfPhJWA/u8DkWyzbQiduRznMie8SRu/h/4aHFZendU
hkMAky+sblmEWmGSYi+LDnf7103UzjsysBdRSdcqA9d8/UQjHe1G0mWbwA7n+LnUpCGvgaEGT9/l
FP9xjM93lFcMi6Tu3a1c3VZzRo6NoVSuiFbZ9PLfDHt5+sYtJojl+QMLh2WNCoVrQb0vg7VImfUQ
HZc95KIl0xSfiYxICDxCnOnKJ6FmLPB7jlFAuu96kughLFMqwcHLusAcy/kb2jZibIrPUsoLnP4b
rdT/uiFQ+JjCjaeCbS6EkLhHEZjFEKxkzsS1rptjBDy/luhrJMugHQN/BGh+/Gvh9igrKSn/2l2O
/HC+9yu/VMORICTGVaObi0EacTiA2d1as5bmionsqs4AN6pDvmS+Ph5QmpdHhGXRhFwXvvQFB6oE
dmikhuo0+ehT1JrYQjMvny0swVJ00oFaNHYdntkEdFmh8DOwH0oayA38OkCFUFHG6kJuQAu0mMdZ
h7qL0DVWw8zANcnFsShX/T3XIVYw/V6cc+283KhZ/pCIkl3KiB4HeU83DT5R8ykZ3a0XmVUhamgl
AW5ln/XsEd62QaYQpjRwzeSr1+pUVsjV86k4rZu3w64nvg857eDGzIEGg1u6rgWq1kS59KEH9GT4
l0kIXqbS/amvZDZLi6kFq3hEOYauTpFK99ECI7Cigz8c/sdP6m7UnnFg8a1rUTPoMhSzStFJsPi8
tEu17LJ8EShvG5USc6P9DX9GIXxHcc3CjMNVDuDc/8DhJb5Pit6twjjeFqyaH5A6Kq7jidpAogp/
6M6ftu0MBl7dDub0QxAHenaNDmI33F8dsYhAio6a8Ulf20zZGKitwg7xBjEYDAdyR3nx1TNqV6gU
poqZop7714UHZ1SS01AbYea+F1FovdYyou7AqnXlU7NnlXHYPqmQDkvkf9wcj9lxZ4GyRzyUCT+v
zbsHjDzyvMEtwj6TDKMWETj0ATsGoMgDusvPd7S1FqY5QtJr0Eu+UtFZxRYUjQunMy9XFU6I5Ze7
1LRvGFdRd6ypmktAgOqPz0rtArQjOSLTShCxVOWnH8FB9KExLLLJYR3Rr1jIIkbl7GxJVoKI1+c+
eWe4UXANI5olS1BNjYeFWFQ8HC+pmRBpsp3EZmO6qusd1C0nOVCkTxle91A1CmZvaZ9/7lxx5Ug8
ToD8jTgWgF6+2j/P1qP2itqw8WtGXEy7NEwR9MFE12us9adPvTgR8KupXJulpKIExvrwAF+ABi6J
mlK2R90D/cYBlU/Gkf+or6QyIovxNrQScEGzo4ryjKLLJMgzRtwYjFM+TpHn8wy1YOPjNDdMSlON
PI6Hh3YmD4Y3EOcXpuax4yr7pLbmJADo7LvsYETmnPBHezsteLXXjfobeN9lb1aWxM5qdO95WyDU
a9togdta3CKs7gOMGSVNJu2gZXtpfYJvkhT0Cr1y0bhsyPJ+Cglg4zbYHjzsC1PTaFokQWaXaptA
wy2lTfb6h/aXLaXajWP54PgMHE7gC7gIAi8iRnkNsGL1UPf/0t1ZmUVtmPIBSK48gXTVbJRpJkJq
KU7t45v9yNrztJbzQX15bSbqHRJyjWfAnmyqduBxD1hCfZr5ve5n/bb9Hb3Zpg5VxJKWl5S+hEql
lPNO1ilI+Gfj68XD17n2m7rQEcc1uhdzj1sU2ffQ6DUsf7jK+yi0SCkfW16mW0M2zJcS0rHYuBf/
Fiz8YelwU2RysSNXkvJOevdTLvbCzDP7eolgfAWuZEIEyrky2JE7MJY99z7jBbozPINuhDDbZ6eX
EG/j84848+lXB3oBTE5gVpuEjJ2RNn1jm7/QviVW6WZFiOUhq0AtmMmIt6C+75leOJY64hHQXNfD
tW8oo+o7uCUm9825fJcjFnWVr4RAKp80f7BqwYKWspStpFx1+1vF/WtHAJPuwrLX6ceMcxV758Vb
WhKB4oxm85gHPbcibQL3CtOw02y4nUPPuBZPiuteJQSYomIVl+yugaBh8MQrM1LvPHN8BZPA5BL7
D0LUFHP5TKNsvdwArwa08T0lTzV1dAT3q7S1vWWpnd6wLV0WB3FCDxjgfWvm9v24uk+6wRDxZph/
1/f/k0s0rmYQQYiAJGLdBbZKMxMRJ71xyXK1yE54itXocUx+7v+v50UXR9Wink0iTRLNCBHw8p9+
/8037NB7Rh2y0oEJwJS5SoCsfKd1Zrn5EyyBsnx3pVqfvmtZV/Oqc2QQKAk/YpYvqol9aXrEDlXM
pVlD24y8e2ccXhQKG5jENMgEmSPYjLEmyPVGNv9ezWRgzyM2F/StouIUn+4XIfePyw7cgJT9VAVj
GCRrylldYKEQ4EcNwy2sDC8rRDXKSvP1JRK/e3+V/TPBuPt8qMP/rwZExCRf/WyxqvVAi5NYzlAq
S64uwV14JGZHVHDGMial5TiHwtO1JeSagRYUfw5FN0tJVH3tVnkEG92+eeqZH9D9WmRBMmCmbS2H
+ixhRPiSx+0g4BfSVUganyx1FnKH+Ktk7ifG4jaAjyxjO2db0EyzTRuDKlNDPCwpPNNGi6p+rTPe
03aokEPyAv87kcHLJnTiQoVy+yqFKMYmoo/k1c+3cZGSj7F1Fn8X8mCp27HSe743/SIbkyHgnkbv
PYE8JKqiaprYT8vm8vTdf2HGDzZykGqiib8wnBRMzzYGbbr/iSoBY85WZ0YXsFe8Y2svkc57wczI
Dh3izqTtkyZ94W/3/dM4OyzLP0I8EnnbE4zTmYEjLAJ+fTbaCwOESSEsBkb8Z9wlQuuyfgcpzQKx
piURZDDvH23vrQrLyFcgBXta6UVDy/yhWrjOtcj3zxaQ65yQOuU+ewZpDHvvzB7ezpIrZ5j2yn6e
vJGSX1UK1nMDGND4fUquiOCchyUrnCB0nKhrXhzqYNBvEMw1jror7qjyYpZCZy0Zi1WewlzauAkp
HpTNvnsDWy7VeTVZoVRrPMIuXq2rijAHkKgJqS5Ff82neAGeXe9Edz40mXM44rHaQM/k6xAht6lS
CoEhBMP0O4wAJlUhyhA6k7z9fWCKRWazDJZO1hl3wkmjKa0Q3cNtgnqwySZ7uN+feXAKeAtmv/Kr
vCw0h6j0QsPrLzhzs6lVtYCh1uszGlWxpMSSiz6K9lw5eIiv/SDftltHVg5xxNGnT3fMHG92A+df
eWZ19P0j+7n/r4g77dO1mqMNkjYvQL7kBvt/FbnV9AlGOjuczRnnRrZpryGelMamC/08xnhYOhZs
xV1YlFBKysSoCNMDN6ewxTpmhL/Q02ZCiGrOOgfPqReR1zruOSJ1zOa/4dgMw65nfuyj4WgpZcz5
QOnn5iCwv8FqZvr30eX+qvHxZVxtcLhNywVHOp2nMZn1F0RicD7CVCjPxy+aIg87tg6IYjbfatRr
sxLknn0yHQUmAa7rLETa+R41mDiitAh5B351/DDn7TWbltg0pQ2Vj8RYN3hdSqzaGPGOKX3BarmI
vB8idEy2PEdetSNpIyod+i+L/E3yOI6GROJ9pmg486CGWPnqjaNCatFLEU48xsfhgN2RmFSN4j6d
Vb4wBQhdtsb6BkQzxo0SM+Cflmgpc/+yiPa08X0/+5hk3SsQcU05/gPmkk1st8N+NNembw/M34AU
I//Q2QTLRRtYSb9cyJh42PMQUcUYdAkMd29wYJz28O16JNWnMz68LERMxpgL8z7XYMpL1Mc6+9Bz
wMkhwcZ9BhYGGdci9EcOPDSdzURvzo8m5kCi1EABmHs/MvjTW45j+q9k7nDATE+Sh5nPJO8OT1OU
bhCeMbWqkOORwa6UnTN6UisZXDtJD2mHmrE95Bq4ND3ynTH2z5jRjDzNV4qvPLwcNJobDspudTjq
iJ0Tmc8D6vBbBgqqC3uDcfu5NJsk+ge4BB6FQReUjMUUaWMbxHaSnEP2WI1qiNSO3ylmwuUtTsxg
cOFDRm/jv6QkUXZq8oWGpMU5FYptgZKWzovVWO2eNuthSrJqj4YN7t88EBp4ANgODfmPP8V6ss4u
pLno8P+gqUay/GrzuNqu4tr2A7N0cLIFSzpFA87/oBFmnbDixo4C7Cev+qd/Fn7Al+oK5O8RhneO
Ru6Xs0HNaYq1cFfTKykOWXNDybiNlptZ8WY5xXqd6qybgDLgfjXbnItd4jWJ1CQjGsg9FY+GCLAu
PN5md3nEqkoC+kSDdsjGsKVG/vJ9kTay0byAgCBQVsDn1zty/KpysZS8UsPCs3SblMdUhOyS3w5+
dP4mxMzSv9ob4Y8007tTykp8SHcWPaMx9ZGvYnwG8JkJF0YJI0yUVOxWU6TSqr3VNWWLldj6rcC+
WC50cfFRek0g40LvhsBd9YnFo0GvB0/O6UKqRUNOS78OIUVgmUHkedpIdsqUOQARjLqev/rhK/ld
RWGmIRhLf/bwO7lvSCCMqojeoAgbvf4rx00iywIvWhpj6U2EtdDanUMqzXhZAP3NnTx/skO7/v2T
aVN6F2FN0rIawUc6d1TrmwZIDEXxctShlW6re+9EuYCXFfQqoHjQthahqNIvHRRXU1P3Zy9BO3MB
pO8/2CUmiko+FKa4QqMld0HgFQIBlCGK9XYiHV//TomJd8gYEj9Y7X87dtzD75cRdMiZTPbxIDfQ
krLp+rAE3sB7pi0CgqPKSDOM5/QLh6sW931a//2WhioWiRCmwzdQtVXm02k6L8Qk9yxsChhXnpqQ
cbx9kfkR5Or/qI4V7Ii9EPmDgGLbMftOBTw7BHa64N5W3vcGFgmAmatxc/jWPKcP4wHzLZh7RIQh
hmybUU3V98Svs8kjv3lE1/sOR8WC6jdnGZ0Lt2NrBWmy/AJIU0b9jaeZlIKa+RRrZqBQ9zcjpLo+
X3TLjSGVnz1Drh7qCGNKbBosbSmMUwFntaEQkGr+Jwc0BNBdC9E15VahuYJ4MCBiHpQU63HdT7Ci
zj7A+X1MP/ltZ2y1EEitrSiCpuvbBt0hYVPT/oSnPHm19Ccxygm+Py868FyOTvLe2Qzo48/elR45
cgR+FkpgXWtLCUnkI9ihFfWjAVlaEJbrtZ3XKUgK2mdcrdd6J+oLov/6AHx0/D+s21/AD4fqGKLi
Z9AvJVYamPWeg2kTinByHi1cmH0LqClRUgOzw4dBQ3OxCgz7l8ua5Wgy1Ya/l9ABkefCDJPrH1iU
9d3hi46S8MntzMrBim+UTG0q3AjnEPNzZy584PvZD8dAlq5v9cn3lFSp54ogV99T9nOMqXH2b18p
b8NLObVUgDwOyU7PjEixTFIjEHGc3wurPeYh11KxQG4oh6MDxz+5GLmW+5wjHiJnBve3J0z1iUAQ
iyfS+0jIyaMeBZqCgS8tf9WCH4WznmIQqQBvERcHy6t82HThBEgpSCx+w/al2QlrrDzh/PV/vKd0
euCHNQiigrzZkEUhUrEMEjhVdog5mY2g9Y3EqHLL1Jyi48MmBTJ+1eVpR2NS7MmFuZU5WHC0FdIe
1brI/k30Rx5mNKEiLh3G/1vwLTGEVtAIHJTrzvtEuddXpXJbkhuKDz//ZEjfVMdFv0f9Wr2emhy1
m06oSPqRoLPM6nSzoaKn3Ii+IZ69kUbSCdsigeGQnHih+ubimGngucZW3CwUjgWnpJgMQEDaEOhx
oVk9iOkLtTgiRli9mLzVoEX9mJOJm6qnjTH1EUGsQ8uSdxA8OpQzyiKgaNXLFsmw9aENv2dQUMoT
l5uaBVkBBpKfO8mTifeT+XNc8svLPJbrluAaQkbxhw8aBtpolShMf080q7HN2WW2mRWwAFKMZQ3p
NSkLIFmYWrlUOM/aE6mudTZ+TSjBqAg4Yan9hbunJjTBwayB6oTJNBnGW95CrAhZAsjK+Cya9r9y
lOnXlw2ibEg7e9uQ0kGtaY+qpe8oRLfkKlZii8xc2IHfq8wdxNNJ9oxNk3IjeeCitgClftZx9QH/
xaDixEF6F5+KOZ2ceVGHOKdAo7Vg+zzWAwyuuBK2gan0dWXp6DHgij1Vp6wHdPEE4azMdEaW7OLa
ynkComqAeECi15VDLbHNoHASFAZtDcfYSFtB3yzakQ4++5YHEL0VGcPlW96z7r3RQ44H5hwIZocE
YfiIRBW5+wY+8L+1k8L/5w9CoceX+MULRCQ95vwPE7DJJlSb+AobUfBIvYGthaxTnxCGTt0ByKkq
KvbfPww63bL1qSkEZN9l38l6f/n7gntLSTd27Ir+6IeYJrSMHJQ0AEvBv7N7Mj4tkpuiz3LKWr4O
CHoPgLj2xHKmB4LhsRosqbX4uqfzFjFM6tQPbK3jBNledS/klQ51vLBE4v7vZUlowzBTONw8K0Tf
P0l+/afvoBIbK9XwxhOthHv6iXA+DffRUAbiMoLVspyIwjaeFosjNONj5MJqx/wMjL897fwdIVr0
raZcRa1LsLNYuBfZYKHka/uTZiyx6QdfXO7R4nVks6xy5OdEcU+qNSnjKAgLPgxvw1IX25bL/zof
obQ6O5eq7EPV1vb/VzvGszXapXO/uiYjsZmi1c0XX0Bz+JjUqIV9RHPc5JpyY9jCIb2ulA3eTWQ4
7IOHsA/v5dZbqogMXxZx7YQ+0zuUkRCusdm380XSj1cCBedRfzRANlSbuaVbEHYCY8byqVeBXCcU
uiag7LmmaTPcenfdIrWxTam22woN5wZlH9+vQUrOP92271i7YkLBx3R0Z0oXO1k4zhQHSpg2g0k3
EErmlBCLgVgc8cucWuPYVBV9SgvBKft6ItBBqlgz1JhNntSBv65UvvEOVQgfYPdYA0L/tm+BWV4D
zQtFvrx1IbbiPyiGy9IH6U75AZeaa6q+wvy58xsDmfR0hDwNmqMDGPjaTKgguoX+VZOxzOeG4cgX
DUFti9+ZdXdUI2yM5WNNSN33nCJUgdxzPYxM81wjCkspD/5jvyFABrUPo+U9E4dlelA2Spdi9bJv
4GkyCVVkSAp4q6ibSTL4Jpfjn6YNMTCKPKi8tpT7JWPUJBuySc0102nNVSlMgnb6LNB0ZIfDDvWC
XDCz/QZ0IcoXyEPaC6VAgoiiL6P9pFSrevUaGJYrrVvDhyNA1uNvkC0Xmf9zxqs1YmgcVfQ79Xw1
fDpj+4CnJYomIrEPFMsEnuadd+ntwCTxwnkMshgtiXsjk/GBfiGKKW8IXJO69A3uGQPLZ5wGOlCV
g0VHFc7sgBIPRT7hzH/YM4coWhgckjbUeyLs2LOKfVWLGDckBvtDye84Hg4CjAC9XWOIMZOE+oPx
uROiJVyJl72ev8H+4FgwvkbE9flpJ98xqRmKXyGGq25jKVm9K1i3JcEKJ17gFSfMV/GOUdWkEjgY
6flcI0riKe1ynwAdCsgg8yqLf4Tf6Rpdz39L9loSNQZmOX8AwFcdjq/BDb1ePWWzQ/4dIr9kXQp/
Kx7e7egfzwX/fsUKxusibDUdTX4s0Zf3jpQPuObdVgcd/eisC5KGIo7N8cVUQO5U06XIOgTa1INT
mqQN9L34hzXzX4YxuZEA1jMy9hjXN/3BnjrxwOy++0S5m1cbsJi3WULgOCfGCZMRZmxUxzHfekjA
F8q1dwwfYoKkz0TK8QWSDkNNfvyuhh515iHVorPGkZq38imRwB6xt43VeBTEelHyPKAPZcB16GUM
wKZtDGPe7Iba7IxaQWWcxRlJNEuJGohcAERhBjeqIFwFIk0hkbkMr/RFEfmt3pfgJzRKq6bnv2uI
C6k3wSUuUzu2nSUKoFSHUPMM6JEvTj7h5vWQ9e13Oq0f9RPqNTi5SYq7W5fEZo4EF6JL3W7kmTBV
yQ9sNcxenfjMMHWMeaaP97IMnDgnNz40RvKas7ZHQOzXcVEK286R4rKvotYrxQXrdYil5Fsqpauv
qslrrJkF394XYeGNGkURB2nnfX4TawIYhbmr/c6rLRTdMgPHCeYCoR4lkQkJLwYjE05xqcjpB4I2
Pu+WOQFVAdLaYEqjzDy0tTEPcJ8tYwssf+unM6XRl4K31mYd1kSsm+Vrwn3nVWJ/OckXe9QEBV0b
cCrSfY13TolZXVcHShUSyPPFhoRvKgpIJUlp4r3U1Pvc01/XaslTTDLOs053zJqbPzrXcapLwrSl
tmJd/ChK3cNrauxUnl0A8TFYcuDO0PUSr6mXTbhylABjaLEu+gxM1gNJv8lfXyvjZ1iHLggY7yAh
lMApP6eVjQHtLi1fR/TVDdffvfB0mcUIHHs+13WdynXBT7Wn5v4JZ70LhNfHIfwOC8qBoOr1/mo8
6WSfSgcwYFqQllpaKR7BjSV+32xpitRYXSwbkUXeK5tEjhgbc80tCCrKlJet2aHAHrCxvl5izXAQ
W0GwIiESxUazoSfd0Sty9LvdsWEKmLG9dWjZcsZ2xIuWz8VMuWSG8ORKDUdqw9sv3K9kbIzQrnac
F8g9uJTXiay86Oov61C7eMgkAVSBMxYs74DTmJO9c4A1mC5M/3rD0jTVvgTvcwvnGNbH86MLf8Xm
AXoYtZW1LNWevNG4+Hpe55J4s7ORiPlWRicBVNgFqq2pxhl3D5qpaIQfcMDR/HURdvT8HEf5bblF
X4NNhqffIVgS/NAHG+Wt3AFn+XZONDJALT3o5QyddOA+IioeKnYCLjFdCrz0semsatmnIYQkidgD
94X7nT1RF4wy04kDOlD/9DNt5ZRd0F3XEDdS7cM1YxbHFeJ1h7EJOWe9vVW8xN+Ks1GfTlkwlNUk
w0Pk5S246nTgKP+GSffqoqrFlTkfp7JYjtqB7r7bhnrZ4xTAQgdKBw4fEe0mGmd2dwu8mZ5Jcd93
UJhaFlKR+KE1THtJc9qPH91bWOKTknHAdBIlkHGC0irOYwIy3WMycRN48P8VoSwZGfiCcbZPeSil
Bmbs/iD6y+cKPtaXdToGBSDGxJ2akrHHeX8qk1pua+Gl4WmwDpMIOgBkoOwt+kyv+COW2+ZIa6Sq
bTFVRtV8svLa9HCj7AN1PYoz57mCzQPJbf0ImpvgGG/0nXQjwlMIYqSGzVV7V6TiU5zID0BhIogn
cQuwpIhTYFsP4mbyL+f6ed91rYi85OPgA6NafTwQVI0MW57WCmqne/CdZIqDTq2Pj+CMUIBLTwrx
eMMtprxuKs84up6qn2DTPhyw319NnP4L4PdvnfvTTtUZ23wdAtc7SKWtzwWDANJawZjHOcT6CcLw
5g8Zji6uwV85E7TqCdPIj1LET0e+D7SW2Hjx5ae6TaES0nAivXQuohRbkVg4JwEE/BZuZKlLxxRE
YD/nZ4Y1DHFtHasuK1JPtBJi0LYDIxP3Pw+vMaFCHFeiyT0qkqBVgNtR2pnxiVQJOunFyBcXhjPp
qL25R48DfiogYXG4W7ZF35GmI8HMT4kicKO4ARgMBgQeFkj7O6tPDTuDpD6wev+iUOsTEN5tKKHt
cl+oMFJFEsaZ81lPTb6maZbdQ4cvqDK6vIGt/W+csDCPWxXOacitutfgaM5sD1oL87YCsCRVVbOc
BNd6B2qVm1BF6IKMDlp0JiRw1yP8KlsXBnnlWQiwjYACcT5DHnIZ7xw8KHR/ASN5QZVGadj1WZ8+
POs77Qx5ab4pC2/28liWNcBknPEQewf9U3nH+XWtKDRdFM+ocAF+LxTlN1oDRD2cJwsbb9DiRqaQ
99xvG33JdT35g1CNlm9b544zPN3tj+r8JkesGb+YsVLjFFb6BvOYeb3NPxhSbV0f9p2HbkQ69eP0
LeB4IYhvPFi6z2U3PROxJjAhasOtxMgt2OtU6g1SiA8W2QmGpZcPLjRKFQ1XfBSKn9I3n2Y15vR/
1Cb+DKxvJiYolxGdWF6Y68cs+w==
`protect end_protected
