`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oWAiulLwHDglts6iqdMUT9Ori/ohV8QguIR1lM7voKoLaYFRvD2S50wWzfOXl1AqjV+esGm+neYh
aXTGcZYAUA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pjORo1VUicxT3KNrha3dwkdkacMgeKv6htW6OBezSAYVQTqVECKGncr9yoRXcs7sGJoZX4VaS8ia
lihJEHqdU7spww8qZeDL6kdfkf73A5GDuhlxghEKWXxnanBE4/mPjb3CdNex8j6f/V0iPwVP8zbO
9xb2L8Nnk6ScRPEyOXQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Peg+7FfXjeQbiaOKxmimfzP1GEfA0xs/a9tFt2w9gwQHX8Ly/Cz5LlJtL5mdZ77ckvdNfJmQ+VHs
rPs/ubGwZr9yQQllrZBHzCwiuRRZU72CLZZmGGqZLsgf8SrxIZGaIKgytX6pCleoLyzOesqXBNLU
/Oyo3S9HGNPh2h+VRbnosGrZKDBWjyQlBWadWZ65Pd2QdVA0z+xxxUPO96CSw0l1/ExlNgleiwoA
uaX2OxgEsUeESaj1JZGYIiMkHilJHZDTkcMK2s3YsyWOqXhwRild6TfejTa2Fzn7TH4K0pu++7Gt
nmVIgHvzVhBs5sa5Fo6vXJKVBorZwCbjGDiu5g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UCcotBKd24z3jkO3jgLbsxNWqi2O9+6jaXbotiZjtapozjfzg09PNDoEdTzj2B303WQ78dPXEphn
GO4PzKGdZAdDgvtFX7h6cCngchutOPNE7wof2pbSw94kWUGoE8qSuK1sO4Z+0LubR7c0IIN9HAZ9
pEoqViQqlFMCXUzLkDk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PIHoiy6LOs6z9eo851mqeJ6D8UYzj3KAeJ9fm4AKfKKarhRamXK6B8lbD4E3RQ3pdDWQccWJcZpR
NH3EOtpAZEu/MkvXzjnjlwMww2/YpZce8bPLwemJFMc39ZZJmCT3SWOlQphiINLNGDVxB/CMtcQ6
rY2up/+ygJWF9vC426YbgHTJvlEVzCe/eGFMA+8YiVMSVx1GFhZK0bm9zeFSEr4sYDaGEOTvCs0G
hCIpAYk1atmrlyyugxDXn8+KvQNZnVl4HaRRFWZzU1oDVAww9Nzcqooh/njU693MwJ2PwWWVVfWl
w4hty2wOg+59AQpZ0b86zzhH4IIXVJ9olmwhIw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29280)
`protect data_block
F0/ac1AzI8udZMEYRTwiqywXJeZ19oc115kzno3hdmHexJW22a4vhLZtELpP6K+oay3hiNDu0IK7
Hn0WG+O4AR1fRDL2SXezqfirLCtCJEWTR8ZJmhGc5rn6LF318rs5zITWLIYmU2/28ipoGMbtO/K3
zikoXNiDstyKzuZlluE1ZHwlTDic5cJr446L+e2XVo0m09HlqB3xyhO7F4SeI7nZvAPgWQZlEhb2
h7iXGTHPzI7/lKtZKDfrgw7i+rWSBvsuaqMkvVjXdfggN025+/c7TKF4b3X12YU/Jk4O9EVwi4gt
HPP6oFql30+YxapNTjdDGb+Kkbla+W7v9xw0HqbSpMN21/TuWSBl/lkfYxp4JineHV5fx9BxakQ3
zvpEmVsKnnSOvwqtBxVDcouNPnGk+IV4Jk9gYwI8btLT68HEgPJYLmVDKB166j1XNhsSgOSBY8ll
kPgteKhcqF59bMnEtVlMLVoJ02KXJSMzoAQyQAl/17mivxx6dJpZu7ppcrtk6LO+p/OLDqVMWhZF
0mpDjKjaHIyYZHGchc9Ug7ByX6FkdJOqckjm8XSPgcZZu9FYLQFVy0Qj2k7EzSMCwz1kkhDqHSWp
1FCMADmNicxdrg8x8F5ylzgW4TrpAcAmv/Cw5bWoiYPyMQZvK1wHpAIoY9AnB0trUTPdQ41dbIec
3scgOssX+v0yLaJD4mM/RpgYGK9biddsN/FFS7HiQhfs9H2nYxA89oRudOS0dvhhQ5CilM3xt5KO
t33GVAJOwYEHBJvDolYDuJzrKgVcYS+jjZhKK2DWLTvt3lTOJDF/sH88TNhrXAbQ7CbEpmvJt000
agoxeWJYsO3eVvK7Nu/p3VpqmJWYNIUPKnNjb/6cVkWE21aVIhoDofwTby7oMX2wbzKx80hqS2UO
La9Asg6I84BR1vYVyohYqRsk6Jl5alwB5wgpJueh+4vfN0249Zga234fbxvX4cWghW9p/txAAN+T
eMododrHA7MmbmiCXofmhnzAraXgFqPuGgehV1KBNhuY0SK10l+LshkA//QXptyOT0A/ALw9bL6y
RvqClhzRv/17wHz0T/uHdk9/piH9+GELqxYlDsyLVv0EUJEZpbp/uFIbt/DyH+A76/XXRTF+yx4U
NjKLzdIqK57zAXRSFhMzkQgQisie0HgSl6FTr/KBOBleufvBQVp8OpyfNrtZ6SvarP8Mzv4GQcEw
jKtktF8gFGHi7WNjILRE1l5tzfZLfTcWU5cJHOv6mWISmZS7FFpwjyQpwpsvo/DuYb2WBkaDzNIK
1LgE54BAj2uN3W1TpfkfgqPMD5B0aoZAd7aJ8T7MM5TzOF4oehfc9cC0GjFa9gNky9vFvfAfsQWf
yfEu5cqQ68hTeQUDeCE8NYc/2Cjz2/NaL43zWUYMlivqJ631MQBP/lsoY6MkqQ22KB/bDs51QF3b
KMHQcT18RYOcjDpiwDcBNvy2RpeXWz66i/CXKSCCfscFAYWAWqef44ybWw4yvZL3vlE0G8OPUqD5
NvTWZOPibK+BMHCcB5GotVr19wWsv9vTso4yl86gKgYihWL3GlgXSTqJzYqL4vBsdWugogBvXhrh
1cSOxJ5ry5rIrjOj4ajY1VgGdmMRxQ7xDFryRC8BDZiQXpvu7l6tbN4Actj1eG0b32RmB1DJxjMg
BhxyADZ8YM38SipoNfmAeRI+QEZE6hSIfkwVSdtCIoJAddC5FrsDtv7fZyTGnz8TGUcVv/P+M56k
dzDOKo6lFx26q2o45hp2II2VgSb0+BCVlf57gB36IULBIlojDgcZQ1sta7j7TTn5xSFLpGOtOcWZ
uzKQcDqos/b+vVlKZZxvg76hHKINAzNTNgQFdgJ9tkY7m1OY861tDNRhuZdakTmwn3OJmMNwa5dl
26C5w0RxG3hHjK/IIdwM/kUj2v0GSFGoairELIIUu7GVc7nNxW2Z7dpBooUhsQjUyZMiBoHRJTQM
MVttFg7shCzIlUh9xqKPcoEs5INShxIaYBu1KHN9++k47JiWBWcixR3M9EWLO+tFHmrBotitXYk5
JLpuo4OtYo3+maDQJKsXeNI56RnBzGZm/gQAyEPFaDR9fg1TPNe6GvSC3RwF86hAaVEuWKLnw5Bf
T9PpE7/DI5qyC5y1SN1DIC7r0si1CUva5k24sv3576nknEsFmaxFFerP6UhbduLScuP4lWA9cjLH
oisbstUxWg5+secb/1dhKVloKsAA3BmFNgavzzYcjtpjWpxW4D0G15z1aRrIT1hWVQXttVvkoPJB
bn+RO5gCLsiuZxajKggnbmjDjSnK0pDWNhbfx+wcB5asEK52Jy5cgzatt5uZTn5aTgnA+RPqSfq1
5Pht0N3DpCSnkbmZTQAwHphu/PciVAQMydXt/u35mQiZRTM8KiIQ8spN8g+hx6TuiKv5ROtYMZHE
IQLg3oZkOCVl4hVsYLoe4HYOacymW/pJ1olaF6zEgkbHr3hELRCL4VTiansALSU+e3/7wIVwQUIX
KSgJGABFcR/r8s/BHaiBSwLbudX+ctrA8jlVDVJsGkVe/cqmhGxnmcSEJLk/jVQPfzJLnr79WQ9X
wT0hOT2T0xM5kFMu+TxD4rS5e82QHDUFhWnZbb8yuH22WYRxtigXRdn0wkUFqK12w5X+/cXywULW
fd3/u8USaXMvJvycfvVhLH+Xxu4NV4Tc3K7b90L/0m2RLnrWBH9WnGkUZAlmYEgRUXyb7gpcJAcQ
sa+WQmbUsYu2BaULET4WOkHXOIJCQYTiTm8K1i3AXL0pg6xcOcqKdA80BgfPq8+NqOxcsDQVKvj0
eZpnqwaXf5gKLgygOdlUDdLARN8/tkapdFemdP2yWnVi8kpaJovosrhnTK98yHSFb/1Hgsc8MCtu
ENmx96PdH5LzoOPH6vBAn3qQCTBrbtuHGSlWXyq4V25tgbijp4Ke0mBh4hW81s0/vA5FoA9V6157
lfhVw4p1lVhDNh0BTMh4H/Ux5IxBbYhwMZjnbLuemYbypWWQhw4eaR/maOEde0c8DWO9CzS35qrH
cLwRSdEp2vFXkt8tQsaP8fIh/gVpXInXMI8dGrjy3YTxPdRyqHKdKPnTsnkbw+Le6Ty6FYmyu/6i
xf41TF2lHGB1MfsOwHKYDpY3uNWLvhxogKvrpOlvd5IqE6FnUc8Lu/JSuKRNCg+ECjFRwX2xKOMj
r+7wrwdVMb81kio8Vx8L4KLbNa6dC1bISXMr1LqRStihmX9U9SxZqa21ae917znlZpVLm5LtWKFK
+7ygN/GMC+zPjhGgJFxt+CAak+gR9aonmskyBevKpYMzyIvCMZEwmIqph7VnscBjsJ2m7yk6kR/2
bQtusmh7gadaiFdF4x5/f3tQu3cXjJzWe7nRUQYLRfW9XhDnfvJq3kiD62x4TOFOw+jaf2hZbEcB
dXGX0CgA7JOmVaMT2kYvnzMQ/394Snhpf5QKNmsAhaS+F1tFE+bhJnWvVX60T+ndl8LyYS5zKPDs
yt4m7s7YiYyOimd0csP2fjRQdBvkKjVTUB08qU89/wNWKfE8tpEOZlzOzS4uHcFWFu6bdubL22GN
fk4iDa3vQQOSYcNCud9EmxFHOpLO/u1EaJq2TlQLhGClIQbo4y8mcAnzcbNZ0ljGzATckfh8EsCk
w+vSDw+KBTbrJenPwm77JYkVHLarE9pQoRh6Li4bEM1ndl116whT/7K18IJGu9ofDVSkcY5SVDOB
goArJhyJQOHnyInmKZrhvew2HVmTrrF5WhKvFkX7hbgmV13spgtQ5NHyQYYd/kTh3Vf6vA/ssoAm
Az9fO9W8uKJX2ammXCvyfWBuTX84Vhie4wepfWJlTOja8kpATHgmqCje/bgUdffF8bzuvUll+pV7
C7ZU3kCxQa1LxK9D1t+MuHCTA41Ow/6Z9gmKU1NPe5RpCbrUAvDTisTkWEU95/vLnIHI+j5kCScC
ntxjTInQUkza+o7/5m1+/h1+gfsUyN5zhxWuW2AUKtZHrBL86l+vqOG30E8vhBP0sHUpqirKpk8P
tkK7X1eEVT7w6K2O/BD9vR4yGTM7MmGH1T7r62VcHTZdj+d4K3Ty+Nds540rsSPhy7OQW5Xrtd5k
IcCB8+lAvRs7YfFn7V6uUa+Ziym7k3ROwoMcFBbm9Xn9s9jqYZSOXR580JdNgocCNKi/edpApJa2
P1rUnq/Ldd1beL3t9Q2mXTMSj3i8zEZNHSi3QULad7mkHeaBxE7lQb4ptBgFS9a1M7EpAZtqrwHK
VBANXQ/Y68xj7w3leWUzYR/a5VJlPqzJRykZNWt9lJJ800+7dKdkr0tjdoQ9DZvu4mdKn0S8Cg4w
RbRfsGL6pqH8ibs13tSySx8FMN1uJcSFsDxwHCfHnxI5PNG45LDH20MuPFnNZwDD+xjwLbK/pxpx
NJews79UOBersxE2f33t4x5xjHTM6OTSiebYDZWZZzGeHbW48LxmG/UyjE926DRC1sReR2WtH+Bl
yidGj1x0obWtD0yimrXjt/9xcNiGqb5Thml8wc6JGU803PxNkGcEKMYE76h+Aykcg4MJP4iyKAPV
rNWotMjN6MLaJ1770VhDn75U+GrrZelNaeZe7XM3fqM7Ug7I6isiKxQ3ZnUvuozGVcXQi8o1dmc5
lV3J8Qa4zEwikCpjx8XlOGL9f0YFcKLFSOOoWSh7HnAi09I8Fwg0KXCdnONv2VARweqZiVwmepir
UvTP5En5A2RJk9PU4TITlj+cSLHDDg8ucxvaCpW+wpJt6eEPbgXjYt8bFf3kyMauATwoHg/As+p4
ndDs7Vdg/rYL0I9D0HPZisqqY9ToBVHX3QBwN8+NEzTosvX+Jl7uWPANJix5lNd+8kKrDWKPR6yi
U8FXGwbSrAyExbTp8Qv9Us7tYORrQ0I05K3gTQ2T+dhz226iMiOEysX1kHUr5qITI4/zmGVj3NXt
hHBgqFZ9PgOLV7Vp5t67SsQdSAuxibfc+sWKSTUC3FVZiab2hVEMi5BEgByIfTEOVt7zA/vP+8XF
BuZUJoVitiQrgekemDB+8qukLUZBBcJgLcWbeAcp7GzG70O66SNeHSwgJ6dwoQ9QAMVAKuqNlprq
OuPIP1hEJjrl/x2LdG7Yqc7aEGHye3BjFkD0CxnGcwiW2gL77MU7XjD60xLxHSza+21OWz9c2wCK
557tiHUpB3h2bGvdfvXuAm31sQYMls8QaNqlK+MmD2KKJO6gzMbYBD2msa0g5FzmYnrZgW9Yp1rh
ero7CgGo8gdeRf0S4XJM+QVd4zRd2mjVyMTXX29kpYl+Dj4EV1Dg3VHIeXZ7D4ZGIxQD27k2w6Oo
eCA94aJKztzBpzLmW6jUs6w7/8DFSLXqLwjOWwZVlCdxL6hPwnQ5QBWmk6qJEe/osEhZW+oKEfP7
rUgyWN31Uio1a1Lx8wmu1fgF02jpS8xaCo3+35ATm5LPVj0N0KPuPeZC5nCaNPod2hcJeOxKcifn
AGxB0jYkwAp8kaVH2jeBNM/SID0hkqzqY+a/bM5D5gSVyQluAKMgAhPFM6Sal/i5UCMXCztRYBgk
Jy0/ACFPwuc26bXJeGiyhD3+bmAAF6tQudb+Ah0Ou+yT0JFNisdkkLohNriQF6WYrYNebNX1IUab
G3ZaJ6z6LAmGuCJtq6p4sCompjI112/DKM0+XoCHy1azNPpuTx6xO2o559ngdKavTBAosi0TN9qn
us/VNzUSiKLExQTXMWi+nzwFfOgQMh9qYAqY1Xcf2+o9/QBufxFxKR7iGr7kfj3aeBXNUTJCf8o1
rplJnbUz6CWyxLVaa+XYTbn5dLdjBMf9uTGRL1h6h5AKsqOb7ilupK8NSiBJx1Km/dFPfrwAgNd/
BHqpc6IbdphsrKHl4lHkMGf3aFdxPXtRurJiBMdjiS9IE/aXljaC7diV2kixAVvxPT4Xv2NDJFQ0
nJBVCVMLbh1Dpun514I8vuc093325OFEAXjKF6d16krz5FslOg7ZdQhI4V/9LW25U4LdFJXeC4nb
Wgknx+KJHzEfzyf3HFiiZiZJ5ltfyOKfnKsalIjDt1w0+vXItZH18sCjfAF8cyL6YRxMhqoqGLfR
aCxJVh20vyYcpO3QGb5N6b2zXp2rbjHCj0yN3l/3utcr0BtWlH/ku1PIQpJtZWueosOosfAV2/Ln
PuUsYQPdYoyyLH1o0Ckwie8BFOD/ZTTDAzRxb2vXdtIPYglyfydXHwC3tFVIg485vjA8pPdtQoi6
C0Ur9cZyZaDMx0wgN9mT059UKz4PunXnDx7Qz2LC25MVwFWgeoXrG9+q4JJB+Nwgjlb8v694wa3a
gGZ91JhJomjtx8VdIhqvxr718crTDRGLws68eMBWmQ3bRgkYiu2bezWYgzrH19LAdKRwDBVDmT7Z
et5e35w+Y1GPbTRHp4t+rTfR8IU/u6+SqnHSEcKK4xF2DFZWbHjlhawFnIRYnkdqYbULsYcpzr89
z2DkVOrHldZibSkOqcxH5SeAzBXt+0HA86zuKQqj1deBkM6KulYC90eD5rRqwslcTJ83Nq2tgS8M
iHeWtxc2GiHjbQx3dOUbmpC+cDk1/ApJv7XMa6VhkWnND4OBi4Pg0XE7oeimA2vpivoclUFa9Ef4
XieMYsT0193XMYbCIiV2dfOFTaOInNuPZ1u0iZQk4irsJHEfgipHAWGD8H824yzKNiXXUvb8qD1i
2YoLLbi85WmxJAidvvPk22ADB4fk2zDSJPE1Xh0D4iSf29NrW6TfF+WE2jf8WZs6qdwQCceSqS2H
otZ4P6WMG5kezE4zS/99ns5krQmw/15s6RHhDcZEzGIlYycOzTz7ziruQQixBV61NoavGyNJoVgs
SJns4dctcm257muOENvyn8oagCuhaTx51d+nDHh0+cBMqy0wYQCkGbJ1hcLtl1C25opnDqohlH3c
hK/AF6s54pzfS3p7Eft82SsMiqFoV9FJLBjYNPfBacBoM6OLPLWGBZzIqJ+Sbxci0jfuF2rdJ/lb
UPbALYhdGjKJi7juoTVkbWF9r4tCCtHTzrAYLS8fzYWMuUNdCLFa1Hc9kPGDLkc8OJoNirWne6qT
R9ZlosH8VWEnXaDxqfezLmpc61IZN4ZvTH1EIbosbYxxdtiR2PqcEHBrWpUgyDO/08Vl1HwPVrCc
Lr0nZ7hf+vy0G7nD8F7uygoBMi41NIXaxdv1vaW2iRfGECTWUBgUdmlaOXP3Um7yiBrhEBtS0htZ
cB++sLXylEvhNUu3PrBrHCnKPLblKYumuDmnjGLunP+8M9153WuxPtGtfxI+2uTYiP3zmzdgCt07
X8SX7YUNTzKNhp+dkDbJnUF0enXgNgoXKFFyxpt5niU5CNKMB2yR5Bwrr5g87U5itKSsHig7sBDN
PcZAU9mYIe6eOQnE3jMQvdYCT0UspcG4ebLmxs+Vuxe4atjotzx0sfBQJIVpUtm/G6nrBaOjzXMQ
aDnhtGVAM7dQOJ2+YKcr5VAZEy3D9G5qKYDqgT2bIzBLLphMXEgRrm9xcJ3ceqCq2YZWWmwy64oQ
0qYc0sx9S7y5owOBSZkr8PfqZQqE7NEajLJzNLTP6Z/I/iL/1g5Nfh8e/L9dgKhaJmKmWlgF0Bil
47XHogHJ/E+OfJMtsNXL6+3FUDNrPBuO5NMocThm5e2WapRbMlI6L+lNeX1QnNDP1dLoMKcY+7Jf
wUIainTG/edBXMwAQcwmhB7RrbEbXymB17ua1Jkcqw8UlUgkMaWCu23O6MOygZlFJ7OWO1gPlCHs
Ea36GS+p0WybuXzPOh6CoOkPwCnkvSJ9LErxOlbIPnNYe15PKdmQG/tKdExiAKkN5O7hVRiEGjvk
6Ckp4eQNYxJyDMcyq10jyqed61H2D6gE5vHZnGAZIMpy2e6zep4ykO01Rv9fVPWyqiTpx+2I3W2l
ivVPsi/PjwsrN9mxQe1KM+6WvqiPjQtAHIrRD0xfzrspOlAT5CjyoP1xKz4UbeEGrw5ScnT8kB5h
+uHP9yHVYj4f0523KqfOgrh2desoi+8zjWW37fuJ6u0X2nsqI66OWAua+yHVNihW4mO209WawB93
0ZAhSeoxJh2sLAuqdJ/YPuPf7hHe9V2C7TQa4QVJEdlcdZL/G4b+c4UC2e/2J30s9ap4CRGad4bc
3p76vr/0Kjpj/kfQMnTgE3c1O2IJexalRgYsaOYNphJ92lQoZgxrls8tWBesYLobfoA1n3y6burK
YygrtYcQWU2OhnmC4MrHaaJfAPfG45jVhzJ6blAoOubDHAfqNFwCO49h3uiGTwoql9Ysx+kt6Q05
VyxAsDWViD0W0RZUrK93W5aCOFN1JTgWmSzYj/JrgTJPe/4KhdX6mAy6WV/9MASHnHFtahL1oQgv
App/EH2uWfivipz2s2b3Sz9Pt8R6GXIxFxOIRV3M3VrztgXxQm37S32s++b7S9gGgo1rpqUSQhCF
QN4HHyg6CEv6MwzIDf49oUFkkMv0dGgI6PPrRyMMF5tco0h4/TyYfloelatOJ2ks3Vc3J66BcUlJ
tRLXq1jYCtAy3ul3ysWg4rIBP7NWni/NhTQeoK+/se7HdA698SZ2/B8M0GHcr34Z8Inqc8czE86J
hVYBnBTtYxDN2Yf7oep3ny5raB0+ZYgFnRSWvuOsxLRX4dh/MqdB585+kc+0PcGp7tDQjc3itH06
yMp4ULPNmzgKpPCYPTWCZ6NCpO9hSFqy+rhOTAavo/QFxrUv55SXr+gqmhlAksK3s87nFRYJW27P
hoVQ7oe3ZB9tlVb4vT9K/8947hfel/RAFTiTqmmzCbLLt3vYG2VzkwfRiALjsCCqT6/a29IqPw1p
TPsrLPmOBvFh53aio4Om8e4sqeI7esNsoDtb0xe2AOzMLMaafy8wqynKirZqcMLml+VFyUWG+u4K
BrOSXZzl+d1VywGkDaE054p0s32KHuuxGYwcVVO4GFFIt4aogokPxBDZ5g7oehsUPs7zx1fU4QhQ
d/tSjHBQifoegtIPH87f+7YmuJXaIGUXb9zL+OzbWQOEsERo2KSZ5+NbULY6qxphWzj388KhOHNO
/pCHwSCdrddafFAZNAVETrjw8aP+ggjrf6Au+NVuWirDzt0ZWHW4pvxb8QqqBcxO03iT92v2NVxT
9yIoaIexX4Yh22pJboZVTmlFmRqZ7XGxQNVbPcn0dl4je1QMuJ51NprUIVZzOOG93UyZPgXJE4gV
c4boVXHrkHLGfz9Qg4AXZHWF/cMOvzT05QjRuFB7D/KyCyFURibFOYxk/8Y8ILZ+pI1oj94q3Iyn
5gktAxqDOKN1WYtwzVDK8mmoERv6gxk96OlByRqCO+OJljgmii4UuytCVMDtg6rWnlHEqTjo8gLx
OyoFzbI91fxpFGNXkiCYpnKmTZOPyNgSXfxVUVVzX6fA3ysSCMWhQklJsbl0LGRfMS33xn12+Vih
Kg4oWFUb04YsrfPztVCHG7A6NKtf+Op8Mq3X5D1RrMWjTWAFWpNekRwXm8flQxpfvryEUAaWcwIB
kaHcdg1KyP28hgoJ51Z0L7GpXJreMEiC1Z95+uEli5kTkDCiItIBo07CDbI+83T/PFzRU6agRrOQ
k20+F8Aq7/ir39vYXUCFUFpVY9SeFAenD0LULxMjhCVPnQYblwfkTwXVFkh0t5bBtoyBDU5HcO3Z
BHViw+WAYQpC+snO7nopWrvuv32igu2RHyGz2ziF7b1HCEIg2aOh4ZsZrw8VhWgTydrlBJmyibmA
QIBOIliIpDrKi9TMDuziab5/LhaQuYp520EtH+2l4JfOV2C/aKKt1kgwu+M+0aguk9JRviHZbz8q
xCUs7Bm4/5FunX/+3ojSHZEc4a8qcwc6GsVxegk0tTyxpzksnBZFu+eV9q82KEgbDYXcZlKZ6aLn
NRa8CXqW3FtDZepDCHf9wAnBBpGuHSh8Qs3Fvp9YP7klwLkRu+22GNt6Z1sZfYGfbTrrZ9XfQ9bA
jtb7xlNAn6lzxzsMc1LrYMv/pr16NsecfLIhwTlyxMXz7rJgr/vKQcyp7b4xFRQG8Yp4rufdGfSI
xzYVmXW5EyAEvnBX3mCvOawMtZFR9w249F4M0/VXwPD9AomtBD8AhpxW68SWwL3vL57F/47R8SKc
Ljht3AUGJ6NNP2SwfBtb1VY1+ixzDDNmzrwI+QZdxqoAvw+1AbxW60ofZ5Pirk1C/qGRUEvDVHmG
AqWtVbhuEjo1jv2KdOTcNyUABQJFh20tibTEn9qNkL+xSgatzcd8oFCDuv7z+LQQ/GCzCoWJ7H4H
cgrtGmHm+ttZlbF4pb2BuUJDZTbcsCIFHhcZlI25Zajlz8xOJ/Xtaf7H/8s6BvIg4gjNBsKsVjlq
SkCaj8u9YzimiEehB9m35JETeNEKB29rMohfDeBU4odPiCDWBDWFFGaeOpPB8JhYk8ef/Vx2o7Us
DjKwZ+V0EgvcUvKWmr7hxgiYzA5ItsXb8vYFTMX019rMAzC0FJZ74s4Y3eHSIRaLR9qV7cvQBJCl
40+MADPXpu/ios7YvuaXpuI5ezRebAk53D36iLrizNnvi6vH8GWoYMs6bhYTQcXv2pdZixVf5ySz
NK9ktDjC4unaNq/3pdo1wqdZkq9JkTQDQD0z+nZ9ZDk+Gq+Hw97V+Oaucl24jLbJHoLf9rYDSpWH
WoBEitESYV7FA5J7Zxh8LG/oXhnMyWVjo+Hpj2E/W+M0WDilyYBqj/6SxotH5Kdw1qe445viUrWp
5IB9VVot2nXz/GUKTFozkbClhjbTaDwYosD6Bi270fU95UaBkAqp/Ce68c+aEUMOYFI6OYoQ/1zh
zqCS9W4JzgtxzyNVgwI1YjFE9LVokWC9jLDEqElaV7s102twqSzpIlFjqq2ALSGtsc6Do7e+E8xM
GyyHpscC69le27KQ7bWAz/LPfI+5kqGcyPzTJgZfXrznC2xHbcvstHUDaogzPhQHv43gIUuG4MGF
599rYQjyhdpJkxQHcI+qKKoZMYmAutpXyldyNM+iSmhYZyG4uEHPwbJzhPYTOc83R2hZVcbeHt+S
1SsRx4T5G8Ji3UHyCo/V3uC+PJ9s7d0HUgiy6C385ym/Yq9IUF8XqhtKSVsCz3avT1RHIarq0ocf
QrMlFEHeXe/bp+yf93FngclS4bDtguiQx9NJ78QfLIzkfOuerSfqR4M3TyJ2yM0oHu8U2bJD43ex
l5H5g1TyckaHmKfCLF9DxW7rlNuPEPc8kX0dfaQyxBx73vOTt4ewxOilf4AN9dIMJixLyaWHEwXv
Z3iMjbHt0mQvDMqcFXs8UDQJvRbnfobRWJWG1gBSdPPGdM9yljqWSbGZFLXTlZxD0O8l85Ge2N6m
C71Mns3g+BEI4gialdKcxwhliLMMUgU5AVndOCNcQqnYFNLlJCDHryB4QMrSvCX+lDCPpYQCSev5
nfeHbb2RtS2hYZUCEPezdJcHNEaKBrJ6aPlSOqKoVJr0sgYRFkiFByxiK8a3pgj0H2JCZqrZUB86
V+kQ4QvkCe6wamadxhoNLokaEk5SEg7258DKAR0cY5kgbVV6qJJS58kuHAE2zSxTcQcj9KnC5eZc
T+csmKnTcKm0lT0jeOUOvrVuvPPE/vtOXp123rmi74Kc/N9csIMjX6cyAMoP7Oci5WMfqjtH4EPv
tUNsk3KGODcnphANZ7JzfumgS0tA/Lx0KUK3XEsk8pX74EG6EvJ7+2fWdpBDVd+sjpD+1m8VIop6
kpe45wDR6gmiAuECiDYQwL0wCz99CJfycSXuZF0PPvf6MT3df/heaXCJdPyygtmvDcY5x+jN9EO5
1q7vjHkoV4VcO0tATBor0S2EzSpwiCm1qTCBoimcW82e9IQ0WQShdDxRcEViANzja8L2tCQgqFE4
Ku62gNWNy+X7MrS7rntgm109e6DA9HxQ162q4bVMga+FFJ2Cp46aCQs44oYn6ah05F21lC7F1lZC
gopl4LWNySyAvBkqs/cQd2uhcLI8X+uUgKk+WWkaDUSB9HIewEISlKKPosC0IK1xnQupbsUp6Dg1
4M45r4EdT5C1qz+A/TcUevQP0S6JPVdDKB6FXF+tvxRzweNBFA3fgwdc+a5aWoLVm2n8SU1jV4xT
f9oA4KlJfjcsUWPNpBc38J3qS8oKU95xfMy9ysaB1Bnl6p7NnkpMuGzw85DkKbqnRZzKVm4oCdgR
rPeLD2Mi2WgzS6r/vpGrMrF9HEqU+1tXfr7k8Er8hw1CQ1nbkiq6cj88Z+5WLQ4ATSf0YtSVZGWZ
S7BLX1FkjKJ6i1mfoXd3fwszfBA01i7GOltYTwJPg2z9M/7HrJ6ViedHQzrbaBBQvAiIlYDxWtf8
OkFWqxrt4PEmKCTKwuSCHBJEO/jx0jdSmhKHeTdEUXd65EJZYzr4yO2A90aGt72Z2ZwITdJcps9r
wQI07hAiMnw0vr4k82TCuOz3THiYCq9QA1lpYBbPivBMr1Y3/TwYjpGkGpz7J1b5vX7jEy6ghBIT
gJ439e0JabuFe3pSw1kLx7+1wqUIdv15yOxmpb4asFFHgoOyg5XIydbSU1W0ixN9dPV/XBzGYA9I
bGezC3sDlSrEnaDpQm3bqf0mAQSk+ylD1Sto61n75JOAKRMVlHlTY4iquIZbPB6pyrCG6em60/vj
+Nb32XUzhAlReqYQt3HKPr5cLvnC44Wxw+KUgYb7GbgBMjriJzbsi4C2oQfxqzc24ctyrDgV5f1/
wA8JFglk5jPoBfJPSArj6ujKTINptarUp4jFdFuVdVmBPpSJJoucLhdYPcJLGTg3t/Cg9QVCRKyR
+pNmiODbz4c4aQaUErLGRu1MUeUsqESBjH3P8Zd+A1Vn3ipnRIRuInu/9pgCIz1YStefCbrQdZWV
jvAcakojZ65UpHEjzVY4PKvyy1Upu64rxr5gyDW1244EtKyyRp//4dv9uBuXF6ovxMyhcg62ccbv
Ms0swW+ZybIaEQIYJtQ+eBZ/Wny6BXjBsMwaS4IW7grqJBLnvgRIp8or01SIE9zQVk/l/4/tSoxf
qyBb1/FX6hhH5yPcfXxkL8Bcphxh5cGNgUc7jbhNt442k2hMDPZWpA/VHABzF7wecf16CUuEq4X5
z8UmrGwr6ZwjSXsvqUES8dAJyZZpLYYUxGCG10anVEX6AcvtBj4y2aMW4aFVmBNPKJaVf8ZMR8Mk
DXHSrSnqZXRgI51ZSUja5sstfexID01tMFCLpRUi857yMKvLgB8tdR2JzrC/CXEXGm+vymLcqcLr
Yy5YhcRu9r2+/hZEl1TVnFOFQGmbebDLKrJJWbuXAKalFv9H4Y1W56Syka6s4br5iRhQQdUmM1Dp
4xQD6u/UWssXEZ3IT29+rj6/cBZIc0M90rclvGnVxnwPqSBsNcLeGO4cWB5RPrxA8NljDKJqsiR0
+L1wzEABKIQoD/licS+pgj0nbosutXvANHW6mfTB8iysBxl0g4ddGPT4aS5Jn4xa6TLywKWeCLNM
fsuKA3hCkyOyz5HG/CLBQ1wyzJ/zW7WsHyQUHn8hmq9Nfb7CIeQN/dGKbrtpIWRqE0UKvtajeC8o
KtMCCVQsRGGscexMez4LZSqopTvn+l7qE/tmdkFchjJqeRZY5i082HSyxhYUDvuwTKPYUI7pMRcI
u+yKWU5rMRr82BbmsJGp4yDcH2B6AgIJcx9yFmVw+TYmzkPLtgLwVufRvV1Yth4QlNGsPVO0yXLy
rF+5yboFgwTniXk0Ef4FbrBDvNLnrCy2wMXxfWk1iIjtUYgs8BUjsVeOFunZabdI6L3uHdSWzg/O
NXJdJ7vNUDX8D9htUS+NgpVAl3oguI+yujVhhDBj9uB95WaOjgPW6ABtSrUpr+BysuMuQZPh+Uzx
Jgq8OxberTWKDuXcepv6BcqT9Y9N3q4KKxA5ZbT3MLXiekQyU7N4+06FRm+IWsD2st8Tiw/coJ36
ffgQOF9SFhaD3P3sT9Xr2sZ35+UpJWeCEcL3CoXta3g7nx1GM36Hao3861ygHh4WRJqD1OezTOIq
6+3nEGWoWb/wP9uF0xEHfCIUEOFg8quYP68ZTrt4W+dVKSnqlrlqIzAMMwDw/1yd3zGGSvbhgWTe
BcsBx9VnRaEAiqa4EV14/z2k32pGwJlDARNtX+42LLoBAyehPwLDoHLoR73nnjeubBhIY/6Mb9Ji
pXCQt1SAd3MRoeEKbmD0MOaZvBDoxT8HJidhaUEnItwuvL1RxJjTKpDVOa2EeJdCI5Mp0286rX8n
puEv8ABvRmV9LPqb8TLbOoo1FCmbrHIE/dspbfjon/04qvXZzxRyCuzqTeU1v5JMsJd+ksyx5N4P
sLqD9EaLntVJT5s3SipG/vIHz3pWKC45yxUQ9lIaDWYx/K7lS+L7BW8wxPSey6bknQMkqz1Rz1kE
Q8wZyojgTZO5Sn/NaS10emVhe7f2H8N96X0iBp2tmLrfbEfiboGK88g0PF5IIXQCFtDOAHbEK0vY
OmlOGZe9W6Mnq840uwFgoypi8E91LvvJag2nAqQwjn/wsSBnopxgus1K6eajd68+rtl/k9qqzaRi
IUw7VK5eHb52E770KtNacxrk/7+bKJZYghGiEO0HO1q6BMHjCGvO2WBTEBfk4DMCSunDTsnf/cV1
WYca422ZgJcB7GeETzrU9fysAsp9pHo26Adnm7nYMwFv+PMLaPqytOP34o573HREWEcK10vgZjc8
GBBqIU0RDlOCYULSrMGEkbKf09bwnmgE/HcpzMayUPOFnR/GkEChTMu48Y8O2I3OLpKkugkMAUCS
+/1gfQYLcMjvxXgY4SxSHZWDj0gHFgh/owWxelvkGWDj4/Z7JPr0TlDv4jkzhqiOjlNwjtvvHXFg
5ozPyYwIRf3Nd7CgHlP+r+/lfOTwS7RBEuB5rJ6v0cmF2WU1MmrPl6+Lua5jNIPLz5nJLL7AA9ZR
DgIYa1GRwYr9zsHOwAdLmW1asc519T1hs+MJZBSOOpuNEs9acUUTEsc0bBkQaKfhcFNktOuVBQnt
Mq1Y3KJp31BPPYuNM9JnHdBCtYacmIH1leNQsJFnFAtSlE+RFiDwlXmTROk2WTS5L+rqu7I1m+Ll
7BUIJfd6PesmQWpS8f/L/CkK83SL9X0HLtbTywGuSkG2HVitsKM25nsBwUwTWrmfEDOQsk3XRe6K
+rA0BxfWikArQaluBIDEsFMQecS7YXC+ATrm/R25fy8LZPfs+yxvfY812XYo4CgIBb4l9RTIwWhx
mVOVqM6KseaewVIP90oOQ8JFHEOwOC9HNSVjLswF9M+4f7EwMCbxzbqLJDfmf9O5pAwjWhHNYXgW
ts2s/Ih0FOSUl/ZAea3IJxzM8MZhoFE+SjdQw030ugw5neIQzvT58qiv8YOAuzasm4D4vUxUPjsp
Wt4nhvTcTu07Z/2ii8NcDYOLbkqFjcWUx/yL+A5nKxdSSbRHfdh1699iAEYme9SyN/CDpUEqWPe3
SbdU7G2CtgWTOcXoHInZgtaUnuYkTsc8IRIACqdHmJsGtRSc99vo8k5MI7tJ6csvsR8wuIgAxAnY
TR6Fc9e2rA5RActFanrnsdj8gNrxGnesQJ/Hw1m8bf1nM5bGUd+y2NjaG+EJrpT6nkwMCd1Nhah3
jDMvnvyadXqx1Nv1yEGD3YJcpa0kVXDDh34wPUZWFwHMGWOviK5ZS2lb56nEEEc6E4jZ7gwbLXsg
pQPci2NPmrpnqtrc9MsLNVg0HahZFiRQmqFU+itRjGBq3U/gfLULMaGpBOxqQJvwdmuz4V0D2u0Z
wi3+N8Q2OWLCxfusxb4y2CACx+a1ARVJtos+5EkoCh4CrY3LMqOujJyxENQk/D3bYpJITyb5C/Jt
VLmP1ont5nbTOrcSaOGKArhI7EKvpXE0jhFKnUdTHj0r0oHsZh/f9+FouvYrqVt8BiXUyAZcD0VP
8+asbDF64sOYzjc3agCIO7HQye9708+bhFyo3vqY42zk4xrYvAh3ScznbKHR4/9mm0Iu9i0LA7cr
Ukz1qFuwv5qJsSdi+l1G42mmf2s/xxWziu78rVB1QrnRsqNGmLiaO2NHY6xsvlLE4znC+TAJQ0o+
uDQGqkn8LITR9Q8gRRBesyqWVOY+u3ODyDwkYZWlbtGvPoEPGgipb98jrfifRusXz09gG+aQKWkj
v36Oqmi+Se4JnNu06mGasJfoXb/OW+A3FCMh/mzka/B8ve0Eed/gs92QMRFQGCX1oUq8I2zpT3Nm
zM+PMG5w6gXw57bu8G9esBoDxxN07vzzm6aFZLjVs7s8Sd31D+y+xPR+77ISmoEJJVaXLedw9mtO
7pvWw2pWCD8tjiTL8L2tCajdD+2fkZxOUc9eBPqdYC7YxTzXrIKdecnn0IY3BZj1c/ssmeCocxBk
MkWZd8qAM40QONUDjTnhQKhdQIHYw4VLCCEBGA9PG8RuGkZHozbiyiG/70IgS/FFKtXJ5ND51krt
vLaYG4JJTiYOvnJ1c1SYFyD3LqlAGj/So07Td87zfGDcrbBx4EXjVqW/FjbPtLHRrzftGQkw2fVW
Qh/3BSf1ZFFFLuBeVp+ArMDnVQiqb/qM97T4tltI70Nzop/o6zisKez7KtAdpLdz4yapyS7XMdwc
IHAqy0VXjl1wlXInrK+g7G4XG5XVYigEeAiI0I8nf9YqK9h4uT1WxO+1SsnxEAV3tXhG++tabPdq
LFkjqEYpt0W82mO9PglCkQFd9z8Cb89Ny0e1q9/MtMIAwV66dFFudSAbItZe0wKHeLjC5Y0N9B6C
k/Hejle9LSmZuafqqhQ81zcrJx79li5ADnJrGZIWqIRLZTDxmVsZQNKIytM13fmP2qvEIe9zcCiL
FPRqc6sfaZeAmTIl++fNUZh/dM+E3lXquh8vUWoVNfhOrDdc3eWthDBVjD+NhxnJTHPohdlXTha5
8UvT6dS7YRxO0mP3hRRl8aHdu9Q2k7ogb0/qMM4JXlMXD3cTUZjv6PNZl381JqT++Kqs7lAbUCkP
diO6RUz4yFck/kkqKB9hW4sBm1VcUQwt2vRZ66AqT5uQNm0jBPfTc0z6BaDrpDxlJxagveaqvks1
bGYaMKF7AZiF3SW2mX7zkp+xZYiI2EYq5b4aG7PJIwIh5YENpLJz954PR23Dldg4EjEUYMl8fYlu
uc31b6/l6Z8B3sx/IHgiCqWm17TuuXnKKKso5YrLk19ZNoR2TD0yUTwmXnf9HBFw76ZbXL33EST0
INV6NRRu+e0aGvLGccfzyhl27RfVBGsVgasBS5XTk1ZOMP3v/+CjdI2O6C0Z7nHgD5sAAIcijasw
h1179xquuwaru2HZwzw2yJd4DEFpwTbx3OTJehIoiRwbkyK+YPcAD84fXa6BUv+/mTnLUe73P4Yw
61BMn3K2NST+dCIDhxDzuxLGIoNZxWyD/RHIHhe/kgNl2aVW9PVgwYZ4D1KTltuaT2zJQGrljrkh
0wpb9TZcGc2mjrLVdmVqaxaCg/iYhVd44sr/BZWvO4Ugi/vbcYPJxe9u17tt0p2Ku0VTCtc5nM+R
RqYOgPQ/kBx6pXnMyIY0b/4kbkOxaRm9dmGXRWizXE4BDG5DjGsvC33ysUgV+inoAt/zVR1K/tkU
qg/EvTOIfbNlZb0EVRjuWDjzPAEI7VBcpSTrMiwItBeO/Uyr4fSD6XPAjgQfIXycQh/uGjPSrZuX
xuVCbcXDndojCpRqS1QcpkMC27BSxGfSaMwtAhvdQF9ARtQAHM5AZZr5icjSP4TbpJcBHtuIXj10
qGQs0sEqI3EHv4Zhiiaena6Ws35Uyu7l97M424eR4APl3lBR74FsaPwSt6M9XMnAX9JtDog2D8zp
zS8Fa2wOgaqUc6+iVhM7Vs8C1mFHVdXPfHfqcwHsCAoY7WTANkskYuSz38RRTNUjruKm3H/Yc2UH
zBTX6qrHd3Pgu5qCN5IIetjb0mpGrvwRIBvzQEFsqLCyz8bBQwvk2PK51Ki6o9R+Wd+0xTrNxvnR
7L5Am2GZCNgKHx6oJJ4cylGLAML/RqTvh9sK/r0pk/IrI/Og3PT5R5XjTT+FVn0GbvvHNVLK8bJa
EXMHAcV3bvny6Pkf0M1+f3fxcPTGTgTFX+VMJj18WIMQJD/IokSrbiWWBVyM4IB8DyKOrs1nbx1v
hIN5QnkpjOxbQiS2RYIdIecuyJdky4IU/xu9vG/w2R4wNOsWnK2YBB7HzVTx/1la+yObQZGypOXd
2/peX17NbTFLxhNFZWSpCqAmHUhPfxSnBSvgH/696dZCt6lO3eDKG6QFSiuhcSuBbMTbEzfDuhzP
zjvPcyfuw2znnE1zzwUCF0PyZrcKRhAQm7YIOreTDsTVbUBlUtsYK0/BOQRdIZkOYPKT1ZhchCsV
OnL7BayyEeOx8JCrIbMqfeWzmVM7ZhnFDGsqGnToSBMYQ2J3pLWJIINn+mLtYSMmTxJbUR97kY3E
7fDA4cUu35iwJqlD/at6DFJ/PqUvYktA4E94b9/QEoijk1zCpZfuJg1IA0YpNNLXaatpjuUCrEjj
XsTwbYr0AarmnBXE8jAmjTsYKMoXPyHCCtFuHHUDfEuosSi2XaskV9WErQFs9PH9TF9n9tjgF5qR
bebasa7AUGxdBBwgrD2T4HYzNPWQkEc9FuYdH05AS8kqIwCdflbwQznoBRXMnTjtKBCbUYuOwND3
jIZgpe8kinUwrcV561WlJduHpNJMC6ImHp6cxJVANULt9NudNLHz7/MwWMGPAJ6/1O0Gr0UdUrDK
H3W+iav5ktq/bksmOw+dora6nhowbaczYeKr74aG7Z/U7bN258qF8XCWnnqgeDVVrJBHx5sOp466
Y/Z0gq1GGJxBIoMk6LTjuX8GxouowVDBZPm8KI40WbS3tcn6UKK2Wwj0tPbYspY1t5bKUoK8vBK9
wQrQj21up+si4nOuiVO69gjy+IU1V2kaj4h9cuqZXrCb2TWLY3lc1fa7TQpwHC/HEQvaHbD+0Qxm
fg/X8PiMiUB2/ugJXIBk54s5Spbjys78WUVRwzyw6RrtkU7owCLKHyKPe7WprZhfxX6l7im7lKeo
l9aNZE616Yh43USa2v2kFO4i6vpIN1bqdqyltxAE3GcpHscPR0qnDNELfk522r5LUHq138unAk0V
nHJu6+Xm0ZBNIKWsyp0syiwUeHf3BtYnD3sVwiLHgegJQlyOaF1xFK4SnnnNQFlm6BP3qIeCGnGx
xh9rp3AkqTALUDNVpD+LLsO8I529QSFbeZno3O0ikq3jyLCzyM2jxlTUyDM14lMbxFlqFBqtZy7+
t2IOfZwa65xQkoXQKIZMLmH1E4vB57g62us8bKmWnlWSROmVPme70FQiATg+/NmjsVgphlZ7sAGE
hw/SQJg4zfJpmbVzL0QzscpHF657AUWe88zvXDydfjqzQGpH9v0hooAVW1hrua7uuOfbSEW4l2IT
vefIgGHEZjxP4vnA4UtB+LjeG9IxCcgq59veUzFStSj9P/ENErNhfuycRE7NCFE6Es0kfs4Dyol0
iiLyD2VvC6x61eRUZKOrrQYQcjOTJOzBskQ76N6BXFomGO5jwgxtNn53reMREp426KUYRzXpdqT/
jNRO7tSy8vrzOgyLQSp0cGmjad9qFfG/dzoMlpS/Q2j8DkWjr3J9u9D65cZyDUoAKpw2jh7U3Xmb
sKAop08CZ9QjdXlJFC8VfXChm9dH8ngSzdAtmSDVML1WR+WJuoablt4CAtZa/PCuprnzcKDWiIJj
C3np0H1c0B2EubQ47cbTMJuIZrQ5AhdbA9QXc3vMmEpiZvlG6mjFgJHJ9QZTSVXyFLJ2ka9IVyhr
leNOaLpUjom6O8UtT8EhG9CpFcvUDxKgcmNcfVGWoB3i0YL9vh9GOT4idtD7kl/t3KT+CQ6B6AoT
Vc07zWO2iaVQqzlkW0u/d7PYWKsXrJwgkSHcvSPN4ELSq/eKj9PTo3JqpGyc/mwqBpvb5EOeIvWf
QdPVIYjPRSHCLTX/OTVd8hcJGiuSPe6afLfiutfSKbpN095D7tn0ZPREhbYe8an+or2UehALL1uO
8Y1lg9oU/EYjJ97dw2WWq6ETLiDKzGVhb0c2A8qql3HtX20BcFhzrL582n8p9q7ZEeVqYixxxLt8
/Rf03kqXw1r0eOc9CZW3pY2llHfxtGz/8phDT8fFCcFKYjomq18s3hZUUseib1Ecvse1ijO54S/7
yPcqEiSWfOSnWVznlYhpsE5oDPT3Na2cbHxg7iKmCm5vJKmx+NX6JwR9TqjAWqhBodnYn4y9wbH2
+jUvQQ9M112ACCDTmY7wPGxEwyvUAcVT47wBrlksw7Gso4TT8wqLX2uAimLBRz2W0vUVhGh1rpWT
nN1iErJxXmzi7DYAlsjewQT/Wqpv3Ui/CBDCc+NezqybWNgcMHn/NbAGh4+rf8YyI/VfHMqmZbeh
e1YUowa8eCfd7lT2P+dpUtSUXwieoAdUwr/IOXp6iMXINo14nJMhDC83/uTCUsfRd2BAp8GH4D4n
RcVhjyBxV3xK2DZYya6CjUZkVyY16uUpS3wk9699mS5VLHXIqNwt2JNcnRps4nRqjJwZygFljaEH
80Mkh06qftwPmbHHNIG4AXkJnOYyNrPXJJKggdst4mlUD92K1Lj9G5kWKZIRYv/ESqN7tXBgRF4w
aEYtuK6X7vKI/8NC0HaKj30lnxJfZogUzi+f1scEw8eodvVwb5KvisCWcZOJf3FXqwOkk8jGKHCn
mWqGVx1KiQSTBxGNepOyMfUCLOAofjJojSxbOuXmOkkFiCRhNVLvHMg7jYjUvltR71KDu5+lnu0x
Z9jxtna+fn+yo2lmJXJJl7a1ifBw6LgERFL1VAAPI9K1/WLf0H5TndF0iUPx8F3HCCvldK0HSh0u
XvZFD14M/WcOLpB0pbpFLlRptniONspiwQRBrhY7B0PwYFxmSeDjNFBmCfu91WI52RGeo4mNlHLV
8jK6TU00zkTABdgqf+r7kC7LBmJnQD1/GPMnlwLAJY64w1U2TXJNTxtimKuu4Xw7pLdlLeNPlMhL
JS3pLFVwK7DkEyBri0FmAQPVzWuXl7zbuGc2wb0oDEIR/B8DCCr3zIx9k0UMyRjSkam54eRF0O4O
siiFh8vPIjVT8L47VywIzNPziu2924agXEAuQE/1RVBVHlHiQzlRNKHyvoibXZfmn2a0UifaBBGz
sO7BT5aL6vdA1D5gSPwy30ttLBLe/3tH2o/HZRg+mId1lNQYU4UYeeKF8ihao9lFBNklk2tzukDU
/nODmmmIt9140/GauFtx48nTWYXeYt0CMi4rdFjuSeAcev4LESqeszPWK2kepoc+aEceqZj3PtqH
vK8wFHaMNUjdjdTUXEKzXKcFrBhbAfPtm5OpVV/ijrSpUUHdT/dFB/C8bXACwFRuD6DcAZxdMZrb
iaH1cv5v1GH0rpkWy6JqsSH8nEK2Rh8NV6j+gOJsdfcIdGOUJAXJfDTSGPBsLteo2l0fNjI1Ltzr
kfACg1IFaDwffOzpl3XXCetwUpP6PK79KmQXfFaB7UXqV4lOIrGhxGocJBwrnk+vwlJJnOhqtUch
Zl2nmOqBLsaJ62eZeCtefY/llOIuuk14OodVG6WXkn8OzC0SqKMgYGOJZzSnRxDDo5nFvgR8Nb3C
N2PyZsLgdsdDFOfnPFkUKAD8u9CS0mPdrgVw81R/mckgtKdNQxBhS/McrcmFEWKP2/ThrF77DlxM
1yV2cJ5VqKmSuxqXzZ+zrEgMfsRMh0O08xsNkG5judQWMkFl1LlI9hEsVQ6teMEISA+SRCeFPo0z
YOlzyYdwD6d72gyGC/4+c45sUZyH3NSpxHLkuXcdVENCLgQfnZP5bcW2LkjmWT81/Scq1XmDM3ga
3ebXO419/fs091DXIwEt4ag8uRdkUe0vThjveludUDels3suO5yKiJF/5+c6GLxcETJ6Brvx6h/e
pWGeaaqnimIujYRdJ18mDNGbrC5VJc7ahJSa5eAGRUWyS2MSRLR/Wkn8qcnq5g/MqbpyKixPzphe
j8rmrc/JNakxS0K8r6jpeCA9/5NHTS51Q/9PQFeYXOo/DlpKrYuTIsUkLvyedYFxnLC4C/THyKzL
HJ4L0rSEOyowvwk35mkaSFEhJomdLWef2GwsVsApZwQTHub4vPFRYVZF8857yjLCxOtPgvVJYLne
VKMPDrdt8jg5V06svc0qXA0sD818OiU1cYZjfr4OdcF3uy1i7fIVahmG/k1rG3vY9WNfFNUbFa8b
3o7guiAP2I1JSisQ7scykUsf3MUD9onyL0/Wtjj//ZTVjBRDT7pJ56YFCKSDHn886fb0ntbKtg5b
NJNzpTjyL6+ngryntiQfzIZ9eU89obVBv+ATVLRwuuoh5ehr9BGOxjFbBEGE4hET/nuHSlPzZG/R
oPX6SbEaeZdhoBig5qYQVMJatcPUPAz8GyZB0b5FOlYREpe9VRU/WYJwJwt6Vz8wBTqy1vf6LdA4
mN4+fPhLIN22BwY4PHZuLP0EflsXiMCGGhDDW+ENydSuc/0bN9/OgvEwCTZVIRHQs/acLvUmBl6w
MXtvoIpcOUDHixbMNgzh2JylNUBM5w97N8+jDp6WDg1ASA06w4W8qo6YaVz+6xcruqLhSLuS/YlL
6Ccv/QCiN/bmWDnv9hh67xoNYtiXTFtL7t/gMydVnxcYK/pAyV63Lk2Zk/Jq5I+brvRDGJ1XagHM
3Wktwt04XFAVs+ACNjzsO1XgdmdDt6sFXtwBf4jhtJGp6F9b+6BO9ynYtNMDrE1PiaOhjr6bBKps
KxrIayXElOBjZPi41n4qTP7Tpm51Jl+0gH95xznIoBTd2PFxu6pni1mgsS6CFpQ7ZX80IGNa1gkF
qR/YkeB8JHR4vyls+P7hcHmAbsoI1Vos5FUtcOXntiJ6IrAp5pYYOgMwW6EIuD5VCGECnwI6KgCV
iapDWqazmdgYqZg2HgTEFvAjfAMN9Wr0kJtepnLeHjdbvA0tOlC19hK3I/rDpk6TcRY0Zvgw5L4I
GErNBXXfsUY8Wp92t85R239ySeM3cW/46hMDbW3Rkt+c4UY5g7Pf4p3NXBUeLnEgeEe47eamAecf
5sPrLQdQPWKqoD5gTAyJ6i0Wn7jd69G1frUi8Q67GUTXAJzUbg+T0xVcOQIP+Ay9wKzbFvEWTU50
YRpeWzHMrD/2PAwLiJjHhecWRtDkGQeBuNE4nQhmSFYxczVes0gLRd9fR7aHmroOyp0C1cRP0HNg
8Vw/p5NvVK1fzbtWmSIZW5Yox14cNQELgUqxsizUyTrUCrP87bPjLMCjd99GUHHgYYLANgvf+FqU
bzXK7IcD+88OpBrZRuo2ksWz9refK8TcyWQ+NMaa32bJtWKP0VVz2rx9cxe/yMlIFaHhL12oMqOt
X0Rf4ZSVNQ4nhCVz+k63i0y4P6PTtkzbO21yDaO6pudlUz+7tntGHBZQLfUJiNr2zhz1f4LZttDg
P3uJtUoW14DHmEAua001W9O7dUQsMiU6dMffSXSXkVnZiWHhyUMc0tiQfXmIDVkBN4xdJJKapZLX
hXXJDtua7b1igFxySfe2TWiC/aMMXvedFHAdwf82FY+VpNLOuctNFvm4s72ByiYlEaaCI2KgFl9P
0wuJnRelHo+lFOVihZHB9wpee3otOhZX9Q38qhUxn8gGLkKS2rzYG5DM8ZVlhsFdiZdna68wUlmM
rLXXTkyKMyKrkLBTTdjEoVmcn1aHofV42A3MLHiXsZIIV2K5CGfBxsC+Ioc3qTfrYixSe0Yc3QTy
wmQGnqkszTAQkWmdAqGmBZ2BVX3AllwMZxipTs3vSOuMJZ6gjNagIpkJL1WRO/9rx+/o/SMQhgIp
N/0FwEQsBqxy5b5LmNYQpcHPjpez4qEY9jbXVKNuVb8d/YnOr7uoZpscgtfqUu+yAi6ZuiBUzGF0
6abURZcsCN0+qSgjqMpgZ0+eONpfwneoTqstEPZyqROl+aGzmetQOpIyrPGdq7HpKEg+f1Dyq8nx
biuamVGAfHunQfMt7bDzD+swLsfv1A9X1GZbtnFsY1pw82YStRaN+KIDPl2izgczSmg/NCmrUU73
YcHgK0k5JW8qiXvwa8Eco2S+8UnlRTnKyARUwWqaP/8rhWdVUPrE56pLlnid/hZh/dQLY82qtai5
wn7x7B3s9a6d/3Cw5WLTZ4d7DKf1GB/7Mfu2kqGs9bfLNyLc+u6WJCFfBI5+w7zSkaHcmhyFWI9m
UY5Dq+vWKJ3RwLt3gGivkelvE7P71JXsj1BcULwkOtQLVFh7KSXAIIDzGaVsOu0ZujjvMXjYTWY3
0PgFZfeIegRKTBic5RlmnIz+f2WinMacf0tXLxaqZwHMLuKN3qBWkvthQMBZvtH9gwrwA9ZvAqKd
dbA1hnJ4dx4GwDNhto1GggwStrnzryqLXTRxbTndk3A+bGApDVLHM/Jsii2gbNuoJVQsbRwnVpcv
XN/iE9OHXna/eJWs6pYbLqSRLkmMhZ+QWBes/3WcWV/aBkY4cUIlHpcu2gr1jtXGHGriMAyMkZ58
dtSBmoGpfOJTS1+zt+tLcBpqCwB+wyGP8cELtr3bwQXqq7Z7Aa6Gd2CpvU4BSxJmdRlyFqIy1osY
IkKiPnhll2Z3O9XFKIEoWYH2g9R6ryJHmIe2xrpc7s4YDoyIITgyeDmWBOOVXoJ5uolwWFEHTu0G
yJoZ891Ejd+Ti3/3fzl9EEDF6G5Qcn4FnIQ1aNHuFD/uirDdGBpDMAS+76zjf8Du+AP1TNWmUDYg
KDMvyGxArv4T738AdiPavHBmse1IcZ80qwCRSXpRj2wOjAKhqAOHtFKcj4KSpkSRJaXK2XmNkmGF
RHSl8aGWwXQZbj2V/Ch3zIeW29AfVc4CqgABGVnAMjSYWZIkhK309GcPynu8+OoXlZqyUrTbi6Os
z56Zw9DcufeC66VgDFstbUSDr5DMR8HG+n4E93/pEoqtXkzbhb0waHyJ1BeQb+k0HXnzCLQF5JnS
fdZ54qGOaefzwGsiczPJ1oEW39bbRQ8HH9a2T0aI+8fAGWdNWCfw7r4zpwWwbz0OJPrr5wXkIYhJ
UI1QS/BlT+JsJ6Mn3IUm2LLkWSDhn5lVWLY6joJhKFWXZHJDFsOoEaI23jMzqaaX2bUPc2LaXhkh
f9eqRQ3vk9AW4F6XDMSv9ouAQGNwNMb5REl2VPo6lDdb6Wqmm7sw+XDSBPYHSsLSJK52dJmjBKO/
O+v9tOgkDpX6jl075yeAaW3luvIF5J4b80/BYE+wQ3dNMvrI+GL7vCdm0xDyc4r6LHUPDzj/kaCL
DmayVQQ40O76EyZX/QVXYc27mm6suaf7bH8yDaRA6o+QPDDHtLEKKUniyQr6d+1e4PxpoQ6CBy5y
pN8kFpvlgPVwr6ocDK9UQ+t+U5Ma2edFPEAQN9yLW65eklXV0CequzY4mf/79HiIHetioiEWpDXq
cpd6ti5tTcktJfFbtX/ZP6CTi1I9N6cgoXlzAOhk8zBnR9yHqSiji7wKtYZqorSsC+nXeT1Zy9b5
PQisjT8QP419tA7kjVjRILCnOEsqEf2AgIiuBcPCaYfWDNsP//VfwWl74WFUpvHFJoiSntrtQeAB
rGPjrqID/loqLUaJe53Gl5Eq4hTjy1gQVfSlofV+/wCg/Xn8e9e3xd3iWeChKX7vZkJUCwkVzLEL
2LHgwsYgkFiMYFz08EnKBV6O2ivnrPm/bedAXcYWqzVqE2Z0nM6Odsbjp6pPAUUhl6rZS5HMDPjB
q944Z95DIR6Kh4zmuRZrBcdMW9+5u2sepCkYZlpbU7v+J4m51xhCq+v3aB2mTy6y6CZAZ5abPkxx
cF7uaN3h6aUQpt8+KW1EKgcHaMZ8qqDwmetu1T9yo2U0H1aGl06zVDCLbOBc2OoLsKKSeFZzGOAf
b94hy4tMtMuUYx6jzMvLlL6tHXq0+P8KzJHAriIDHUntgiFpUVyg1A6wIT82EAW0ShNz88CvYKOA
HSt9pmQBO3sKLWQjPAEPXGcA/92qe4D8XjoHHHL7QUdm/3mQtPyabVmxhZWSvyxOdKcju8Tcs5Rn
yLpZ0rFPnsOqQhC31FkiDmu/10ocR1IP41eXnwBQwiir+b8/O0M8dNc5g+u2mTTrgKmJhM7/lmSi
N1JQAlj94KiFjccEZR9bzpQANhHTQv7+cBaqZPYqhY9LZh2Ah1hbKT1XW6H5PJmBTQvBzfyhnEAg
r5vv2MbucOXPbPBE1o6N0z71IM0XhbIktCl6A82ZPNpCtcPveck7kHQ1glfDzMWmlOy9nUAex5ZV
PCyYUjxXvXQ6Vc7oSDbAYhg+dODvj+G32lHLjJr0eBzpFEBLqZrxacNmRjQKZBow+jxHT6gpPJuj
/oII36+UTBxGo5I2Omfk6GrH5q6eqbFzVmK7deVZCfk5pIXY+3mTai/enFm/1sdLvHpMQlrF8AR9
a6ddmhLVl8LtnUMSsCE9OQkiSm+Lw726OTpZBd5fjugy9/qxvr42stsneYPty6K3FYMEHKLSdO1Q
y/jlapJBRwvwTiF6tY6IotgtvjxvPNyANdFO79HJibOPVJRK8xSgyR5AG635Ha4bwbmIdhw+/r5V
WWxXugA7HwkGyR+/2W6cVOcya+lxuNqx/HENN2qaViKPzMux7LOpo7VqdPqjnhPp57/0GpowKCwn
Md+ZSTIO0a0cm83YbNNyZHosfAZmxKaY/3uNEI6wb4dAGMxVR75lgnXS9ybQtPTvkhDNIQvHlL4a
sk3czrECWvDAjeoXnUgNVW4Cz7BM+S9w2H9Iupuzg9RtEr+apX0oQwrhTOJ+J8RMnHlIyL8Fd1Py
4mzmucu4vPemVdvrSxWaNspqyoccLsKx9yaF22DMAnRoewgfYQKpWeoDdnSIgKkJQcFmoF8fRuyj
9ON3uVXcVqLytgXEPf9YTyIjmNe1Ug2VtXjMuEojOsKzipwAEo9XC2S1vWxbem1ynQYmjkowAC3v
BbB8vyCTdRd76uArtZRWRdyMslgLQIrG+3dMQspUIolcwt7ydQM2uSRUDYe62mW3ZPCg9c7ISBEt
39ypydn7ghp9FhqAo8iFH4Ti/DUXbkK5JgkVjPTbaftgHRY6bcvEM2iKeI/GHaiUoqnh4XFH6KXO
WhBqz4wdp/AbJn2INdZS3lgqbV0AFGSJcWM9/k9pzmM4agMJ/wOPPfNu86WaSbF2CtwTxqy0dQ7U
RzMiCxr6FCADdyD2WqeiMGW/RY32eeuHz9lY7aPM4GzcE2pr8uzKC0Iy6dqf+i/CfMI4gJ3S7bQs
8jpstepySWowSLgl/OnnsnCH8nL9J30MzkAkfwePeowKL1nqbfAA5dmWzV2cf/V5EtRdrZXigQZL
u1B0MXdkn6SNK52WZt20grf1RG+s15LODAX+JPAZj2WdxBCNmJ2scbHdtvlIJvL1FPW6qi6bRNuu
tfKYFTiznt9x/PqxFnwiaOWu5hOXvTfQDSWzaGl75/n44jAkx/nN/qw1tVhBQ2no5zse2rRnvQMW
OmFIhmuCT5kH0jlrJ5lBIMGt2nDbpsL9lsufOhCYSNGkRNcYMvvm3X2QwOQQwhlKqadlYSR6aoRL
K/rkVyXkD3ol7LiLY38IzTG5i1IDchbpzbURbmjXvuFmsV0f++bNHP6SXTpgZvRN/8OrSdBGT2VF
lyX2FORjCSuHBjUraHyVba/XHRE4edLOJ5Oh6lcWk4vyMiUKtW6WiqNYkAW6ofYGiW+p1GFKtA8E
0z09XR9zpOY3rsUwIn/VjAUIWRmP4TNyTDwyVdTLEqJwvfaztnArQOjM6l6GeuslaDZjlu6gFj2d
m68LXMUtkMBnWtqE9mA2PsfzI5UVyVtFBP9ekAKY2Oo4eRtI72C1IsH8vIuT4bbfSmA3UyyBpekB
nDjPRnUQr9tKAJ4ZXOv3LPAKuaVjwMSubkBErfWi9QLEAcCosPPcYWVwMyh975wxBmQfghmM5Vbf
d0FdCsjn6GJpaS4z2mgS9RY9TKTuzkpbv02PPu1WAHrdhpPzWPHM4KAT1t3hI+9bD2u84qwsbVQP
nyxDdAr7jmXnq0PcAK4cfE+EKA6FauhDBDKhhtC/7/8RUPxqGkIjZgPT99YRbaSKHGW4r74+mJJO
9iOw45CAvPT8VbQ0+sr0vMPDkTXOPsu40DwiVJG9o0VcjpohOECQCbriHxqqL/iBaR85Z1OgoWLI
nHmKy/EIA04RATY328dlWC8XhqALCScjFBdbHCRPOl2u/8RfOC6e8VWNWVdQnlmoaGmRL1DuOy8u
gLmbMHnGnvRiWjWhGGfzTlknWGADY9+R+UAgvMVq75H1ExgWXX3okDKjoNlvDk08f1GKj1L9B3Ax
kogRFGDP16Jy0MXKPSrJZ1K2KMJUIg7fw6s572nXFv/muIjLFnDBDoniCuTGEbF2FbO6HhQ2JLiO
ZyEBXxrjoemqtxs6tOiaJy/YL5zLG2kJ3NgIipXJSMoe1hZNQAsThfawLhNcP59BogODrzFWL01M
wFKkT4zr9psIyrYazstB2QHHqkDF4hMP/9fDYJjirqeI9SQbPuCT6n+cGlVat3F3nqq6TTO5p/Yz
NGwTT37+JPlRRfkoHf888uPnQmIgftH/Nv/kQP6DDEfFCbTWyTSlk4J9pS3e5B+4J4CIdBhShtbh
QgKYY1FbvdPfccEB8JGzAxTznCjcRUGBYl3+TDqS3qetQZSV5xmioxzWOAHXb+dZ8Tw1NoclsceN
5K9SloBiPYmQf8cnw0kw6NFrrC6e2Z8T+lJaniGN7Jn51Z+9hRJm7M6CnvzUeKef+27vdaqYOIbT
Nwxmf6bCrHUuUX5DdHLPEU8Rts3VGSHkBYHXD5IMG3RNFkMD6l1zIJedb/ixYj5kAj9L4Kmxra1g
ynI7Cf84Vm7jj+ncxn4pOIZmZnii1Vk+sos4Wm66MivM5LePqo8smMp51VKVUYsCBLHAtUGATncU
7qOxf2DkIhUQd+Kgkl0/tABnIopnI7foJowA3olcV5IpxKubQ8VueMaInA8RT8SFy+V1CFI0uS/s
REzayzTyoM5/XmKzPTIWkYdYxKkrHQUk1vR7l+SoMHgKMz6tvKnPLtLRIRuuQ6OmxnpeUynDj0uM
xtKJOj4w5ttYdhm7Hq7VtRpuCNnzTLZmCT64Gn+D5BrLbEZePJ7CdRemoHUrJM74lZVoHnVnSDrZ
ieza+wuMgdHeIRA3GeBxezqp94LSSogtLBrg74ODPsiJnPAZRtOXJVx8KseoNTVDWLNE9MP4smvv
3uVfxSs7HtVznSoB9z3gE7paTM6TFK2jjGEjuAyPvzN9zuO/siwQnfQ8iXcyF6oR3gtJwwLqZxjr
EAneQt+eovI6nwQQBPgR34w3qGgoFnCDAPDti9UmO5uXH+6isnyFZUGd7s5awo8hvMsICAGtgyl6
vSV6OApJl+sZUNC2ctJ8i3YZvYhB/+S6A5t73zxG9R4UUWyrQLdgWpZzGad1SjlJLtMqOGTr2/OL
n0a5TZWAKqNSE+YzasBQzGL9sW+dooso29JcHRRdXlP7nEDy3eyYIRFvnyihEiAbMckBWd3ZaLJU
gbRVcCXH4vloGJgUBnESdpmLO4KOsp5HYQNLwkUjFsDUcattNigobWS7Tt/8oz4MBc9vTFsH/STX
9O2uqjbz2+XDIthWy/AkD5kWItQ8cA/SBB8BrVJ4gvZV81YPi0/NObFSDR6meQjOxj3+x4zDUJ3K
TbRoS2xvgsa5LdF1pi8XmYymEAym+8IkJbMDvjWBbs1ytOiaEcv4SW8pzsOfbbvWixKvPTy/pjq7
H2Ww35gMtxWREKDRgJSxW/Ds4vChveIpVlVaQzxruyLzZiyxI0lj5bvspHFKtBTIrOFfNlHY9N5K
ZIk4eiTvO3lvYoOVQhoZ2Bam073t19fdsbBPfTjkUfGzIkuKM9H9QR+b+cL7TQt7EAOy7NR+dh6a
HbTUv72atPn4ngafNOv3MK+ZAmIzIekr2/fyZRaj+lDidbIGX7LeyS54Ilh9O9ZRPYKTZ6NMK3xV
5CCE+zKtUM5m2bcb45pa3KKE3DUaHTrZTxRmB7xrjWB18E8TGeMHGzNN4heWnHvdd2O0lw8DEeLq
mdUIFyjM8PgmU1GCaGjys2gBiYjDotnsTXCWlLsvR6Rl/Zu1bgemqXVqGNoUA48WZk9GLfokPi5e
9uEFu1YXp9qMkO1GA8hzSr8/8cw8wGsIRtqfexQTN8SaNLHPs/ImshC3gJaLTkCWpmr+ZNDiSlYW
yeMJOxAkOs9/+Z9sHHXRNAsoo8kHML4HmwnjZgCYmcKDOh+lt64MkTY4l3e2+fz9B64LeeKw/sM6
7Tb3ecxkdWOxB1HXtKuqRoTCL5ulLeAXr7Cjf+Q6ieaC/93oyszStJD+1VjHbwnNh+881llzpWoB
aLLdVDmHMZ82Im0XDYbvRkqvlB85ABMtJ5VryQmJGVzeYznqfqFwfNSo8D9Rm/WXhv5pdWTkkdXI
WtZrg5IZYOUCTJXUpLAuEUUEXNQU4YAlUNCVmFOXGakAR4kDfJJUVj+mAsoDGfyqaR+aBwItUwFS
GfyOrjztarVmooZ2DeUMBV0/aSMlinV0rJpOaQtdSPfqXgrKJ6RkpKhHwyoQJSik/xDrXmiEiuge
gROSrLypY4vHvVJI114vVy75se4mNO83NskciiTvVZyiWvYzz7bz9/3CUXGQ5C++b5thn6L0BZCs
JeYX6ptQGEbzX1ZUxPrWyq7BywwLL8J2dj6+myRo9tvgtPYnL3O1qMfYvAZ0wkEkHoM4iKb9uI+B
PPMCsSy9aMm13fAAYLKaADXAa6DC2flMhWg2Xsz+NWBNWGkore1TErB4BBmuCt6PLh7qGYoAzzKQ
HrQKxkpCR/4+W8exQK/5ktwUTTOvKPln1YTs6sG95wbEPkN9U5Ab6R0xCVxwdf+LXSA2eB2d1wCN
D87me/sJf4yF5TskeDbt7XSMPxKmtBSfsXu5EKdofyp1+4msJBtTHRoRk5X4w983OZC+/2E6u9CW
V3wcP/ByAv0t4NwJx3HqMNL9gb95a1kFL7ycN8iXj+6yHJPdl5TpGIOKBGtYInPLr99mrss4prny
eBO2I8GwDq4YRivLvVViyHnMRfEC8+y2kwF/41axwR85n+h4OLNzxI0MnI4Vk1lObXteY5+jJwOT
77EMbU8t1KMekcL9EaTztCdid6Hdpjg1dWJjHMKHDQJ4V7A60r79q2qDrSIXRqITjRL5qRVcW9uj
77Xt3qVw6/LUSOKayBRzAptxJq6kx4pqQZwWRrPE+bn7Le4K2JWDYxyE72RODQNpNcpgYFBdMq0m
nUhqgU1NumNIuR9vEbPUayqcPtVEiIq7vbOBcIG99kd4gi5gJ5/Sgvs0RRAYCCZ+FajNBkM2nq6T
K2BQ1CjVMDCk1Z1jBdTjIJgfQsvBYTAeNPRCy9lifqXEfri5bpxAJci7VOUJZzQKdUr4xQdCyF+k
bXlSny60ebHDw6K5i1ngOlrX+5u3Yw1uiWiDXhi7RWrOzyZ4qHMvYbsOR31R2dRnT8Vk/H3zev/O
gZOrEbTdPfJSKzi1Sl9l5AHMQAp//A0ZF/hAaTkzHU0ET4Z4ZftPKsp4rC1g5sx01JXr1E8FEM/m
E3g3SnJBQJj/O9FWVW9mklbDcfE1nJ8GrhizbhOkA8pZXNuwv9OfQcDHc5jZIDOEMFKham3JbdKY
qcNyIW2SdDpDqIalj55cbdw6a/c0eaArLz5QWRfuwPxJjuX4hO2fFl2zAdwyuCAWaqfCegA75gTu
mpuy8AAMon3L12Q9zeyFqmzSwloO/wdr+LEk3Y+y8sviyAJiFq2R3qUUgekgdX+ReARKQIFgL/RO
+/90LpgPHllO3EpUdYyHv7onxESFycaRkk/0G6RizxO3Kg3IAJya1QY7I+KaNm2gWQiPH9WAf2wz
mNpGi/f6UAjkya8AzLsU7c5adg+f6ZjBs9JQkMYpbIeXOPDpxqAT58oznt0esefMM8xhC/E76F0E
DsF/ZE9wxRZzn0HUNl7LVRsrXz8vAyW34g5GjujxPRIo/duC/msz/fhnDs7fbXk0hMZg1zCsXpR5
4T5JKFBC83MIg9xOoBAdwl+bVWWQ5B5hYK2y7l0MMxHMTI1NRSlTshrRrBFAEE6FPmKLPwF5HE4Z
rh5L6+YbFZfco6Nlk3BttVmE3oRzlHl4LvAAhKcAILk/EojnCnxGPOmJ0yUB0j34G6lE24E9u9m1
z1Bw6zY2pSgjugMhJCJ/I3ZTxFLFjkzrNyvbxj9bG0VV8e+JijlpNzrU6ulb/9OJ/0nmxUKggwOP
ZRAGV4g+IMkjN/cVpfjwNurJqiEGRTpEeE5TG4t9PPNHZih3f24ishxXdXJhO9tTWCTlzeFv1IU4
jv2WHQF/DbHNAhO4RM6FU9AHGkgJfaO///u4Kdafkw2G79CGQWlImeaiz8QHQUzszD3dxewMxCKK
XeKg3Qzni3jVIGgq3A1wvKz/9YFThz0lks9LxTfz4T/tFEm+bnZDe8MnqRY55WaBhl0DuB55E4ec
4y1J4b3LE6NMz4EwJ3iirVSPkDPJceXahfhPzt4Y7zOviXbrOt8IXYY8EUpY0AvQK+MmqaLMH69L
9AOd2MAWvbe8M3FV4i5eKFQIijbdWupiBt6f8x9YnextIUmqHLvyc7neak2gX8I1BkDEvDYKSQoM
uy9IGdARvBsScFBgfxW/xSEFZUzWQXf3jbV3C0j5LzaiFiT6hBBoztCDaGx12upWce4VNMcu8Yto
/evUqNGMuxjojdPu/n8OEeu6j+2NAI5e1W6SVm4DWpnHvYpx+mimW+IYX/yGSj0CtgCV2m3S0yVp
3l3gtQsMS4vyO02V5WIm2+N/V6+gcR1WIMlrb9vzh1YBSt8c5v3AFTnn8sU5nl/HCp7Z9gjxVzeU
LAGULBsDez/YDwoSk79fKmlrg1J4IA6gLd3Yc2xteHdgoxvM4HQaRNP5YOqJOlLlS/95wye4mWHx
1qb9Cev+9rbvUsj8FmNx6NqzzSq40vmmADYZm3pTW70p4HGy6Hb/y2g/TSJ1aahuY+qdVR5wQlsq
w3Sty25TYsOjge528FvdWhP/xXRqH0SOPQeAbK5HsjQb1bgmfZR0DBmqwTfe9ScU6L/GizK07fW3
7vAEWOn8gnpAHr4guZFeD4L3n5ecJPgDK1CuFKihlBgbTWjyX3uFh4wbodQXAdP2e4b9TPIGFW8Z
t5fpA4IeijkQ3BgmtCu+rYnTmC1c4biGkJZJVe8P82BWer/bPTvQBMjGDO/vFqLE2hvF/Sh8yPle
U7U3SYq1sCn6zSXEHjWuwt170og8aqJX2QsuUjb/CijTJcy7Ilbp+rFetVu/sId3aKeIgVgpDO2P
aZKk+fKQuyG882Fw4X4sTxQTRwtXQX1SfH1mz9e49q8IjgI3hW+834LKoGOinIqayjlcpUGVjYs4
TiVhGUpNTtV4TsmvUpBuwxrZ8RHTl7y1Jk1/P9ev+cyS06Q68OphDJ8+AzeZNPjsMSDZtZdU9oxt
G/4arbFdchYfbuOqnOelV7RTy7do0Q1CBPw6q1TEqZiBOnBEfeY4cjtqpWS9xkYvyOk8kz0qgqpR
Vw20b/HfVGqduMmcOoT9MtqsAUoFHD9i/NF/dMZQF6qsSSA8eldu19xTIU9lG5p6GPVjeUUEbjJ4
v0+j6dnnMgIq1xMIenJ8KDQyEshGRQI9+024Ilsl6E21jlFF0J556qDatEAz16giaZ9AJWM3DHbk
a8r3uakvRGBiSR4HrdFTPn7ZNoXs/mYlSnTqTmmKIK732rPV8qiiYnlYaXPhI9P+OoEORzBnxSU/
o6JAF3xagWOB6aHyRWZ5U+yKNLu7AqW6Y35377MLCkTKrxxUdn9EByvp/0qdWzWXQ5jjmdwHE/ME
I4llMKL0QEpP2Wanmea8OoMf7+UAIV4UawPRWMf5OAa2fvSAXNOCxctMbd4F4Y/0G7R68vvfoJvj
cyNWfM0yHPfuNuxp2ZyfPxy1lswh0R4tQ0nLDPlv9R9KNlBmLaUVlryhGrCJpszDjShqG/AcK5tt
Ng2TAkt2ANdYdMjlpULeAi5DA+SAhiAv/+sw9GvDjOHOy01CV3wC+cDPpJ8ji7H6u617oPIdSyIL
y7GDbQAZVNY2l7fL2en6EyG34euDVJZDos9XdCBlnDQVcUvnDmZs07KY6qvymMXtLPwisUlqNg6L
7up5ffxK2zeDTty8+y0uMEeZ12nd7haSThUNkC1kBejal2ZzYvcIzHHLXI8gkzWZlQkwYCBXO5LY
LXfBJ0JITSawpH/wGJj/bYfPQ209vJKhmyXgL9btLqjPojBi2w0X1LyTDJ5Xa+u8cdcs26xg0cQm
Iju0FwJhAmPz7yBeIcksK4IhRHTfqqvy/JIq9vaOKdz8dCdSRmMR6BwHD3wqi02m8lf0Pym52/Zl
D07LKTbkyesy8AsyABenfJ0NbIb9niz0KYKmOfH5O1OZ4BEtXw4ymvW84ErSkAV4L06PCaoKLpHa
AyG63gkpXbGaWPSe383Ou2Y4o3oI/cZ8/j8OQKTSBU1i40jzCHKh0eap5zzbeaLsq26id4o0bHMF
8B4mIggZXnf//1ZCoPV0uFi+wlcKW8zff9Y5pr34qsa9PIrouhUZpfDRjHohOnNvsnT/ZtWpGCPX
ylb0dIR/Qzjqoq4ONtSvFefIGrj7BYovcPPjPcOovSPZhlzjraC5rTXxsdCCqfxxmmEgOFgMhLVq
BP+6fCoVZYFbhNKsfe55XCzJLxCdnaV7e/LfqdvIMYqQUhAFu4hgXKhIQs0GXMbGJn7Rc/41iNov
Gf2BwYaQ6XNvH+1jRsQ2wNbshTmenl+N2cIX3H4NDPtKhT0vqgSx221+tbKYAEHZzGyiEGL8LxZH
0rBrAOYNjJWtf0w15/O6TUCcN02x52iW+Gjca6uEOvmXrbeK93Pd3WZbu7B88TKK8RhIU1XKKCxd
7RIy3ty/MwWnbk7swVlPvC+hp1nnfBQIsbUA/KZugC1J5zkRqKZZ8Xkxk0pmmBKoWk0AJdOesZb0
4z+3X+eeotAcj82FnPxMRyHZ2bLPmushlohMti6fwEGtnt06BF5UessR6qHpIqkgwRZ/xm/4xu0F
674kLTlUseNM+1WHajxKsdObRFY0S2fDR7zbNv6N3gQyaokE2pxrIKUOVwBg4oN21Bz2nCldcLBB
Gu3l/pcx+UQzqc/ryWS63PfKYNMi8lvc9x/CoFZM0oGUH3dBhKf65W/Mr3Q7L6Oy2wK0nIEQLWHC
FGZvcKXkZmAoUImhZwcMiZQoBrHscYRvUFdkZqzRtbLnehOO9Nukr035zpTEPS/QsClL0jTEzYEW
gu4FcYlOsB+HwgRNuUX/iGLe70otrBRW5jCa0P1hSfHiubspllKvkbnrsyYbTqsJwNaTaQICUQcB
VX/53A5/blnpmsLYZ/RE6MlwF9sYiFhA2CvkvrsZkgJKySAyJSu1SK4yie3vfwKwIwE+OIBx+4If
KNn2o0CkuvHlbDQbN539Sj4De+S32tWHsQgOmhbzaRFxzjLEk3T9KHOKNRmslcV7TDISn7HW3Piv
uvtCGiUjHHb5gXDJl5Im+V9aBQ+OCasyfm8v1oAMsd5CFZ8pnjCjdKaAsx6PlOzg61HSf0kf/Nmn
cKcQFzRkzwXkx9NWF/FROBPpIO6KP7IzvAyhPBGwzWEBV0icZ+mPcENEs2nWcKLoev/RiCou+ARi
LFBiG+z1i8MnmSl2TlLA7sl5W1SSfPTaE6YDOdKMne1c1cgjysGc+G+Yqn8T2UPad3dK2ecJBYtl
EdAbwXAiA2rwZ+1ICCSGHgpa5PD/eC31COZigqsRxPtbKfpSGKoBRtroXAYkRv0Az7cF35q8g9nV
IilytclV4KaIs2POTpnZVvFKxJyCqY7Zt7OSJFszpJKRPeoqzz9o0ToNralzn7RKZXwWoe7Fmbvb
m3rIsENFmhTWI+Vdec6ye5G7QkmBHo+tk0zaApNujyQuyz5p6hlmELpIm+/4mDEflOtPAPRdmpub
UnkcXXE2dZyUJ8qUeV82XSRkoiF3ATWig24EboPAkVAf2hJorm67eUepvGmTg+6Tq26n43ZGa4AN
mopSQEcA/uqxae7l2BH/6iI6JNr+5XZNw73O2IdGvEpxKiquPIHZw/nUdLRC9AzZzD1V2pn+mo4/
7ZaO6/TOC5RRsmcyb+esh8JyVACA15su4id+HqWJhwEgsiyGwXxfbiHzonZ+POTNKJFG4A5MjWW8
RtvzlOsVVmP7v2qXYnkA0EnIzX1isZHmFUcI1KxQHniTSdR/7t6iDFuh969onwcU9sRt47Qky7+l
TYhg26aFDIKohBoX0+Lj+RUPvUSJ8qlCtWA7KAMejW4EoaKXXFMakyxwu1sKqX2+0BOGtbE+yC+0
jg7Ym+/rFcOheDmUkdJzK5Q2Zxn7ml/xFuxcQtNXrqu6cc3y/xwnc2udsAOEoZa8rI6/pf/SEEMI
XY828+vktg+bdyZLVizTCgfPbs286vIhjVRirI3+idtjfGc8KEIiNYOejaL3viX4ADRI41VLudTD
vsPuNnWre3iwCBS9cye2ztt8SSqjzKTwu9MHscTZrd5LXpsj3U1ITzQR0NTZ+iotukzH1Fa1oBTe
ASnF7qWSInBYe9rygLNS2NpuMa94IL3IYaNPdRyvBUn96DblZvFPjbY336SJmulrBD/qndfg7AjO
x7XotgbppbAzlpUEpizYNUuz6PIVnaU2LCAYGCmiOKTVc06B4rbtrqFoq5nidgKlC3CsBDtY4lJn
s+n/Q18Sztmgy8gdz9g18IJVUIj3dtoA37bY15hDjlSYV6XM1ELyxvY/vhbSlJqPCj7NtqYZSnxl
gZ/0mbBiIV0oXs/iFB/1F4t0b0Jd6yAofI/CcKOeakyRnEpAfcoKmB2UnehDCHL1aa4o3f2K7x4L
eOvfJRBfAheBx204UfmtnEpyycRKyJPm+Jr3gG1FNMkeb3jvxKMSmFQnfOEDo0QEZiCIxjG9/Cap
ueAKBkSoLrN2mRj3dhbGI171b8egLW/4czsIDMTEEKP7msI/dZOFfNaBLIfW+WmoMSBEksU76GkN
K0D0IzFXbZpkzthdEqpNgAyaEZ2Cq1eke+3NWCiTm0Z2AJdzekTESf50bqFe9l7woZ5HgzEFJziz
8i2kncPMkox7XHNOeij8RVdOBioKbXJdGJhy/3179yUUugV0+ASEwipbZR05idaHJjEgndP2E7tF
qbrjiLFrNuy08ZhIu9U9LCQdltmQb5E7IWV+w0mUGDUhnGONWlONwd3ie6PwIVrqkQE/uUk4Tv62
lq2+kT5H7pmV+8XOqPAoI4C12mTrLlVc4+bJ17F23wtBFyIVYYDYIxm5ayTbTPf1/BObDfVwquII
CTEWDXW0raa3/mEf6lJy1irJC9cIca1AOEHBwMeI96PYk/sEnnUyBNhoJu3MvKI32AlP1/OQknYi
8nmKkfIJeK/c93VHm9LRNWSZxuKdVkzSVJi9a96we/wp95brMZUdsokDsDtH/kPQ3A2LlNPJecxJ
qKCbvU2AM/Fv/jDmk2wrjSVpuVtDSHHy7ktFX3Rxhz7dNHgi/ZPkw9D1byc2FLLJXU9zAzPrgNnm
A+6AyOvwBdjMgOgFfmdTPeeuyEZC6UkQ54EkLzRJZ8IAR3ci6qrJyXa8swLHDnMhxX7q7TAAKDCi
/MKvZbNtxuShycp3ghjNNyxfKJCoBO0LyRHyAkR59aJaKUrZCkUKNDstdoqLhcC8mcEj5q034xtv
ZXP8BtHWRzCmHLLydkG2KTonmuMwS/Scr+iEaPVk2j5zHBT9ZjBDNhHoI3LJ+FJ2rNpslnEi4d3e
1HbNNj7+fJoS9bvJzDwdrMbIuXBf17UBe+Av1lYmwi16dQo5agcGUhvW2nW/vD8lYkcJhNfnvYGM
da9A5AZiTmpZaClMWS+h480UIolK2gJ/8fDs27qaRZWpYcV9OOffR1dDJllRBKtXzxhWWPXq/MpT
e+6w+AcsEzf0vWXJokqID7mzMZ8ukQvwAMIYV2hvUfInyAa6ZJwAVh9FGcSQXOyUxJ9CDYNYA94s
HxbP8gigiAVGCw7LQ+ZirENtuIYLPnd/ImzPzy49sQFNwUHhO+wCO2kAtL+qALfBRmemHlRro35e
YXMo5APRjwcVfnxlLX+SB4qHzWMRScbLrEHqrDCu3kUJTv7u+N1XlitbWKYVvM7dctBM9ewJM8/P
I4/0Ao1iA6Xs/xa3aItw0gPih+iZiPUG9pEduVfyU6NJn43VNwEeGPdabvyh4XuZ6t92kNb/pELp
zPGjYAH6ts8y/q6C1IXDPqHRfN+urK+2oYh2q3OGc7/gs/nX6ooocbCRaBDqf1OKocU8irKgLLdA
s4tECpd0iwGu05nqDP4hWiYo5JENHd1XMVI2BG4HnWXWibrZeN7Y4quSr9DZG1aWICoNxq+7gBHT
0kNAyvgHcRq0PfM0wkGKmo4qmZCYUUgTKf6n165/wOYBDjr+Pupb0H1lHrsCSR8SIAlWv0l11G6D
d8PJH50yqYMBB68O51X+I8jL3j+eh+N1NNB3d776BK1EjYPp662eyic8OYykrbkGz1U8MjoDA4lC
asENOC6k+xBp3RFp9wFfmqH8XDedrj9m3u7dlGzaOUs5VRNCtzKIBXcK8MMPhmgSpboeY+Sx5UFO
A0Ft5+qZiyCSNbBq/2O+e2eA/Q9JvwyzmenLKppd2p6JNlQiV8Ns8ObLljm4q+MhYtzeyGJOmKmv
nQCWoZgAtT+ktnIT2xcYWmg8in/TaxOo4eNNjdlZ+kkGqRt0B1ciic9XOhcRXtvjB8aJQ0cr4pV5
5loWc2XkUG4/vOU7tiK8UGSo56++6jXOgsydXLO7/XBnt5G6KZKIAXXHbCt8rvP/yTvLrH+t80ad
0LLj5NmHwEuvhZkT05XiHuvAW6E3bqarEsotO9keAqVEa+lzXIiDqHchok1OdSeuKGX+KlXzNCyQ
jIbO1jGOzve85jwdzqWuAvQ3iM1mnXsvp/MuYdmB0juTKXDCcrEx29sqY1aNiV6AgdH1eJrk1nUb
51S78BmxWM54zT5stl+QVhFq/3D1qUxpNWNWGU8DGusJyVbPERJW
`protect end_protected
