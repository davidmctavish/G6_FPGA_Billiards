`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f6Oty/eDcaGLsYq7HUHaI50CR3KddeKCWngOPrYzxgssq5w1cJHPpguHxHGFdy9EIfCRoyTbcbsJ
kzGkvWDMfw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a03BS+f/GVrEwcrmiDY3uOfCIEA9kNUce+93LLKYgIl26Gpdil8/WWz92OplHD1bpM3jrixYXHbd
BnEHPXgKM31RhVzuk/5zfTmy3nsu+VOf0JvjM2HHeNZ+jgbmWrZzt8xEvN100yexT3qCgLH3sVTa
mOE4p/RZ+r3F8M7OokI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nbUiSMAPmx4Uta8/yPjtP7MHRMUGv9u7CIISzhQDrv/X8gHcnpa6/8ubhCkNOCj54n3b7Bn8UxBw
+F7p1GRc4oCPtwT5LTsoeOsukmuqS930j2k768KDUIqcoGPiZzBIaNulEraYDQiC2kt+eRpRPxMo
JQRN1ZPr9DnZM5uZxeQoQxd959BvgqoC7gQakDUcu/tLh4AGSNRqM19H0DdzEj8/k3/9oepcPo0I
DJ54cZYsEJmPZHTsPMmu0U8sU+8XKnOZkHerSO3cg6Ic2LKtKM23HBft8jb6t5JpiqGR4UTN9aAV
zrcmnFt8zpphWudQkN7uqB2eI0Is7l/qdNe4Xw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qvcDy9pMQR5dFHlKRINwzCU6wJ4e6PQXbV8+MnmLuLNhgau1fKZnkFgiRwpyf0UnKN1PEd+ix0Wc
qmHHsPasKZF45LKqdY5LDM9mD1dWGBmaXOk6fsImJSTvf/EHa6SN6Cdzv2VDXj1RTDAt0Nhgm7VD
vceZGP0d8idcHL1sHo4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ORJv3ey9G0h5DSRenT9jsgEdHTJUq1G3USaqvu86Um6q7L7Peke8GnAN5JYozuD9HwaZjtRqcq/R
VtP0h+69M8H9yD5YTEYdsXkqq0RUXuS655hwWJ/uekzsap8YiIJRh6d/s+hDPz9jUHvu3GfIlNIA
mg0YXQw2enlThFsTR2ezx9Rp1MZYGrkGUy/r3GbnT7gmSNFl7X3Q7VV2Sa2uwghsGojzMo0lHUqN
4LN2HwSfUrpvJ1/w8mLBRdNyHtTBXcqqbbbU/Yjq0lilXdnIMLuM4UwG1F3EANSbK0hmYN6o0gOI
EQZrLP80jOpIgS5jgO4vLdGh8aOLHOe6FIfyIg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13712)
`protect data_block
znQjYNS3aAdNPe8VyLh/OvkxAa8F8tNwXWMv2jEuZYf/kECndfl7uAdCIVtS8KSCA/mTIYh0PWoT
TT7LvrdwX17Y/QvQJRFTXMYG4z8h4AqkVV1AictktC4kUiSGF1ELVXwcXZ1gWLTzFmZLt+kwq3gy
laAcwTsO7uv46nLVLBJN4N7BxfXKy/8K6rKEJc1FzUIYw6Kia+8NCgAucD37QawSUhfLNuUpm4wm
aE7jobK7b1LzZjkEVsZrxGB/uj1q45YiTSzQM4VgSDE+zxESxqGLle7Oa1Flxvewe5GGMmmAqksa
cA2VfNDLkZpK28SyvBMBU//y0+kn0g/NKmNESV0QDeJRc/GJffeVFUzL6/xwTb+bmO7xvG+iqEtf
1sEke/Ugx4+Yy6FV2szBiVXO9ByCVe+Yej1pFF+lT5TTUTNWe57BqXgzQNUTQSKCDMuMjiZ5BMfL
6VUZGPol3I1KHHDjlLyyQkubSb1UPykHiM4phhsINxAYnfWiZgvlNgY8lGK6ADCDlK7jSLihM1la
Ghw6qOiVLGRA5QutLi3lzC5291eD2/ViUxeYVRpE+6L6TzPqgGsbXftqGChTL1uwEMXYoOHit4Oo
JJgkoihyDdU9y0CCtWrTOBOVjrFhHTBu7c+01KsjWYMpi7MsKAySJpaz66sXgkP0s7uaKLNOOh6x
/C0QY/Lyo+D237FXTI7hsD+6t3dFrql66vbuDoDGlUXCgroQ/dmR2t7iA7xztvQzka/W93S3j6bB
sh5n/DMKWbC5e+lJbER9cULgXQOQV2o+7EvBFoNOFsFApdx0o6/COMeeb6j1aqfrTz3ZsU81XpJX
tXrTVD1q+vyX55hw6jbjok+5usKji53//6Fqhaa3z8YeKUw7sMUDuPFsGboAdiXzoPpz+NKHPrwq
P5tEKsgeb+/x4T9CWph4tDEUdBIrf/uGWu5GegJHveUu+flp47T3S1Kh7+VWotMTlokkmUFvyfcs
4n0AlyLaenFpsnVmztkyg4k50tp7YqjLLqLxWLTEe60nwn91DV8Y4mPeCfFE+9FRbt9c4zIHY5zR
gpnWRQOBGokcP+yqQ9Fh4OPQbkb7JCIpAgaZL6TS3wMUJFHrdMlXKlNIqVbHw10KGVhhEUdD3QR2
Z8EfGIa8lOxSa9Vew3SrSSAyHbUcZe/HDuwJB0BHsVowcFyygyFrRWyCfknF5RY2lbQKwif6/+BS
lDveW+vfy3BmbtI4ne7U73xC7avRA9oaXrhohC52o6U/vTAeB3+zxjdbuni1Vg83tSs/JgYm7gE0
sM3rUT7bvcEnTHRVwDtGhxezl7KGjGdMmGVUMJ2Yu/qruvXjK5iDOI421YzYw7EsP15or01f+2F7
l0eOMdcTKi3DIV+9wFn6ekq01/mfFh59XLsnomMkMNQEmVzXVXHYdh7nsiDEbIY6ZLHoffD+bBia
bxpRRL8jCS2Zo72/1Y4v1NYjMSNOe/2jpOTCl021mOqlCxZW2/HJdJtL0yO9FpaM5bJkEaarqu7t
F12UZ6SakGAAiD7HKU+bx40v+xnnvJWnWpSB9TZaDVVFaQcJFtZQTw5VY6rhhkKKwgddoYcAkwuO
GKdthNz74UOmYbbUChnMCALA1UM/UZWbbcMdL7JjtVqrarIDG7sepxLsFktW4MBcxpteHsXQAg7F
uEYr+uqlFqlavedFnQy5Dj/Py1UO9GHV1YNWRI6LBjqLShPMSRTgFhzmQmWjgF8DQBeb5MerX+4X
KWc9dsn6MbRfYHnZmz2k5tHiF5D76juILuQfATDtax0vV01k0XXNTNQHDL1lX7mhtGBuUFleimQs
q8pSFGvQO7U0KkNsTIA6/PyD/MAA1V45uXTb7oNFE6yR4oyAPhGjv5BGfFAkx5yFgacIT2PtVrZV
OW6DJhULGuI0Tp6HynOSOWAUCUrep5GUv9vaaCHSHVsOyCxBk3pbEjeCuf6C1fX+/4OmGqQEJHAw
D3/IfE5cOu5+o3w6qzL345zmHLdL+J5oYMkEHZm5nFHkT+UZrJPhbCUbUR4xxm9H1G0ppmm9NAan
JiBodA5WYe07u13suOnaQntQg3ixYoJ1IjD2QX4t3z3Sz0/gmLei/fItXNzoPyYCcYl+n3WEASIf
ZEScE6mgg2agK07RvCIgOMrRUDUigL8idhk4HcO5b2J4YUcDVrJwNUpfyzVXjFiModBvqyU6q2kl
bclFPHL2Mkju3v6yLN1l0H6Sl+UIbLjpAIQAsqmQuICtCXtroM8MpFKULNtygQbimnI3NCV/iDEp
kQ5XqoxNrnsVjp3++Smg13E2KDz4hnyV1QNImGgaZSKbhwBYcvQp2SD767ox0+fdyE3qRzN3hcBa
3PkixlX8YRJZNxJEu6u73hN/YSOATbxSHzFJppkTcFZHx+dQmoKCZjgDzxWSPIIQXEou4PI3JOgE
POK9R6aLQdswBxzSy1MSNKj0nICQtE8X0zcdRpj+a4UqNW3ltbTwNP3bIGClDmdACETloct7U0Bk
y7Ya2Cld1tVRLwK/Ldrg2fKIag17zcRXNjMXwICe+f57scMzEvGY9tTS9WApy7mWJEP2wWeodicb
do+x7tyAVTBdrW+WKrlctmmKuZkA67JhoCFcC/IGI43UBcQkWipWxjc10YVDNOwCnhN+shANeGts
8NfBp3nEzuKlMNL3HD/QOmk5OTSfWmH4/GQ/T55hAm0gH2Fvvli99Btjx7+MhuBlA3kPL7ANxGgC
barLIrYT+L4Zl+exStAXPFM2uZbJtdD++wWk2eB5mJOo8OZ9k6NHfMKt6hdRlq4PD5WQ/xCLWXht
4+2i8TAbGlb9X0KxsltfOM8G6KDJ2zZOhORRD4iJlqmfvon1mRQiKDTiOFiDSaaoFuXSoIALKW9h
S0onMtnhjoOOLD8oQDpL1RBsAK1hSYgyhTu7lBZ//4XWRcdG/pHXLpNgN3HUYU4FH1ZQ++KWIRLH
wXcIEBUD3lXeGicAGTTxnNuzvkHqnj62Ejt1yP0U2hVvOS5bPbkwJkDH+6ldkmNI1XSDqsD1PC6y
UfBOrj4M12PQGwiC0SnxcfN0x6dQEslVniYgTq0VMRUf9xwX0Ze/M94ReKliPO4nM9JW9FdJr2u4
iKpUONXDP3uiCLTWe5G4Ph66tk45wtm+WOt2x9qpUOM5YSEGkYlcgIjRd4Qljhesaumd4RySr7oC
k2VoMm0lN9ESqFGPTh2F7polporSK5Jezi+Kqyp9V9j8HesZn32nd5INBGc4fchCDGyz30LNZF6B
iI49rLloBgvWjsoi4FKuPNhoG7GVWobHuGJ9WI3ojHr16EE7xKyaekeF7jx+5mP4840sEgnv8KuU
G9ESEjcsLbKkAPXY4pXvSexegmwblRaECLnNXfRu93LrRMLuUGuRZizrAZQVO4eEZVkMelXIzRdN
TQxO20IRBToKqWkQPsFgrhs7B9G4bCslYq+5rZkeaGRv2+zox3TYFCeJc1crQ421y3alTA/IaHB3
Exdr2NSeE0AC3QfB81TiyIerrLoLpwNngHVfPbXgq/CylG45va8b5uBMqWGuyhq/6dm3rb0fOOO4
CQX8PLtQuIpqLwmlQ6gOo921qqPuPmuULfYJST/e3lyZsr9C7/jqMBIJ6w15z2h/b9VV9NSiwavb
V4uWLJPuyo59xWCyuMGoCXMp3gx1Rzp0kgTkQCvr5HLoLE75qimfol582BmmxvrEp9ExUfNcX9Lo
eOkZtG5msxxoQK5Foyt+QObz5nHCOlaH/pzUmKaC6KgX8qzyUcdd1qOhRDtbm+ayKgKnMViWPR1h
GTl0rG8r/+5hwa4Q3Yh5+6Q2je9T873L7twjyN7RXppH2I6y1GJvijRYXpkEAuNxMB5dfXqTQkiu
qlw+qeuqkBz+d38h3mC00ai1MZMwU83+xrJYsfLbUv09JZ9pfvk1CfrgS7i6BCAueuO1/YygQB1f
4LnLqeK0Bzu/QhkMy7xNSucVRg1a9FXGLSmodfc6sY/IWLvwNQTC2WAXf+7a2hgeRvP+eC0tj13o
yD1GMOkWcdGLd58I3HKyzN3xFFK6nHVnAbCmB4DRKSbtGvdO5wSVea2nEMrBLPsM/+ezL+A5aFH7
ngSMn5aiLfo9Gjive31QCU5YlziEGtjA+J+awGmhmszDAiBDaVKQ1KbQWTASNPGJxPJToj3ooemy
+tcy0FIPFsML0W2hhrmatbfwUIxIkGe5N4q65CznyWqedg3ouWpsr9kXoTMM+tK+792RM6KzJRpA
bstA4ETO+PtXr5KdloqW9yv0KaCO6FRE/5fuv8JnWKxvcLilSMle1J5YEkk9fSvcUS/ONQ8/evV5
UPJeafvTGcqmxyj3Hjb/xoqqQZvI8vCmeRISS/H1nImBr+0oy/bJomQy8vl0bNxqA4Z6JngOwvw/
LQU+boYj+okE/v8wST0t9ejzEd+0sHnskJXobmZuiwFFjmjvNl716hyfqfoQ5twBhzWWGaO7Fy7+
SAC8QtOW46qnTPyqenJdyO4Ucuge1Nv1sxoEsZdccYtFZu++PC76RPd9XZTSIOkO06k92X8z1Osa
cVtzvam4qh+sI6xFvdAnyjkzmz6tkO/Ce1sG+yE1kd4y1hzN4z0GEECjq4dUoWAMR0TNIKTBmOaj
87lEZlesGDZ5ITJ0Xow5gw3kL+U5a7iWQB922JZjwOdckeAvFQX/4zy/FkzxGCiQwP44YCrkh6nZ
5Mx1eOD9g9NXxoeIKYcBCK0BNWqClfs6Pd+sKnIKXg9FHXVqS0OhX++V56h98/Pyb3ZU00H+bhzs
U4ZBwlxFLC42XYTeLUb2KGfB0m83swOl4eGmBxgYQhgW0/5DKRZns03uvuyxwCHtHg0eSw+O5ogj
5JUR18uakkki7xCgEPtqP+ZW3siIMsAJNkLntFJ7WLYkWOMfFfLAoQ7Ys+c9GPsy+oJ8FbcLuNjm
F8joiul1MSXcn68jRljwhemJ0C+d1IeQSTyKbgaYJnrn641qWuIS/p19Ez2D+vmqQhopgiWAz459
nRyG+l/2Ktc8BYFjA78jQM0vsvzihLcT13ATvafeBM15i7RkWO9mB2EgGtTgnvjerzaEyvqTv74K
yxPc/0AsBNHZ9od7aZDlmPgK2qwGsQm4D1rnlIWx6ZrwCU6YnZY7okWf0VWOLyyJAU38WIP0eG0/
NxHslh0/GZjEPwqoqM/6MuB31d9NN7ZUYUFBg3JRX7vaq5hbNSxur1iLH0iGEUY03tOqwUwdHSFq
p6LD7AaK+iT1Dx4qfYucpcPYAPZAl4DWTrAgORqP43x6rUHJJ7N7tnCDMiwCcci1bt3EZy5paLik
cD69OFxgYbDLBgSNhpvp27MHcKvDHu0ti2ALIgqacsd+7jPYAxfkkog/KjMVnGNb3oirS7KNLIyP
87TjVTnZv5J6v8TDSWWqhazv6rOywn933rIt0upToVW5QU+PSSMjlnQuPOkLK409XEHdYzDG03fx
6oabCcu18qansSIibuDFFriZiCdScJ/pPqaNDpXVsdLHfq4ZDfvrvcZgtCAKKAbJw8U5aqfNOJ5q
y/gqTrbvWR6HdDy9hqaAY6nfBXpXaHqd+KOqxXaWopvdXlJjQsx5qRIZJz2Hc0MOTDb0Lx7nW9sX
6BYodMo9EiYioo40SecBtWxnmoLW2BW9PYTVtBYRLRs2Ghfdi+4wZ1qDG0EtJODD1StLEPmo2TQH
FQ9GkWAkEoUsntNPFIH4ySO35X7sKCLocq0eUW1FqcMUInNUUPHXUJa5ePwBlZ61uPg4qq9gQXGu
YDPHU4EOLnCDyxoF0+zse4FkMapd5jLbP4YYUzs1cObrvJ21QtMFEIuBEGSU9p4bFicKoX/Gajhe
Lblh4RZ4Cdb3jEKkm++7WSwcjo5cTX/sxRXFC42vC9HXveWuhy2qcVUPo1pkpEg7JYLo0QKtL7Ar
t6IYxOa7RPjalA7JG5PYAoXSqdG0Zpzsn3MKAUJXP1UaJF0GyjIF8HVBKddBDqS/24owcS5kNCiH
9h6DL4dQG66JZ7AwzLJZ2Xs9JGu2EGL9ADFOKpPt43vIJX1tDvUY/01MtBp8nOVHkbWjGFPgv1pS
++51AJePe9Q+mHw42RigXt0dXPRRcWiK4MhGmTMHAq6AQ4chk/1SeU5tK0Jx69OINYimmlCfhDHB
iuP2pQmH2cWrLT2LFK4knk4AijVJ/7pJVzSH7sCldbpv5Y6F90dQPAlC6YahI3r9v22VVIymBib0
15H3G0yINeoFNeCwpEYZNccjgtNz4qze+jHoHyZva6LgtG/7w/A0l8N9Rw0wipmktwLuajjrlqDh
tIkEPTbMmk7+FrPHkzEDMDsOdjz1keOGKE4ByHNgY29GKuz51LOJZZ2CbfZDf+ZfRdrWuCZ6YRQD
trqVjmhUiVH8JRpUgxhIMdJgIofM/DZJ/4Ce5Q15t0XXtMg+tl/t3lTqg/os3D9JTyW9IDrAF11l
AD1m7KuF2sggTTe+mbekMOpQnSacgyblCoh/gxMuZQSPPMg27LmlExS9VGUCcPsq/5O25PAxyeZs
WGfGtNumHyzoO8I2Qwm7fedIrv3C935zm2nO9AG0hj91oR1PiKXosYks5t5QDeb5VQtzkbYqicMh
pzxhEqElaOfKzwYDb3RTSmYjIXR6hJy1/Q2ykVfh7CrxMkbK9ClnvE/JfRkJprhzjngNm0pweCAt
2mx5hTiiXZOw+ukbwvwQTqFIpNgWCJUmTMnMYLY1vdhF2LDbGa7c2B/l6yKdKgiV/LlgQRohPQxr
N9RMN/0PhV6FDaPPVfAMrvx5oQ877uCyBEM2vJBfCpRYGbT5fwdA8V6mo+GSU8fVav4p2fbNrzZf
4dSTrEMq23zmd8x2rd1rv6H960YjRgctUjwMkG4AeDMua12I9Mea9uF2J2Kw857H9NFK1scbs+zX
k1K6eG2T2CRiR0aPZYpobRO4JBt+kRB10yCetpSDQKJ7X0CxMgbu96p/mLWT0fzReRoGU3tcYTaU
ofQcZJyGajmsg/itfHtR8gyeZ+pWhlRQoUxaVv/OZgpF3DDFT0/S0Z6/osF1hgymnH/sY5kw6Wfd
nOrOR5G+gh8zIAui33kSWZBzmJoXXorjkRG7DysofJRW74QUmGJUWF1SFautoQTEHWuLKpzO32xL
Y/mTFglhpbFB3f8QS8xhsl4B94uU3XYMgbzgkPVhHj5XOTBeJp3YA+nt/44qhuS2WcYk3AMXwq7B
nupuFFEa8Mf2Fn6m3KJKDzFr1qre4vmMeAEn9bjPnBggd3rlgEbwO8LGyNVHciV4jbtJ4fxbEOXv
Nk9Gv0avpt3v3ZfszE8hQV4lYM+5jRlvvFamBKUnka+VTdHqWuQK9NZuCeN+HoOCh9MRAWYkKrO8
D5f3PfkFnhx6E7LVrg8AQeKi6gc4IIlZByPQhpw5phj1XDdwETrPY/IcXPAOCHZxK47mg/T8IqoY
5b034tgDlHQHLar2v70/vastBwhroyWYReXM86eOp22aFjUqlkF2b/DD4SE3xOi349V/swW1JIEa
LEf1cr+DNmxT3yg7CiYfT788pe5HaWG4+tznBNOcUbl+CLjCEFXdP4UN8aBBTcVb+q7s0V5/Qrkb
rbM7hqUDlblWWj8AprR4Jfi6DPoalDbabB6yNb2QG/4bvjNUBWDUtjdxWl1cVd1J8GG4ItYrdA19
M2B2Lkf19ouv4J5D8FHPYkchoXdErVKOwuirNwzX0JSewTXyvBbkYLgImFsmpJKMevJY4VYwW25t
KsWthsONph4M++Vmo2+ydiwh8GNWsarfOTHpku7VvTthnLOin006rhk/95OKF1oU42Sjlsv2ST+A
4Z4wzxdGDvPE7R2jzf8Mquy4WxGsaJKXPrbaMO/91DJzlgkTe1MMfONlmVv2f/EfMxxJ3rAC0Axv
YNJqaBZqV5X6VuYj5oevE1hHS7pI2RlO1s+UA12LltHZ/qatlxqGbYbta6+olbp/I0R7bkyNoG79
Wc3lH1a+1z0Lpqfvosv1jKCSKfuY+ZkgM8NeHzOfZ0NS7ydNijmxaGG14cHkWbzQKOkwMZfqMmcr
6uMsxSfyEl4HXASx9x4Y77gQE1Sx+wlL1IwYcvi46l2FOO70WjXvhH97CQr1X6aV1PsWkIbvm7dt
zbqhQDaYGbrTzxxvqfl2826Zd4ctAIPO1dJBEpkmCvOxE/jJnIFkoRpqkqybfs/rRtEF6GW2q7pc
+Ti5pyC7n8OhHC9Aat2aE7jUJZpNODM6zNtU7EvkeomNBXRUEeNv1LflQMxp0r4U/fT6ty2k9QRo
0PvmsuOE5kuzacrMu7h4agOH7lspT2zO/L1E7TZWtSz7HRSOitKLTY3tCbMjn7MgxUFPdpPt1PmU
VqB3R66IO5VnatPPLg7fD/ynemzfgvG0/TPntamAW+xaEjX8Qu2+ntWiwdts/dcwEcYqzTUJ93ix
dOHZdlYP1220MmbYovb4Ol5PxneNFNQz1/d1rU8zNg1f2Rx0jKzJ28ux0T3Ieghtex3EGkvLtVh1
vLWsyVMymelmwOAmsbyxgZ7vLj7n+uqcdOqELKXWt874Zxg8YNh3wlZA7p/MgINJ1CI9fT6DpZjn
V3YKsxPpsepYwLsbMmoP5ko6tadbYwT6FR9AJJA9KUWwkx40uS+4qap464vM1nkN7AxroLAH6/ln
fR6PoYYzKxo6/lK3R8NwA/CwHJIkYpcfhfnWPGpp83OXfER64xVAuGmXxlNQeLgKFScTmV9vIj0/
aXTUk3jUY2VNK5hUrFGvXPhN6HBHxNouzU04fXGKyJQlLCt/RqwtzeuBXVm1B7Wwas/i8kT56Wwn
aAF/inIdgQvCeT9XTLKQ4IQYetk1hPhPcUFiiUZAzk2iy/IQLNtgCd6RWiAnGaLqiwRhUuRKQpQ/
liFExfwfwP/xzmw85UMe9ohqlnH49fHcj+eEo++4bvJpH1CFZ4rwKmesLZpA22QIfkeYuWRBsKR8
/U5yBfbeGUfoqn7DrUcMuV6aQq6BlfW9U5YD04P/NJ/5nwC4K9QIJzkS/h4aej2SlWVdK1zdipZX
kfL4JgJIB4kPjXnzNXR7CVFIJPSU3DlHUDxg3CSqp6MMemeP1nmUYknqly1lm0UAX+za6Mn045Mx
VlsSymoTdCqTyz/PLBbRaZyMVreP4u1dAqHwwCuORM/ADRCev0WuEKf716ezRMdDLX9S9fTqGVSU
AFr5HpgYnlSDpKLh3Q81uTPl5GSxz4wMwT1kBeiKUtSHaN81WH95JWekbp/ZYJzAiwah9EdYHIru
uyieN7N81wpiJJgJYPXxL4+I3Ms89rb7JpFW/gOyxBp/i1suA3c6dw5+yiNKMa3+9FVVwjX9ZM5i
Ox9Zf29uryDCK9eslWdrg/f3GjXgCuIRgxNnms/HWr7ctKMauqF4ckTXYT8OPUf52ipVgdUjYPKo
ww840rTK61RS1gQU394bASUOKePrBDyg5RZNpLwz9HTPxNFEJ5Qo9V8RCjzgfiURgwtewPJrBGrm
y5/50HUKxxnElpsLWHSsGni8pWRWw8Smwmox+RWm7jahKYTolxvAmsfl8uPoi6FHYqKBhrJpNN2j
u5+34DYjVgsW5lRriT6kKbwpe5ZaLo83bJzOrkEik1G3lGSko6f3cPlMic3H+0UQpFK5f1kKH1dv
ui+FmeQeTNAlOh13LDdrl2PfcPf88+YMJjDMyMzXXk5GVILlajwxJWdUT//um6yYp+jr2hl1TO0k
E6XS2Dde0Qr6G9NGzl14npipmNEGqTi+MDRDttBfUSlXlUtFJUwUsn3/nbJT5JT9B/knee3mjuB2
gljrkzv+tYMBSSZUIK5MhtmSuKGxhwzPHfK4LrW+EgYGjzcNh9c5mDZHhVD+Odd31lIJVX0hQOQ9
pXV02PF8bqvyYWBu9b42adpKo9OVsI9buzNaFMPzvOsuvms9OkzfaUTOpa+vJ3fH4HSvggouo7PM
mKHF6zN3VXht0oR1ZYQfMom1px7GQhwkl8TR4eWvdJtnL5NRFBXXj81WjeWJWeXU8oA+vPd5swi0
aHwqRxK0OmCRkLk5c6Zk0D/TTqS48RRoj+yG67QRzeVtqUNer/hrWOIYN/qm1EyLBuEPsfgLibn9
s+az+N85CLZDnEsphFEB0XmO4ijCSBJagvBX5lYpeeUaoyBscYICTusB/CRoNpHRH41XZIM8rquN
PKvRsCoJdtwfRnVXdtO/ZIM3WBaZ35LcHPJrbAL1Dizt5BGkxzgq4oKwoGeqZVhuCKT1dMc8jkB0
YyTpGVEe3FHIvDoSU75DR0c9SH7r/VPh8XFDbRvadup1LiPeHeHVXtEQf/J9fslXLI+wIb4RirzS
ve3d2vCvavZS4VhhfBHkspCL1uFaCOdZZyZG0fVJ8fQGx0hd2z+JmryS3Et42RPDDNTpKjsvBdg+
yI6BCUSQiN0QFX21JpDIKJ5hXOyiocUIHgvC0jsTpsPJ44XpkptLZ20TvdtaytWCgPwRPcnCtlBf
CXeCCw1sRXgcIXp03LPOoFvs37vbcnLMNEqpInWSYrimqTlIH9oeIEqoAgHKBG7ZS0zqt6EP9kCH
ISAEUoWJ0yuH5AYZ8m1THiaDaHfTyZDVdbF0OnmglTA34wmfJcQt5jWmAqOY2Fdvxve4PBbjh4Lm
5+aJjukGkVeYXpyq8x2wq4ljVCeLNkP33qbIrzHJQSPoDdVy8yLilhkaygvtEDbtZ84b9EVn4zQ2
S24hFVXV5Mg+nsL/byecTV1957DbCUBNlbDkv/Ru+r4FC4ukPs353RoOIvtN8RuzrOFnmoS67+FF
adfNIgNoRBhpxQp54amVzR4s4twor0aO418JqlOiYfA4qdUZ43xulTTHKMH4d69C1qV0OtceVvWp
6Dpm9tu9CO1JYEjyxE9hWn1AXTWYN+h2LFeEjrsuECy3LP9fH8Uji2K3nCAoSzSTCNtDgICsainf
oKkKuD0wOPlYx2cpaCQ26G74htC4zMCxK0t7BwTcLHRc+/RHYsfHAvDfY1ZGUge6m7Rn9gMQgWjZ
eAJKir5x8R3uutZmxaj7zCOzaOHGmn8KLFzZIPjq48zXXGrj6F1842ddjn+bztKnoIXX09fP0aDL
8jHah/8vAtp0nEjswY2Ldbot5hC/Fy2j6PKiw0HsFxhIOdOzpfGaRkKvPqv98YlR6B0bulrCZyHP
BUC5AAr3PH5QcMmBucXHLOg9LdovdNQz50RheKGbknpYBR5NIEirJxosY3uAMVB5WxSxvMlGgrZd
OKIcPik2kcfaMbrpRcoppHhCaCyujyxUAKJ3egT4lqxwqX+RA4DFBQxWMz4TDHjMBlQwwhCP9UbN
exHWTWCR14HUibEDRT3fVur+SQx5rsQ+P41Rx7h+SabagaZtUhOdhlvnDE4TVA1e2qYrS1RnOrXi
b+5veBYQRV0eUDHdlG6iDiidiA0OCXJsedhMxjVZl2w3RLq+5CjAv7Yoz1F0NkQyfURqir1LrWU+
oczanhYU4u9lwU5Ekx3k9qD3BMZnfMPIuWN7u1wtdYlpxxgmalQIaLZ9bQxYBMxVgjpPqcoZ8u7Z
/EPob52hKhTnWqLx1t9xL1IMfI+BNb16ypz8NUlYTsGxRPa10IEKFck10TEJbjqm3a2u6kdB/BtX
dTbTA1KKvi1reEoJM7pzBmBgntRl/YawAcnHf6Gn8hEy/DNsg6hfkrGk7TrqTnHrT4ntc7hgkYJI
wpybdgqR1y8gWiMnQMUIT8m7SHCqneMnxyze3IRN9b5HPzQyGTwbAXgUQ5qHWEVFYTOqtyxlcfiF
gCuKUULrNeCxAWzBzBTLO/sUVYjqR4PWqRj8QmlwtyweDbBDqhIMce8/18XbD8C1HS4i9L5vTVwH
zppztpukv0mbcwKQps9CwnR6Qt1roTFCKCZyAoZ4peKkifSczK8E8oY+eGh+gY2YAOUvUY3WmnKK
xNfzTwc+en3BGH6FLt0fR6LnRgcQdjsKmuQfBd7jsYdR+y7mqDf3bnKDhtnnxdr46NcqGN90TBxo
3Jm7O6/mpF0WEP8+sxSxky/vREc2tneCln30BBuTgWiIVuBsdbVvgAvJg8yqRkTrS6Fmzjh397mZ
6BZaBgK2Iwj+GPGz2mhexLO+DQP4fwSXdJr9E+yoSl3+SE7MaAGfarD1hCbsdV1HoiiPKyCNANQT
PuduIIG9sVA6XaZUszuBaEa7lzYInANKk0EQ3G0dc1Bjmyzd7MGb+MeAH/Tl0z7ECj1IelWsHP9s
8zJOUDDpXtO+wO6FQIYQYdBi5h9ETlxC5qwG59qx41QaOMGaLaPTfiZnq3xM3dL/+lPz4a6A9l+e
0G6wCAKwdAGWbHIkGEESLM8rAjsiPD6ztz7mTJzMpr3YXA/lwpz0i3hOQyLSRxRIoS7irGlHLhOs
perA3d8lOoKGFeA8RAYrf0WD3XX8Bv006eTDqgYUUP79i+Wnd9D4U4aZEcjF3eK4Hqai6pajzMp6
90P34TtP5afcs5LC6Bc3u1EDZ+mD+l1PRWwpnp5IjiZQ3VHhEbuWMglW2WD+HGyLm3m1ksWCZcRl
ME4CatHz5MjAp3RvLve+5G2EpsGZTWvFR+TNWjJy+xqO4Ix4NsQ+d8KSePKlinMNJr5eRtqG/BO1
5nXn6SlHHeB6cSZcdWsUkwEMPbtzVNW5UdbtQq/0OB1ZDRAWPacMMfNW4E4xqCfiKx8vFra4rVeV
Gxb+mava7/a1W/xtqbPBwYfabhOdwKDtL2pjMO2oukUaiKo2EaRfev68wQSfICO4p0n7uNapp/rW
g5rx08pJNMzrpwn1nN9WZDxZWeh3h3WWgeFrZUMfA++xpxJwJBFiR9u+UbGMyltlgOp/X0J8hJWF
3q3mP4FytPXI2klMYu6IYOv2W3eq0Gs8Zb93MWQBqxLlMGLtvVZr/N4PLXghtoWkDCrTnxjy3DHP
mLBplk8D0Y3xkLQcsNimrfdiPMQsbk76tf3csegbfPc8nu6zw2Q2htrVPDIRczJffeDsbA/mydIe
1Pk5N92npW2zctyHwFkPcd9YVKuI+YMcOGF6SszqpE6AXPLlIrbpIPZAx47b+54+dW3CaLYpq+C6
mrYxaFJhyV+lyvVZjP79pLjXp9+bZi/RcuNVKJRJB7EOwcQH/Y6ArinUB3fptwYD/t10atLMOS8J
s3iQ8mke58HejszKizMSyp+NNrHN2UdfuLbIcV4PH06suaIRUvBCcI1Fr6fG/iO/w9WXQiJW0OvE
lp5AyMaTFj4QH2iRiIrmI82ZP9yTRcImWYSHaR6a9Sfyq/1tn+Dc5+yhcfpQsIRLf4mtoMtOv/Hg
uOZhstz45PswqDMcJkRlD4dkPcZt3iidOQYjj82TJmxTAXUt3/B/AN3bj+B4kVzWw6PNYWlEcq8H
aXcwNMVBMPYu6MEyqfMKUFRVz//sOtpb9qdrUIIsGPIAiiMMpYyV1SEhtBZdxjYZE8ZmKStDrMGB
4quM0eJNxRmg4JuLcJeZZRi6EngPTpEfCqtrZlS9jaX9ru+TDXKXQ72JEsGu9fzdjiE86ufjrvcd
rxNlxV/IE6z32+r06lQfZLK22oAP4n1W2xDrbqkQb3loGbJABHFEsledqH542yv4XWV4zF2HpMzN
1wvczO/OyrQKGa0F+SceKo6gGB0M3Qwo/RctoSqgzBGrxKDc/soSYPnu1WZxSPfpi4oHmz16dLmD
8NzYp4zqEb4IJu+LWCYe1AfJHeEh5F/10/srHLuekdhVFbaq0FzY7ehVmcF7YoTKQo6l/muFjpdd
AVfKJ3wAeVeMTlYTxO4M6/A46mWiQyyenMNdoX5kwXdRogUfrbRayfStgp6/OevDq1b8CDiJ1sU/
mKnWP3PPBz1eAZJxLzu1k33Qlu6FcZ6+I2yIgRFltORRj0NBbMr9jaCwiSNpb6vtRhYA1O54OYpF
SEYtCjAWY4obbKY1CdlNtXlPzTr9+ps1d9U1xdTEzhTPJC2CWelduw3TAVN1ScNpmpFrda/nyXii
VmlGd5mPB9suzfhSNYC5HLCWX+mB4S/CBfuG5kmYudGzGzaEUlDKoY+UcFjaglv5ruxVr6J37UHK
C+J5rKxRByT8kWld95YPZrT3c4vWgGZcyQCy3XdrFyrzb218azXCkHo2txg7R0rZM8v793xGlLtP
jVyluEPNV77qL1T3e/2uAZffxoMdOmHajmULn+rkXWAXLRY4DFtvb4GTb1WqCK51AQWkU9el2sen
q8+KaeIgm0B5V3Mv+xazWjhIaGxh1vuojG5+1Hf5beCyI0fnEBgrTISogfWEYLAvRrTwDpehqxF4
hdxCpi4Vk7cfrOLW6+b2qas9r3l2a7eXZIt9onVAMYntevUITb9+wtP1YaAONDBC+Fa9g4LCdm2e
xePVmpOypX5EUM95IGjzCF1OOEYRxdKqDGYNpSZj7t5YAO/J42Rxolup29PbiTyrdWfo7+eaTr5j
38KggbBtxCemCkl/0UMyM8oFJRdrcvp+EWejPONi8KF2Ix7zbrShV9Wv4uSOUv4bY5ixTMLCBkeu
90oveSXNzzX9y2od/UGxWdk4e6DTNke6XRuQWnmL8lj9qlyUbZ9KxHZjMpcWaEH85sJQv8KZOufh
EHLT71um6SFn0uBSR7C7J3w3rXb0ZV7E0136QfqrLA2L6qnsoXPN0PkA0PDLl7qggoTC00Cceqet
UxixOYqtum/CjMtC3IwDveIev09qijq4OU8IKQwbdi0PvQYLRLK8nLndTPGgae9Oq1u9yJLFz816
fezX+6AhNTw7P9OMwwHjTHrxYmQxND9sYBsxrX/RFU+0wO/nHR1jWdrFVQIYW4k1sIDWEPEoDI81
PgDVLoQ9E+AD3t9fggPEcy02ZOkXBPpmzTHOV3vggX96+uSuq5yBH5uyhnyFmr+803pFbq3BYXnH
6zN/6myXsy0OyRsiuSzeRj/OZZGwaEuPgz34DfvwT9ZVMdsYwn+bTc/20St0t8/987g4k//grRtr
gP0/M1bptIbM2shk5ysoJLeEV41jBklJr/2l8DArmJ3cinSxU0bfEi13IPDt5rfnHoEGPBn6R5rj
A0iP5luJmGYgZWXGLecFjNMJsOtbpEqhUVm6uWd61VXiZGeuCd5OdjulxN63AJ2VmxU3I6PCpqpQ
ZzfRC2Cn++TkCRJmGAi8oAXwrv6HBqrHNY4RQErLxzn2IUD+Row7XvDHvKWaPYZ1T6r7Bokncg3o
LUHuln8OWy6z+9bqka+oTJgrBYDqiKr1Y0PZsk5XCJwctf8ZmgGZd/GfZBw8VVfKN+vyRAAk4J8j
HJ5yO0h00jV/IV0Kxci5yUQDokJronIwMeImu+SogYY2nnh/N1AGFEhf2fP+ZZAb6r+hpGBnnD6S
ac1qBGuhHY2mzk15RCn0J9bD+2cR9w2q5DLK6JvR4DpJiVUlMBufoBqBpV2TGwvNSWScw5Y2PZTm
1Iyqx1vSe42n2Zuvh/c82pk/qhtRD3jLkvfRTIFpFsgZJikqSewWTqsN9WHZrcyzaFuuv3pC72do
BTdCLBl7ksiH/kOXc9pPl6dfOy9r0kdqEbrLlxIK73LqMl/totbRkKDyp5KSBRCSmjHArTkR3P2V
UMSHnJOsBIVbf7b2fzFSBqcTynSJTsO/jMvoSX8L8mXy1gvV8LjGbPINnb566cE7ctwudwC3WZRL
rOgR4382wwKBMpigTwvwkBQk0ypN4xIWpld+ndl8KBnN8tKa3/kq7RcLFJXiyhmAdlWQ6GBEv9tk
Z+uA+znPGFVp9hmnuR79LkkOg54gl61HjaqQ3DuM3AL1WsOrL8feSXqZHZViKLvgGStg+liPdvsU
1tc0XtWH62A9Bq1qWiJ3l52Q92KfdmdkUVsv/IYAREoWhtXkV4dytdb0eoaNdqWExr33xazv3UUF
e6GL5HuDliyRmcOrT1c7t+S3Krg0coEfgU1CRMw7ZXsFgEwCO1E7bgC+hllS7nUfGJGtXgoHqJAs
uw+KfMLe0DCfbCT2XGU0H1UteQ0KrEAp/cd5Dp/qbwETS6z6qsae6j8wbd6tOVzE5Z9XSrqfenIB
50EB5xCxLTV/1ji9UNJIELcfS9SUdCQH35wSwV+WrfS/YgAlVOhmj4+M8o5MGHit+/5PfSE30GLS
kftN1BH4F6yvlgy29B/fFecgb1eW4qdsiuoD4oX4y1YvrjfZqxf8bCAO2lcY44CsJz8YjQojv213
4qq5IAa4Dp5UKQwEIrZYKrNu8MNWUD+0O0JjgespSt66v3H5fNyNqiiwT5zeeer3j0rXLNzemWYk
RZTYroWgQM2BgSGYfA0xwSDecH3wkCZcwpUKW4tFDGI6egSgQFvmfLfBpdng9AhmWZ+Lh7FNNsfo
OutrbqkCX4FdPsy79XR0+oZVGSZviqaUJN0FFe4PZz+DiSy8fiaOKZ69B0h1+ACKx6e4at5rKMS0
PvaNcUZ0FOvZVP/cjWxxzVF2gweH8BglmfktVZSL3Alz+Aia0suhCJjP1aqDbpLzVhJA+ZPMZKVm
tGYNwNECRog8XMRMRMIuueMlMPDt6nczAlUSJPY+Rkz2p94MAD6MSOsVVLsrqHYRmIvzps9uP5ed
bkIur57uYOU++62nQlmqfGNo+KDIcZ3xvy4z64yRHW7bbySUhS8HdcvoRk8wb4iRo/C7NsVVp/fe
5dHOawhhsIxVm246QkxRfvQ1oiu6Y7rRIhsWGVYCCJ6TSc+wmefCvqMTQjBjxE8OsnWphedGgZx7
duvX6HYFTeaVtlTtZe7qGgwNO7NSguD2dCA+epBq7eBvvOT+/jxg9DjbcrZfBq6I2uBut7am30dV
b3Rkm09jesGqARwNn8VKnDz5mkq7/GgxwTmw1T46MaX1w54X/76MneZzukSUaXX4CrMAuXAtMueH
Ba1Qx6BFhcfzE7g0f9LewZdL7hyAe4LSqNT32p7O13Gz1TGjcKYP2mccjHJFnHM4NxGE7ZoY8PDL
vpAmOc/9QnP8onCjqUKY/kkdwTxV5bpv3SHxnvftfKtZm3vIUMyThxJhefpHZfJ9odlAidTji9iP
7PuKNM/A+/zKufUlpNx/E9RKAhIq4lpULdmIbcJx1WGacSg3Xt/q8SPDxxp9LpResF7g7yZ6dvio
eGiK2RXuLD+YhITpbOA+hcpjwNZFrh0fQc7U/9ijVr+CDTB76mcfYIivGwKFc4mzT+PEB3MZqD0o
5gS3TPdvSkXq5fCnT86XOc2S+CFwI9ulZDAkOX76QjOVI6NBp053+3zkZXGGkPQXgtmSBRLbOPPu
XD9/MAGlncxBHX2+phXqZJiTBM1vFfGds+AM4v/n+TvQEgPKruDNRScypzSMe101luiKKGOWeYW2
MtxoreLtN/BKqGYC0PCL2OzFPdG01UYUX+QxMgxDogXE9X39npHq5Tc2k4KeZ6ghzTH2irptBZ8D
7UhcRnxHbTDp8ApPamMvUXjQBdgLcbfR/g8bqkPMd+EbdzHs+WwYxz91KFDIOhTKkB1n1I8osYmd
NyJdBXUn4957DKhMfEnisgocuNg2DcSsFTr9FSnhQxMP0/5YJgPx+igAVIjQaUz4js27FFtPS9F7
XXOo02MwhRiutlSsJSczoTIO9WaOUlD4kXScdvVtcTIc8Fq3L3O1HQK82gVVLbYTJsQdllvZyOs0
lC5jM7CCf9hrBsgXPUYBhWC3LNJ7PU7NpCb0t0McRFVqYwulJXn1gR4z0Ry+ahTLP6J/xDW5WlJw
wLX4sQQ697Bqr5ab3J+GldU57m9QXaZIU1pD9X/7RksTLg94Cfs/06zWw9SNps3sQvMK6ePR+N4E
1J60hp7bHyzFP+Y1pIWORl8LkT+ixs1tXF37J6cKxhewklgnZ0MMHylG5nlexLhiF3chL827FNIg
D+rH9QyeoFyO0RFakmTS1V/P3rM8ULlMSIT8El07CJ24TFYxlvp/OF8i3yExDU+cfA42rGY68Itb
dcugluX2SkrMsNwRqtp9dMXBrVgtQ2Qcr9cKfNCIIl0KfAXWveWAiL+4NTt9ibUqRxnLy03F4qVu
gCyudq/EclAi7JgZn3B8n9YRiEvURVqNMPjump8EuPQnQgCUc78jx11KIFrzdnNch2HxdJ0u41gK
K+xAEaK+CVSBaNs32q2dHzzY0jtfFr5GvpmLgSIPRRI91r8pZXuob+t3kmxGE6zphDlgcWuuRn89
qGs5wss+A0hR+/SiWIckgX/KNQvNGmcQzLuu0DaaVwJlWueMZH0WqGXwvkxUMnX400gQvLQT2740
wfwP0UMldDqHkkuA4LLurGnjWNKeCaMVLDF9wbp1C4c=
`protect end_protected
