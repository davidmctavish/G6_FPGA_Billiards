`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NDQmFrd0neS+znXO61WKTkkyFwGb30eUXh20zauYzhPq903FnYFn6iqCfTDu1wsVs1hZCksh7F5g
EojEBshQ1A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJ/PaNr1NekoGDX+vDUbgtS3URjWvctKH2UkONT/GQK0btPzH6H3UG46yydTijq+RLGJ9iX/g1of
OVDALbvNr7Aoklle5xtvtHMNm0LXIMArCDXig1h4Am2JkY5YZCcLSVAma3FM7QH5WE/V7Whn2YzG
1YzVtWV12G3BZMMhf4E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gcR7E3poZ8oa6Dr2ZZ7BOIwu5tYNOgLl6aZ4ctyyNg083SU0Oo0Qjz11n+5IxuIJh2tbHP9/8X/h
37a0rCcmAs5zTtJvzZDNTOAbDW1PfDrBrG/P1q0Spe27Bz5KxrYxRUoRG6MmwgMKhhg3/8AJYRh3
I+bGagtCgRd80hbtLr7WvTX4NaUMxZFgPj3sdHouUKjzVL+MSXjJrkPA9xDbvl3EUFfR2cJ6DoIW
shhgGPsgIoUCdMfag3uxHP87TaGqiTfcDTlZDC7fokdVSjWkui2WcMfywXbtt6zaODdoIjIu7J03
7tM8nRu8mQ1SUSEPGMCEoH7BvG5TSqcB8Gl1Ig==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p5eRvn291TVqeA2HIdI/H0PStfMNSKqo4XDrzymYYz2V5CFdOVe7WP0Si60DAqcRCaFbqYyaVAaP
p3RoKXCZ+cq7IvmwGgSLAUb2oks7C7EqIGMW2jgArk8543VluPVdQRWBra9HelZkjZ6jJTEs0ax6
j0kB9VhjgkYQdA4eTbE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rC7o757DC/fwdWNjyT6Lcxh5xqXtixJf6NXEKvS794D4knEVDsZT2Ne0JCAiHq+BEocAz5tkVwac
Ikm9nsE+Cm8U/koLV5h3DOe/oGFtvcw5x2QXDe4KjK3STXT8FHCIi8amt01f9UPregiZndEPCNeL
3kJipW2+MVIhKyVwNGLIcHe9LllgDe+v8m7EchAkkO3woUV54I+p167+EoqqyFcESuCq1iNzeQFJ
9EqDAr5MyCFGAhANhewPssWlul9QFHwy1a87DSmHLiGK7w34/L8fbH5K+F65/JxZemIqtUnKIc3Z
RqgVpjwyNUeGO/orqBAmoP2eu21qAAd+ZDumnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11616)
`protect data_block
GmPD4QWl0t1kLUYKVhSIbcxKCezrc+ttdn+sKIyZtURT1LFTMZjSkpgUC3HSlEp6zwpI24p3jRcj
EA9KowIevwhoeXtXqnlKKerdHpFrU5YqnRUL9ZmhN0Au4xu0RFhIKF0PVEB7SUo4XJ6Eis2cos5u
iqKmd/NHozvQZdaGpMFaVXcxK3cCvsLOgWcuMiObK0vvejwiSH2ce2KU2kCGoGkrxxjmwR+GTcJ2
CJJzO+/5l7u4l1vgv7cGRihzcotVFkmo1eGVG/sm54S6aPy+UaoImw99k/H2mPzKf+/i3HAVCtyN
yhdVXOC7kCgwjVhz6ykGHsWDEIwBzZyqZjX1AtfNXfXpc837lR2+B1uFSfks0Yh7gPCPo4dJhStm
CX3fyc4KXDAfy29ztJfmSXMExZHHIVrIJudCBToMslbA/8oD4002MnyTmqLzvBL3e4T8Al+CU6Ta
+oqmkOiO+IblUaWqd+RIGA4IF7yvTgZ/4wB96FfgjualtJXVyY0i4hVzdqpp3myPnBFqNPzzTTB8
Dsfu88qDZ4yuhZN8oZMqipS1DbysrSOYkPIuc4D2qe+i7poWyC5C6BgWf+UOyXvLeoLomz4g5qyO
6Pk5YcuLGvreLdJHVUd1lTZ/4BQ9oUTCCeFoQp2EmxtMaatfguU7ZTd2o4EQh35kDWxQGXmAuIjh
RFYymXWBhoZBvy62uoAZsc9WnU6lG1OE6gsjR0MdEIi0KG8t/QdbJtJ6erhiCN8MrD4myks4Jck8
UjxE1BfqkO0QCekCfxtLQ0wLtlFarLgRUHOeA07UKYU+1HWWeNfKEoqhDAl86p8MTebGyLyxJgrc
ZbvJK5ogS+gUlc+5ATXc2enG6GBHRSvlLrlz+4h7+b7gYQQq2nChZWXD8SN7q+F9I9IuhUuJ+Hd4
xo8GYC9M9ymVHI9yvs4aspyQfqqT+wWCBnxPyP0F+q+O/gBKm48Nu3YHmVIhJTaaRG+gubXsNXca
IuTh3SpVRm60bD/Tj7oGqcgi5etbRyfSWQnEqs/ia79rRGaWoL1Hnn2AdOFmzjbkzmgNVQFr17DU
/smgD8xAyNxDpokxn32m/wBwu/WxuXHMLHmtMmr6xbpz43YzDbwpUPNeKVVljS+tsbLe/buRckjh
8TVDHXqXBrouK0539UVveqBzo44fHe3W/WAB+SpREcPa2eYDg5FyvvFwCPneNCUSVU4Yqz0A32ws
XY2eNULM924NAb8krDszQDBDv+7Wuq/VVQcNC5WBAQZ5hsXfyjyDTjZr35wIgCL+ENw4sgdtQmM3
+2/HmVBRrwuphI3vydxSre/TbmOprmIvqZfE+06UrIlyDncQkL5I+26DzTPLODmAK0S9SPfdLMxk
cCnxHEUQ6E5vFHPPbdmJQrJA9NBudrUw4oLSctmAuxJ+wVXit2R0bCt4Cy7tpQ71ZEb22lq3eYOr
opoOaH+GK7m+mMeZ/PMl9UaiZ900l7TR30OLQ3jVKvgY/okdyH62u3pEyFhg6GybQ6IIa9szbln/
qaNS32Pv5DXzlQUnMoCXpl2Cww6RadSmtnhx3GmD71YN547oNk2zm3az+r4Ocf2u7mKiDMgvg/Bd
L7KntbCec2xJ2G27iuuOFZCnq14ns+oP6r5SFuLYwlBiHGvEpWWBZRzM4Y7uuwCPxhx9TgqP1T3M
YKnzdA5bivFfYziAZqq//n3w7Ek9OPNMKd7LJ4IKREsAYKdS5/nlKAmNj9jt/TGiudsM3sXWWGMI
WO2YXKuwXCY85zBEXBJcr4Vg5HSYZn8M3DRYplYNMfqiDhp5fnPX4fMgzbQcNV746ggOCL10Cz74
1Zh05/YPHNwvn1yMiE+Pzqg/kwhXoYw7x0kHTz9BZwcuGrt2dOqUKos1Usiy1UxT7iCaumfTQCMC
gn9rIKkLJWJeZsQ9/c+SdNZN1uCNvjdl5CJh5igiXseX+Wu6SJiG57zrhCAAvSaU/gi2YYgU9faJ
sFUsbb+mkxOQu8SdbEZpmEzYFrswSQ3oPCPhfHeUcAoBCtAKrztau6nYsNnnp3MHiVK2jQy+ojpX
lEoVNe5OgnMqI/zPV0ZdGgv8C2NAO2ftD4zVqdZ/oBG5adyCqDKKR05bZ+2Pf3eVq2PqgzGmLDUP
0BCSOhdwkIC/RrasNLkvRaMz0qc8LEvGnTijFx56r6s92uxvqIC9Wh6bOuWVD3UfAo1rqWDSJHg9
6YvdGuYujnZQB6ncA0ik41RhkJsDnzctmDqLtfoJ8mZijEU3nt9t3gA4Ma3fTle/ow8w236iaxKM
fg90qqMk2i7kWYwzyT+2WmhYkIkqKhsr6XODog7wTmd961yi8lpZ7AfjK9zJ2aQtMpgtMRVtgazw
UqnDL4H4YxozPHNcHFJyYoC8HCJrx8acBsfBho4B90AJb/PAN7atXWta+b5kSj5n0hTYKnbeEob8
YGqgmcRiCP6qs5JZkAgEHA9It2bREfwSPcTGBeAoomtE7waJTlgwH19xp3VuaLqd3RAq/GFAMRYp
MSdkm9GmTEfKZNR0y3tbdDUtxT8pCb9wldEeVMRCAY0D5Rtd8FQ6IgsSOcKv1xwrvciqEcaANTkf
QmkeVjpUAAnCcaumXjbKMQwntkJOHCo2mXo59koTMXjzdoCbwNcvn54LmaeMhZ9aW4b8Wk61pCkX
nErOt0zJbtRVLnYX7W9QmmuND94bqhuljnW5+FSCQlu2/GtEVQa+/2S24RKs527FMzgoj1X5uYwY
9A3v0OGc+ldCF3TBv2VI6AusDWB7K7KJZikEpZzA2iefKuNI+L/Di7SQFzidQTNb88qlrZqR4vBi
1//IfayZvCcg4tNICgs8/BfInrqk8xfMvXYwPU6U4+nPDI8Mu6YwbkSK5T0oj652xcUtQEjAlmdS
HZchX1PewLxkHKp4ubicBT/soVFPUTrjmEklxKt4hI5g9ofGE39AVafvWwhoFQYQRQ/wHyikYT4z
63k8qWzOQk4P0ZqV8tMVuHKbuYq1qnwWIb2XL6ZcmEj9IF79C1O9meSOapG7+oItpI6odPRZY9+g
gd6yqR1zatuKv+YpX66AsmE3vWOTNFkyuUmtfBDC5GemhiMbI6IAzX3t2VUU9fac2dVwV/n9i3R+
0+tNoFgyHG+3jlvEKETDvulER804/mIBfTJgZZHO6t1g86Y0XGwBhqNNQyYMo+vhmMhm/x8lt49r
IzOoO5zXhaO4I4V8nGCHsXdHqKcyl1TRatN1oATt16sDKBtzHDoKsaKruFA9mLD3T7xegwb8vvVt
2D+bR8hpjAK57LFxk4ILyNZiwieI3t2eUzTkUurw4M/9RAQNu4v4Ks4KciPcfj7pzmtdC8DQxKBH
OjpAJji58apQhG7Qm26IDsKVYMquBKEYeZudhIVIDFVhy3Ah8D1BWA2t47opLSYpWzZacx8jbRte
oJ/PwQUKnSQqmX4ka3c3K2VQWzw2XU7i4GZK4XvJLwcXxy7KRz0CycUCPpmcKX+Oqcb4hJDwYYpS
R4MOC1ijcBNLQN0Occc3LlB2IfEhjeKKcTCikF5ssOztWcMphPHfNWkkwoYIgTUKTYBg2DAEKEjK
LhDlXHsEOCKfpkjtbIKYG0wN/wxB7htLQpGfRQVGnt3a+yKNfGYZ4zEa92PwKPgYXPDwJ8AzjB19
OR6DgOjO2bRocVFqrnHnVuM+uUlgOuu9Obk/rhhtFcJGYHgr8VZMqPbdLKjY/fk51hJENnRSsmHU
4yR3W22C5VzTz7+KdKlhecBk7rL+wFoca9rg5s+GDZPqF8sxmlQJ/GCd8XMbxvEDU+63bo8xTdW3
cjplbyX0KSv9KyTw98cJjuXupoKqZ1wkkhxd4QU0zja3ijQXIl0xoC9RkKj6pWx6qcRT4yRKURaq
avNghMu8xjdyGheeT6dLS+bTY7sZmiaWPKJyRZJ4COoAV8gjv7QHrT82KJgFDLG8yx1SGhyxjHz5
Vi2QysxY25RGqgnnhKD/QThBKVfIiU1lKd4ZOCte9BY4qDdQEbSca4hpTNnK+Q+QH+4A63tlzIIR
NocDIm/fzHvl24TxqfuOaiFNarpnHO7WUv1pETF4btSfM0wySba6jn0oE65OsJe7Y/tHN724sK0X
umcP9KYveKlFpQMVWYceFgcpuHzxIiwd/bW2n5C6kHOzq2HXlvjN0rrLNMiD4StMlmvY+XnJ9gJP
mJpwJEzu1DlV2gtB1ftp0xTkO5uK0PZr8OUFd1HUKAyaCaJp7TZcVw0EIOZdnOqTp/0CiXCZqB3R
jEsywkIhVO6B3qF3zRGTNHKpXKGB0OwM/P9pZE5BBHzNe09ijXaTsdtdsD/hlVHZ0simHY/nwhyb
Y9hWIphrqj/j/6rSP4wFKU0JhNYPNVv5NVHjVcuGeOes8B4jGag7USnSxV18dm3+1PwvwOvPpVR2
DJjMuTbOWClbXhpZDXXilBfsAzGG5M8ZJAgxnoUBG8o5cl156EgiY1CgDkK3ta3zihED+vF7taj2
AMNAISkZU+2k1OGnRdCBY0lLCOGF3+pXkkT3scmIU89/BBfXKdUdCcr9erLDs9njTn2Czskz+o/4
noW6eUXZiG2hHOsA3IrA5Xe5kM2UqEHmzIiy8ieezx5BTXTEBz5JYcVVt7P2KyMJSGDwcvZh1Cg3
AKXsikFB+YdyLxCH1negCBfslvBpvhoQegCKAO47+revusVC3B6INiUJEQvfPftxKGEOu1bnje2z
RTfEAiSok/y0yjBGA1MQUk/BePyAvQi5hiolDCrdg0dHo8TR2Y7HeDgcNP/6sJix84HElQunX30s
M5C5w3hAe37OrFwmT8g8zEJRkEhmcuSNQ/eu4e0eYByHYk/PvbVCBJeeb8knyt5Q2ye7M1ofBYni
fYxB1w9RPDYhEBNh3exolmehSp+dbTlJE7yE5BVZlm6yQLUSqBIB/DcvfVB2Be23P/WZ0X4wBuVP
BWg0DvbHHLNvR1klKhSrJkrZ77R/czi9gMPaveeFrAfTN7yoa2Q0/1pQFEwAYQW7weDOj4qmGdiy
WPsr9YlVTkrW+OdXYFDIpyMXiKbYDmMEtTG2y3gpozrfxa7vDhAf+o4IkcJFgVmeTm7QoG0q6DgZ
dxfRuk2eDknyRKogOQLmuVpQqnsvGtdCXwO1AaLKjS19gMBSA6qKhXpUZ1V4+XeYH/f+DjKQfaeR
VULMS+gHfsrQ4jk15oLbTA3mXvodxRKqwm6VCy7LKxFK6t3tyUhvR2JkzrgvxDVzFTnM00mKVnD3
UltaSKNJFM14Aa/bWu09vTAuyK0A8ZjxxefmLG/t1GYd0SE6I103q7IPG0AqLxKlQHT0J17X33YE
g37SbNk4NwMHJU6txYoBH7P2/0j5RatJrK2Zq1Lg0n3wSgYL8VSdrjSmMMwBzaINrujJnPXnOzaD
LBPOxyJyF9jD4GWJxhJpxYGbGwCpCgYcOUjs81GguutTtUmxupThlmCA+sFY8aNt6iNrXSBargeZ
Uxz/+GyHPeCSIEqJFwGHKb1KO2FE+N+PMWvaax57AtdJrNcr6TXjfEROWy4Q3KqLp34RxEUX4n3N
ySNWlvB2Lzgbqk8ATM8Bj1MxjgJLLDA/ccI1n1bWn2V80JCOwPdNGHSdTyyno373tSoIN6EMKpeQ
kGkbtm3K1+d3R8NyeBiJqxEMm11A0ECt0MHNcBf4sEDqdLXCG6kXAYwdEA/9a6Tc5umNwQ95ccNZ
Ck31iTSVDqMr+1rj/hMhuPyewLNJuRRe1Qr6DJ3xcWUW0UTzOaVvoIPYCAJhQd8mHxbjUAXNtRTt
BmCYiplc2QJhdaPXb43QztwMYG9xm9RiWwqwpG/4smmS/skY0ByHNOA7iD54IIKl9EQXbxj+BuyK
AmRCk/C9MRBDQMov2BxdXvIUnYlM3B5qIp8FijGN0YrudmsGA65s6tg+0HiCWl/LZ01HLDow1qUO
FW9b4GEve47SJ6qLWy1Xk3z32ExB1rDMxCD9hOPLjib+3yWOHIq6hSiwDcvQBrRkw5bDeq6iDg0J
bJ+RPSMvtLTliWrk0XG34giwPOw+mEtyRj9l3bodTpQ29gH83rmIS7CSSSDRy+XCdArmsSnjmH/q
7vyFRFhuDQqndkScmeO+0x6ikq8FoV0wVHSEZMv4zmL8Dh2ZQd+GpPlwUSnWyqb+8/+qEaHFDDxd
1HlbHA7KpMu5VG79PJInfolrbuEjdmjMtkQ4eWubZMO/O9Y9EeIQYl1WGkhI/J8sWjZx5BG7IEAz
vg+FyMtz+Gn2Yu5y9ncZCUfU3VRwFQ+sAzourb0OghtiUo4fpA+0yS6Hmm5dl/w6bSCz4UBBHale
GQBj/aPiIb7U1cu3akxptC2hRav0CEYhGuuAFwCMkS6S+N+wgFvGAul6w56gqQERzD2+LrPqXKnO
xzXzmCaGSYcAXX51mmbtEoL4gDmcxwNwDA2halWLBxq0yxvo/9Zn7La30LfTC2EjflipxJbfIfAx
u6BWKh6ZdeasCGjvVgffMmmBt9hCp2FrBb3a2NN+4dG/YC3k6MchF0CQj3QBDdsRDroGIoH1kTEQ
dpl1RsswMcrrGi28scKBYZKqwtV7FOLkwF/NUISWpqHSbY11CMBz/zeMBKY47a1OUn4pTj+C/dMu
0ZwO8ExKmJI0Z9r1T9Sq/rRwlCPrV2VZIfttrTeFFh4gNdcN7YrnivyRGNFM3Q0lKRYaOjnTgpfO
8w9CqwvzDfasdWEPZcG8WDGedAPAPgpsFaKk34ZjaSKzqesfP/YGMffi5rO8/FwgtJ0xnOc000ID
5T6ctBB6+Q1Zw76yrfqjb2SjsEBX5BCVZ/PhvLwTkdvLr3BUIsnKLDTiNOseREc2eMiAKLv0SM/I
AKmFRx0jbZrHk7EIDUglMCLiQJKp1VDBU6kE8rSDVca2iWDfWQuDycPSlKoWDxsG6xrSYSsk6Ocf
+UiKeStM3v49eatsFpllCPO7PPJuuDJOFvqZj0sNe3trkfHJW+OE+2OOB+dF7wyDDW7A6N8jU/Uz
s4k0Ro18veQXf+F80LoNH+D53LaEt9m0RdI8RFkWJfc6woSN68RJIxSvfLs1MNHSG/dJXrS0g1HR
RgXRSIkN6EkAkQ5QKD+evoljNU/YlDLCgHblAYb+i01rBdhGDSg2JmeQB1SdliL0Gzj+JxZC8GYl
XNBhRIaqvIUEo0OB7QGXB8LpO8qen9wEo5s8mHjsjA/wnIIsrxfNSx76+z8gdbCLsnQ3N1NgeVJO
WcYGgB6VFaRyMFpur5oirwwa7wVk6hh4KSTwJvpULjdHe8r8c/2Cpon6Z9NWJB/6BYYC+fyOOEn7
6Mo9xVpcAJ4lUF03TyVdQAt2Wy9f5MXjSIwv7Z0jJV+rypZJHektqWApY71hdldVwOManlOL1gsb
2KignHReLtT+fqPbY3LbMOMU5faUhV1ksK+86PdfXBRhn3TbKcVPMtg3AqLaI0hf9TaPc60h517a
QomxKDS4FouRrBWq5wre2d/y1FnbuvnTtZhgdnGUR6GUdSULkXlAr05wSfmL3xMdP6TAAeFFW8Hs
VHgVPKc7LN0qo8z8GEsz3KuygZkdNPttrFthyKg0bHZIArKWvNF918NN4kw1EDjQLorsYzy3bnko
uxLGdviJFMp/s2SV9bPNfXIOiOXuSCx2JxCGB4QyI5tZiyymq0AlSDgbbc93vhmH3i6wnTmu5+6C
he4rkLcH5RV5PynHoATjEprr6gjaoFpo83RRrj6oP0Qa3qcCG0ZObazocBpLU6gi5F1QSDIP9C6a
NX7Z2Com+amFbQrIY90gx6ne7CMzzEzyF9qBrW+aI7tKhSIn0Pneh/+S1fruF6M72j1WnJZ204nT
lidjHZI+c1niUuH4lmRzgJ8PiibpU70rGQdD/dZZMeZNI/5+78yt1jBFGMrQrmXAaXcgfL+UBJ62
w1B4E1y34Q8ErYkejzLAtdKQ566C0S1VKvurQPJVoOeQP07wyqNMiN/J7GYHeRQ1WHKVxpks8ZHl
OvlipScaWOO1NRt4iY7C9+XzuITEiGeemJxbhf8yjMqUXpOeRaI3tjokUNLf92RyULI87KIf1Ji6
GDAngrNsvaOzipob6AgX3SljiHOs3Sgv0tfJMkQoFLIGoMzQ3U6HfPAPROup8CaulLvVqi+Mks1s
JL24mSNTj0gSl4QZ3LZ1GfJ061mWSKGeDHO2m1qcPNShKW++XFosXgmcYYME5WuM12L4dAO/LUPu
uYjhBueNFVp5Zwf9a++QeoQk4UaAkb3IxC6k6Y2LeK6yBzJX0szZFqe7I2x8YMRlDUQ/+/NBHSVO
WwQfPoJ0+FkCQTBT0AZHZaxFyhxQAS0FRt6rWDjkgXCHq5rqNtxpa4qGAskFWWCcdeteh0tlNxTj
Jla7t/CcwSUpXlXUeVMDkmCoXjicoBZzehhz3SQJRJuiAlQU8Cbiq4SKEpDfuNS6Ih5Ato6AdBgN
I5/0a7/7wXD0HCV+Vv1cnOnrZWQoNllUa1q/PSRIeCbcVOvigMyQ27zLIQGW5hI8sBCK4YtXASaD
PL4yHIPahbm2ZfRTZaQr6zDxWGEzjnY8g63z/hmp/z3tyMFWNyp0sWTBcpNHlREEupdslRB4lbkk
rGpSp48fTsLUvU2XHcgQnAPht1oPTmxoTxy8JiYeXxEUmV3qbmdn8ekyiqnjD09fIopVvVPwte0S
4i/6RwvgiyxHv7YU8botaGXjJ5MWs54zZHD+R7TwFE8gjAgjLOYWzIUEAXpvy/3+P9O2QOZpmRx+
GuR9CD1kTn48NPR/DmoEAzuS2fo0GO6HuwIl74/a8lWX++eT4ZH8eBvZyVa26+pnAU+xIIeCt/4T
KFllDYjWqq/+arjGCvlmJHh5RO2W25Wrz452Af0zPX7P7L4Ey8zkEygWGXlkZovGa9QQkh85a9vs
E3/BGr9YH9cunisi3wSwIn3O2IxiGtWUVojnaoN/0sbIz8OZ+l1fmdRGa51nUjVc95mX/HWsZzeP
xMm7B5Q1hdCbiqHesDob/uEbiVARigX6UMEOizmL4+IfA+rp7/Si3GMNXfETxRrmxTn8dsMdS5Tj
WVK4kNLuzBst6Rpvn08TsYlMRawJ07+rBSftWwDo2zGvie9oQ1VTMvbIcHaBxR1LgPjGAwUnwUj8
oggksYZDSEiRd/IzDHf8i7OPpY8wbADOzeUDeKoyLBSYpM7hrnunDq+qa2RcKja+gUWUp/KplAeK
1025WHtddWbBddQCxdq4Q8bjtxRyILBWkmoeiTuEf0NYu6gAyC0M4hDbDbEwIcCPNTWRjr8n8xew
Mdnt0uPuVecJ914+DNJPeeq//DchZH2gJXHcLQYEYU67hCdbn/OAhfSX5HPgl+nU4OmCmpWJ4Eyp
1Je475SP7iDq6B1Sh8fylc9Kq7RlZikTH9Ti2T1NJG5tj3z167xyg23rqQ97NXfALKiREF69e1Ph
W3vA9nj2gsZqibtcWqiqxhFSrK3Olf5h7w/rHKoe5B9DzdNjQfBwu4vhhnd6wrN+3mle0d9JJWKr
QfruCBuXUss04AAMrPHDYpVfnGhJWcRPnjHS8TInD+ryXX4ZsB//i1xv4ztrvKTAVkXIazmwXPIW
rfaTYCmgACH4NAhFltkJgt2PIwiCrgtTprxKVE2YkeCNPvpTpB/y5yQi3C94JMoRVpcnFsuqOfBo
NgL5kFEhyy5/P6Jr1a1PQNo6PVD3TmkURM+/KcNqF9HQCcHgu0NjCzx2/orUmoorWLzkb9NaUfty
LCzpPROQSp1/8pOsttPCohsjGwMOeaRFKr2XqBH5M0fAXkiJ31phMN1jraaYPTQJO9Br6Tg1qkGv
HbjLiSX11unX/vTW3BTvTDm4fVtV6B4ZbLzSg4vOtxBvlUk6IA655tJTR8Qy+VSGIo0Z65VxAx9k
jgqIXA75r1fdnvc505/AweZX/pnXQBpVEzXRHEZulQtbKqPxYJiqahQIhGpuqspTfYVGpNE3Dm+1
qLrk2lE5b79TWI6jOj8feF1rCX6P0i7RDs9Q1H2xldvwXHgo4iYY0ztfi+idJnQ7vzVVs84wXGnI
34rzwuADEltO/zLRtQWDDOkZM72pSnbxQIa5kNReKJbTG6FCea5beCh/M72mZauOpDNiWcRpcjta
IZqsubsexX15ox3eEGBA80TqZQlMGX68QhufKHAMN2BzYFFBm7qbhwnI2msT1eJOnzaj7j31X8qg
l1fwz0wXps+ZCbL0udVCKPDxMumCGWu4PYcsfIdBVPJ34egnWlNYyWXn1kv+RRoHv+NI5ouL5dfI
FOQLwall9vQJ7PSXEnujWw1SkqYoeJYRuKGmaNFZlQv8+YCWXO0aO/dCJAuSS8ZnVEZn6O4EHOTu
TYyMyvR5zRv1wkwYIjd9B2rbwcRrk7/nSXkcVVneNacue+3c667UZyuqx349DOvtaR42puMfy8hp
JwYj2rIK9O5r9124ZDQixz5aYJtjjZneyiom3i7/yg0wYJ7meqIqb6jWnYOywE77sFexzkClmAtt
e83yY9YvNQCuvzj/lMuQd3W2VM/U+tJ0Y5hZHDmSFQNXF8ULkN5MD44J20h9MEHGOm+h/gN9KCax
AENMKSRU47Tvo64OrBTCOD6YsDOdSorkKfUKgxQCITHCaKklW38e57tKTQYyirA0otrvY/uB3GPw
4Xcjgzn699DVEai+2taKQxFyxdSE7uLhT7kTdOsiOjgs9CxwmLsZh4fScMbWT5V/lVnNZ7q24uRI
D18d02ZT+ZTZ690ryDmuPEfDOVAGr80cy1x4CEagf8SrgMld3GRI1bju5wyuQ3l0gJ4bOpsbB6Ag
5NrriDztnRoGbUH/PD020eU98z+9KkxSbIwhiCJsJuP6dkjSWZ2dRBYf5+eeFN0Djt+vVnNFegJH
3UkCSbg0XvKRCMT8ByMTew5ojlwQ7Km1pk4//8whBlpJakZdQ/WS/YDBRKM1Fy+Iq9iieweue0QW
GeVsdSV3+mDoYMaEpEEzF2IuEV7nvNthEiV7sjPfetxWKTjGmb1Uqp1xlmzdiNjHMd6OxyqFdGTi
cmHRmsXKXTNTlJJRixdf+tCIUIj0SBJtIakEAIv3AxXp3FS/DwCJTzPjiNQmIiPi5DeBE1AYq9td
ex2aP30fn9EyeBE3hXMkBvb6yoL3eP3PL9tZz05hRRlFRJyp9Lev3EoXO2WAM+aR/CzwwvAudub1
wyqbqcc7JjRDshr+bLczy7ezwhSH20ABDVQ8VXQy0ArA7UrTOCD7WFTWFCLG9y+1H9gbTKbyhY2a
EZAuKt/f9QOgW8tgxMQcxZtqbZgnPIR7di0cb7h96IJZ7Rtv/YA7ICDy06l2VVBzcb8bh9yeqwW3
aLhPSduOSDvQhIxd31n0ouZihrZ+qKSl372eWznG28Scv0iypXNAHvdOKCA+r72UN6Y54nSqOSka
EXiMr/nDZoaqcaN/uQ/OcnPxIjtqbDOGlSpXq+EqXhUCOdrjvq04+PNzbxsyZPwxjmL6OqzAVveN
feez38V61QkvyvqmEbAQCIFU5Lf7uprrCenYk19v8qYme8ev1GB7VnNuPbpVojh3GuZcGMcZAVL2
MRdBwOeOl4oPdImAoz3fMWPPLRJIshAIhdROVhxG2oFrSMyH2PNZ2hKF7slhUj8dk1s6q9uIY6GF
tJsi5UXlEgGGrsglflwJuE7C5g7nqXmce75KytvUM5XxVTCL+70+Z1+8EfI5WxATnW7QE4DzADQB
2QAj7DHijYAaCVzmoT6PJmjd0IETO71yCb9/EoJ9uFdNUQbz2K+UOFdcUsAEkHdRCINTP4+Jts/J
lbQ7xhGfMSCh29+FDRVOdjXpE6q8zfD15/EHuNmewisChRmYzwlHtioLPiwK37pPNSIFj6G+O5ZD
tuk4jBjXSa3dXuhFiuFqU2SIT51qkBJJYIkEwrz4DBkrGc8FOpaKbcKxq4LmQUEkhb/i7c5DaSST
MuWPnA/9Apl1qh6N00eVT6sujQUNicx0emVSrYDK5h3Id77nzaTQApoEL/YDhv3AFaS06pO51/V4
c7tW9ILwvXMR0g//eqSaB7Z67HJcUZPsn0oRnK5wrLErqiTt2BRgsYPUXCLn8QdneSCKrVoykLjk
iE8J61L35Xav2gQAbdmJiVBDOV3qpe/oxuEZkc9ecNiYbzQbP0qBZ/0gfJkITqn0pmj3WW9wC+Gp
j8hmfj4ahwH9Uj6WgVydS3Kmt1de9s89z1prnNAmhGKhfEV5megXKGDVjzvqSVYwYoIoDZAU/Yf9
8GU9Ggk0inV2lnTfCCOVEHuHR0yCsYwtSs9TUrIbnguvCfVST4i6TnQAIoSD/bvKreJ/5HmSQKf2
hwpvfC0oSyajcV6ve+2pDJt/Hr7BvD380k1/6PYvKQhzwI3xLo5m2oGhwTwuRbmtEMFDuQpAxQoN
Q5oUO25xJZSwNm6VOngK05klgEBJIcquOXsZfAGFsmtU9Oz1TfZf8oimOCqxng/PuR0Ge/lcBRN0
7htt0+poOKf7irckGBNDnPGqw8XtRtC8Doa46W3msmchta6H8k2HPOMcpJzw3vZRwSlHXMLExKZo
4WLdzikJFkUdAYGFxJGSOhNQxm4+qglBEMkdUtx1h8b00E5FnSBn+woJuFs7g3mXLDPUnCBjAf/A
B6CQxmZjvy2ZXemtvp9Ki77qxBL8lgzOekOoP7XWemM+JcOu5/Zwde8zFNscap8SiphmvwocFA3w
WI6M4cF5SidOyz7/ZfOUM8o1DZMo0QBXmLdq4lVHNS+1k7lkSG3bD87zjfgL0Q+RKkBt6/abQw5a
2S6otT20ic9fvT7sk9a3R6hY1uj6mnZTdIc3d6X0xpTL8pf2HGYn6MZ8/rh/UXEBQut15lD6gF+K
uRW9N6uvEFmprtkuoz+GBLmKzyhq/AKMXU5QGe13/yq5oGXIPlNJ77f0bccD9PcpaO9Yj5tX+At1
lMjQms56yHjKthSB21rAZCalJ7rtPJBa8q7Oex5XHeqddffzi/4C/CCiItkm60jeR3U2SL4wlBrU
EFaIJ8BoODsqDdzE8Em8FKDJ/QEeYD+buFLQL1RcdmbZoEtVEzsuKMtYTfhb77MivNyIk+3c4Jmk
yNgne3imf23TCyLyxmziJ16Hrp6tUnHs/H9uBcZ97IW2nvLhx6MF/3AjyxdZwwqxMGFxFLktCSPC
g0pTYtwgwSqQ1FoTe1Eaee69Ru3rJuk+EVJwMR3HnyuBq3Jq5n40Z9YqU3zO2I9LUICwU5nyAIe8
tx/uS70qhd0YWESgwdvY2oF6KjL4YpKj+o64mCrafszPkudIf4XYJeLCE3CSrtBKowIBp7UwRvfV
VKVM76taJsTih4pEAIbu1riiO/BdMds0eG7TT0Ek9SWVpan8RGsgOSGNUNuaUnBE/iNjFZcvV41g
G5xQMuBfk0UwVZIq+BajTm30EZ5c76+BqV5kliK+7gXX/1E4laPbTKeLH4W19pWfNw0QrwH6sqTf
Sl6dvkeJF785TTiEf9HJFFcvSCq2tSWOac8UfeahTon9KVIjpZTd+pKy+hp45xe5HB0wWaj5LVgh
1Aw9RdpKtasQUz6vps2N02ZkXBpyWFJMIRCoeYd0mFO6OkV9ff/Ii6xqWY4ZLDjQnRW0y7nhaA1p
4V5mxHCFGNUCJ0kVvwBTwThzmNoAammve9AfhAujF7l599kgXnr8NCQfJtcORbgEFS6kB0VoLM3v
SJUdHcnFmbHZd+n/ff4Ju08EfNN9fXt23csB7nA68Vfj18OqDhz3WXJLxOwHfLTU0M3RVSMzBFno
Y+oFfTOnc5EzhXCGi8bqU6NjvuhfkbuISrxTzyViDgJMotE1iw5pxuHDZ216INrVhwU7mqbsz7/6
GI2ws1TVtcaj0w9w2pBwfMbuxiHiAz2fWXwNHs5MoFG+eOGyH+lBj1lY+q8a7/2Z4OXUjjdWMShH
/jfIjaN4Fdx76LCDpNJLJxQF7K0J0WxyM/Tgy4zMtzzOlZ9NJX8GfhHr+5wD1sJK8PGtdWlT9+sc
EOOJ/3PZt5OvSgi1zDxVU/XNragdDHCoiQlDONlKGAtyoQhrGUMddcKyTLPfWdwbcSFfdlt0oPDO
RHICvl52dG/Eld2O2vM/6ZzPepdLKKFipdtnHeX9DX/4Il9H0FEJYecpzbqjxhJ1G/0Eh2wfCJSU
Mm5Fv7jY7Yzo0GH9WFPcCXYBFihrFYwrHzFvKRWJxpVX777zMuPTRFchR76lU4DFt+t42CsuBUgg
jaCqqOSfbBEWeN/jOqWkKSpv+BEcrZ2gloMxY+pNpbudbAm6dDyRvHCmK8SRbJ3NPU7GpsSrVVyd
ye6ZEd9sL78RkFe9/xSAiAGKGUdOUxUkXXivFICizjDFsJq8rRrRdYU8/LBkl9blsBpsEGlJ45WN
78I4iKRJW2DX29Nh+zNdlbvdHJCsm5QGsegOgXL2vMNjQhQeWi47oj3lphOC3U7b5MBz/CDkEL1A
4WBke5CPU31A02Cz9DzNadmKJCCLIczlBdjRDiTigqe8JPxb0iHmli+Lj9I/Es5u93PFSprd6Eif
TU78uR2eJ5c6cY2Ax3bTtG+RFlcay/8U3RK55Pj4VFWwy/ATiMB6UKiCKfv3b0vcxgsG7I/RdFBX
Kye7gaEYsNorDPDP79FIvol7zMpVP6mp5TvkWebNL9BPb5NPGtpndOyUw6CndxatgkR6B913wSvV
rrIbPcR2piuwQ9EGFkAQ6+fJmoHf/NGVmvYEdtny557q6Haruvds9GjFuYzQKNl/OCayelAxiAGP
TzcBGe2vE/1/y9MEr0KUfJLUCZ6pu98Ss7pQcotDSCz7a00A7nKasjU7JGPxRqf22BhCoNPiIkEt
/Eq2r1snLfziFtL4Fi4aw4YAPoXKKZR+KrMuoi//VMNHojA1Zy2t8LBrGr8TBM8UWDzUNgzAZ7NF
0P08JzWo43pM5oXcr2OWXOyujYn7nBiyNuRH/xQhj8uO+PZs4WTW4aAZWcfhy+dK3/iG8Gd5eFCZ
KXbhZztNXzBZSXpoIG1n8yYIGZQh1zXUjivfPz+Tsu4FesZA6cQZTI6LRcYnH/0pklIb9D7OHruz
HR4K61NRjeHbSRMnPzmX3cS/Dm0PS5sTOUBUpxunx8dAZBTkGkURR0s9OcPgGaX46aGFjMJYFsDA
ep+ciXu/h2rDowoNYFGTo+kmyM8T6mt/KCHIQWF3kfZgTT8p33X4FDZoW0gZqCYFjYvjyCXCEO6P
LDadyEdSQHZIejco2HfPJotuehhsepIjTSVOqHSvUItJZuOpXMFy2dMQuu/jE8aPGpxzzP+sDPEf
J2lhAAcxd4Mx8COls59qJobYL1xWD5MQ8d83IKhJUVN2Du3+Iu+aZ6j86li8SGHIhLcvM6DaV3sv
Qtj7oADO0BcmtTRrPcHnJMonk53IswLZOnOF1M2siiz1FDNelYA0yfhcjqdeN3uXGVDq9TBmGRpi
yKyYziN9LIDOu/jdWKzWAsG9E7dBrmn4EsL5zA36Cy72DzSimqeUs5I0qCFp
`protect end_protected
