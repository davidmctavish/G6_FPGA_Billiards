`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mhzBm2jqBKrF+bsl4cRzZQYBjZX9Q+pwcCzrps+U4bzTbB+asJPd8vPVhn3/loahOyMMk0fZ/ezN
ITDHzwqlLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BV1BYjJ3npWZCLFHXtDV+Qd6kYSohSmBGd1MFKi9lUBXhDVwc11czLcO2DFG/Y0PUi31756iUSf8
YqI9eS1cBBm1N41q4qzfycSTw9Qs7K64IjV4Z3tWvProDN2PUJ1BSDWtnL9/nO36DnWDDcZY4uAo
QV5B1D9XPZRfJNOBGp0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T5hroK1ySmIp1ijj4NC25zTPvG326JZBg1A51lUOeVdHyEqYkDqmypXIZL93BD8orhA0LJ8rgyr/
We8KatrfgOz2zuc1q5GLpo8q+7CAAoFBg4nMjZpQ5uBkr/ga1lIIgZiA3cav3fK52cWVUnPpD9Y3
7AI/Y7wV1qB7oq3FZUEZss+EeM4bgD2SJfEjZJFYrznH2SqjZsvH4/6xH300bg6ReMQpucoIX6yM
qniuvbEu0p3ldpjMp2mqcRSDlgZd0AiDzrtTBosGzvUh6nRIugnsqXhBwu1jTlC49rC60BehcH9k
Fz97XBtdjrTuWkEygciPwHnLbIO2/zMKKlDHpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
32NRL2ATHjfeoLmY2DdgNePlbV/Eh6zPW09DL0fV+gMrTIjKFHnJ+dgOALi8MZMLauKzOVJTZknv
R3/vHUI9qSk5wFlcPDBFYxnrGogVEO66Zy+701a1d6qEGg9Acq0VdaSfEK/nZ7UK29+K5sgSTeQ+
I4eNpSEpoyLtui2NV1Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tnRzKq5Oyxo1vldbDtWHPqUX0qAwix9kODEDtyG91DBOCiL+f9AWzd4J3OfPKZaeoInSUZFQu71e
P8Y6welhQbrBxHT1zywJ1aWJjuUwJQ5IbQ5d+E8AD7Y27ftiUV0szxVnUD2ayYaMYUJPMHPW3VMX
oH8UFW0auVByZ3T6OXxa2G4m5+RtdVm1UgGrHlpGHU9HFXtayLwEYVOUdaVOwH6Yt3Za5Mx9AyIp
vcQdD2W5zSlPbCTRelXJpG/Y5kXEc/P8T0TDTB1Rp/wRYFE7VxnJPRF7vyU59+4AauluU+y6yUWb
mhQecbdewQsTTmvmiNOfxqD0PwbV8lTIDoW2rQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41952)
`protect data_block
pqQS2C9l7IewXxdLDpjf8VgZLdBSPmMsucB4f1nxqCNVxHLIfHCZgbt5z7NfmylRAwcXlJER6Xk0
qRcoR6IyyAH0cpqqUkDQ7UTaaqAEx0hbEM61uJx9FQ5SJPV6Syx4es8hffCQj9+D2hhekyPqKaFX
ghF2Lo/E/lbeVqyhU8YI8OvSKV0CwRkPM3OAmptmMTvVS3wRpfAT/yffsFRcUK1hFT/jf5YpTiVv
c9OJyr6+w0o0C/YW2PJUuYtY8uEMhshO9fOwhIqUDlYh/3/LLxESY07089FbAWJ7cqQIIm29X8T+
NL/rsHnF/jxoKsltLpKI9CT16NiYG4g4p4Z8gd8rFV2kwIc9DVSXjCLD2rsI+3mYu1IiNeTSaOFq
Uvdo95yy/Ksqfd5Q3VQO/0vSvMBZ0hkydGMCtnx1Fxrw1vxi2ptNg113frVF0pkrKaA6RO3WLjHc
7pyEuItNlDCelGV+Tj36eYRHbLhZHU1qsC8xVzjcxjKHvESRjpb7vnz04iEMLt5SYxOTQ8GzQbed
yfqVFZAG2CtcmVuRFJO9r8wqmw3lJpAcVKUl4FxvD3qIFbSM46mRlTYk0y1acwiq2rXT+WOk8p+K
DvX+KMgOcSf0Eq7v2DwMY8c8RsfVIDizGIhsTkzciEJ5qyI9ZdHOyUiqubRLgpXVTtkS7QK+clXI
AToiw11rUdoP/2sW36NTOjN54cKGRPmvfPDY0jy0hT5K7Y2bQe9SmJb/O+0bB52C02+bPtKpShHW
OjsvDZEVz8boz/xenvFvw4LVn8wGsmiPMjga8o+ZQYvZRx9F0d9FOEeOzlKjxiRiNp76wAt7ih+r
n5ne2a9ki+5UKIOXnqWjh+inZp6QNLFq2zGX+E6pTFGvNUpQAmkk9EdHH+OWxP6yjeW+bupzXkvd
Q1tFs3RMlOCtFeTP0z7U85uxIefkUaXlcC2Cf86TUp+4eBu5FxM9ORM3C8B87hHah+B/rezrBlgT
IJ457ey7UoSi8EymTkeNTFryvyydIH5mWEMlvNlSA9JN8ncvIIiIPatoclYlSTV3VA91hkV06UHM
7LfDgokmHIQBpBPvjhDLiN/PTCpf3sXjR2AeoBCvwPLurHYjTinjigt4wur1usRxoTZn7GFwTpxq
deOdeYX7ZtwhK4nE5hdMiwqQDMKuYBOXZszm/KsL39SgJU+2v6IDVDCfz91GLEroRWiGLNNgscmR
7Y2oh8E/C62FRzpJQFE3jABHee0wHe/dgWQZ7z5NoTcpQGc2rL2akn0KaPgsTFbndOpWNae+9hrN
K7kyfa7o9/ySYA4+1FX7fSzJyEZndibF1HExnrTZAa4S0Od0IV2D1lwxjFRwta+Z0AMaFyC5Vi7w
TXbVFytcD/nLEwvhDgk/M3uaOxm7r9zMvSFcte8TIccm/80jtPTk6+Cd4xT0fh2aY/e1s6aNGWOe
py/HoxLRZpdJLuF40tzt9ebdxJZJL4iVN03Jxuv0jeA690MRyBZrBQAXNn1mxH1fLWFqjB4Hi2Zz
j3Q6tBvwnPj2uKxsFtX2qxuEjMbEU07CZBp4wGWP4RBZhWoiDhCHzMn+yBKQI/kR0OyG0/xTj5Iz
SKEWbyqphrpvNvYNRf1MPLwTS15wJ+PdJzpv+mHXbMyPu/Y8xMPnrW3rU7X9Sn6r6AzfvF1Ob73O
rhPsrAXrQHkFhejPsRyK6w8QN7qBmm/Z6EmZuhBXvNBmjn38smwjYcJecIuRESTTyU0Hda9ejnIr
fFa2S1Hn2GjoQV9p/Snl3Qj2GUJfiCFwu9wqkHQpWV8nbMGL+asvxh6GVTcnl5/WPz5xLXtDXiB8
3wxomGOX1MfGsfIik9ut8Gpc39XOqCewCvuVM68yo7b/eVh014W6ter/vBsqED7vwUOwhoWaAiOS
A6/5eZAjcIlbdIdWUvXBLsyiA6YXUGqd8SZTtlu1zpQWoRLrmkB8pf6ikeAkkzlrDtmeuY0LPam8
7wJzNPvguAK4X2I6q83UwVGL9U8uOgU5onlPlCdX4JlsiZdkZAGbQUq6yjsE3Z3qpAn5h4Tiw+4K
VLCtSRqRJHrgjcGHYUspCks2S4MRPpKgJvw8evnRA25nmsewG39DuAUcz/V/8AX/fbVql9jZzZFj
Wuz6kZVuhV6fMaKFQ3KkrKU0lzuRL00vsgYQinw5lc0WKwGQPHyZ+LEYZtiq/z4YPjD4AQLBySRM
fk2ejNqlak5SyCOfNeAOV9dUUwS/c+JdHJuooPf8uoHRTmEoZCsEulFM41rUxCcyIuc4dwdJxxat
hNBWz1dtfr8EgjiswrLFGhK62hqojzf0bbtq9d9ytg5x0zZkaTi6teymdUF2+mXt6aXb0g9HaikO
P8rp/88d3VSFyOMxfUEE/OFrBz2N9vCvGitO/jQi5WGGatldcnQhJUE3pi+I1M2SrgKkTTk8+HCd
aI+W5v1xVTtI2Fz60lKzWaOArCBBiPI2x+Ivyoh5VyhTckS2AMyPqatsMREuq6kZElmhgKxbw504
jDBrc/mefCEJ+P7JQY0OG1ZybwbjjOmHEzSxcP6M+M9trEJkogg8aVy2D+/KVmVgOB+Y1tChdzH8
8CjmnXKG0l0bgUBvonPqjLn1zxN9qondUk1OFhJGI77a5fyyKiNRr+9wr0oKxc2p6EG/GQb+uE7c
qufnQXsVYw4m4W50qTDBaaN0qquDnxXWfpds38sRDh86a1bfBq0czPhBDlB4GPG7d9KNrIasn/UV
X2EmCJAZ//oNZD5LhOYf3Hzh+DpeXK29gztgyzpzA7eZ28rT2ULROwDLN4T3YSbeyqN9x38Qhcmc
YrW+FMHttciAXVjQI/H6FwIHVdMA5dc75HcUFBRVuufSY0OFboSfGShMFCqYL4WW2MeThG80xADx
noMFzEBrxJh00aeLDqFfREXfdXcwZHHw5+zJ+5Umd2wE2SznsHcleiVVJIE0Lw1lbKJcDfwrw6q4
4o+4aWeo3Txgg3/D2BR/XAV2iVN2iLtJi2w4MziEZ08g9XCGl5sExzVjcd5awBlaNIBCMM+7Frdz
5HKLkKOudQEI+r3GvJETtsJQ7IUJ10ya/pSvVcekFP7ZgTTuRw0nyKjdsrurTvwPIJ6fWS98p7fm
7wZilNjgPVWQ3EOKJ90IH36LEa2Wa1F6nvhKh7MZ7851m7ZIVqZYICnWpDvv0aPteHCJ9mBbEHE8
Mox3XpAzpq+nyMPviCRctIdERUnRwuPhjindsSLIKDuWSnxXYXLh2SFF2A5oqwxXYRZrIAhLnVOu
p0Hwc3VnZ5KOaUY2Y6fLkXej/+MjB7XmtggGdOdyPDb/CVX2TbNEN0MzpfFeTwqb+7g2MSliHirn
/mX30iv+JBX/9YwWV1ijBJy+cUDkJzwS/JtlE/VhDlp961cROwkMHU+UX0h5E2kjs4q2Wpkot4tc
dVXu29fzoAULuHQTsyVWdp2XKGXB+U0EcvP+h6AURPIy0fXU/eIan03dfqjhwoyvLCXfqduznJyp
j89iiM9upBhNxmRgY8/84mHHU/dA5l/ioCWzoIGalZB3h5ncIr7IvSmu5vqajNlrl49pkW4oleZK
BBUaJPNcxPmbwCPIrvwejtDWSwCguKK8DpMB0f8EJpHtfWi4j8v+kQ7vtiUk59ZgcwYSGzQaEAn5
BnqqmzNfsBx1FeOQ9SnHEQn4w8B2dv/dCuPM+lBRp5OvD00EwZpdyBsvH9KHORyZiP6iwC84h/Mw
NVbZ2QYosvYtX9GRWylesXt8Ke/+xLnKjeUdl/O+9AmI8j7kBR36xAACsiMNHNv81+89EdpOjSap
5a1KWtfL+WIn7HXfcSnvsn2hBXbnjWXvi28nzLL9C12BrhSsMj0V6KFwKelHYujPZf7VeAUwvi2C
I/2RZPqxHiqaAxmtq/V+vAuDWwhoBeBI9Mp8GyJfI/VxM0Ijn/mZetjEbqP8LOCuxnEH2KXeb7B0
CDibzNPl3VGTcrTSTUNdNH1dZqa14o7rxBxzmPsEFhyJEivY+eWMEdh5h3HqsxIUjZQH4ngfeS8z
5xwxYzTNKfkjjIVAx9D4UnOeRQbc5xGVUKmJq5nYMBqMgyY2oZPUWTfEw0cm+B7Ikif5LziR7CQG
k2NApopVvj6ougfNvCbbiEq3MEtnkLyuOQAXnqGbq+iJ8uHcMuBZmUepgG3YiBG2vyxe2UBtJGB1
nMY/zJSQQFnDK9WUq4Yv4qXfwlY4cKXoPO2l7ze2n44d+VMo0nLnXhjCS8RE4DQpCkl2LcREsyNt
Txr+TvZDzyigPo9mMrBdb+61j51s9oWO5EhGBgGwmnSnI1coqcvn+quUsXi+m1cfIbWiGGuLyEcn
KwZW780DM2jMXdEQu0pQygCo9z+BqTo6lOONBE2pFr5Y8QklzZwtb8gOTb5r1Ji715U7uAnhB8kK
t9PtsKDiXdDUw6UHDmeo+NHFr5/Q74n+aj3a6H12OHFu3s2h5m2t816ViI6un261rX8O45HbZfno
oqKKgA0rSDTWVo1g5hun/SSHQuLN0uHbl7rxy+purfSoMgFLFCwaMRyGsEEYb+S4g+yc3PXZDvQQ
SHTC70M8WBpg5g8HxyUzUfdoN+JiV+AB0g8vZdQLNxBimAeOWisF0qVc0HTF8kYNrxuIYLtwdNcg
Kg1zpxoK9yFeQJNjk53oqdT/Lmnl2W+2FX3oc9u58gWxnin0ye8O+NKa/HEV7TQ0ZYBFKFVMh9v9
iETR0x6/nD/LuzmdsazJr7q/w1iH8I9b0tvY8pNcoRZngYQNlqEP17qb0l8/KQINzfkusWeuFUKH
ghI49qDjjV1nyg3I5djz96rB4+N/gncCrys4tqg8ibYp5oT2H0+DtCSWtC2m2EDXM3jEmxtxlXC3
HrcFcMVPjy51T0MxCpw6z32LmnvbsXH5bQxVa7rgjfwObwvFTh+AjplA1PmysKYLLPqJjLmeMlra
69gagD8mNHum1xkxskXtDy/1glSN9jolU75H1wuLg74IYemt/fDan1FKjvqm6x1TsTHshPSWIfLM
YCf39rrYYE3JvoPlQTdijY5Ot3XsssopT7Vqv/U72AZTjZD4K3aNVYfwoVzguf56NgNFXZG6bWqU
epaqe1CvkepyZk9RmmEiPd2tvjRGDPUpPFwjLvPngcqOCnn5dxGyrk02+bVpnkDVv3fxPKmbTVfw
JPTHH8VMGDyYmRxrQforTTRczSFGzccIteokqRbmeg4rqr5qlfMIAjmLcQGTadr2mwFEqKMthYs+
lyyMZy43ww/OBWWBXPzWXLwfUKsbuK1cUfLIz/P0HgEKiXUHFMsBZ0XCfJE0Wkvv7wxE6nFMZXw9
XfycQV7L33HVUCsnDENhZruAijM3b8B8GoPDDf9DvyTtZt3Zbq/DlOx1frx5F1bcZltNGE3veFb+
qsX/xSbZyCGMZmNhAyIl+rU98pCoOmYEm1Ww4b4OTy7CeyMx7Z/5K+7DZlkbSjt/Ze3gLe7fflSO
Sv6P1Osk+pl5sCEyJN4mBpmxQ0KIaS1S6NL5bU/DAr4ilx359q2cv/R/GnAgDkQsa6DXOe1ypxeo
1UAdeer1C+p531ji8/t0Jz2idtfA66YJ1UJrhZ4alNTL71aEPauWYE9vXesg2suDZWvbp/eNdsnl
LcKRKMfyrdhKB0kb6PtGf/MNKTwQA5leiMqA0lsw/vDYAOpmnVO8W5GxYEPZW5O+1+DDzb9q/kl9
YSkRMAGIOsZCljAwWfbO729yvPY2Mgwj6fFiUdZqHrshB2wv6NT2PP9UWd8cLfyX+c9JL8iJpqd3
Urnl7EZ8gMjei3VBHLu+nAUPjnLchuFCjGDWREgxXyjj5IcmluEh0Le4OaAxI5if3TcC8gPdiOc9
7SaWqR7YPV6UiV5YXue9Kc/87oBMqdq/L0nYEHsu7DnLKQruhzeYK7jHaJUv6XOx1Wf0ahIeTruW
fSpV0j7A2B2LZpkiDaLLvVub4Tv2bReKagXOpe97HR2TSirCi80QIkGMHRag2CgCLsPAbV9zX757
XXgllwuY3smvIqFizSOa9DxXy0ROt/pqmhOM1gJJjT5W+5QgAqMiXb+uiAib6Q6oubKcQY/eaqij
U0Of5ZqxPNHmPwEdu6S2DxVDbvYHkvcE5qts/VDZRLbI7xyYpMgyaeRjONsYGN2bIMpc2pklGWhc
0JVcWF5F9JqYbhDjsIbka+pRIBWoCRlAQ1HVZ55L/Sv8UnlDOITMo+vmg+BSEV5Db7V+8+s9F+Ci
4s3mwkM7GQLjsh9sc1N7/2oOouOdPJ/tyA5q19kR1D0JiSQKFSUQFNMIgumBI9M+UqLWjquMp5lZ
go0O7MCu8+Nx5hfWuwihNEqXMYQAKs/IWxtDMingWypmIxjeojknZAjGWMWoX2AoUD6u8dGl3MFS
8oqkJM1CU5CaxrnuOgRKBkYOy8Fjxgjc+JePGBy0drrIzBTVQ2B60sMPcp2EcgfVR9JYmRHhlMZ0
F+mewSvjYG+M9eDxOlE3ZTG7Nsqb2iYnn7tl0Lzd0IJ61x/+QYocFrEntS6vKo95Wuenak79x3Mj
jBokeEAE4TnwFqtsstmV52zk3IsAdkDINAFF0xc5yDuE35MrxGOeU3IOFOLqSLHWse2NvvCuYqs6
MYG/RPXEerrjKtfv01fgT31pCg1SCXpkLWuswpPXIJK33xv1hT6lYbcIS7HdTfKecUuRgDMIJfWi
vMjyn89a3cPPI/jp6hXjwMWd4UafVAH+M6ddyhqQe/Nnxv68rQLw1XaSD3R0V/nmBR7QV5L7ZbKg
xlsxhvmxa+mhREX+N8Qb+7JaUpujP/RExLQLgex5s2MKrEpxD8W24CsY2KB7NBRtij2Q2NfWX/AU
/q0EN8JzFfjfnsp7VcngfxSih8M1jvHXxdUzulJOY2+DMtlOy5xDgY/TaC8i5NdNfvqMjw7K0vVG
V4NUi0hW+SFtzb0MVPVUUGmjGjCR1eCIJJJ5Lv+ldGCBts/q0scCVEnOAb7uDd7S8+BJctV22n2F
0jVm7L2ySXg2tzo0CH824R15nShSuss0VKWuDu0T01UO0xtlcjdF/UVZFnV4l/f7683CVaQ691HB
e8HNdkWu8YHYqm2Y6MfDEs3AwV2dflD8EZUg/1XM/szs2FyzfadH9c+sYo/SXdbMLK3b5VhdG3yv
7rHlbMB0fOKIQNixu4PjuiJ33/8/W3bGTXIyAc4lTgKz9Evko00YLk14zzBUkAW+itXXS8L/B3uq
LQMiPJvZOumdHTVTQVvDw4WtFafdtHVYMTIQsvNrve5iCQaRGmAECAhFD3Ao7D7xr91R1UySsr5x
hSCJNnqyH4YeSjdXepMuqY6q03FDxMwgScOOJh0jSSDqSp/T7/o0SY8TdB8GiELLj3lXEEQrUII+
yL/0/ivnDq8z7H6RpSE8OHBfNPdDvYUToEmIdIdvR+J6ubsoDxuM29YTG3U9vaJHwY7IpTAkNFLv
PYW4XvIskU63mm6NuvjSzmhq44ubqouloJqoryI9urX2s61KNZjQQC1AyZOosDvvNKOilwQdrtU5
U+3f18hgnNP9rgPKuGmm2zaqeFxh5HA8n1Nt7lfm7BpjIyoiKjCtsDBV4JJbFS6EA0RnUidQkc7m
Jx+ZXATn5WmT+d8vo+zxpb1XMvm0YV+bnyEqQf6Pjqz3SxofiPbTl3no2osv5D+QnzAzugTrTKx1
ZWzi86TYXCCQdM102HvP8/IcEkWuFnCO1LYVI7mVyMPg/HMcfkKshSAhwJevlTlg1xfu9aFufLiQ
FCntAf4qdly16GJ1njI4gnnvoVPJHwoylR9JRQQMCSMvPfVqTKsLhHNkTn+LS+MvYHfkYXQAjFCc
8UpWwzDPy2gAYLHrL0u2YuFZAC41oyFN9tXH81+kDYrEg3fbJxI5yIUd9Ct1+mfCz9NaRfW23eI8
n8iAwlwUYEUK95UbpPJFdRsa4uEOk699Ug3WIuMWc+iJheroOKVzs/sdyIeHUs+I/YiPha4ITXUS
w3+j2rOQbkj0hZLQ/d4kLZG1UeRSvPPL8SN1EA/Ndr1mctiY1uhuGLTlrvJx+PLeTPZwuJ991esM
uUVvCPHAW3p0/hM6Ox3tybQ3zI8svUZzaZZcT4UXkPoVIq5wifag7oq2Gl/PnM/7CYACYwc1rQQ0
S7SV4qmjagZjBnyj/+wheDcuHSy5MyJPyJF51OZBsMI8iGgQA8RW/9Jz9da7dDgHu5FBt1evzDrE
WXFlViECHpSSmq5We2PUkgVSkrWwz639n8jHPuZfLib3cqFs+fQoY0Ris0Y1+/22MVxhceCdbkLL
/7VAL2NGxHf6/8rIshq6DZQA6tT8pndd3mGDm1n/TYu8dlc2tdmar4I0B/m91oea10cArNi6+mGT
Np7PlKZjBaKgdEy+tnAF+Pk9NOZBfrLCT5gs5Dx92vxpw4rLXSAhEVOwjbndDZ/juAU8ngULNRBg
NyxmX0qFOHMdPB/9LptGROyia4UJ6cTKjHR7PW6X0tElwL4Q1fCc9ziU/O8oCOGj/Rz3gMYs2y1U
VirK36FX7OZAM8qIi0zMHx4a0UBeeh5M0qWyWyPAvoW4AAlDNrZF5N7WD4SaDMHXE2U0YHSSL0AO
BoSmfa5jTGtHvGLo3GoNw1zhCAzjrc6r0r7D+cSqP7AyeKFmdXAOVcDKH59k4PW/VrBXkkHeAB8z
nrSbfcBJ7+wr+ctL/zwP20pjXsvZG4am8LzjuSs7SgXLHq4tPTFFqMk304t18LF1/oouKrdXh7Xv
520VgFV6ZJo7FLs3zy5LL5mZTZWHeRo1A5g/YHRb21ezzOgsoz5h5k20BcYfiHXNn0blUOXcf3Im
JjDvtyuO6w+ICJ7DCPYqSAY+nJEjr9pl0Op8Yohp5YHfSPwcWCNHmFMxg79riiqU2E7+9QLXLPt9
wec3geBO4ureKfeTTwtCuHe5KOLkamHJk4Ikd1eAH6UA1S8TJrLdU8anjNWviQjqTWztBmcS3KTA
JaEHIEL5ySs+M1unwmqVfsQZbQbs/OnO9Z9CwxK1I1Ro2o+eeIBDjWshZ/2hAthqDCSxn2ZrX94b
XGUZsbc6lvsMlfudLD4DJD+AYoXhCMDRhSeRLIpzG9Jvnb4VXLV4jXZoovQ2EIEczPaEKORZn0QZ
PZQLDB7yeWLErc8BdInu/gflvxthSu4NmdQK0oTwKaMY35GK3B0jrVZgZ4XxkSV4NBGJpbJ6vyi1
D3zswv+xt4nsX2PP4WwW2GLSq35rtjrxleGMtB5pd9WPEHN15mfrI3GVNnccO5uRefj/CsfYFXIi
KNyxjtUbXZPM0G3vjOniDmPDYvL2puQxjWhofSKM8OkE7lihzOg0F6At7ZpofRmKFqAxFk8eq08n
7j9lNSPRZ0YqpfdtUb0zO0gu75kCGxIc9SnPe5AVxFQqwkTIQOeqYBnxIsLI75GctlKsS3RRShjN
1LP4fH9dzLZz+yfIKiu3fKJFm3eLlHF/WsAYzdGkA/xHB+97CEcegbcePEWyes0WAK9EmVKU1snN
FTDIgUSNVT5Dwn2WAJbMbh2GMbbUHIrfZGnefpcQ7snGyY/+iz4DoMPsLZyKrnvNMmWOblLhnFoE
0a5E0QfktaS3ec8+pZjT82ISEqMwWG3GoO/Hxwhz9B9CLvHn+OzhUmKcdHPZCfhZkGwrwOvEmEk0
vaVkFeP1yvJ9Lf1GNmXcew3yvBBXK9bcpjmsSn/hueB253vaSYUPA6WtbeayPsa15PB8uFol/vWG
/bCcDIsX7/V39rD/fAB6wb/G0cF4Oerfp0hMTk8/YBQaN43RTzXq7jcWHrJiD/iN4+ma6Jnvdjva
qYUisgro6RHmhW5Il62lqZ02CZY9hgIAPpPx2dwgZhSenGuSUOVvc64gSVcLv3PCCYvOecfvigOx
y2upwb4iuE1GuSGX2QnLiuzuv/HUuM6N28NnxXkmAqxuGG4eUqp34z6zQlEShdHLC8vGLjXRC5RQ
wJ7dJd1btcxyCSng6KieysxUid+5cP2ZrXg+hr/1Y99YtY63tfWoYUF9EPfOXKmdXXAbtSKGVJeO
2tELorM5oH3WQCP+zAJLBhin+LetnaXkXSyScAhVnOeODsenqQsHIwX6xd5nUMIpXQWEA3a/RDj5
nALhMJikedsEs0OwtbuIX0kIN2awFy0h5Lqos5pmIhRhgAe2XdpJwzYZ26QqMMJ4LS9CM2V/IYb1
4qD0XMQlJYinTPpURWNCX6RrUyWAuY9XoAiEQESCX6s2hO/hMSQHSADKAvfMadWJeDLrrgTafvZT
vPaKE2Qn/vfKzfWlavLoqbu1eIi5mESMRG2pEQghZKOaCA4T2nRdhE7j7UwcaEOE2PDh1oMgItiU
CnrLpUp+fa+erB+yZz1uHYG2NDtAnXKlEj7rd+nRl+IpIcfV9SSQ8XrQeOs2ewizSEHvCT7w26r+
tTBOVKmjalTTwisoPQEF+koAdfK2+XTlgbzaFjY2NiB+5q74TUZqf3ee1uN0GH09kRg3PFKiX29q
iGoHc1+0yGugXV7aXXL5RgpKide1PEWlfk26APKHjW5BhBnGOYMoU/iZmweVeatqYv7hgIfpc5M0
GJjUjXoQ1JuEnmNSbIbAGZ95LvGsLQdY2PSoXl/ZjtKBhcVUze0lngKUPDWTUo/DXPqkv1DSDAEB
qoXUMH9U7eqcIb6SE/lkKvPOSR57NxwbbA9U7rZOqcMGwAKVaTJmVMIYm20x4/ukeHkbjff9Kikc
vUyFvDLKPvKY6e9nJ3kS7F+Vc+r5wpux/x9j0Rhh0ZpDX7X7tf9fvGJvmTVUAdpEk5+bhB7uNCji
ta0Ox5VPF7Fl+qce+LudahxcJJHMF1T8nvw3YGvWp2GewHAQWC1shSph233pwwlZNCIZaAKeQNqR
XwwfX6j7rwz8ucfZWOq5+4SVYiTZg3Jrwwj4bot+j41jlf3wc8lyqi3LZzdZiDuyXoePeVRiVKIU
7RNxZKG2PDpBGlbtEfDFNdAiQv0wcLGymcq0WgErTvIRsbMFAGNXHXdE6vXX2tewj6bG8mDchP3f
zCx0Knvk1OKl2+L5zSqFoiM2kUx2acumZmdh2+aOuwB/5cw/JWsUXaUWgxmqPrkNxeqCp7Ih+haf
F5Vyl0NTt1r9WpzB47YuvvP2g/C6+G7SmTAgSrEJeu5TWek+pGKMEBoVGDBMFS+LgefhfUNKsNbc
WFGLGB5YK5aPrGhYZPmInMwSEKR+SdTGqk64gSGr8bkXAkAUhZlz27xNb0CMqcEwP6c/jyFUEJOn
PMxQAhVy6V1a2Wfg2XzPaXLsWyM9l7fqSa5gJrEf7DqC1dqIhU3COf+phNSgMYJ0QUbgGh6LGWov
hMRteJdIN9RAlBSbPgsqVl3AhJuzXZYc9gBE6mt7xU3VpVL2EOuVKgRVeOUGEH7VoLjGp0YBxWI7
Td5bmP5DyfKuXEPQ35c2IyuKJ6HMLARm8sHhEabhhl+pWz/wXqYOWqTai9m3ucCKOZX9euExTb9g
fsr/JVqaDdsJjgT+f9/4lIAPlyCfzbo4dXt4GCRc2tGS5z7PihoItIKJmAaR73zAxyajad9nZOLK
6uNcP3VwOzvuBb+xkTZNhBDhax7FeQWek+rTRU1m3U5Th8vYSlGGuIARF5rLlTYRz3s6vMKQGzqI
x7uoT6LuAWBkc+uuutks3njcmIuoB1AbDjQbiPVZxwohRFlIpee/27qh2z1TsMMKwiln8zrlD9FR
owtP/4seu1yQcX0e+SOeM75XVTiUOE/TMRGdWTCWAqOVCcJbhbiGb5DawINeOR7N8peK50aPQhSl
mZ6ocX8jGmOPFZto72/ZSZYGcl19IhPe8wNlGiJgT4aj9auD6fDFaDFx9+JtKJzUSM5k0sLdoDyD
x4tbwVi9FcFMFXsMNgRYZawbNc7ZhhPvb/5f25P42KVWjf58aiW2X9wqjOegr8NPapDVWxv5dBlJ
QeLDVYmeNInsn7bftRlVq9aaaiS0mnenBBv+qTpiHKudebBNlTBIMrpAaxQQfPnCcRKpLkP5wXQR
Z8XrJLJ+UqCNvPP/B+QcsYAMPeFKZBA4J/fOBu3MK6y/IwHRUzVpBAT9jXX6uqozrKjuHoT0SUfw
v161DH98Z+uIHMfGHkF+YvvlzbvWCETHoIrGdwIOFFed0fU8kx+TJisAKC1LLE6nMqjtuhiBg/fU
zV8dWCEkKBZbZ7iX+vXl3QN4MWQT6P/SX0YY2p/xzqSWlesGQLO6ke1S6+PJ+8zfkxLfSn/cmoSs
pZD4k7KigJ429SG+6i+6M3YaeuHfWoCG0g1inZ7sYjhM0EmE66b6M4bW+fMTKo7AGaKx8t0355U+
GD9GUATkt4UaWmXbxDEC6/F5J0U2r+7Gd69B70/NFG4w8lfdEvrrKCctCwSKllvLD+9QUwth+oKM
Wa0eDt7i88xYmm0VhbgkLuIUqaUvU7cCzti5AYJuunwkhOJ08nJl2rOExejY2jGPdYHok/laTQAa
YuTTIYA34AJpISgdT88+8muGAGFAtHQvdHbWtulVA3hjKcQ1QSWf8doOzq8wH7IMcSA9EvoSgIlY
86w2zfT2DhRaM+QhOQZv35ALswHkLD0SQ0i+ut9Hnn58lZZCfZJ0+5MVDIcItknUu9rZS5xlgGjR
WjImQ0BMwW7vMQJqMeNdLQO9O77Jhuc8t0PGJZEvERGlHBmlVVPINlSNZ3t0bC5iSGBizcqWa3Xr
KMYIe68JG8m9Ecw/c5Qwrh+GwVBc23MNLfUtZfj8c/9eCKuaNy3v4m+2qW+zpycUplmFbwFDEyFR
cLFQvcFeXPC7PQ/zRIFbQ4yee8e3npgcoOBGLz3ncceDMsfROQSveS3QyipxdHBFGnA1sniZgv9z
vV+Uj20F3nekIANJ7LJiiAyMCxcDxbf69wjETBr8+VM2ji4S5fVzGyGiNeU9bU/lxmjgb/w/kdG0
KeuzBCoPxeXT/V2P2q2En3Z1rfDokTXYn7DfsyFh8uTqe/NIdq8Awun09gkEjlZ0DehJKqq5qJG0
AENa1qgBfLiOzPqXguZKzaeqlCZEwSdX3KsUxbT6FhiaC40hqJ/11rElAMMZtUOquP0M5susP2Zy
ulHDy2n6qOUBqNzd0FZK0LXxNGTv8nBfu6WTJ+S9ttqg6ed88fq9mQ19Ak+1zP831/u2JiPz9Zaw
LwijoSkuqgrZgSrcgObxgwV9NK4lnVnGWOblnDfp5rkxmAUAb81Cq8mw9up6bhip7TR8ahzISX+P
zJJvS+3NBihiPHssA0gA6dYDm6V0mstOv9j4oSq7r8H9kExVmFNPXV1MlG2xqL7WhMitjb0Ppmbx
QcySnd3rOT9hxZZig392W5IL/Lo4wjcERV2tbSegl/FNEha7ki9Drzxe8H2zo3Eh9svR91HCrrJ7
S44tbvZ5xyIHv/BeNAEIb0SfG8tiV1RQ7CREZp0FCepnYlx6kIKmtfOhCtWTW+YSpOSRNrtuzua4
wxclGyrtYt8rEdiTDvrb11wqgkrZ+gJyC1oAJIVg6Z/i8ZcYbn1Y3paIR7lPr4uZNY7ZzDrT+4y9
Yp+tDFFU1coDB3VsN8O3zEot7BulTHz854psRMbDzyRU8SXV2Jw5AA+yOQYHKq4ntUmBkREYw0Yh
THU53j3YAz+vCmgOER9wwjsUnFKDWD/U1G/swFiOx4puF8WWjCKOE2kYJOE6ni8/5v/+DZjXRq79
k4rOj7aOiZgKftaN1xe2dvOsLWohrZZYc+inxJKKFGbuuATwtrhUVMy2LzApGS4CGPtNszPCF19v
CjSYE1TfyPnmpMn5dpo4ZlxKn/LmLykjg32XN2RvTglsqsjxzWm39m2OuvYL4LfkOolOV3RynfEY
FRs2HSF5hgLWgNqKIB96a35GZQrBTHNic1CL08R0HD+KspT0X+v/fUjXgJzuiC7NH+Pz3dLlfY00
MIK0vbn/x9NckJeVZ4vuIen/x0WLQwaecGRG0rplPRS4gGsDA1trbkc1AXY90EjuNVafYCEGeP1P
4G3jWe6jQtd20b8PAM5NIXXkNNU3YDNr1cdma/yQU4MLhTKWbT2Bp3GTqytSd1GVgUdLyl0/wD4R
uTLB27n/HmfLzZePT9tfXuYAQn3n53nFShx4QSJlCQr1BjkYNXl1MbzboSEF9kAfwbAV3FYYYAvN
xPm/xq66pqXpEfu3pL83o1Y/9UdCxBn7+f+wTyQqJVFiHIi74aSREcQ+IIVezCr8GN9YBQL1wuNW
jWbABUIyCIP5Q/CrIHuPNV7/VXOecEEQ7qW2Uz8uwUkPPqjs+HS0arfDinQ+F5jTVwVKl2oiDz5Y
MWrzZ2SUkyNdsBIq80thd5owY0lXk+OuRKVoPVieZawUNyzt+oTIPKU38E+y/VFfDzU59p8aQQg3
g4GHCvXPXGjhWslFQvn5/7VaH1oI9c8rnREtgnU9WQAK8prNlXU1Cad7pKy67bsaQowEEc8d93tS
G9BFwO4AmVklB+n7Zc+jLI/vGxnJzoa1J0pHU3l7Q8Pg+523iB/98oyvSeifK1xzbrnE5qejLaz7
ZOcj6n8nOKXzaWBNPxXfTcdykv02WxnW4yTEgtNz7WsUPEGH9uPEwcPz09Xn/7bN/MbRDGd29l5A
R9JNir1q02xw+CBDOX1CvDibFZxBop/jV63AyMcjzkqq94Vf8nXMd49kRkA4gRJRXTpyYt3SXf/8
4F90Q7FpgcC0bsZnYzHozUaOhHIlmB5npfhFaiW2HJe7suV2cdC0C8WlXfDi3CJUlgqzVdur3GkO
ZlQgS3IjgE+M2J2ldwOgg1UxFkxOLkdiT/iJ+T/A/kfcVaH5NTEIRtJMtuAgzPX0YCTqvZG9xso+
PHr3xrF2IOqxrhZ7NyrnRerp1VP1bPZ4K+L/Ky76xU6AHI91sigXvGh5IU6dh7DgERE4zyVSN2s7
/ETTO6fQZQ2Zh3tQiW72ZGFa+z5fgEFuprLYevywoyh4uWmB5MITzAFjEGm6KRwrVfyWGNVM1iw1
bBlMtu2Snl2PJ3SUYpSEuOF21gXUVK9NqPhz/NrG6oK084xR40u3XwSJpnNmntaVB+Dek4f9/iRk
9xxXW9Q7IMXqt/3I3KUFPEgBp9a/Uo/6H5++jH26XkPByrFK02uPQ3FANX6CqhRKyOa2WxtAcHXD
h507lNGmOT7zcKOoEGfaCdAWKfN+v7YkY6jE7EvTLUe10/bn125vkJW0U8rLepUEhJGQBYFD9Stk
CyjxDa7kclK/jdpmt1HLA8dOWQExCOZi0z31L2lXZoN0v5hFJpUvBCAoMj1pP3TJFiY9NjcT/fH0
fXx7PiDgnJFcC7Vu40S9YhsJyhLjyGEp9eOGjeoxDBp5K7jiIAkXaVb1PGtcTFhemmOhnia0HJYR
A0YNXlPxDHVUwn0UcIWtPYDJ6ev7KL8kUxYyg38bBE9A+BBeSk6K2PjdE2SoUQUv+E0aXoeERbEF
LZaMtWGwVxp+CRThWxgWQqtbOCDjzRcoP/QgINx5ksEKENG/Fuseq0vugC1GIgiHJIrf06sllBGP
ejJVWIa1p1T84X9MOOkYe02XavzqAyg+ICCAmF+28hSR0XCTtQ8S1DkLYAUiwiP9g7J2KEwI/wLg
3ylXz62cAJsROZDwKxrlDKKFHqf85GQzb8O+0qbPgwzBKoCuXxftSrbUDX5tj5wmBFQw5gf11k/U
sDe/u6BpsqVi5v0Qybijw+6vTKkDSrqp5KLlFczOzw2U7fvG7IFS/o+KsjecONqgB4T4x0H6Zeac
mnoElifIM0rrIvqlHsrMtTrDjYZ6wPiimLAFHXZPrg6G7X+OQCloZcwjVN76nMsSJFPxGdySyvuF
5V4I74Yjywx5cT9e5bgLl22uB3uyB4pqy4MKeG/no+2nAnCOwynNjGPeEZLoLkbiRSDSHpQcNTg/
9VDJq+64FTpGI0C0whIqW3tA+QSzJLgX45ZUrJiMT3gFH+UV7ncNhIwUbaiHGQmNGY4AOzZAB70e
iNpV7anYsDEdWY/ecJDYMEMP4Cv3HYT33XnTRYVK/qnHtL+E91rqhjlZ5US8jUdIexbtwHncNsO7
FOQ7C5Ob4g8U010u8eQ7L16un08HdEl6ZjALi9zNar32lzff3M8ky3wZynJ+Wwx6F+LWdEh++0z+
H/WD5AEvm/TN4a+ETB3BWr1yVfn8cZqjSKbqybx58jg3+rr239WM0w5ztcuhQb/3w4Tx/3l8qazi
kdWVJaBz1PSsb5po7ZwD5Gw30zujTGqlnsZNyp4FWz6kxSGYqayGRE4JemXw+lBrzEjLo9scbwHj
zftvaPf6SKIp9yVWAdBOC9JiGkeXxWiKWsUAiKNkrerxDTQTGT6NOvXJ4zkB4sLBmtqGjOpcMXas
wW9BEG22iDjKbPB3UPGgEcu+Cxr++qxUoy2mhACVGEyIKuWy8z4UTrXmIZCHTYwFtiKLqkJgK2iW
SLo1UGFooAzD0ywErr29NHtN07tfRKEq3v3Xbl9yrWf4/pksarkb+DsFJxFzQRLP6vtA5aotcStz
hTmf/OGz+8QL0Eof4ILauPxs1MDqKq70P01KKT5lBKz+6tnev0jTz79aZSlN80umQ/N30HwzXdAo
y4/gJ2ocRU5miDPK2Jijmi6S93xhjOJhr7erKp8theS9yWeFIT5chnS7ssPPf9gj7oSk4BmgkTbi
SLBrKXhcspWb9Cx5JFC2ZjwWSXOUa0qG9xJRNTNm8V1LzX8bMHbT712h92QdN5CxV+5LO0+Y/QhA
5keHm/S/iNaft2tUE0XmQbz1aCGpoEE35d1bDsHY+CmmEBlHyDGYEwMZt58oC7dzH+op0aQepip0
EQIpvaal6FJtKqNNQfDvinUCj8ZkxzCLWTRZgIvB27H9sOcTXQSxwiGfHaso/FMMUExU9kitoZrH
TX5eldSxA+pq2CMSzAiRLlokwd5/K3YCHrWqTwiCt4dQN0jb+EQfZl9fEtX6N2829HYkMQlgVwoS
rL46leut7EKj60XKz9Ad2nybFYD53UDYBqJ5+5SvkrTF9Ag8acVKaTHAzyV8gIEHL/jFhDXwaIrh
8kLclazToU8BUzRNrRcoJgattRdob7dMH9b48JlAgUi4EePfdrVPA5fPJEVezmNnPZ1NJlCmgnSE
KeGCPQL7cY7oXFUbPtNtwm3zV+8qCW4aPXn1aHlrbizWZemx7ssV9valKSJ4fX07eyGHI4ZH7FUF
xYS3IQTQ35S0Y3rM6z2cMO9mXdf4xkBBTJJfgN31Ch4TE1PJH96tRmpxZB1C7B2ioD24aD0UlvB3
BAnhXn1MqMyQNKvX190hV3fMd1ZZbByEqbgGz3SJLkTQB0U+Kq1WdPNySNzk0iZFS/atEinJOjiV
4nyYw7wueSDx9x3cKBK/wB4OL76yXFO7u4GI4rS2GvR5+lAxhpzV8FW0z74HNrkcHuvYPgGvme1o
VzSUbOnKgW5FGX7rhseBxmzri4mcNjIu8aCjofRM8EoE5XFlPPbYO03h5Oe0rgURnE3ELd6jOKa+
ldY7dYbFU9PAed6CviPZpb2n98/7sBjEqsdpimWJdng6KdKZKUE63zuJ54bY/zB88uJi4GEDX4xk
2g8M/fhfTDUAvRUH2WODmZAYKRQtbG995sWVpl4AeUTocZgskbQlxg7EopPsbUhulBA/2u/Q9mJZ
moovLuirrfX0HL/6lGebaFy9Z8o76O00byIfZPalyIyOdyMNkIKZAoFpXUJuzpn3EqRf5BSCZ6HA
3X77R5bhhcHY12UoHsZjXBPufd9zAunijpXfthNbA/jz95QvLMWLpxBlfqSD7rL0zYv1YGQoT/M6
BlpYv+gv9Nj9AL7adVGltqf2uZJ6UiJ6/vlCk0ZBEmJTq25XYRRHVgMhf3lZlZfsgTBUjN/I+OSl
VZ8pMvm4SPUeM8F5vkcI2/tHJu1SATKdbwTph1mbZAl3NMayU0SA4IJm68o/Dsb+KXi7dPO6LPjn
+YObQypuk08xJTCsMjBJY1CpKWbyTPXpW6t5eFm0fG0zMtluI8qLQTnCweUZtzk7LGFmbCf9zrHx
+IAcoSIiybvSqWzpeX9eKvBPaHGUmUr5NeXLh88tUGaaOn2J9Y3lvqPcPUt0W08N8fwNYcpb38JB
spWln1/HqlipSkk0463rTjD2iGBEMl4AXugDoSEbdiisZEW/HPs2aBPh7F30DHQspuGHw7vwbsDk
oPLLjZtWgBxjcKkMtSzNQSBx6Nd6OLbo3etWyeWXIBlxITh67x30xFiDy1Gb6is/wfWI7EMqxwA6
Aud8rZOFvOOemQ2mmoYiV31AnnsK04C+HdBRWIYjmhEnsk9rhp+DqIv4VtIkpA6P88vdpXygN7oU
q3E9u3pSmAJNMkKpzJIEbYWVYUwLDZ3B6oiEwkuWJcWnIs4nETZHZmZCFPwUaop+i3+vJOS14B1B
tNwJnzVC9z928ACxjEU5lOCm2bUvodXgWWj3HjdEfK0FzfNE1LxLILwN1EL7XuBj4DRC+tJClPdC
9bkqSiE8d9jgpFdSqSIIii+Qc4u0urVZQnsNC9Tsqx7ViMAjb87ymiywDSLWSYE36zkiY9kRD3fp
iec0/vSbEYGiwAOy+dMPjaZdMvx3RZsKreBIsOqgcJbPREWnqmtwPpuHPqepiYw8aVUP0bRe9Vo6
rX/NdDaORizOHOo2o5qGhS37bphvs8P5CHhaUH65S9OFO7d8DxazvQv+ky4CXmjmk0EWUv4hIh0G
gkoJk1IbrXCVGYhWI63zQcJgQ+bk9/+pbJv+jXVM5NqI5+7feudpzNmJpgORxhBfiMn6ulMeqLf2
GrnLpQWzFGHZRBUWyVSCgvE7581AGnSicV0wg0K79jHmA2ni3hKwY7CTfbYFSqSd6RBZWsiXLP/p
/X+posZ3ItitKbmTShnGA7P2WxJkKoKfWctBBpcHBEpjG9nbXrqyH9usd36vGeV2KcjB/Uh7ZGAN
Vyvl/pGJGJ5j4LZUJx+boBoG2BYaJgG/hOXnOFzJecZhidiENrlGvLmje1DVvvTk8Px2wK5nQjIY
LWekxYPkw3x8yQM7X3TewQUO5NofHwB60xgOaxOJSlEDe4TcCn12cCduQE5VUTuFFACbWoZt6nnb
Do0cA9PCs0m6z1DJBTN3yXHIFo+EAeMRXiXRNjiPGv7P36btMDrgvzcCmLLKU7fkcw4phrIAjduv
3RqmpG2L0QKHP1LDXnNiuJLlS6VuZ27SLbKjHBL47pz+GYKAa14/PEqa+JRfa6AXqOIm+gfLuv/l
GfzQt0HUuR3RwBztlcnY3TagiTirbRxMuErDqJgc/qereVKVws07dSN/bGfLgKlglRtuaBUjhun6
I+lNVUHGVikO+pUWyIB9FnbIWbvXraUKpHc+xu3fwfD90wN7y6e7DK4mo2jHjrHXnb7tNcYC1XDn
ayjOTnm+kj3w6BLz1MHcjaBhelg7moEuktLsBT2yfPj5JuoVWQ1IsA5LhkkwEvvQoM5au3lT2rhP
96lla77chG9CIiildAICmuizysVOBJh9kvbtHHLGaAP4owiM1wD+woJaeUg4F2ansGVSpk9cgAq5
JZDIVYUqHMdu9EZOeo770IGpKdq++7CksdTasXf55x0dEjutOB2pqP8M1rLZFnT1wB3Z2UohOziw
XAUk6veUVUTcF8vTCi3VWguTzv0RjoyN6G8IYC0V2X4fc+iHiyDzUcKbX180fYp4xCFw3EoJ3PdJ
O/Ok1MDz9MVwCXDI9soLTzb1LWFRLf0+tjbG79743Dp7o2MA0efLdA5M51XNbLaPMOJnK5pS3aS3
W3vzG/9dcj829ufwrOqYue9OuH/k+IkN/bQf/OuejNDfnr+VxmqW+6gQNjzgriy9Z8jzrhxSQm4L
bCMG8fMfrAt60ujITXJZa7mTjLaELLUbNK0ChEHuIR2DoUoyOvkY8Rx1fIjgieeIlJWPhflMzGm8
GnZQICCkvHRtljdvOK9tkYmGQSr0BeK/OJ/X6oBOpxw+FV6vKtBCKq/w6Z4/j5RGcygUr8oCJe7l
RMYhl1NOdjMy2FDtbug38Y+1VlUPA23UTFVEi48vhvS+vnH0iq2xMGZU8BlQSwThOCYKK0nUvp7J
qd0lN4th92n9GwqyGc7FcoDFhuM7DuFmCPmrAEeMDnxYHpPgUuzFFwXiw0r+ETa2U8DA3lXRkhOf
B9/erS9sZPToQMpyOnq/EAMLkQDWmfCK+nX60v3JQm7SZjQa2E6kod6w5SbTv4nhnE5AzRNTs6FW
QbtEEOqSx3YmkGoCZzrZSHQ09d50LdvmdIiLfPaVO44diKIbFRJwB8h+uBhvdGD2JTlju435HarJ
hmp7uLCM6QCJT+x2YBOWTvoBqq/kPqjDAKvuowXywj7kuMxiFziWCQeJm7/4QKzx28XQf+9qO0OW
kRNOSyJBYr762Xp7G2vwVIu59EmXlQpQn0eWXPsp79JrRiV0Cr8ngeYELK7x2H6iwvloX32CxQfu
t8DWaEnbeAvdO3lsqCPgRXLQfc9hXdMcL2UCV/2qXSXJJVnLmbY/v/4Tp0Sx2huhBnmhZBYlvtCW
CB5zZEbIJUS4yVVPE30dA5MmLfAXJfjM7Na5Gd5VoSjlFL4m0yMBIkE0sJt4yiBzXRkhzdG6bKhR
QqoDHP97s+Jj6KEl1/Z9KyJlvEVobuf7Ityby22dHFPKNjCkaVQCvVdavsEsWZIedQmPof93A4ZZ
M9tn+El82nMs3tOPHkgPen29iSZI1aYqJ4UNFmufDYNUEzZiqwEiq19t3pgXR23IMTj2zcfKig9h
DdM+VddsjlhKJRDBvrpjrxu6dCrZy97IrrVCPy3GrOH1NDhF5ag7Ou7H65XGt2Hrf79kfRn5m8ll
hQeECj0RyQMijImWx632P7f0nQZSNp5hxKygXEVKiAojDfpigf+kX9wdOAIzEbvoF6z4lLDsNMRo
A2hUWpSlVX+Ga9QOYdyPQvDdMvPR2RK9gabTAdoUgem2YR1+Iw3iubcpbaY1nRk3jLA0brNvgNse
RKOk51BS039e6Ob4Y4GBNzpuzWzHtzx9+QEfNpV4DydboEy+mV/9sPy8M53qfFoy+osoz5fMw2Uh
DUmVRGrTQ+0bW1ay6N+kOYO8Hqf3Fm4CcwmIB+VoD1M9AJpSkFL00P2G8kfXJBr+t/hDPEG0d9sT
AWsWCQHei2Pbh+GVnHGVQzWrZ4PYs3GYRNpWFJaiurPcQED4lP1oAGgU2ta/gdcCY2AXnZPrpCY4
vY+J5EguLrYFUvwM+71/yhUB8vbI4Grnk7+XgaJbKtV0SgaNAQnIVDKw3OmqZEz76VaiBWLvwJoo
zi87wJuonQ1b1LwQpOnJ9VYrj2FoKfeF7CdtIPP8uPsuWsvirQGHp5vPcAaLrtWtSZ6h90g/WRiV
+7x9Nu9F3ARvdZv8oV77Y4OwqhOdpfKEc0TN4v+gfUUFdg/BzvOcdQkhGcbj0zskQHjI6pggNSKb
bP5VAhHFv/tJELgESUKymlFLcqH0f06atFPMUPmf2ZKoHxJIeALKIz2tr12YLBQvw12DADwHtl2N
4cWU0T47CNhOQ19U6pJa2JAGxsPhEZfVYJduReX7oaoFSaV84N2IegYrcerkEU+4THsEK86spXq4
nPueZl+SS2OQq1Ql92SB7mZ1slBcJYKveWXrumiFP7aZt+snarRlmdx27dEZPqD8JziWKzBpshIC
sr7hea+rgx6otfUb47Ss96L4kvWNjYJXP8D6cBo0O+Ndb2+TSnbT8iztaTWXCL+viKPubf1mZQ+a
9ZGxF9gZK9gO9gVoqPl+/pHLRqYPBxJi2/SJz+mtm1RYokxQtdHpN+vH6licz1AxXs9kh4nmxRX/
yyaIUmRRz1krXamJboNPqO3USoJltc9foYik7BD/0DMGCANXLU9K3DtsjYmb0Fxrb/4YArpVkk1S
tbv6LzrLPouV0xoB4W6TM7dM4g2bsJ5Kk80oqkjnQftDvySNJRvcbT3ixF1Xp/+XT/fq9QbcIq+q
0b2k+qn+YH2jHxUnN677MHxLzX8TPQjnbmzTAieT+n/df+QB8l5c3bq7kT1ba/UBrLDE83x0HAay
SXcnLZgmk817qZ9vCYx/FB8AIsl7b4Qi5Duu1mjCrXv/hq84NJA/vyxIW6UDshmW8j9LWfKHGFZW
xfb6ILnWcXMWPi5p7DKOUpOB+vgK1I8hFhdmCr8GagEpZG3qb2CX2W6mFNGDui95gjs+DBo1NLob
e8a1Kygc07gp80hSd7TJZz/+ncIHMUytKhsDX5T5aPa6FkrkcR4g3OncI08IYHhANRr7dHD97kSS
JFhvyyrrzDcRMBivPht4ZEZuMCD9HNbHo3VZbWkNtRz+RH3UotT/CNx2+huPpv1t9oNwO/M4W3EQ
KqNvsB8xkSWVyEuAMyVefy5+g6fBAapS7MT7wzUVP+LQm1fRlSNYmummUeAQokfNndBWB68UDY5k
48Ekal9IGwl7XYpRPw5QFZ3Vov7Iv0SYXL8wIKRue25HGa/ZUCFJmmWdfnsKFQFdXvFV809JlLY9
n+JVqjOTVsmFBakP4u+PdZEqNksDMw8KgN447FA/Ad9puSuQY3pT1f19fuBXS99wMKLelUvBGq7X
mnEBc4j3jdItOvvRDeJuERQtHAJ9GnVajPndoFcVnnaBOSgdIzIy8ldMQXRKutZACE4wTm5oWNye
J0iwYsfabi7ME8helDXNJS73zYGPg9josVNOGOC0vfJth17jZ30RvpLttWSZCBt1W/gBCdpUtG/b
aG57Dv5GDbPp6yOo1uwAetearB4gg1zS6Qw1CWo0cWHopqcde7cSWvsjcUVdFtwUNtSrnk+Y8TUc
8H3DGLiRED2h0fMyY2jQUOu2eAZ925CPqu+473Hz+ydHbDBTOILPoGe5oh2FsBXcVF2dPHy4I8sD
liOhtx1kCZi51hPLU7gU7oBltI5FmBPuFEqQpId9g71FtMLH4w1zsEwZU+RV7lbpYy6jsCgtsSk2
svttIptpZPproRcK/AoraDlj9f5Lf/2gmtdnf3qy4gZrDFxsOkXhwehDXJxFFH0ZQJFbwS+T5CWe
YilK2CzjdHzG5oacnF4pv2/F6YwRzhtQqPvGMHiIJZOc5JidOVS3nLg+zarjg+0ZIc9mQ2BbOS3L
nUtV49nYa3Ura05N78gIwTo5zgeMkQfpto59atY2gTHkW7gTa8wgyHYLC3PrwbkEY+tN0I5aZBqC
sbTTUIFN//vEnBfec8QUGhhZ9QcVLwjZSUKW1Ve4vaMqutApcJAeXsCMK7LFIyNbsMirxWCRKmYg
kwXnV5/KoJLV6L5hOIANh+SxdFRWZUvqrTl87ouIzsMqo342jY1dAzCKlR6vJ9luCkiLYflmGCIT
rt58RSxJTftYkKs7P3UysPevIQfBDjoIHZZ4EsGK474ENwtoDfGUgbxPp8n2MrveFV8Cy/GfTynY
LQ547lMX/AJLUGGxChl7nBTcHOaLH85LOOSULeBFBbS83w5w8jSiroKG+FTRKWRcKWlZSGCePRm+
KETXZs9EaONNnboX67kUqxy33A531c9JRkcEkK//FSVX5O3j+AkDX8H1DxyWDY6Ez8JUNsSO96SP
GftMAmccTD2dtogGkWDZTEAhG9datGfJ4+gBAvK6NKR/b+twr1yvDxjh4MoKFdmnGzMDijwG/+Pp
O5rO4RTHz668ewxmDEd0SJMGlqT4l4jw76DdgBrzAV58EY2ngYKdvcH7MN/uuFKyS2kOAleShs59
U5JmYD4Ecbd58rowBM/Lw0Dwi68wlo/ldvr47sC//jdZSNXHY4Zp+HT1hGRZKAH6fCJgW09P9OOD
RSdCGpduXR1lTbOARTt3Z5pNN0WY2aEWV66WpmJa+cq0TFK1EwY10gIg+xJKXWF0a/bnje2dR6fs
DfsM0W5XOb8zAEwezkvMDzk0SEYZTvjk57iQFxNKhp9eAyKBlVsaUKedSHGxsQ2At4DP/cXZyyIv
qP1wsKUNJGJNHOloJWlxlrWZwUYbRG1mgIAnJIMlrBeV1KkC+UklHzOJvRNQ8a26mq5k6pmL5Jli
aXVkFlmw4kAN3libjqd+p4JoJzK8Omc3PTWlBPFfYjix8C5+tsctOYBJMJ2tzqKywLkpTA3fSeOh
jyLRdCZT/wNmwXvUgz4vq5wPAOAROumwN+RUJKvuJ2EdKYkpot894BCMFO7rYjD0+5fbOM4IAF0M
I2gI9u404f4LKotr0RmekBIsAH0ef0hDv6QPp2ObCu87q4Zre2vIubVqyNibMXZPUuLZtaG6KVOx
3TJbLJrq+tafJu1Pe/qjJqas8dW0IfHc2ZP1o+LSTEhbhFBViwC7ksex0bgotyODQZ8XeTn5Uz1G
nruQqcBetvYPOgMxF99N6xl/DUKdFkuy4AEjMfKTYYVt13gcD4ay83IDie6mO1lvJGxWBmXlUXIf
pzVFPSml396qxeunio1xfVkH4rd6Wg6yS5CYZpPUdhkhxnk8eBz4GMFKMXdtMiVduMvxkMdIQhHO
nAVrBCrMl6HWT8dnIV6WqPncd/OwFAADXTvWrLnMGP5ipbVZpUvwj+k8iADyXjP3yA700vi8FDU9
4TfiSZCof1KzHHRn9/9/CbanPAK9tfwz3HizF/KnhOW0CEIUGuyXqcLNmTgVELERAid3i8xik51v
ByiYZ2AimnLNqesXQdfJn4WZ5nA/vhrHuP6bUWDA9qmKg7amWdbYvKy23EmMwHlFfGOqEM+BXNkk
UW8jz5ANbZlTXbHLYnHhMGt4bW3WOab7MiXmsreymIOdFRKa8XDJ03CqMeHoqbTEPVEIrPtWxjtS
chXI2dnIcO9PPii1ZMJ8E6fW4ZGIDk4arVmII59i4LpkK6oji0Oul+An9pqKD8yoislTH9M2xYMC
KKugNnGmkReQUHTu/SLSNhuFjasOdqYliKecGHBguUKcL+U8MLktTEPH7gd+JAsMeDPAXikycReq
yyhRvYzQPKc0rXk7acfxnoNYHgVqy9mXronS+nWmuiMa1NV9zwGC+ITDi+5lhe24u3ewJsUCmLJy
cFKNGxPSgPys9A/U01wmuyOHYk03vJSqT+0LqFaLiXpkyBE16XgjbtLlWLs3yNgtS0XVtdRJInD9
kxj2ApIdSW9yD3/MmS9oPlweu76/pQBVE129L1CNzxbhOFbkctC9phqutbjexWOQmCGwXqhgepYq
hhHCSAJQwRsZUVKdpoNBvYamplKIpuQJIkPq991actFEQbTupMt2xSVixXxZD+raBI9G2sWggE2y
l6ndR+ce9VOxOv0M1L+cDO3/s63D8WCussHMkhRIfkc/ergNZhO6L6scOgCkjZkmsj49zMcOi2Ca
CIYXKxdgw3zhWAtVzIv4plYRrMicX/X8j31+X3Jw3bYUSbKpVMCPKlIyKyvsxqVl2W1HtEX4aT/H
+6/G6hZughk1aADszu7U8PquIWsILe8/jLOewBVG8FWVw4/zgSXM5fw+aSpUvlUk/hod5LPnbUcB
+TZRx8mXM3fqzyqsGoDsiTxA78qt2xyElAhxDbbgQj2+ARcVW8JR///t2XKIMfNkTFdkFbV2gdNE
qbwlS/zj6qsBc97EMPYF3/87xtczy3aQgtd20Nh3d5wNMiDVLIgENfHw7ZtVK6JqcrB/y0e5MgW3
pMkgLAu2Drq0aBSCgpEBkPa0U0Qubzv/yXBtKnBAGnOewYnO86w0Vy1kfHLQN7PD8+yinf0p9PX6
rzpjHBFKNxAMHVp1vM5eUwIHj2u+waZNgx3qb97kfzcEg1b6+6XdGp15ehVLAPpL0sUjcHIrRmNA
C/SMvtm1XUeXmz4Mvztt6ePjZvu5QzD63aiEqHhbDpRviCvVVWcuiGkzbRpDLpY56fMn4WHehbSl
oAxg3ra84ivzS9H7mkBdNSAzHD8jvmI45x5qgS2zxp6LPxN6ESMaOkWCMJ1/2KM+GTJtBOaJMVrC
7QO51qaheP1b2jPXHRYDQ3IZt8o+kv8fzf3RIB9y+fOiOSR1+KgI7RIholHXENnnqHJnPHPtv5gI
9DQcXDvkN4HrhQxDHEDk91CkGMOIpHht0NcZxuDh5lrC1gc7vgUoXxMEaSYZZGbx6C7fghC0gzGw
N5zlzwc/HFwAxcBuhmOft59Fv/Wk/4rwb9wHsNuguWA33hTyRLFE1lDDWbowH6yrciqChrzGchhs
RISoV8lBQTxj7q8LuNPAGAyscaEhV5XMQIClZAg/dmLXhJsF9ID9K2JDQdtj3OK2rANjqvufJFnO
hE8VHaAWi70UWmJuM9U6Xko+Vipkho+7Z3BINVKbVsy65nDRVEHWQWayAYBiP5Myn3IVaGMXsVFz
Kdnd15d5c/5MkQs7g4lI+9CdhPRCfBRTKqpV6Xw1zGuTJq66NFrdFgufZUdx+XNXw3K7Xs5JrWG8
mMh1JivMwkNjGlPeeDRvR4WJE2ThS0386Yid1cKkshCdnaxOq8VwAVN0QBJNIsRc4tlsvpCWx4Gy
DW2I0FDSOkGE7MstcfrS6wnzFruHjxduRRHX2Ml/yBxBAuEDrrAt3Ayysw/oyQuBUbIaOtM5L7/3
x5sY9PVBqG8iLVm5dDN4dHUQrWFiv+HBZAh29i3uodv33+VKxZW0p2S4ACIyJOsE6H6MgABYt7P2
4X4ae2I9cj4lnCVpKn4tjg6xKNBRxfuT04zAttMdzEmGIGDuxd6KKc3qFNBOKd3G+/8czmtckLqY
0Mc7freIdaxB+Tk3Ti27DC33cqbDZXve0n0iJ7S0nwHLyLdG6ikCi2QVDbHxUV1eDliujavX8Xmf
JvDljvDTaf/moMvCE5SDnXfXAASKkJZykwLxihVdbbezUnl6jdPr3CKDQuuS3nq9OKoROvrCqyoP
Hu/qesPa8+Oc2/KRmYalCpJxhhXirN+KqAwYs1I9Q0VsBJ7tKiCpfixftGJ6ywi0PdbokkoBqXOJ
OJQm63VXJCKnOvQ/aZ6s8auzwK0tK4TTTJCfhnGsDajUBxqVBm6w48A5qpS6QxXjLaO/4w4RgQvD
cQLPmJ4jpkPtAcqCKZ4K5k7jRsE4CbnxHhrilBRc/IUWN2+NrJb8EOGvPGTI0gxq+nF6z6ddnPz+
gpEYohGtGHRwLHZ8VijOJpbgYCl8jU2bGC2h8lcaj/AMsaehCe2dcYEWlgshSPK6d5MCoNIwEZ6q
pM5zridwlWGqH0wzqVHnfNIKR0H7agfoiOlpioh0ASZU5GSRoymcOnMk9PseCswoxSimCCOwa5Nn
rshZpayHORFo3PwGppJcDfVtYCGKHihFNWc8TC6IFNS75fWt5U26GibS3H5h90/M1jtc6sUIw2rW
EGtH249xxte48x5KNvieDDE9N5At089v6MUGvDwZ8Xy4PSnlv9sfiNcplTFK5CZw1NXDQfrsce3h
dxMHXBTMBmmxbfxsFxs1C2PCV3cSbP2zVCTEqAYGvBOc2uZr6z5doXe0v/q6cubpdA6maSS1snWW
PvSdUSirMsS00zphrtG/qe692O6toGdUvV/YNpKzuDIztMeFhXRnOK1xfJUsczfUCR/0YfeBrGlf
OExKnbCvNUUrOLMw51wDES8VB1GukUOspHWPcPkxG7akK16IHefz4WgGJnrrfDzy9JaSTwCcypoY
nhTOPA5y0u9NVWH0QEwwnRbAfDkBnxrTdj+ip/zKGUeiKrBUWlI/jQtxYFnVfAZZTP3Gx4N+0Yar
dqEzpmyUDDzFQABbDYBhTf8HKDsCBWdxVo/p7W1SI6tlpZAj0rBK6lsIBB3OUG6IjOM5eUf/Q60I
/5ha8WQOL7uJCYIVUNP14vhnx8k8LNUfl50KAbzpUqKVZVHtd4T9x1Ziicc1QeO2zukP24YZljK8
weU1hyujY9BATNDsGIjbIQZaOQNG/FeUHg/6yzmivmFI0p1PTR4AnmJSmwF65kpFPf6dYwswgK5b
h0RS/31kJrgtCY7/U9jaZrV0yJKVaPkOdEtIOfJlQmohzWHPz7VOZBX6d9EhIoAR/U4oIKoS/snX
AGZ25GLmztmgJcSCuZRuGiNbcVLsrkInKXrYAcItAQ1txNOUIaGPDq1GUXbwyEKZA3FGs5m/5rqF
UENMVPrdIHWColNtPL3W5uo66+/XYmzwYgDqAs5P8QPsrtDIdDkLddTte+wWokGMeH3Kf8lycfHT
g86n9D/GStvV8z0V8rhHe3A4bCOh+HnvCIyQnKKOjWyec0dLlc6dYg0pEvi7hM8qrMs7Hb0RFuPd
QSYiTNJjKK21qvHtuaukSNj1m3c7Vn6b6GnnzcIGrbcWw+g+xc7XXe4GjD2PQfag/pLH7fRdMiNR
fiD1H9E19Bmi6ggnPcE7PfR6FHk1sidTXE4gb46ooDonPTBYeU2bmuDmpQEEkVGO3g+6NqdWkuZR
tFW4rMFngbWSGnqdOlq57yJWQ7oAdaThItBw8ZC0uBrqKt7lDH9a+cR6RtSQCIXNGa8Z1Jnfekoy
59BlDDo2PL22Ht7b5vy3gJWWiI1fVymneu2ZQHIifNX4gvTTCKk9vbkXZ9jg9q1N8ImSwuDrjG1c
VU2XkDvMF3N/M3YY875cJWVzZC5XjT61ysIdHHGQa5JzvcGYXau6qbMWWAKELV6lci8EkwDbSOmT
mqVhdTZMZl9JkME9SemeadNsxz5p40a6Zq5KyqZ9OxSpeqYiaGuHSwCg/LSJz5FXl6ay+sA9FKFW
A6MhdP+v5QbrKi7I37hctqbmGkmfsii3+OviPFvv9NwY2HM8RJbzavOSig1lWpNMZ5ebbyiPQ0Jo
CE/PRJ1h7q475/r2fLTiHsSY3V5cr/Fd/j65gpbdq6IBldm+Eyq7HbUkpxWGbAZKGj2flFDy/ymE
/nT6jFRgcA6W1ouvWyI3RwThNh2SHF8pQ+OZKTFm3jySOUAnWdCVxtotUEGrkLHwTHHYyjd40c/V
lc3HZ2UCSnyAsfHe3XfuDwhk1NIZMTWGOHzB35M7pu/PF8bbiM3nzY/2urOQ4+rp0UfY/76hKB1v
GS36diMHE8vGvP0p89UsZAAWnmjSo9qU9trBHiFJ3H8kQl6d1K7PIpbEOef16TZxk9eaKJJ26tc6
g4rsXfusPQIsh1zsOhSG/NrKhKyfoo6p33IqO0KzaOok5jCSQN5olBRsQnhXvcev2WgTF1JSPfRa
x5sAMXWzwuzLtUqeEys3e0COR43SSe2c+jgCIj+XkMTAWO8kmVHZGYMXxSttdi0L/Ox0U7zF0Qn6
3qFz6Mlb/p9v830bELkdollg6Z4CYKMWXgxqUjTqhxTJvMoAIE2mSsEIt2IhdmtnfGHtsXfT1udO
NM/pHkJcG15hj+6TE7N6Labm72RXdCtHX2V527Wrtu+5y8214CeOJgb/aXJqjrm2xXhRgBucOz05
WjJUF2Nh0jEx2duxVxHNzNeZJh6KIOllM7Y29ydBye9A+/TArKpEMFAP84OJG+axU7kEefqaB4aC
yPhTDkaJoJIQNEXRM4cV5gsich7iHRXZpYTBcRdE1sjhLkMZgjizeJYGyUQaaMQCUQpdKdTaj6XH
+jzrQUQcGXQSZqxjrbmSrTpN5l9EUqgeS3AHtHS+KlL76WUI7r4iKim6gSWkkO7Om3UDASjehG3l
oaW4MB7niJfSrLNUiKWRan7hhheqq2MEOXAPdPuDas+wcN1ADMxJ4P2/wChydQB+AeGwdF5wb/61
zwb7ojXMyt8QJLrKPVwZO61LVBTadUqLBpqxG9Vd9lW8qwCBE6IW0FTah0IeAsC6F/sDDIx5lZ93
jLH9fMh1IfTKAgibSLvm1NQHamHtqlMUA4hR+7HWm+8CSqz0aZEsAOTVjV4VS6efnH3YVqesluZx
mfpUHt7+XNoShI5FosjDC/v+CdOVMGx1Jg0esDL6bPI0qZQaU9l4uuESEwWP+v3vnJIwqm61fG+I
f4blD4RlwRwm72Jq2sKXkVpIEll4OVMqavKq4lYAMB99OleYr3bY3CwBMkR4qYMO3zt8t+qX977e
6doBwjd71ezW85wjOZyzpR9f2tp0oz2tvBLMv/v8rylN4keTjEvVaWFeukK8mIrkmKb3WZJtr0Wk
+CxfbslPwx4SUn7I8YlZIVssbINRdXdGHbnZ0cBRC1/ozEG+uBYWz2Lxnf3BiSPdhd2i5WGnjGRU
Anotv9Mz+z8KDJSpqi/9NEu27s6FP+DZfDjhPM2MK1YQB+Kgcd9S96JXiVrZr6/pCL0+9HNszK8b
KRl3n/RVsz84jwoOI+Ogr+JpQ/jNDMQ8+asS6kRRL0/F784qQMZurCltwaUzWFb50gmlR27b0Vvp
t1LztruDvosSGsLQVBK0J5L3byWiTZWOsehjNTQfmWf0jg6Tx6/RUiRM3sNfzTVN5HHdZT+dwfhN
y+3l4ma2VXRWYpa3YaE2i6bbrTfFflcDUf1jvRcfV618WiVJMdWB0/i45HadJlfbuySWOHd/kfcP
Hg25bW7OSR1C3drUkwqPTFBanYnAPPFyxl/hzdiaUusPLFtYQaiTN/3k3IMBPP0DB0KhzXGF2KGs
+I7+jF4vD4W+9X9X/KB3KEduDXbeU6XOfTD+9VhlDJ5QDDzHnunFej5bcGUtxmmAO059kC8epKdI
apDWQE0SjAKfgJ8GuHBRd51LAlaxiMoJBeu2Ta3vU1wX5EoNoJfv3lOSy2R+y9S3EJjciUkLBHgf
0x+6tRD2TmD6hDbRnIAnUNw/ctNonzY8huVayTF0cgcEp7pU3i0+kgjwg+PytWbbwqiQUnqDXWfU
k70kuZeiYWTgue3vxi3Q61v4kY9lcXWGlr5TVDQGJjwb+tnggQQWvUe1ystVN7OT2K5hEOWkrYmT
pVW5UvJTcNDsOs6gQzOOTMBN1g7kl3SljN/VvOoqGf40Zmuxx0CymyWfEfDVWwWrMBoa1s11L7/U
lV/X1ONriNn1pfvhhoYPv54Mp5q9LehNXEYuMmqvgYXwcjrb+QwsAhZSzheYNiITxEqAzRUfa8XM
ortsM4SNu0tTfTcWcTtkEhSX9l1OYEUZYrVz/vyeHcNBJq1yF91O54ZxyZK1vQ4Q8hB5m6IPhfE4
QKfRFCb/oTsC3Q0OXjPg+gnXgJAGMGePz43S6mMM9KMTzhqBSlovOSz5tRkNzluoJojv594Ieqw/
oHliiYr3B8A3LKDhv5u/DK3S6WGlCWrU9H6iNELqeBCRRt3lEfwHt+inx9S6TsWpk61c/8L4E6pd
pVVYa14fhwMVTGEVLT6voIDpoes2du3N9osKONLUZNl6Pul+RpL54LL/WhFwiqm2F6Dym1gaxNhC
tmIE0ccvwxGuUuJSPzGZMoGMC5HiaNMgF207zb9g8IeU9gi0FlX91JrJ1l87pCKErSq2AZzVbNZ2
CL8QKWyWGF7v6aINJoH0/5B21A4cuGGwiF5ez18gVgCT30LbTMVZy4pl7II6X1CjOn19B1VOb5aR
pVF33sWM6uxImDCjyirjACIYkLhQixwMPOHABI5peQHIPTBCsOS3zXktceez/Ka0ofxLzSYZzZPK
aAKp3pyoEz0Mq10f7yQICXq0neDkKc71Gcv0I0/KgHCbg3mZdCtPTo5FOiV1UybE5QCM+d/6HUb9
hyJiRnBulQVnLhAICRaXTndXb9XLxSmE1Q4c//OVdB400XJTYw+ZH/DhfjzmZXaSGMDVnhCsHG3d
s32WSoYgT4It6ajcDSVfNh6NtR2bRqkuz8ePIU6h0bM26B7S4MxHfLIbdsnhZjwEiLC+0SL8RA4u
5KthgHWaS1KO+6fK8Fh143XZL5tbNjIXpPKUyqnS4aeGvDi2z5B4urThhwy/38FV7rt8oOhJTUAR
WoDS/G5Ih5hgebIrM0vERdEAKfwLoOWk9QOkDQdDCIKkRGGRxNQa7wpSBDdUjy/I7zS+YetYsfiQ
j469CEc6J1fWXtqUdkjawxpPi8pbU5XAzOktLnucpts8K8Gfi8TiSqwzOq5/xlUcPUAE3rU/PONG
7ID4h4RLDT9ilodOBFBITBV8eLN0CshaRktsKCR/qRlvN0azYNqfvAZmQYw0bknknPhEICk+nOdn
dYdYUWkaP3i035Ei32SZt/wiywV81pDK+3erA17oJt0BSDkS7TwIqQKjDMXYX4XDTRUG9kvVbU0h
S1mJ6FaKSYGbG6cFkuGtkevEqReRQ9e2sg+KmVCozpPqhAv6HXwRRX/i1ryZJ9cMilOqg4ssi7G6
Q6+W9yaKM034/s1X9vntJxHopIJowCVuPFsCuRfqNI/8gqSZ70jr6uZc3YIJqYf5jp9Mfsff3XEi
0gLAy3eUh9pDZOI/AmG4M0OsLsbsAKCqLPFtq0ZnOZxNfTZeq3ROVMgQpjkCppaCeKjHwuSJiy+X
ezE/sykfVAiRsFE5EiM7WDw9Nwx/q3Qew46XuKSna4pYAtPso+l6FA/U/9XIhbRT2TlLaBNexWGh
TbYEwQPrLLr8akjLzw65beaT56V7sBUBkbQtnTOlbBFZvMKzzlQrSn110cO+H4ag4dd6aQCo6obh
VGjUY+rmHNlytXZDox34wU2JRZBn7HiY/Y92UUjv69zrCoom3AQ4UfOr2I7I3gIUK40Tkc3OnPsG
0Tw+5DZT9XxTpcVZPlADCCYMGJTNDS7j8Tl3K3Gnnso0WPZ7Ol77B9ZEKI2e18Uz9IPDPruD4zwO
ryFGwn+uJCYN5bGweJLs7Mg9kMzKiCL3NyyKQUmzS/ugpmvoX+U5BWdgO1mH8/TiNg5dAOgwQqMH
tutbvG/S+aotHH+0h0qLEeMDrvyTexNW8olSfM4tl2lqE26z+7LHe9FVICDhvxZ4zMDgCxVCf2EK
v7yxGb8q9e94beagKL3afz6KuPGDWnUdFXACnDktrWmvzwSmTMXmCgnBEd9kILawsJRRqnEROhDC
y8Q2f+09nz5mL3qOJp3jum2Str4dZAf5iYETiwTXeMc3kTi8EjGTesLb3EPf3mDlCGuSCZkv2FXZ
dJqmPcVekHRNYLlKf/xMthau2m4X1F9lQ4JjOOcarSjPizjq7cv1jdbxh1PsnZ+hSm1yDOnK7Zek
3r/IXsYCROkYe8CJHCGU/qydlnZy2oGzZBT5tHyZxtLltQsPsOpSgBgEFqehXLr98JfSFk7VSMQC
S07H7p4p27xZYTOFgqUBDgHzcvEUg7yK6CtxhW7uMlHi28Ngm4BDkLPkF7xFj+MoiexcINSmOTO/
qdaEmTVH/vsuD8NKIMsaRGpaTrngmbwwZHZCFe2k7oEewXK926OVMTOEn2CIywy6rZ+S4ZjbDZf8
PDQdNkdwbozlxnBpg24q/9uFVkwOJBN9X7PExTDLZftu/RSyHWjdOhSsodQ+vJvmY+9uL/LqpOEt
2EO19hQUomwoRLMuPN8bv6ACX8sXcwKPDSLv++xHmNnf827mxJFdUPzNk+8BWTwWvouDH7tja4CE
odLFzyEnJOv6f3pJ2A7IKN/wyIJIqp+xghzQNRsMTmoUZfNYx2rp82FO0ckVKUYM2RF0f/A6lEAZ
oNzx6OvRUxDcWHU34sMaIOB4NUSWMrGNCtIektvesBK4wU5WA7PMvyxB4VOCHyPVjfk1fOWqCsrd
Y25OKPn5s9VlW9kXcDpl3W65s9ZcaUGuswoUKw0cS2XQjSVQOqWt8jNVs9lQ5yMaveRHufdNxjAU
BNNo45WF8ffut8iySbQhk4QWNMMn0wOX3uLPuHsGbJBZS9U8dO/DIzmvIgxiGRZJ+mNvDu7iiC3I
OJTgkSaKZDTaaVg7lZBsDVb9on+iWvJF0GLAuS13ZKgk7VxzZ90DAkGr59qSuJ6+gXdVyeWez3Mx
ys8TYX8K1o6CML8jTX7UQioAsgzmxOWyouRmlr4qIinj8Dhk+QkrEE1dGMmSApNPFPMPKF5rnR8e
WqmN9cZEqBkSOlvam25SQvzduMpylpiZX9F64GdG/r2rZZOGo4bUFqBgyFOK3dQG4oJAZcJ9S63u
6EFgXWrz3Dh6Cmb9zjTlZxwlHwPq22eOM5FYVlxSidofO+FNRTaEGdL/r6OYL7H5593vkXgJWDzQ
HCQ3S6bLIJPm3gNy8aPMMq4u14DcpyNSbi97YrVnQJPbB5XDI7JddMbLZM/95f5m8xvfrzynQf82
uLDvLcR5ikWXWgnGJpKA3SO15xmwghnDAbb+rqOh4im18GgDNfW3kvFlZYjlAJ+lDXR7CkGrsR+Z
uv8xbemttf600RCHOrb03sMxPu72vzeNnJ219WvoXpbpwlvR4bGpjeI33abnvz+Qg/NiAukTqqMc
YwmLnAzKYSa+NSH+iAvQigUMMSbDn4Po0CkXbIrkMqwQuQXqmjKdOw2SGVnE7IvWn4E6TqCM6sCR
DY9prWpSgDiEHFX032UZk9ydMtzf78Svxr2o63fOweZ7BRohLX+78sxDVm4qgZ/WMYIX9gCkuopl
8GghEk3hyjvOaswlYiW5caLTR1+2SVRm+pWxOH+fP8EiL0sdu+tzf7FZPFgtAU1hDaAGj/uaYEEx
8lHjImzr9bJ529uNj0LHR1+hk99X2y8S4Fa2LhfrEWsBLO7nGwFF3R5UoMyjaIdrAFE+U+ZYHj1m
50h0eVwxJnWe2G6/xJmApmUZZznD4ByUaqUbIBXcMd9B0vHOJxdHYmJDiotMrmQI2UAd/ABN7wJi
i0BHsGhrqne8DGAshQizMBPLLdYP9zLGaaFvx2de00pFxTX33SIUp/qcgzdmUktRzoHWpchOJJUx
ZxLoEY/w4Pe1xRjaCOg4cpF63Axbybg4ojCJNh/8vKB23ad5ABx51qNdkWbGa88ETJ/KPAuMdOBu
g1wbDhutYd3E63TIP94Txov/WRLMfmAo4Oqg3IRYtna+u6LicycOsErGHmDvgbDT/iE2mq/TfI7X
LwXYVRQuezqgvdRwSlC+oSWXy9ncj15CeAaP25EtwSyr1HOFsLddj0rWTfsBuDhtVcyiSsWOJs1Z
S6eEnPld2p6Vrrz9jabQ4vj9YQArbI96PHSaV5f5heCkQ3crin/rG+lixfyoSOI7yfdnBvFIEocl
mXOy3omCEkwLp9c6t5ll78UtFBmFP0Uwdq/cfMIpCqIrzlp3m1ANTpauD3y/OLBynS9oaGHO9wlB
YRuuFwyhqALtFqOnEXrFXaRK5axDaylLKUuGTA43RkNn8k4M5ru2Algo02ql+GmdlHyb2oI3ge9u
ujZ4WSlkYeZh9VA850Zt8wHlY+to0wzBZQ4LYTDZ0B2KkreiBw/xMuJ1OassiCK72B7TrV4BX9HT
l46NLyVP8WyHtjyFMcF4hsC5psvHXn8rKfoq/HKCuH7Quvp1m0vtv5J53JDwYi3yjenc2TGN1syw
H/VXO8XZNlqOIYRiQ3uOQN7z5JP243QmAczG8mgOi/8wdAhFCsC4vvq/n1PRi9Xf3B9EZZHBwEvb
A3RSx2WWyF8XmoZeuHP8X0j7MJ/CXRcVfzrjKj/apJCS63ypw7xS93u5QSgptDkdz4KyQHOKOsor
CMSLWm7jAxcRxLbIZQRomeKkevp5XOqgRBmfQ3cOhTuWPrze1ubqSxFQrF3/RNx6oyGfa1dFHV2z
J2hxY2zvdAP2OjdfV3qfq9Q8JEyqdFrW9+uDR/Dme2bh48DSL28rKrhNx/Ze/UkXAktKRonMO3Cy
GuzyFSUpjyafVjsBOwtYhGs4bb6R7ZcjsTtNGtm3S9rbwb+LGvUb4nC3RnJn59uwA17c08V8zSRY
ZgIt3eolu/C7wBqGGOviSUNFPFrGt2J3avBpxLNR1IkAix2nVuPy4gu4VLQM2fA4WSZazUDU8IJr
RdXu2N3mKQKkR+BNvPc8jq65Cgh5z/qWfx1kGVQkGRa7je46BQ52NHFh9NfMdEaaySzRk0njtvz3
vz6SEZY4hLzlAvLxlVhiIaLttCHratqSiej+1Q6Em29B8aesp89SnN3MeqVEWYZAvjNIsCJijGkJ
+wF4+x8xj5qPKnt5jO761rvxhbYounlMEv2njEDo9L05AEMWCJd313gHoFXsrsgkPrY6IdNveZ0j
onhsY/qJ3suuoXIxafRZXKQZdGFhiKHGveNbpxHOY24jBlCarty3XXukA/2yagODny+YfbXQ7cho
jOMEkllFnTm0E1g5fjuQrRCFYtUyUbprMKOhY5VomC+O/NYDEmjg++D/LxgoUHeOzQJA2QNmY22r
1UDX4Tl2hxZSB0FeNc6SOk+8wIdgqaV8c+vFAhghL2gn7g7smvPAMi27GhnEEu+Hlc4puU7/gU47
/UF2HUGEt6/JpcwjLTH2T1p3pLz6cbERlBYxMqusaJJM/5ptk7zZLKM2P7FAs3kFe7jMtf/n4kA/
bdLgUjG4RyB8tjXy0baE3TC5c2T4/bb5se5zPLhBM681cgqljSDHNNR8SuwNfrFVSijix2wdGLyv
yMwhUkfylnCu3rMZDWURPyCmVakBoE7CQRd42Y38gJv6tGB5sQGIK01L4Xw3QNZ0HizwMG8pR+qM
r1NTa+aKPjjPPimbV7x6BunZQrOOWUdW1vBRVAWCcqBFIHiybQsimaa+Jwzn4C98XqmGmQjaEKm9
Nmxg4VEs9uEPZB7FxhnbpNwjocymret/k4mLZX/XSefQT4ciZ658foaCdZLnGJ/l8TN+CJTUQPUL
kpQNltUhJHlyQ+fmC163OM+I3pgpvGVHovZDR2RAw6f9+IY1Q7qchwodlSnjSz7aLuLz0bPLT2yi
EcUYjR06/IDbrwXEaInTSCn6Hs1pRmK9IHnmxKiaWFH2IpwoMFi0wB+oVmnxRZVtj9c6y0E7qylt
GvnBB5kPtbNsyCh2tfTlxXpChPUCZFnUIm2w6PRVA4Glu1qWwTmbwgViXS6mgAbhSNO1lKz89D+N
yLTFw7S8/u8ezvbxBIc5nSu00NHAtx/+nTkd9u34hqli2quzliacJf8xTgA1ujSb5DdlXq1T83/i
a9kYfGQD32Pcsk8N+sQu23BjPtQENhhwkvy46EQ9rlZV07L1oSQZje/6gkur+4MaMFxmMudajvEK
iPCmDhrf1twzMJoSJ6jgPjEYqVBILEdeUMuH2LK0F0oIEKyvTLMyCLSIVTeI8WyqIpOOxa23n4lV
2EQGBmoREvV8TdUedZ2ELM60HSIr0jlgFXJaD+HfGM5eToOjPq3NmoZamuMVaUHs3kv7tixxbPVi
1CMwZ0LuLCqfwNMrQtkIoYjava1+aq06Rr6sDEufyJ7Ych0N6SSbkIPioGon8UwNO7kqaz2fmaz8
lUrWiJ7dn8MC/buY7y/qUiPUnQ0KBBkLGPJsjTyOB19eNzmNEAQVkgnWkLigyLlfZJQj90NGcp/O
L9hr/ateJl4PAzDOX/zMjBKD6t+/gpc65PUtgJdChTknqpAve319VxZY93twAhw5vHEDrWG7TPa+
URlk+TuEVuN5TZPj3+wA4ztX1lKxGiKg7eKxyGvuX4h76cyRQZPcNWQpI5OCEw25clm8hsYUMVr7
70yPPlCBpKQG7dagjkKFAm/wCkE385rFbJIutWuOpo2h+7pqpkSU2DpovpP9DRPvmqqNoUxmqEBu
w1cEp58nbUad3R+5ZDyiI/euThe6JQ3CyfMYNjvEEyvIHHRHqR8QEwy54i/DSHQtjYNCxdzjGwch
8AVYTF/tpe28NVOMO1fkx2V5RzqHfgIXerHb9CBRA05WUmLx6qNIl3g/kWaUxu+QpCdGD/FCyYIq
jvVn5P6QkWSRgeXOYlVL2+9PVsyxhyOlKqL79GUk98ZsG7afU0wg36Hl9TMkfcvYns34zw4NxNKA
pKiI7JEPn3Hz7YNw1oHEuITKobMX2ESa8ggQp0Y3i5GT9gV6vtdJ84AGYjYGviQ3PzWe7rURVYLL
lp7tc00YdPGITXmxB007yR7tepvTld/S+3IJ3lAGQ4b2G5u6HgbO4OwwqhaO0m8R6CMywhRE++mZ
c5guzNPfzTALrlDjuPtLzuC/kycTwBsmmvuQoiP1dkpyfsPRDkO5ZoGaarIOkJBkV7b/U+UChOp/
+WuQq1t25dppgQzXrIkKMsDzKxLjlBIsEle/yrneKFDdv0tfwK1LtzajLd4usf246Ws5YPVPsudI
wg12wSjCTwY6Q9vCghcCSXhyJakTEH9e2m0MDGJB14e7qcBRVNv19JMGdhPVpbr3ohTOq+eR+IFk
gehStTIJ63+vveUFuL638sCwXiyFL8wgAvRONXFHC6nncwb5/4dN+lO/VqqD9hxo7fhyLJiAeYnO
xqzPy6FD459S4zGLQyClGFeBr7GckmZIPu++CuT++rpse7g3z724kCcyUlSNTVe9jQxuSycGvwOB
OT86YTfGM0VzlZkAxpGrU5T4OZXzVMnG2wD1fsslcx25gzfm8XXNTi/97lwpaWUH05xiinoCTzDp
xuxxtajATFGGvB1M3+JkEiQ/vAvWKU1lfGpFoLnboGGIhW15lrwjucIOc8zEVKXxPDLyPxKpRUH/
Zvax8HSCU9f1MU3YOZhUUb3IlewcSVl6mlB1zj29vV3XUxIxIHggED2/3ROcN9JlRacu69W/wj1/
VtNgN5HMjFk/aMvDDDawUyxhmJjwKbJQLc/9ZdzYRyVx6OEU6Hhn1LG00UsTD05xqPrPoM6GbTvt
dqvIM7A2ZniYSfBDg5Jgdx53UU7nu/pGzREMXlpaYrcaINTps/1BwFXWBkqR4p9tcBoTmfwiPZA7
gY5Xw2oJwZ77/m2Sg++mMz89hBces8tXwpmz+Nql6GRhY3y2cXyVwQyZdhigvvUUSOytFpCkZyf/
pAX0+sHJE8z9422QXNQDN2nUmjjyKHdFeIQUbUEnst3eRUHNTMtuK+FdAx6GJXdgNECP/wmiuGE4
vuIFSctwsY+cUdfRS2X1d82oAik9K2ZwVsbNrQRhObsJBOWswfmTTuq7gXhDlkUSoFsgGzno094p
4SOtM8q0VQCX36hNPgGCWzzWIKzokFk9D43uei2dOxwWkBrJUcEjAfndrDAn+0TnuwqfNCyQ8HZN
GLyPcvVEHJ1RJqg4q6BwpMjd1dbz2t7st8alN0vD0OmoRjLwb1dOyk/ncjpvdDz1nJ7RbIM4JET+
5ewZOmwxgOpzZRFt9+VmFSz+7tVULwLLfsya3RTr55cc1ZelPpCXc/gJPSSY5zmb2RoAFIc8qAYX
Mnc47H4sOtq3YO6dubJfuJ9+U4LDdCMsjqcBcMiDQBrXnuN/sTDQJ5aAzg/wTuHvO1JaWVMMm+1C
L20DIaEEvfmG2kqfPz+hhNecxah1vaQb1cT40dPaSmepXcwkHCG7R0pGRQpXdJuYpRJEPjkJ/NL2
SV9yQkV9LEkQdxL3Wd0sxtAjo1RvVWqGzBALoQZBiUsK59orvVtdEuTkr8NDrFUXcBACOsKRa8vE
BCOO1KEEnTnbNuMHWKP+WVEL3tPQO00/9yhyvOQsh7RnUw5+i4X0sRe2u6Eku/4wSBrInW68tdbX
w+tzGirrvhw+oXOhxB4HqTEBFyjwHhw+ikesg+Wts/Rz03LyCGKtiyKVLJbnCCVUfUyUBhjK0tIZ
FSD7LkK8OHHFPVzM/p7UUE0iTh4hAoeq0l0vthhxUuMsjPXVy5wt0VZceqNtjW4QcjPT21FyjHoy
yBmQsyh+3evJyzoXLrKAxjXTPA+hfdmb885W1MoW1HAZumSE4WuHvqUwwXw2vojdd1eTA3yrnB6K
FxnJv6ptL62C+cUTcaPuvtm7cIq84ro8/I+2m2u+xh+lITUPfBaQgC6jQgR/7RQVD9x/2cUP3msJ
fd3CiMTiYo9upgYekg809jn8JIMLTwQLotHytrS3xsggRutG7/0EbY3N+Stt5escHvy77PKyfUz+
60qhUg8l+D9yuYL5TeGG197c8YxUjH2Set6kVrtMSTyqsC0Lhornia+uk2aL8Gz2x4Qv1BtNvIX/
DUYROKOYkycRg/xGWCcc8wUDjnAJNByJygxNfcGJwqw3FvgKqwhLh4awEpkrFyrgd5R81Yi4QioR
/BpiTDL5/iMeYAf3GEC7ns5/MI73AedqIOZ+RsotmNVcQw+X0VpNyG9kaPns5ckD9QWgjJB3wk5g
Efb7wDNFLe+kIGIoVDlyphKNPqQD2gteNS6ULZKnzzgR4xr8C3Q6HfpnsHDRDGP+87q0zwVrgN7u
mxUqyekpv4ZTwb9VtHSAybnvs61hn9RsxlMJMEVDHmSH8cNTl0bN+ohdrpKUQ2uLOupP2Kn/3Gib
Wx0Z/xBab0JrDpv2I2ntzyX/ui4ioNzkXMUE2i8FWbh7saXGcWlt4E6lkpVF/2yOCF2JCXlNkUAB
QlxytInSlMtztM3YjBnSKo2qt38NqlAZ+YjnMkGMXkwKmsuh4gRoUStafw/jp8qd9GuNsBdLAyHc
XqXX1Kdf2yGKBQRrC2izxFVp41O12kMRXf6tfFyjv0HgmEDYQY+Uv7wBGBIKiuy5bWgmQd1FocDG
Wm8/kA4/nF4l+3TCP86Y3Sxso4FmhA5yTJ4auSgnMZ+KKDK1wQ9vBDlk60/4HORUpPWfihkpxpat
aZ1RceHbfKDmI5+cDI/BnbonM/mLxaNwTgpkYuGXxOfZJ31fN+r3qsTDL6hHfLh5Ah15iI3YznR2
shRY1aELd6cyN7Eo6RCX+I6GoLKE+ASgUSI5a2vgQSuOoJuo5OH7/QdjyWj4nPaUzpCRyDY94uzo
FFjpcwcxlwdcYlMZKPHnCnZ8FmQM+7sp8ypkxbDsZPF9W8uKvQqqukphIbtgqOuOhbuzcfDwmWu4
8HqgrHMhX+xpneCQS1GZobBlokkaJpBYa4M1MFR2C0nyVYlHVZXdIoF+Bp763WRuFLBXmVNT6R8j
n2Yhwb+IRtDP9ccKQJJ9xYVmyIN2x2a0P+yULAhNh7F611MKHNiXiMtleu3mJO4CPqTVHZMhAnIo
lZ/SaVL4oAxkgXNg28X22VcHlrbzcgxcJO70DXj08nQJSJKiPrTjnVZh43YnNrHw52IUYcfm/y9s
HujoCVd8Wq6Ys8WHsyJrb4RBsK1pxc+H1iQt2yL+noMAy8xj2ph5paEMN7baLv08xpWbxIg9Hp3U
gJfJBPic7s8lWU3ME2OAD5FYw4QuV2JBuEjDKSruHFhgk6Js8ac5rGWWXi49X13JnVstPDcg07k7
h4W23KAOFNq0ciTFGkeIcxfWxIwyTcAUb+HKx6Boc/wOFSbHdDJnd/KV5XhEhX8O7e7W32uNJghH
JztovA6lmNSTkp5F5qCTeA4EicJ3BDQKl6LNwAT3+Brbp4ibI55XJlH8BhbRU3uKdWmMDklgv9Sv
QYvnobYO6HvDX4Yd9XFLtzV09jhPJ0/ah/Lcy/PK28xlVXGkQo8lw8Gi57uBvOqe3vqHNz24UpgG
4hL/baskWLN4xa9EU5uMyErm+lLdCQVSfov1K+0Cr1/DsFSrjw8NAvY6IdRvW/6vr8AIY0w2m8Cy
/20HmOGEPIvrKs8HbItf//OLpTO2WYwcNGt9CaT6zcdfgfq04tKf+izei6q0RqAggYzj8zfnKLtZ
tj8ABzFV2VUT3CiVlvMOBs6TiWjmUVMYeULGEJe8Nkatjz6rxvkbxSUcVNq3ZqoLKjLGbqjAUYYf
LilpAeukczXHRB9NmGGc93ueDYR3Xu8YVl4MV6nTDMoDUR9n/nQPcn/C4rTjpUGP4ATHMkY48KtK
RRUDTEhXbTLcgZH5mlxmMUXgVMVpMN+Uxz2LP6LjFHDaD7ovDbugCBlf8eUljTPJp35CAInBxpDu
YTSuBL6e0nFTHUR6mB3Ms0Fpq0BCt88B97vAhRx8VDkYkonRNiNlKzO4V3JTelkQe4pbunBInhMz
lEBUQ8y4tyPmKtVbf+N/HFk+5nD0oKRtu7uduBqTatfDAH9rx/hdL9nt6reTV5DeECLXLLe7Ls7u
4ce1OaHp/QM9t79WXS7pEmarekJnOEuBkDtGL+7gnqba1NA08dlBtA2zPtblrr7y78r+dOpvEqyR
0Sp3YlbG+tx2Q9csCCHJmS5C+ORoUP4u02/+ExpWXzgmUC9Dizc5uGJJ/cEI96G3CFVCj373l3Uj
b4AzI7dFrFEBjGbN79QyiIoZ4JUSqOinl4v422XffuZKCa+A/CqPMtsLAdNYei3YuwURnLQlSszD
M1cAPaE+YqX4gK4DWC2sCXjQTXS/+qx5hl6+I4cE0/jDF88WgdcnS+fKkpACOVXLuHvGo2B/7bDp
dm2v1kvZ2MfU8V3QUsXg+kd7QEOcpohHTZa1JrKi9bSAnSJKaX+kWtyo2or/8nX3gch3g7qIbh8U
n4UCBV6cguwGxlr5BMVBcYXdV/uKsGIFORJrZe4oUU2vqHNDZEA90qdKTOydgu/HO39PKCjquuL7
8sVhSmiZPu85REOGdxEeuZCwASrrkdbQxu8PTy8JE6RVP3VjJLDV4H8sZNStMm/mamklhkKUv2RX
tvAuqnnBPjBGk7tpRnfo3H7Zw9teSNhcaSBSeB475v2PKZosLinQ58skGBFbSWK8hpHXfyQ8xt9h
CFMICcLWNwqXEWYaegUO8r0NpqcJFUaRWP5gX6neSv1T+jOl5Zb3dNcDFKO2PQANxS9z/EYZkPNY
XlKzdUC6weDhDg+u8Ug/KWUm91rmiqjmWH/8LnODCKI6bsvbOa2UHXslhYvJKiIpiXRPa4+HQ2FB
Ymz1Yex46kR8dOpL0GFwS0j3M6Jw/pzPheBZi/b3L5kNJ3QLxmidgPnS3aYM+zLvfNzM8mz6z/BT
xPgz1IZljvu1OAzhMt47X+tbyXd6bceV6pLVTkMCKYw2xyV7zxPJXGNFrAE3VBwTN+EY4JanVkm7
e9RUVcX5XOTIvlMh0g4uLL5EDtZDsZme16SGhDU3jx5nRk5WyDdDVaXFu6sysUykWCgFl8Sy8Pcf
voSKb7EA4JjIVOpmiS6uUZfZ5L2cNUCxJldN3ck+MhWEBtz6T5BfdVdvo0lP4OTp+h/B9pjrocqx
GtSCnORcAMa8goiKYkRQBSZXu8oMXrXW6JQU0ACzVcW6pRrOwgtxbCDcgfWKLjS8gYQ9M29+BqN4
i47tRC8sTGF9l9H0QxIzJ0AvmGTHBWFnRRF/fmkMnFBwhuweREDUGHSkiUn9rRsv+UVVJVknEXGP
f7T30gmPSsdWXJJE0KqwqbNrZPl2z1toTIA10Mg2EWfkMThO5vK6eDIoPYmiqZk/rgamHjEEomJ3
gnPaaasW/cz39zma/GoUJ4DzomUqGRVBbipwiL2wu1I8FRa3U1cLjL16dw6OdkAfDfU+QaI6VInb
Jbu/Um0T79Arfl6sk5IL72StFqJuQhOvrMx5JKDgPkSKmzYzX300XxtHM0stZuJA9MuUm1tbBmRF
32LQwhOhyFFQkkGjYHM1T6K7zu/Z83Ci6m/XCtiqpSwg7blBzD43N1LNT/+vFM4H5kGh/WLoXX9X
wphfdATG1PYsrFGguMcWhexyDva6i0d8D7+N0eavXMPzf14SFNKB3Evo5b32zK9Va/bzYj8fTcVm
LwcPx31LIPrVarcYX5ow5t88KuGkevUOwa10ptT0Dl1nE3zS58n5IGh0SyCHtfB0r+8tPMS76VMX
5Y1IKFFT4ZHvm0uHBjSnXvUBX3E3pKnjgobhUmaScycafta5v92kH3yDXq90lLElR25qzYam1fjY
XJP0o4iS4E2Tro3luIHHwfcKaTF3YcxNI8sCPENsAh1nzfpRHfOzC0/BNGkHU5w2XXDkQgc/nG5n
UHcg5OJTkF7+xeaLJ1XV7wRQNVjvsqSspaAn4EJsGoCKMTOTU8chYNL4ikzKkdD6JnC4HBuMzgrJ
EFGXxKpjed/iMxYa8Dd3NIx29Xf0tGSuSW6Kqy49zdVRuijo4yP7jX2qgKVfdd1fNI0OEEiLlkmz
Qalf6GI6CLukKA5wxiUIU+j3DqqRbr/f1pYUyOIizhZhyjfKymhQeRHpUNEZ9Pl82v3tovdQOKMO
e6AeO/WvKlLNkuAA6H2iUpnvBsfdSpIrKvMv7WpJ9pcewPcCRWBMj33SeLSL0Rq+1HKEaUIBhbqM
FziJWcPETfT69rq7eFBkEER1FCF4SYFoy2h70mZpRG82e9jBjsLHFKQNKtbltMGWdD4Pjc3Uk1sn
RKk8UgTr6YZP/G4qTqroElqzafV5fEsYG5qzXSiWqmYRBjQnUgKmk4+ZW+gqgGTgyAghLq1zcMUl
9Qgc8aUDmmTGU1eJdc/tGQ4K5+JvvU84VkmF2ROwa/EDSEe0SbL7F8lgaTgNKMS2ps9WHrTcK1ZH
skrnXq5+EzWKjjzdQUvjvKTq/9InrXJAv+1Yiqr/0dmjAyKYGnspNkdAsi7W7Tw/qalmxl3Tyn0c
mDjFCYpUI3mNC7tfc+lGZpAnRXd5FEgGjoMlo5UO6oCd3qWSSnSbiESVQgtLmskrwscGQ5jluznJ
AGCmf8RxSdiwrSpACq6KFvMPFfj7iz1XA0WLESXxdYINOsXzF0SqjtjakNbzvpKL/hfPTZiMXFna
2Co0dQM3HOi61jcPZsuzxT75LhwDWIeelxA3flWHIPTZwTayOJ9mDPWFgpfZvGHxSNUU/HQLkUEG
YocKSyFd+M2Kn7AVU+Y2YYqdlhw0eamd2b/xuIm1aAictGuNcCwuF92+r31sdzfWjhQUltedFZY9
wRblo1MLqtT6UotMfMAYFmOMYbrhTSW9ErDnyBX+IWmCgvjXsbWEY5jlUqSqOwcWv9U8MNwIUmsO
BRkja7Z1hP6Lp49oOUTEt0WQjWFWrprFAMu8qwvCkoRoXuE/6YRjX/mzhSWnw0JHYHC1aiCUR5UW
SFNfTRJEDGyKEmrj/2F39v+HIT+xD9I2ufFXFwpB96vqDsAeKWMgbkVErwfZq0slZy2KR4IYG2rG
yrcZa55GcJ82wS+cU9jjeN1LJlAPRVXb2uqXnoIZokyJ9NYtOiO+4hTj4wZCfU17kbZ+QkYIWfDG
9EnYSzigP5xxnVFw6DOTnk+VPJT1PrloRO/L8w5SCn3v84Q59uK+FKri5tqJp95gFzfebzqIPENI
OCFmDEJr4VWk9RJRvuEAEAeX7wrIzm+fr76X/vTjzRcUU4EhGD2r6cTSjqpCAeGwXVcdlsUnlm1q
qAOaGPM1UW3Od5V9ZhFuwa07zB3AM1QIyBVBuEL9B+JsJbt91fLR1XRH0OaBpIL6KN7Rp4H9i99Z
Qa/fG5iMq+1iwAKg4eJUSZPJ4Qp+BZnMDlUcqOaM4tndU1VmSicVupKe0Q5J2UwUd4w6TixIttwd
H9k+WpHABPQUvbmflaFPHBW+JD70HuMyWvfD+E4MObcADMNg/0XbyyJSF/0bEYp3Gs37CBPQzD5U
qMAVX6xAutKgmiAJcFUgyCu4BI+GkG/6KqBoXbKqJ7lATz3+8BA9dFezH6AxCM7NoX9hXYWNwgH7
tMu+EdaNkQmqBKb/kEoyW+SYteaMUeH3G2L65Vl3uKE2QoxppvK78+u67knL8/QhOah4v+mcsH5j
WUUHYg6EgTyIBenmJIwQhsx2buSZPb3B22o0C6JzMvi9En+QaMvQsD2cfwuha4fPcIkPI5MsIIA8
EkWvQ8LOS412YvDbTILVE6jYddQFe8mMZ1Hy8EtDmj8e815KC+FSpi5UEGrFkNnOwl4ptBPPgLgm
7i0yk5pBC6I9vN3+949hZovZ5dN9Nzcc/6GnK720ZuUpgJES8SxSYPnnHdyJP9KDRDIIYcA+zNJG
3VK/wnxE1SskLsUOSA+1dxktBDW3i88VtreCo9OHtKLqftSSleT/HtZ9Tej9b2dO5xQVN0evDHt/
FYvGbp/Q/cLmdfK7aatV3CTnZUXhNud3UlrRwoCMTnfX0X35WIbbZgguD18UBkp5Fg0/+83sZZCW
e5HBllAuzTvDB0V/uMuJgkblVMJZhgDYi1ikUbT8TsGLIJrsKvqQpbRl0+YSEz9qAs/fevYPQZbQ
L7CpM3lsyAvSm3zSVBOPuV+bSONU+hj9gkK2QZi2qTzuvVctjpGemCGIyEsVNTiFPcwL8x53MQkB
l90+/9zU1OytE3PbFC6K1e6cYmUXNktBnRyxlCCDY9sWS/DvjJWveiHO9P7CWshz0Ld/YFmoR/Sq
2T4gbCos2XHFpac2kcFhYXP7JMGfr1VzccEUbO/Def7MWwLPwqhlSuidt0cSwfRZIc2CzDBPfSo8
UQAVJy+lpfzo5vmO6oGpzLWIfRHpVdpgMeTcP7uXr5IE/4SEYSwvOuFmFeNPea+vuOJA/EO2xcyb
r3sk6uiOg1VEBWF07bwatMmxCWHzQmHVm8VuQjSRQDsvbylJaRG5TsEdKPvudkzp6khMj847WY/y
Iw64LV9OEbYTwhfqpHeh6PFv5DyqjcpRrJrbZKM8K53Uq8aNbLWn/w9vBTrKdITH68lIeUbHrDpI
/b9VLfe4a9jPCJzK2vAIjRZo/IOhE/R6rbl9CMYlkcdu9DAAkDISLxOIb4Jiz7Y/VP1eQux/cKRw
jl2Uu+j0SZYfQEwg6lIaulZSZiZN7O/91Ql9x4hYBhB30MEaKyhpgyFiMT4NVCRfm08nKr/F6I5U
BmicLjaT2Se7Rg5eV0FJea8xeEpfc66E6nspo9XYPLDGMcK2FATB/STHC+Jg24wF4TMTF75SeiO1
zuEAmpw6KEADTJ52rB1PHNFC4S6e8nZtcvmliP+OaqnP2nmcUB8ZhE999WZtARAa+O/jPPHXcSL2
bTeaR4OgGJ5BpyNZ2U+SgVwxfyp98HfEhpUvPQ17qVPmNuhB28hKSxCRH4g2BIzziiituDC2wTdH
v9sR/NLGkdgKy27W/8Cvkrd0/8jmk1w6k3Ce30115dhH1o/bYYXGkJFK5FZlzN9d1t1uZFgKhB6u
QM0Ubpa5b0XAEJtuFukogEvkxa5OOyaBmp8E1FgZz1EtamI3wcqOSuy454/UKUL4FHqeuDcU7loE
JjCt4I610XWRxPweMxvePzmqM1O0UvOqndm0I+Ofy8fililaIEcqVsoT3mHTmh3xd+HkcemQ+avX
8+cXHwCbhB1N79XC6vcYbc2YpYNTBxy9nB3ESxW/eMiTSmgNfq5LnxzyHumy4Fjcsb7nkQIYKqZW
rr1+BTabLNfixElC4P+h8GFhZzfnyt3CSihLtNtdCPm6tPnRvGGp8y8xorCTZB1mPU4dnX+NbWOD
4+GS2dQjLNkZsgxy3WRoA7X4aNVsBNAXnY6uH8p7u43/5aOW+/Ps8D/63FLURvHOceObx4LuXykj
tuvgYplgG3LU+ObyFqyeJiIaR2jSR3oxMtkqutmco74csyrlbyE5aNEzbG5rP11B6TQyrfYiwtAE
2Z0sV1F7kX9R300stsLptOvvmp5LixzzwBrItQfROb0DH5Qiissh/BTVGVV/zEEOLhD1chb7tGNt
OYZyIghE+P0je52CmLwfDSdo3WTQiWGmcQ3XuIXdVSRRvQLEmSWb0o80AyYopvdoNTyIPlUFStPG
938Z60dMZjyK9w8RPwKlJ3xvUamFmMohqDhOZQkLyu/sGi7x0eWOZKTQCFh/MHyqGOdtTkGyVB9k
pNqb3WdfTuKx7gSvej/5ImSCGI2ay3UIsuVAyV4EFp5mcVx7tqNodwNS1bkRtpiUr0ABh1z+x4zu
3Jf3YDMP2CiJmc3ar6KALUM//+rBdIHcuNnx3M0yg/qgSCHHW15IlrRL/X6uys+0ROAKxB7tyQ/7
TueQ2bFfPISszXjG4fP5x+uCRUrzewr/mHLGcHHFCrirV29kh++FFCr5TH2fVuevhcphqzIJQK2X
w3JaKDOrqLlUr3fDeanZNFDI+VGTtJVPZD7+MCjOgQA3uyIio32d5U4d9qFRXFnH77Mlq54hAHqO
ZxuF4pUxKbosV4qAai2jDklOWwikgs5Ceo0v+RBxCsldiJ305tjZhfHqdTe4svGFOjxiFjPaA8vd
uNyPVAI08+2WsBazV8GPF8Rg30E2IaLoPvUCfm+3GxaoE3uNlmq1H6/Fu3lkYwv89X47MVawy5io
haWXB/+/SrcmZabHvBsVfK/tUYlHWgWy4yuzMb8O9DhFL16qOvO2MIBrkep21dEzd0FbovZya/qR
oM2lzE7Xh50kNAY8DRG3/LKdJQhosIqdzmw3DPC/GC71LkAQnQpL7YXcMAXK9nkrZEU3EvU7Xdch
V1gmxu5MsHkTvNeQGTpRNQAnMG0xAbo45PAd6imS0D87r3IpTtxwxIijbnXHUZKEtm1v1YdfhesC
bh8FzTn35Y5pHgDOpH3WQpvq7zsOYTng4GurQixAkQbrBjCikrXof2UBMCuWTRJVF3e9eendazAx
t8T5fLYo90onU2wxhpRV0gc7PnEsq8u+XZ8Lc1hk6QJJ3H1dYQctXnu0ZWkrzrmPkvMZOaHvX56Q
hfKOwcxWz07qTEIV7AfXcbIZylx82iyEz9T9YKcHnShB4hFj3UFdb+jbaxVssMPFoo3UxLmLSAi/
JiSzsSJ2q+m33TuMljFGigDiNIda+UO1HfkpK+tocd5ovgfg+cac3AxKEGjOuDQLJEvVL8yIB2bK
A953i2ZNZNLDOvvqDyWFPGP9MbY0fCZOaK/d4qOxPzxFzk+jJoPwYsAST/WvA83R4jXaagq9Ae67
ovP+d/q97bV2rpqunum96rPDByD5sbsUFTkFDa4nx/8h67Z8aOCVKr+QnY7LLLYouDkYg+xVHVHT
9E6NDIrN1Mh9Ybcev0nMwzwm8Gxn41/nKPiIDN5kPpuAS7/mwXmJigS4qy0PAXXfiZIonR3RYjrG
6TaRD4ZuGUs3kvkMs+fw4U3hsfNHR4U1Jl69DgOQEq7SQbYnO8ooTplCZmVdltvW2rQfsdQFRmjH
JB1h1pB/PslFILr1oOEx5o0QaLvCzcxOy+I3CTjEL35aIDiGn9Xvt8kPhuCAV874Ce1DJmjQ3XVO
+MXdXJJZMiYeHgqvw7YSuwV3uDXr3+OpEYjey/SK1r1drvC4J4qFlIg6yudywRuecdOUF1ho4mEG
hH11HJDkHk64XPICQvZwdU09HQ3X/3hGOkjdFBQ5bNZgQZprAbrae6VPJ7fjtfPUqI4nzwmHFLbh
wmvZj8TnHx+En3AQhW3ZIP62gzYlPrzN8emH/byQtVKX3SINj7s49zL4TdyFOg952FnE7oAXhMv7
971gKJ3hZACyQvzR7VIqMHAleq2UGcWmwxllGBTcxUfM0kMiNcJ6O0ZsqAbTLLAsLdB3tAoUrLVx
2CebHh2d62uPZcZhgG8zXJSK8GLHbBTHr4tiB6NJ4rQxwKJuxPqXdgt+AIP/b6FdVJp1P//sy6ZH
hvt3R/iSoMDs1FCkIcPS84V6IhC5X02gk1Gzj3xDy+I8KP1XirAC8sCnAkHr7KN7cJmqxpcU6fm5
gmCzLMrgV1xqUxdexHgy3g0Cf4COG3Ut8T+ml9ndMnG3tSZGZHmJX/BmM/05IeB3+0+XtllsFF3l
jwK1Z3364udweZGkgGzQTXqUQMwXC/35bh0PJ4azbgVDfEMIbPQoPsGXgUmgH7L8U7s3OQ5TNaVS
zY6kmbIEMUmaOc36dGGaq6x/s+yHdr1riXgymY/iUlNKpp90LuLwc0SIM6cwsY1XFeTXV19Plh1g
sTG8GVsKg1BCOEtcLl0/QQSJI57vPJfAU44xoW3D5yFsKeYWQiHky0BtnAJA2MuDHlfR8o3FQ/KN
sad4Zq6N3Obak1zXNIQ0abcKOa2j36GK5OL+AEdIffs/519dJWLwMmKaEIMiuzChg47GY/ZZxjmz
n1MumNjLEWndhBsUuNa20ox2aCx1bYoAgNCyjewsu/ehYJE0Nq+2bDZGImKKGEbLLatHu6ciIbGl
dTddcTfSTEOk/GNCJzXtxYbNb87a26WtNXWZ8AQt6KxyGnC589sjQhfHuM+M6igzeYPA/2U2IokU
0uNKrRn9FlN7d5JL7X8gHzNJcvXBBm6BKC68CCWMbZLGi3lpjl1GD+MqX/fb2ZlaxgHjK6iqQsx7
9TW4fIA1FVq3eUKHemD+BcLjiKfhD1OnRTp1GUEsqyKpUGayGbIerswNc6NHn98G5/qHG7ltjhpW
SCbWM8VJR4A5AFq2lMjEk1vaW8//IdO8F4vb3XmvEB/a2bF52MRgNwX5Q4HJy3FLyVaYNgzkpzoi
WjabIH2NaR9qPN70543HLTTc9RtEi4Nwaa2Ubc6ehp4kW+cERU8vwvfSrC8HAqHpo/+MMb8b9VfQ
/4HwYQvjk62nz9f+3e9eqivFcJaOkU/rPlBPbk0mUNsoZRV43KkvtgjOJkmEKfCA43GBD9Sl9Jjl
8+pMvtoLjxzGrvGRDAi3ojsUa2oVBrndPKbJcHO6hOSwnf36gKEk40FwwHX3uKcaHcl9AB75csiZ
ygHrPWDFUkszlG+fwVV2WfIQ9hzusovu1KLN4pPs4qGsaUT8OYbUBPnKAbwJu41rIvhlLkcedzkm
aQnAs6XkvuyCmv+ITk4AXv1cWQTzh5D8TGa5OAghSBdyJ1qgX0A9OPXwG5Nm3zAFUiTlrhyG3ZK6
9seiWLWOL3vii0hSpCE56ZmGlPyLuWSoY8CrCDiWTx+5rRWkFveJr+5XfAs8OeTG7w+39SdH0zVk
Ww+YlbEi1BYrrLRN4Mojy5M+tZPuo+lnSQHRuROQm2EvqCQQ5AmQY2s5AoT9zoFz1EEilv+E6gSz
GiX6vU+mV7GiQbgu/WOH6gUJO7NEyd4byjj2+a2pE69ngiAVhVqUJIlnNp6kgcQ62KwGPSgeX8gn
wFdgNu1T9oReFubC3cHnOfDVGanP5dkUbr33eIU1XHMSsgOmGap4/17S4HSO4BcQUDYUAL28DjOP
FbVt8wjWMtYGd0MIIfkZ/zx0otqiCWepAjAuZCOKQX2Ixs+sNVuPNLD3YwCCDlxhS3NP37rbbN/q
ovyAlc6TNm6FNgKCgShZ9uF6n3hQ1FnotQRsElOgJzZ0IsImor+gD2/NLgzqqEMq4/q05Mq4x22q
GCfZ7lVfeQp4/eV5MD4PDmRpNsb8COqQmjbEgHwfsc0W0CEGBkZ/hptjRAb87d52EBR5rD3eDczZ
qzI8//aSyzFlh9G34bJ+URndCiXyQxebh7qDCE0B6dNZ2GvDRpnH68ndWFKzKV/uOX9WpPYC/qLc
SV/Lnb43BMMqSbtwiVtm5MZYCBXAIrIeWxY2CNqoK1e0HCHhxLWigOORNwIA12nF9Y6W9C2EttcB
++fREtv/ly8Vi8STAJ7mHPicjhcxJ3dBNvd+07rpk+7hcKaNpNzYmUb7WkoEIYcxUZ5x2xCaQ1gV
pfmDaaWLc8IsTfKaqg9wjO/CpiP5JBjpJvk0ADRC1rlb5hJRxxQjaJD5euPGoCEravqOOnAxHeWK
CQFcPoQ2yDe1sIwzAU6Y+zFD/YvOunXeTv4j5unG7bCgOOJwMdNgv30oiouTAxDWSniORzYTS0Sc
mag+XPj7Tqu51JtJRVyyaPzTvurWThMqUQ4RQlTNOh+lQvBlT+PnXuNionOzwj7szi9Gu4ZuqdqD
aaVXo5wg1mcJSR1o1yCIVJRfvMhm+pOVLi7nlyajs0NIZmaY3jIWUlVkeoZ/7XSYu1td8+iQ64ke
AYToePuNlhC9peqqPGxz3+wsJdmMZ6XmCbOiA830LgjNhnk7EzC/dF0CGugwdVtch3uD2akEiG90
lOl1QQEgAcp5lw/ZzUR6Jtu3mC9d6d50avic26ZTCfCtais//H/trza+WwJt2kZFO43eiRjoNFb1
9oa8wsr8dLgWon+KTFmU1bFEUwHeoLXbL1dRWIPDNs5KndFVCvDHSKIkW3g/nHQbTpDp0g3FwHIh
BUesAa8XletKv3rrWSVNPTo6AGyoEUV1a1LOH6BFL/rseezwUMDHV3/BQZPXGH/ZMeBDIeqeXFCF
B5yXhdZQvp1TQ6hk9Jh8/YbNNZVi6+eqjIDdtmGWZKe/bP6iNLTL0nX57cj+SAHKqw76uGztAJKg
78Y/6LBUENiesBnKCFei1RJw63vZ0jd7Ra8mV9stdLaLD/eNOr7x/IvPMAAorUJIF3XW92DD2Gfb
lA1eY3FFypYvdrVx3s/mVlHRJ5BJZS5FBTJKIwrnt2EwmCASJeXWxTT+S7N1vcl6intNqgvMAXeU
It1UJPN+ESjY68081QqgZVIMIWCW1LDSiM47FleVsCT/FNvYy2KO4XPDjBtbC/xt07i6Yp4I47Zy
T78yi7ZO3f5/CNz7s9WAi9UXy2uRFmipQe2gc9GiRRWwFF7MEvgFy/S7KI1F7AXDGPkPy0gUSJtL
RcTPU4jtRDrxqb9PWcsdgL2FC1zJ97zL350mq6nXOyMAoTeriIKU8+G7ZsqqEPxVV6MRE793MKc5
/EgTSo7bLr+K9krn7gj6NtNY+YhQkK93EobQfoH9q0W3mPFprl8qRj+ldU3oVTBxmKArAh4CgszH
nIqJ3U9yODM1GHmB2Tyb65QROLUCTJ9wSMunIznyJl6kKFz8qtnYUnroQ4b+6gfit8LtJzHEp+O9
LRoHb2BFDpSVwQwLVCLsE8vyqrcdTAcj+DJHHKYgbtM3al0jXloNpv3H+bObUPIVCx18pIozGppj
apC7gSFpVLKGjf0R5w3l50uI49LByjHMJKha5J7bcpcnOab2io05ez0lS0LqSTl0bQVgFJdnDqXq
Kmko1Ygv3idOqq0T2A1YBF2FhH0rvzC8fVEBPZbnueWmrNq9wMwwoO/czVRNh3y4S8nDuapE5Nme
qLODoH1kp34QpUWfq0AU2vHaUrXk+lKcYdD7JKQtLuigrPW1RQi24QNxkfaIlebkNz65VfWEc20y
OKdAWr5RTmFV+nuhrhlBc+zxeQ+2+rUl0MT2gycW1Et55lEEtowWKCQgBfrQGKxCYTvAASaUsJ3U
dq79Qow5/+ZPtvvhr+kv3PZjdQyIl/UBIvnuLA/gkHgxtGr/XgQbPnIOXORGUyRUnU2/xEbUB7Dp
Q3eYDxyNo33Lb3JLdXsuGjlBLcsbIqK46rk2tJcgLzlSHzpJFEVKzcbcvWTZg+lv3c497xey+jWJ
x228Mp29kkWeYL4jvU8mYn4LFZIqzFg93goOmFA53MVkdYSKfAKU+quR9D8qIOA2M253+TbYDNyW
jDCkNZXkwEN2eYUhlbGvMAbS6iGgldFgIb7oK2fg41qDbX4Nfq7vL4T0CZsleiYONYp6h05SoI4i
iuEigN3vNIFVJEb0yC6C90ZeQby4zyLv4oFKcavKEB7n+Q6hk3HwMpKS1TuyeemptQxGkEdbmPxg
bvostPAqUhN6H33teXFzTYda13nhXcpPCnAL1x3eEHnfx7z3P0M7Dbmi68Va+wMhb4YirJE2cz/D
Z8kILYohC8srJdNxI7DnuEsLvmAkvbNePgJ7xxAH5D0IcksI8HcqtO3f5nitr3sfS+KpoBd8MjKj
IScs5B0tJTgeBwKCsyWwWh0ramt4cTNKuZKRAmAOkOcCLYyt2QEaBL9rE3RlSViq2RcDo94zrMvi
43ZZlgvC1MvJfJKF93FYBQwEeSBvHEz0CIjIAtKIOfb8jKo4uHjYDBMakcpWq9jBoncH9XjuJutW
95io2+2nfgMJtxjWeT7JuHlzPXs2QfMaKLp4giHQ8gn1NNgvbGzD7UCqBgaCDTrRouLKhTWdunsP
r94DO/M9yq4rXdFNJhD/GTJ2J5VTYWeo4HmA9HALeFnJkBTC0xChnEC+vfKsMlt86BmroR5buV18
Vl37xd+VfJzhtCY7Trv05HbWx56SfbsBYtV8pwPlm5vJC55XbNGf1CjIfvZRJRZ1kS+nlEPyA7aH
bx1mWh+2ZvTU/Mbb/T6KJ2V4DkNkcL1sImp/QOk96x1TMV1bmBvN74XWm27dgq+vNpPSIcjguaJY
dCUVcYXVmdmeSyaCkshR7c9QeFH6RArAwaXsDH2/SnhW48EIHf6jN/JKdkyEPAy5JcVKHCE1X1Vo
ckV+NP80wcUspjHgy2Qfx7HwxJhsrnx+tFEXSVTyJkr2cpvgfCVLbf+zvRhX8G+Pl4IIEGDPWFtc
2ExXr8Uap0XvQWy/ZI1mlUq+alWgxtG46UL8UMKewx3IXzKPGtVSFGECj7TUmDxGBU8zcpt/zQxx
NzJY8xA5wQfmKal8vijFqt5ylULFLKybHYuUb0uQkuwGGX5e1V0tRZgJIpazAnVa85uDlFtuQaQZ
5ApxsxUz6JIdbXP/b18RGNRffxE9pz1ewm3X3BLlJrmTTaUUh4tBJjU9twc7syg2qP1EvMpmWJ4Z
lLcJHPhJk2Fuu5J8IJWsoT/mViUxvPgmYv5h+ozcCnIahgJiNhDIu3QPi7pIDfSISYBWyvWx9c3Y
U0761Sjr1h4qKpmIBLeQJshTUkYZ3UA9FhpZI8/5J7mi8HeB2ZtD439lDekRaVDA4M5vqsz3otzP
EmGMTsVSrUgc6Zy1lg+QPYMyEAJKBpk+6lhUMgCMT1GniVg7HeskfsVqjZQVS0tOYZGWUVfLHPhW
U3YSu6QW6zyUZM8zeuZZLoGZitBczUBQPENWFPGb9yJhwNZVjf23hfo6tL3xiPZhxbklBn9DokVi
7jcAYXvZ8jdk1rpcuWi+lYzylzhXCCw/8EMPR+TUjpsP3tgWykfWw84zN05IySDQHy9WfKJuy77U
3onY070mEIOBPNRyuq127CnBnVvQAatOdJPjoHuwE8FEnI2/QH5y2U7SNrdMFe26v5UPiW44Fp9c
9L02abb47C/rE1F4NQzyLeIR2Myt3M4C5GVXRw1vRfaTd0H2dP9bgy77sUCVV1dQtGkGFW5uQfiM
YiGjnriL3au/C6bRFvmdnkfh6YXAFxOoJBd1p7+Sg6EADs36MRLD8qtwyfTf5kUNSXOZ1EOOLTw/
Dij/Hl6kfH20Qk2cYDD42NkyrQFQJsrdUhdp6yBv3B6lbFXtCZdvn2AmiIxOAL6kPUcTHkHTutmK
brFyYfSD14tm+tmoRFtNseh5eIENyqay91kD4+W4ykRcaCjGehN5udMYLgBIaCCIk+5EHEKrR0eY
aBi4fK/LZCIMNTfj+6EC6h831hjTreEdZk0kTePnDskRtAsr/n4+m1hd0ro1ringow1uaWTKglRt
HEYJ3vYpX75lI03rzVz8a1hQpdwIkShqnW5teJu7RVqul9+tCYXlJbV+1qt4ngRcPA20xvbbyz92
ApAxo2YcSa1kCEXIRIu5mtZ33dYSareH2dZya/7KfUUL/NbEl102mNamq8fyE4g9NqjEJF9C0kRZ
1qVt0UHLpeltcBuJiptsGMuTDrPDyJIui/XjP8O0hW4/UsZbhy70ihikMFw9G55tlTli/p9RHenZ
exCKJq+CY+uxLi7KoYWll3AFHXxRsLpu1j5kmTe/dCnrwMKqW5LA5l/oDygqMyVSSiVTQEVdDDfz
NYjsFxhi7MnZ5G8wcJ6wLS1W0kYuiLGsctB1woa7MsiuqyDg7g+gBHOlOO4Oy2c2EGJcDGbnILk1
p0CbiAFmbqT00E1VETTKb6rs8EvhI0a8aQDeZYTKFt0ibkGcV/JWNQ2KXq/LfNJveuuwWf4Wclp/
3Lc6oum3yDGCbCeAsti2pkfqkLdjmI4KqQvnQD7LxtGKBgBHKbQoIFLLgqlhPKIyKRQrPXnFC23E
tBHnt4HKnnbdlJlFsDI28A2P/3lefiIzvXExekVzFhMbrcgjbU3uwGzJU+Myso12k2tKnD8D5EBM
dphc7ne6hCo5+r+58GFA22johyxtnyar01jCmelR1wGffB/AtAMtbwOaIsm/6D6gUrF/jpj6LJ8p
iY8AHL5KjPAlDDNgJ4jPb1w6CJKIPFdzgdc3Z9LnF3P/cHcbPVkR3ZaNwB1bKYTVLoII6n2z8YH+
JTd+EsAidX39PhYADl/pwQwxv6c+biPEPO1QsZXFbd4i51lm2Pfyt8BTMBWqyNn8pJ5C/0Rdl0pl
EUghhxNN2imgynIfmRCnmXM7OI1Lxkfy5ltzRJE9bQrEzH3vwOlSZgaduu7Cao1xU4vMJIAobu3d
V0JjCSWt4o8OAt5CrJv0JpRI3GBNw2RDdjAV44q6BSTOl7lNpdzn3QYyw+RQ728SwBkHenEUnJdx
`protect end_protected
