`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kMVQtO40WFFWwORqlrzHTh9jiT7vIuTxrisJkQCigS0RmImuWR4uL7ruq3Pcd4oWBXvBaDegREIz
CDN3u1VdYg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XcBW2n6WkrqVHKuSKm0k8FVXodvyuUkn/4h71DtxO079yveyFowRmGJJAvA9E3klwlct+mOIaBlx
Rl0gRiYT9ci3386lPMo2fzTJiwqmrLncCyuX63xykg8r8DptWrG3HTpGNUrbiF/aMbKfwkDl245e
tzjapboWzaaI/Eolkgw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRJgR36bUbiZ4TJSbWLudf9pl3vHpvdvi5taiF3xEM3ZRgb6HmgNjhssZFvcgNOA9ZtN8qcmNNS3
wIdryjdhnx4O/SYlTrUF+mCWXVe4rye0kpPM0Ypor5M4x2p9ejTCj4GBIlID9Juc4DctX+7MlVXb
J7ejoQkgh21q5p75O9slXaM7xm+LKLvE87fY7z6GJt64lkt2HqydeV3eleOwSpA0cLaa8bRNu4VH
06vJI2L5Y6I46Jjo/EOP3ipLbyWsemPg/m10phoRrGRjTSLKkOUe2YcNPLx7hHGQ+obc5ncu1IhJ
u2yPxSqD4BhC1xI2Qd7bXOy854xMHAkuAe/44g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4UinzjZfrH8KFllFmZNlujUFJ6JXwKqaqM+vTBPTs7BLruyOm+DV7FTDvQXz9Wfu12XXbAMJjNLF
EpaecpifYuPwikapTc48I/8WE17QGNCy4jsouID1rkfOFZbhl40q29+YDIn9Vif1mY+i7iUV20vL
AOUqn/t3PZtSzt8pzJE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NIhHUz9KmdaeYt1hgT5ZM6XWOyH774b44B67T5S22/6UouVLl3hW4iZRVbRzFV6rpQIU59zQqbue
EyHha6jXEdTgFYsN/j3El1YCLBtiFmtZZJQErvK4EJQ1gp+G2ErcRUcN7mpvuoFpQMPRd+ADZRHy
6gjhZJtwSWg+/eNBKb355DhfPT7RSFe4IVELl+8vPnvKM4vsBlkLnTX1EjlW3J+dZAHQDXoWx59y
66j819Q63IqSw/rwC47m7zdCypmKqb9eG96RCd5Hy9q124ScExuLQjTE3q/257lkgvw4LTwLXL7V
sONL28EhwXt8i/Wa1183oZ3Ln58ghMJRZsmjbQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16496)
`protect data_block
Uwamr3VNdfbdv30AF6flOKGKmP9TXILl7Qs/mSIQ8MqzSXAlnl7paOXcZOTniVRBNuXzGuIHAToy
jWwhMWhwbBCbZoYyHJE055rYxACqXiFGVEQq4IwG2W6zGKBStAjdxBS7O3oDVd/rj34qOh6WJ/hO
JPnRm7oV2K0fkZbHgfqxWdlaWXTjZluF3qJ10KRfCLw8F6UmLPV5Sl8IlXnb8GrdegBD1UhOfTvQ
UYHHkMXTj635iKxcH6kQh/aYi193cXKfzB0xUVWGP43gxaAP2xPY6dDAF9t+IeDRsdDCckuw0HsE
nVmobVG2lSpQrWTY9wZb90h79IDPVMciFMeRRGgLCJKz+hN7HNatKDrD1XmQAhe49KYaEBp7knTR
MtrxriThIwORmliBdeo4HZetzXB/GjOljxzrdoRbwFSuECPAxOqmFuJLcrzKHHWj+4g8FeV9/h9N
SClmoUts8WHb19sKMM5ZSt1+C3upEnyEg+ER+y6P5u9x8aETtR6hHWsXoqYof/GSQ/MKYOk65k1w
iAWgLEz5W1mKX4U4oyRt20dR5YWRepc6/NYUqgy0B79sTw8QNQL05phzh7dRBw9Jm4wfZkzgqfi6
Ads+krh7UDqgvLCmW5qg0Ah35jz7kWQUr8PahiH9VQ4VKJToeVeTiNHCiMrEi5EtdFlV08zNABEK
pUgDu83qUH6TBiUBXxmR1q2NKSzkx07TMXvTZdKKPR7Pl9wa7w4m1UHKjjFsmMJScm5i8+IYKunI
uKKKMT7zEgmQXz+yTg4uPNfovrW0RermDWGftjfsvbOBAhvhkISOmIfEX73ostC5Xx7PrnJfzLhZ
U45+NqI4Pmt7fP+ud5owOBB4e0Szy3emoMWj1UCdgqxKXgp1AkyN9ip/FhJbiuenT6sw4PqLPob/
RTBeWI+ai7HFrz7/1f+ytn8TAOilSyZJURPcYv/UUINGC/nrJW+Mlq8mQbz0ufhgChWrR/SVJmJP
rFnTU21yFoVNmhgRgdGN3jRW37fYJSZRQQ7lG+zT1Xm2w5Evci99F76UFTiMOm/RUnD/l2bbG/dm
b7dAEncDwWEvXwCn5xS18E0vFrrFHwbk43ZN6FKs21bDBZxmHQhLXBrZ0Xp4b1dM37bVj+t5sghs
NM/tiiydwwN7yVj5q8JsYXahVxzZiqfrVIfhv9xm5jjz7Lsi9BNZ87SBefjOkSuAtUWBq6/C45rA
t/UkcpcmJs5T9v6N+mVcaOBwJ7hN01+yeQoYCgvc+9q8s5QVPAS3/wgHQXY9ywrAZM44tmsfjnWm
j9+ldWathwK92QmtGrue5sC6bl359bN4n73DmYPovxhz8n59YSV89p/iMwynCGpzzbDbnN4Z7omP
NAoghH2m5oix3zI4D52K0SO2B3Ggh97v8Spx8C/LIvSGIn8WuZ0mdbvEyp74qVLwbqcKQ9ACEyVK
70bbELxcUco2xcBAYqF4nUmYowfhyjhLUr0qEyi+lThkb6yttwb4IJDBdcF+Xj2HgtNf62EQG7oD
QEd3IZAOqZxnP23XFGxoI5Q649pAaFHtKvUzcSq+E/TBKoQs5EoryaLdqN1srB5DBg3M0fP30gPq
WYAMeiqC2t18O3dOOpIdFH6YkV8JTrdkECg3pIg85g6Nl8RWCIgq2PJ8EdWbdotXHQhcokAXdgo0
nBqRo0t5gNXv8Su7WySNcvwDjpNpOOiAuVanzydSnOdVMaXb9hAPjXuo9J0ar8SpU4qOCVXfQNEd
Fq579m+AomtD6GJFBGItOlos9FwyTbVSaBQSdYbfoaJFvNPUdz6fScnw52Gi5SqV4IeCS836r89M
Rc2qVBatgl+nMoymMeojb8nHThoXO71paYJ3jPjSBBqEpv0r0P1VKAThdYYKIL6GVGa3Z45y9CfA
LbYH/TuDaQRv+GDXMxF2Tikh85Vu+iIVhcFS7RzBB0ZL/0arWHhZ9SpbpbRwvp7aO4HVCLhJw6hV
/5avQJKmF19pcr04wU3H1VcmV8akoKCujqF7AxjZr7v0YTH0KZYdNiie7qhdIZypviHh4tEW6gVC
1MsFm3r3eS5trhznLVa5rCEVBDwt/hUD122WiDTL0yU+mx24nJR/tnZfieqXIPHYbnzgc4ZXmR8r
OxsCKs16Nt1LvdVnHIhf3LtvpnHAhoHC0ddoQX8fm9QwGwtk4ghir+M2CNR0pwN8lnmGW+dG0h1I
dyFMUDsSuj6RrtOEU81NZwTnFE7OuIuxHRmjArXYWB5hSTxTAbyAZOijaFIF7CIRt6VFJJB+DKAe
+7d/2dfMmbUd/CneX8huA5eeXOuDgDPa3aLAXp6L3rKLHiRvOtJw1ovtjkgHe3U9k1WMC6qloZWm
8Fu5c4mrqf10GfxT5BE1dPpqd/2XLQ+ctAhvZ3Nn04cI0GJ/0SYmISjASEwtu+ADPz5EdyYCFhh4
lee0M/EaDAEhWM8RaHRWLMlhFbKB2jjH3+QT/mdDLlOy0Mjf+iy9W31K7GVTaXUXm2iN0IEjs3aa
i1xeUnPJ/qmYc3xEvN+Ng+TbvOnMwwaANelfau05S363nNano3fXCKVjxWcyjCLjamKSl0TKZXAi
ya7YTgM+6Y1Ykf1GBLTSwC/AWOhYpIpTwWGqlmfSz5xpDYq0/fUm3Cr7iV6WsndE3d1Iou56oVTa
4kS8uDUm5K0ZII2/wi7rXrn5t7/DiwoAoliXMcsqlyCPDH/GBQjsogmulUabSPjuLxae6yJFuzPU
2gWKaqyXuXGUIHKD9yf7n6mlWirgj0upiEfnDCUWMxUylEKNJXUwA7ZRP9Qzqb3HE7P/x4aeo/gO
KoEap9VtAWq8XB1D5D/EbU50qZSGi5hPqXDQiyQjhgklHj8tJ/jXEBl3gUzA7uwJ3dN+IyZCvs8K
d1/d2UMlHlYIurOp9z51uUYe0d+m0yXiUo3QVDeR3ez/FEuJuTwvYwrin9R26VwYwI7kt1NF8XNM
67TsFRopWBJrwe4kG//aOuWl7BhDDpxa3IyrjrwodUakgChhIi3gstt3UtPz2vqVcrQld7iuvnsb
eUhAbdKbtsTfuK82py3xHqQMnJclnOvdxfP8EYe8lbA5nVeCt9YaDFzg5BzGqXcSeJYRLDtV3oYA
Tkx5s5/eXD1T6R/lCIEhIlxN0+lNg/5Wf1MVPJ/rzPMN/1ZyqOHZJ6XSBIXlWTnmvY+XwNhJzi9V
ulByEy/PNQ6W4HT1P4qUYU96G1gzZWOUFo9IpY00FdDlGz2r514NGOQhQgayxQYdQmNCX9uB6s9R
gbUWGAIhhbIqfxirM9EgUy02aZCRzeMGdJPIh9tBGUFEeX5D/sUOZaxEZ5OqDeZbo+0/FAPlkdAy
iQ8R84c3Oz4V1m4y7Szr/u9GgjKlLtjnIX2L4yDMxTiLpOgspgk7B2607uOk30wJeIBbUJf0qkRd
f7+E42hMsktZTJKgPrUitSF2pf/0GG3mvQxaWufvgKYKjpz0P2o+FMKN+6yj2k4Ocm4nNoOa7aam
UJ6wWXrk0Q0Opax5T726IAkwQROeRh7EOVhq8CujTRP9f9JajCMA+dXCk6qcq8vHQuq/mm8cCiof
NH7gW8ObDkXBSJHmhft5PIAvBR16NzCDf7qn77tMcp6KQ02n5A34pmbB7kk5T0tlcZaT8fuimY/b
+js5nAXlbTZtj2vXEKw3eJ86QS/4f8SawdXqBQCLtWc1GqLRRObxTZpKc4Aq12g3aONbSy40MjPb
98tOFXM+g1z/uvV/11+oqvvCOEDqlH53iB0LMzlF/sZm5g4mbP0NzzPNRJECom0paRc96ZH3kdEr
ZrcA07D4DnAm1i8NYGWZOfte0Hc/Sn6FZYBqVc625DQx+kX6oL5ZoGa3XZp6wsQInUoh0Gvns5P2
ZqXd4J8me4c/gH9XUPmXunayZI3qd2j2baoz8RUhc4WdVf+TVt8I/73jt7/ltcOJ1J0tK0S4gKHK
PUK/pJGT7FdaB8bAp3VbJzmAtfGSV+r9EDuZVj27jg3894hFXMJjchtyBYzsmlgJDSlLzjtDCoHV
QT6XuKkv9kFdbcbFTF1AfCE6UmMY6ejed7gXFGLVK3NuiOS0XYBCaFKeIpc54IktPxUETX3r8ebf
GulLXga0Itsw56g7hveFdvyZWjj2Adn0lC5nXB/hp8bUfEsc3nFcomkhzZkkQ74HrssWKeThxB0B
4up7GpEXGMNE24b29NQAhPV2VGz9H7DhVx9oghYe7Je4i3WiDhUpSFs4MStM3SlzLUERI3/O+5dt
iHwij4xFL6QzWEfPf6MOvhOi04otFvL8EvvZQ1+mYztdLUcp+YRqdJu8ytcFhLtSVgQKIqClfKXA
xuTtr9hFrhUbtiSBBxx03upl7f54dppkVZk0DKtpxCsn+OYbIhJdxwxA1FN2/Hv62CRUq39CCFWB
kOIqG2qV9VVzWcftbPlweS9nyUdoC/UDUQM+Ei7Zq5o+XuINNV8qryxt5ip1MMUv14wVfmZOA1I1
RVjmwIbuVYVHspbipaZ5CY7wm64EiRIF5vGCxrX/i3QqRgQdvoxcojpD+uO8I0nla2RCN2QTsK4o
NvSJqYbWqYRJxeCa1xA8vYevakA6KlT569am5OTUYTFJsbazk3Q5/lu0dpGuP/mHoyZJBBAWSLS2
dbX/BAafGOa/N5G2d4DPOgmZBAmz4jaxtu64HzmH7ity0OqMXWImqHm9q1VvMr51CuEj6rBXPX8o
yC8jVvG0hiNKamRhTT/Lle+pRrdtPCaIi6Dslt3HBXB8PCvjAStAyjAJ8+8SV+eH30QaoYd7AhWB
uICoGPd1d8awHcNDR9OppW1bsl1HcbAeveKFlyJMNLXyStWr/JlIvEiEzi9ayLzrU0uYyk0ZMHf+
c6kuEWXzSHiNwAosCXKFPtcnRoR6V2osMEs/RRNwTOaJJwwcv7uz0cusHiHd+lLOppnNlnsvuSp3
ZXpkLnNYDK838PC/L7OdfOhnVVp86MkDZTlP43Tl/fpMDTI4XtPDvpcEbJxfcRVRnDnzmuljdFz6
VbzttvYHWqmDj+Ji6Ku7dLmJZ7h9H7mcPpAkpa55BRDO4cYnxcaLL1VnSfdKUPAs9sy66UkytR2t
pXZz/AdH/ThwHodnu7Uedwd5DvMA7Go9lJ0DhN/+55agdkcUKaN9iKQBtiNUy/Z1NuUgqFuREGNU
7cTnNBpuRWT5mwVYKEjwYm3OTX2YK1jxHzlf+zkcV1a/hCSvaUAZGZnrGjcJ9IPt1EHIvpMDHQ+J
lLEqDcC9+ue0S2WdP7hEKOeOZSoTDlfMxs5MomAedM9v8qTVYwoScHApz77v+zw9kSoTCq9+Nnje
vRk8Nvv0RoaWFT1G3tkiGbsJpDzjPnCtuWoVO72Oys9HTgZ1sI01fg0dT7GAuP6wFaNOUVBbOPN+
QPN8/8BrUekwPG3WUUYnHm6A2+4gn3tBxXkUl1kBZxp3z2gzm7ddvAHsbi/5tLsiw6brCsNe5CZa
+N9uaNqFoHVFMajtI4D5Yc5RCBOKwxdgQ9FJ6mGXZWgkP2zgbgSJWBXJDbapB0ktrggpOt+oD7Gz
ekT3BEhC8OTD11YSRgonAWrLVtvB8iQ/CDrI7EknzR8cguD7g+8I4dNz6+qmNv+EcW2LUWsC0gVE
gQOcwhH6+hdE6JKIabhtBqhwmrkmPtS2fhHmWXEyctBjuoRd3/5iZkq1OoQ3aRT17LduFrFMyokC
z11fzUgtcTaOJJe1B3ij2ovYMY5iAUP1NGSncPOOvAqt1wMUtrgsA46Q5V/IKoRixkd73F01yLwT
pN8j4VtRIoH/cOmDyqoAmWC2lV0m20iluREASAVFYjsZ3NWFhNWvgj8hRMk3KKY3D+F8c1Hn1+kW
4xVPeLRFY02NO+6zel+wObwGFzSiua9vUKtlOgyNMm0EIzUmOuke2UEyO0dpKAgirdshrg8GTx8G
W3ROn0oDZ9dh6lM3nH2M2K0BoyFW4DXzOcOUBk/EdsrYFaLodeF2Ozdu3hMi/AvTkMvovyl2//zJ
RPJxg7RbGnK7bH+GWUsxDPd6iajQzhgARS+GahtaFWbod1VdopfvMYEenuaaA9CDgy/1u2TZl6WW
3jX96m0LcAEIKms4WfmZ6XZ3TbGQtw34qK1rKqfg9BPJAOoZI6TqNVLnLLOZiI0dijQ8zlm89n88
mdqJNG/BVqG6OTFWDYX08j8NIEu55Pt384mJr874EOaqv1wv+oHJSKOXeZgc0nUganEmqBscpdNR
vW0CxXbHQ9tjnaY9znddDD5WodVdyiu9LQydHk+pn9v6OUPuFJinHmiSGlOrSFGSm/04rN+5WCFC
57WWozdu3KXw8gbYJuvMDf0gqH9SZLuoRqTxNEaVwIfu6SZup1MbJnJrGufE6L5r4f4zWlOFWl7p
K4pv96NrcTYDN80jilv+cfvzpf01LHbh0ND+zAI6jP4+IWm5ZQkAEvg0cNCwBMwERo3uINYxph5r
RqC/DUE0Q4CUDRHQo46xIk1CJbbMf0PmU/o0NI2sncFI19LpjLOfkujevCliu8BC71nGL+i5nD2o
Y2YBahNAy+GVuKUDYQqq0XaNe6i0ksgZCLLYOVW6Xf7NSQ+IF0rkbuVOxY1Jlf8uyK80pYzgVBE1
ccj5KgqQicRgJUuCAANPDD7fYNb3p5F5EfY2fi+UIl4h91eclVrFyHzJjifMbtB7JfLobenqRQAk
YLmqrdrhoGuJRzN3nyR4Qv62GzY1/a2qbjV1YXaqWdSzw/4uYIR0Qfjo7TJeji0c/5wYmO4Xboo2
RoiUPiAovUXuxiceFsbQnyjtUWNCTneio3SkAxYtopkiJ3EzTpCjRsauQHB6bNL94e/feITDkMEF
k5U3gnBe7UcdXCXfGvMH/cShkBr7lfbnOa4SCq3KL9jMB5YCM1AfkC/nbYkQwHn3+210aPmFCOVi
xrqGhX6aYm1EoRHoa2uJT2SsImZEIphmeJe59pAD9USETXKt+ht/ENO3RFfH+JySFA5DAhJi2SKN
eDkfAHE9cEfWsHxS4RBf5c3wbY1+pXv1xNhWAYA2prcbFcfI/yWQEr/3IVPe0LrlSk9n/psdsdvk
0ekV1zpP71shaUrZIes2IKFkauJMcbMucgYs59VCEtTah7M/GObUaHtHoxQ9Ke3QOzoF07PisA8j
/gry7+Kbc0LrpzZITFhq8hsqzw58IWWUE0zHiyq9pP594jGOjyohN2Uv8rHVXrnXKa32Nh323cNB
y3Rrs/5mQkBhDfY/uufHB+Sb3LqCWa8GboG1SnLIPvZZNg3vhUo5tJ2Hy5frkPlcNlRSgYJWtgMO
JHNhJxMYDA9umRUUzimnAlfx0QdSk9v639R/94cC8reX0firYXz093mUJdYwfR6fRd5xr0W61230
5RwEQx/kk354RKUaujcRwTMHn4W+DSoVtspQ8vfd4Yzmpk5/eGK6ClYEtIt16QoWeFB6o18zy/Zc
KErh7Ip1tvK5JNmpkI0tFYyvyF7QWvyUZYi5Dw/PfXHggeeiLJNjL2sfp9fNl4hiFP9d17diozbI
iSEbhxCVgVw49bXmvSm6GrbnPtsPhGc96Yd1jHcY99o21kCwFqbOtTEh87kdBjKoysh9P7hBLnuT
yJPAUgvz4t1xJNfJie4WlQqPgrVeizgj774Gvio2HjR/sG5RDUtx03Ap3ZdlQXSizqXWZ/MZSZ0q
xxtcdMdq/CMlLWOuKq8l0rSPhrw2osOheWa5DU9aZZ4yYmhNCXK/bs+G/5AIBJXkEpOFBKGOgMgX
wVrC/iJgZ7Fmwju71iBN9B+PIiQz8CRNgP/J1Yzmec+XAfMRSGdXsYLZaHrtpHLfm7JcsxC0rjQE
Snzf1mfvX4MUjmoD9/uukH6669iftNS6PmlL5Dtrq3cQYUOeL5dqETZev8XkQ+XKgNK7v5zgwg0T
5w6QCshxSFKbMwqBp/3HJmTdKnE0Z5Kx7/XfpH12Oz9CVV6Wkhmm8xrzsfduH2l5yKB6hRGn8AAC
g4FPt4crdJRwwJR5Z9xhRTMnPmirtvkx3o9LPBt1hoFaWlt2pkaUbWdaVlgp6pmW6s1jBqMo4DAk
NwMqry/TUm+8m8/Zdphwbn7IEb0C5Ej6kZ5IN+pczXqp94wAI1fmicmKje1IPQIqAufBXO6M9p5Z
6zgUBfzb0BqH3IAaMx+wklQkbqkeHQ8FDO3WY+/iLZCT5k1DPMtGYrHkdIGgboST9nSFFMt+DRee
DC3PY/mzdghJO9KcA0VuFdsNrmuInq/m/rKzaGWnHhPaCbaEakNYcClDvCH0F4PYm80yyCW7z9rs
5iJ9dTdwERZn0u28RjDH/YcTy5jJ4YHXfj1bNB4NbbdinLvJAszrQI8upmsxv+e/6p+oxa2xuDR+
o98I03nofaDXyLBVfAb1QTE/tlocdu5Fpsryuamf26WO9F03fk2+S3AqpX0mJKUU+gMakAKMgobZ
TNZcry7dsVN9o0EZ+Y3631225u7VG2NWJGe52D7HKdwN4U0IUBdrbyTaFisavhHv6cJh7BItzvLL
lJB0KwyAMNBOfVYkt3cFm1u1v/fY6UWDizVODbJx3ZW8NdVTsOhG3Vnk/xwGokqJMz2UYWY6rEDL
uDQPsxnJNZ5fKz2DgIVxz9sT0WXjpEMdWXw67bR9TxptQeoiJviGBlQP2wcEdeRMdHXGYbjSs2wD
QHR65OJejyuprC4sjeWigwKfUZQjd+W5ALpXHoOvKE7lFtB7O2fopuRgymVcjP3n7/LCSBB5hBJQ
WqvqLP905S3CvtZZiF58TLMB7opbDwbeb5I9eiKT2IvNSvoie5A1pMhiYXNqQJlH0yk5hh3CJCZ4
rR0msgEnsnOsEfkJKD6xDPCzMe3QShCWgDG+K0DsTz3Dvh2fPJmF2Lmgup/XWQW8zhnIrDDAkldO
X/QUSElveb6c799AbgL8MdtYvRwfiCAWTs/e8kKd0P9dbisqgcXoyvpfU7RNgnd3ZK1Vp7d/zegO
VIzCJ5efrfFWgWka1myLetWYCZH5zu5KvjIG/s2Q6yU9c8ZATNxhc9/n7J6A2WtHKTnLdAmkJtZX
WXVc9EO3LcinGuHjJnMq8/Yj2OPvH3mnLoeZTAVsjmMGbNIUcRNxdILECk1TGQHafPK5UAqMXRtv
xTs2GbqaJPNWMWS39yyyRTvIFI2UEVB/Ohqrte++nGVvXLCKWzgGHiOdI2AtseqyaZXURwEHnvy4
NPllcp8fJZeuPpFM/WVjzUpWm5X7nUCMjFChJ39Q+EYa9omHddb3Uw4oY/1HLv3mmPdE6AUK7y1v
OATnQMQmzSaksYi7/UNfcmP0IgLiqoCceCU5T9hsjmWo84/allXasjeYv1p7H23VpuE6cMGLTBxY
4x+DcjN1h750G+RbnozJQ+6mMbEoYZlfsdJ9UmaK8jGpNQuxIc6zFcNSAifDkvW6Y2IB9WPZmSKa
IUqFNjWXjyoo2jCn940D2glCQu37e8IPYI61N0sEdBcF6ZWxBXYU29Xz+0ZL5kZqW3nPa6Y5SE0v
FA4A8vWfiRWWMOQ1fKDNDYY4tOxwroPzvdzPryQ2ZIK+1RJ7YxcOISALk1WDZTrKfzNAjyNTLgo+
aD0QdGxBeLhQX0la7yiKapWB04yCBC7iSTk8+Hcz6OFgfiIWnMMf6EVs56TE3GwOP1Iy3h3uW+0c
/Zp0t94Ms0MvI4ycbfzm+cSD06j6ftMtFZu3hzph7MYKbJXq+oPxCIBVdBAyIzITfdKV5tC9NIwF
FdlDeJkpTIo1XswgSd8b26r9IfxU4h4YFJAXf6cRSUihAIO1Szw8pdOuEQYshhE8CU0AwwEZC4IS
ER/xCQjzjCpyJi6bzCRfcrLL/TpCAulv5AeHqqJVDADkOp+kcz2YyLkDIjHIw6G2fLr5AS9IM3S0
Fd9YzcMmtMtmv5N6nAss+LKmHchbuFVP5SZ4CeK2lJmlbW1j1r5jBRTLs6hyrQRCnSmHaAoYF2Xo
8yx9HMIFhijX+M9NtMX1zmz8kHx8WN8c3c13zyjHM9ZOdMncXtHcsJ3MNTxJdikeser8sfSB0iCd
27fPl3BDe2SAuUJcslAb7M/9X57egeJRI6fCevRe6ZlsQbwxzadL61AVTt9Bs+soI52OWVCtcpni
ME8dTOJqDjcjVWI/RKBQBk/eylD91aL/Jw+3Yyxc5guMFz/PuiMF9IUmygKrjoyRJ3V4ryymXJ22
+PcdLGEAJtzkmuK/7cWFcz+2v30YYkJ3vIW+P1uf/m93rE93SDuN01byFnT4B9pFaR0aVRbPJmAK
TjXuiSLxWDkOSX0PFEJEwFSUSlKN/mit9ExO8jyBntaYIg+xTYcSuobzFftZ2PxBhNLd/9kQbX5d
cZyzt4e5wLTi64LrqKkc/3pDx4E6YpKTnjQeRgVNKk73woHw7cey0rjhPVNOUJucz+/5xq0LX5xF
K84gOSNfdo+lWpj3lLJmMR0F5Jo2cTYsYVtSkFPIjb1BSALDU1bJitPjqFw36sdcXAIPWknVSEHm
RlrvONZ+0PCs0yGN4hFpdK5QMRd9WU9njq8qa993WTule5nwuxBh7YJa/ggS++CDQbh3b3G7y8+v
aFIl1hFZo0I0fIIcls7XaxcKIjhWaw0wNe5q2JBVBcy7zSl3M2YOLyWzWV+if04lEt33T3Y9SqJF
+Zyy9/3ytagraddgV/jX9qs/Zk4v8LdYExPPZ2eZ6HnW2Us6jvhFhhn0EOoiMc1HYlVgWHdcLIpP
AM37D4iEHcEahesDNiXyDIg055cezJfppbG9g5ysRAiL0oDpvd5uA4sIfV4Vs3uv3aiqsfVysPjO
8eMzp8uaOYxSuznO2+TTQYhgJtbvkx7qldtXcH/i8Yd6JJ9QiWlTpqBZZMceOE1dLMDrsgedGjFl
Rq2+atMZ9KTlLqrt5tF++K+AJTwEGu2ABGCqTYCKjfc0f2JMII5G664SCce8HfJV5uR4FSwN9DDp
Z8S6VDLA1Fv4N2r8RbB/ZgTnvZKclkTwD4lbdlFILTRrw9swK/5PdhiL9lLkzcHCGxvr+7trUiI3
26CvOzseCdfKLTQVZznP7cyU4NB2OMP8sdbKqi79XTtOlmnzS4+FfnnDphHDE+XR1BQHAO8BMxDI
ZwIX/XRuTudgJrhIKbGdd9xNmL/AnrYmJsm5Sm9Hpw8Jl1AlZUCsSu+q6G5fpB5jkXuBaGCfZYRw
Mgn/BZKXJFrIuIgiBpEYNysaHYdDXt/zmVfIhWZg+9zXy09vx6SieH7rlsv/lGQchT56HjFGZeOu
5S1aApHuuhlfceLzfdTZZztQiEn+FGTxM8bi57ryOmUlSQlg3GkJ9ZQ8wH3LKtIek6lckaGhKJve
sShvF3+RglUSi3//ikhFWW/dCHtDV2ZveE2jX0Pb6yXS9MpMu8Dbvf1WM7GdYK5VMzLTVCYpdqPw
VCOJfTjHcWEz9+UeH0JMoDfLn4JrhBznQGTLRn+x2ocWcvSZZtAhln87u/1cGsF3Yz9N5kdsZDJi
jt2wl1t229eUm0oja0j5eiM58uUnBHkwMupw0NBy5VpLz59hsCFRn/yo2GZC5G1sNLo/LzE+YPve
TM6b1V3Fn27gBahNC5W3Tqalrj3FIM9MVroir4Efgok3zAfN64rLJsYjOfJeZPsMn3NY6XoFQoN8
WHc+oP820aNppXkfbqKTdMMiaNaDTJQtixcUZ8Wtv2cIYOdaGHZv1jZ3EeyxpSyG2rJ6WrAtSzt8
FQnjCXqS3niWCQ1eKieXJ2QV9kTxiQHKvfqhskV/zXYFhrJZzxE6+KlwJ/+b0e1RadU3/krChs8S
VnOiSTTHN+wfealiZFWxTW92Rad8f9jCMe+UA/l9/oAQmY/89eKqkc4d/NQpuO1vy1D5aNAo3oUA
YDOqqZmBZxOe01gukoREMGTlLhESh8DmGgKD5nhQXZBYt1GGJ72qTVOJX6Ppr9xlRvhlthSYtlYR
vM0arcIn2gz8stn4m4F1YqKLZzSzfklCLKXdKDSoYLkPWDDf/xbFmv9p32OqSBS+029piFNe6Qc6
CfApTLULW8Wd4kV2ZVpzWTGpmhRGs9pOkRMsIM0q1YgPYREUQ1b2tTEPs1leN2P1yFtxiXDO8CMn
103sxgabMBaSHwTSeT+rROutTM3SgAbzK6K2RZEYvqx5kOx4Iiolr0bOlMdhqVeYC8xkmqKesGV9
Z1rNCxAxgMaQPCdAhK7+W8yWg2uxAObFhETdRg1RgCbsjxdQr1LaPBxdsSi1ujrWW0ozKn66t2N7
osF5nqJyXq7+0jkNYTHSZRmYtwNMUDXx6DZrDjkCCfpgoJtGyJ8VhGoM8MYJvItq3PNSrrEPzDp2
iHrhdRMx1YvRIxZzJoBG53CziWnj2VGP+6ui4AxHdA0T+CV8YeStnvCfre6KQNBJ3/lCw7sFKglm
yVvMZAQ8dmSbG0bhFdwLQslHf4kiA9+Zt+0usDBoTGkoLtg7GVpa/3THf1+TDcQK4x2HACMt/kfe
MHPZd4j0kiVz2gqK4M+ADj5gL1U8Zuj8HrQdk2uN3b/sv0sk2xTp0NlrH4gYbcS/4ttRiCI5EB7C
dA2LWF2n6N1c3KqWdMVytQ7AgxLjmtSyT7OF0wZ8DNJlOzWwDdWlYwdvx/eugbSXPugqZrERRta0
xvL329XTWxAkBWLF5gbfOZv7us2ipeKUw2qUrDTszl2AdpbIjnWMufwwUZCTOOlR274CRqjfJle4
aQg43l/zszWSqOXN1ACPe6ISsXoGWbCMVRo1WEJ2SJkaWsBMFUWyTFdNirAvPdbATRhOxv9J65GL
I9StoCQxahu8zzNv0N2gr9enhceU2dbtfLCMRoDsvgD5wSCxB+iulZ284n4vE69DnRX0dmdzn8YV
T6QrgN6rdCZjVILW4apqipR33XELm1qCHRJxEybwBs04tnFYiwsMjwGH4xJugyEe2zfbBSyTVw2b
GAc/jdQcdlz3NVGmZsOP9U7a310H0ewfB+mdX2VPg4qZn42H4jqwjwAEJc7xGHbKuJyOGOsHf1hr
rdEwc0jRnZ5kUAAIQhbflC7e4HGC7wx0f+deK7xgsd/hGcR+V3qiI6nWIzSK0DzWTJSNZvmJY5tl
ABaRFdSjPRuE/nlS8bqik4mxmfRaIccVfEIG8b4955oLhgypwBfOFqexju/xU5osvM78s4l8vt+Z
i42WWBgugh4F51D/NhIVTysmPbS7D1z4Vf89FKeWtZ7EmamEv8tD1g60f8Jkx9XQ4UlTe4lk+Z2Z
nr2rWaCvAMapPgeMl6TRbA3jwr2PvG8D4L0pQo84NCWN4Ne8YobwJRa3MxYJgG8qYeRyPjkyP+hs
S29GOMqVp0CvLkwZKMVnSCR93xNbjCdd3HtvnbW0WrGicEFLBDqjIu6LHI/dqMx3x6tHMGj7cC2N
TJfiqbXB8zQtcF4Ea32/0VT9IIvjts3ERzRPm34hKTjS2BtaxaR2zarrDVw5Dv0b0AKxn9mZ5RXD
FuywHtUovjNQbRk96GrqVzP3FYFBUrG4xMW4pN3M6FZ6gVrW8mfT78q9sV5WlO8qIxO9b5Xt+77m
skWRYk6dbKhKW9W/KTvVuqWu/MCh4vG5mI79jspu3OR6SCi87BU/arw9phipsiaKtt/UIAN1VosJ
/22cxwYLjOj9MVtusxDagJ+KXA4O0C63kfrJgTz5YAM++ZJZVlkSLhBK/B8YjXvn32M1NgkWjtCy
Wtps8Y9pqjH/Utwy4Ib6hNP04EL51ztDK5eSz/ZE6j6ZCvmcq8GnNE3AFI9i8v4tgmzqerFVNiFu
4gsbP7TN9LKKXwqhrHtX/Xb96HiZyTrxH3Q9yYvf7jcWEZGbIoATPATmDp7ZarqT1MC5vcvgmD7H
vFETM4Wqe/oFPVFpVLUb4oHTKpuR4z76dqhCJc21oDYNeY01QVZNQwbh3R74+ZP4gQgYe4mAGjxA
XXgDxvGD6ZQ6vxjv94LycTS6BZgCkNWqNgbGEMS2E4gqgKNVoIAhCeRy/q3nBbARJXf1t4O0pJmq
gqftvrsqkeowmKxaa40Xgul+BS6BS3DejiBvjqyu2O8D1ILnftrOG3KIbjoxOtUFoz3lsXLMn1QG
k34OEtYk+ACzgG8l0Xh3wt7GZ3dtZKyuFGiztJb7OYW0bBjqml7JK4qCEHq13EcGzMusN2xDVhoV
RuXdRAseLWQffzXGglFbYoFI0DvWGeDhYfxX6sDI6slA46mVCXfg6Zo/2zQDRht/GVLjjwvJrN67
+/9tc7X4fJ/7A5BF5F4fhahSt+BeRTA3cA7L61OsZhxjQFiAzMpj4z6icqsplDzJkigJBbrvwNak
BTsvKEcJNQ5sLZc9cx3cD/88BAQplEQlpZrJm9kWRFznrK3Z2JeMmL/sLDs3/01KWm0qbE1OR4PE
Y9jC/lZK/1+cSt0Duj863nYYvb2NsqYxEXQk5sEN/gBRB18dcF5wdUpmQEkja3mVNAWAd4zpAF26
LowQAw1BMrMRv6o3eEfOWvBUUUEc0/cFU4+V/e6359aGeMvS57ud+hCVtWu97nS03w921D++VCIV
TW2SZkOYxxH96twMHMg8cZFe8y12fSV6kZgU6yOy322mv41j7HCuYu9fwkyiycIQk/gqY4nsD0U8
5jPMY+8LKEkxVHshlImkZNShf/JI3v/ybGiW8BUnXFnpXccs4krtceFjEQRqIl9cyry8xCWJ6qzO
sv1fTKnPMpnH4MKUhwS+dQElrUtLDn/wekQpueOf1HThhYxMgCG1BBpza47ouP3U0esM+iOLOuEb
2QR+RnZEz8dwNFq6n/48bh4Wr3783bcDgRsdA07vEg0sCYWJ4x1CUoDjA6/q9DD2/Bw9MnzOvkE6
kvWPVuUSe/dTX/E/sWxaDzxLD1SCpoOn2X4NgWy6hkwc7CbM2c5BY9XBlrzOcOTI5RLOknEz+iTt
xFNI6godbQmh4hFjItuUW65xh5NyTblkTi+QwN446Ke/RG0hrCBkiz5tMqbFaoNBQAXR2jDOhMdD
5KEnH1tXqahOYSQis116XK0MAXzeht1Zmh7evJ54XjlsBvRZqmHXOOgNb7HMKIctrgwIpy1PZo5C
egvYqmzDy3ttNDsQjgkG0UMyAi5wOf3Tio+h51Ldj29EyccjWZhuY5PIeTnKB8uiHAiASCR9jPDS
ukhdYF5ibT7ws7W36aG0C6b+zEj4I0mCCJh1BBJmVhjzZnWM/UJVGUdsLGcc5lnAYHNnN2OdVrxg
/FzQG+mByIp28F13wse6sCpI2tN9pgftJ/XCjXh7wpW5dn7aGUakwVwauG82lD2YYhT1APpgNZRt
0IZqOp9CHj1nDsmwPemyDCXfaPmvBmb2DgzSIueDNYEfVkXG/uAN11x13p91L4fAtsSL5n2HOQEt
g0zsut7Mg1Ms0ho+8RrCABOH32+lrd2yUqJKfQNI9g4lgWmw2mOGjXHcwNgLgzHwKBitoyeRuQuY
1JjYQzk4aJWQ7tpPkQ6t+eTDnestiMFWdOuRwB8LzM/0m4/LeBOqimHa8VXBgc5jTC1uEbvv6OMb
vbwrAVTUWIiA+IFrL7I7hS/Au1T9P3E8YvzSPVDRWaQiyRfIN+GPVksQKbrAyOFuG9rkhSAlXcXv
hrlCvUvKop+gqThFRfNMjkxUEt2LLxvQqCyF5iofg8oEzMcZHDHKUZDpciFOKmpnS7P+mS9HsG3K
DAnHncxVOT4yQZ3idFUgFKa7QZBc5FpuFTTrW14CxJN7Dgwnfj9GjFWxsOmY8SZu7ekW2E9r3xHb
L0t33PE5zo/PoBMgca4MLA+jNpJghdOnn8sn5yHVru/qewMZHQ6S4Abx511OmNRvWP1bYgln4BuC
1femvyRncKI10ZkllhopaaDm0PcrBZoDjpDj7/ZtGywHlMLgxpk4Y62duyEnQfOFlMpbqITClQ2V
PjA0ifvk2CoV2bYQYO80qr2e1inMV8Q9A4tBlnIEoBezViLexHYiUHEtbU8a63hgMcmvdTEKINgF
izQbPmLh/7YssCeRA0FMAHKwJPy2QBoCrzZuA/RGfbn/FAvbDBkwUoPvW8Z79j32Hp1KZ3RTh9+M
1bkfEj/LS8DXbrJYS0Ts6O450cAXt5vZqSmtLSke0l/0gD8p496iBo2b/DIQqfI60qWldEv4rcYV
GQKrmOOG+fHi959fLwMKddG9zs6PnCrCe7H155DtX/qfVOgSOKAEpLcjz0dQezqksSD9GwQJrSYE
lbjvxqF0DPwtylBB9Bob08Tsl+wkewQ11YTKetDR1+el0hOE+3jL73rUiSDNQHP3xTOp/fx1xWUD
fPRCr+DScjenRr4odUjDGzSu9Xc/eeZ3/vTPaeOYc9/y7sBz3ww5MDYdI9g0dgziM4byHpdQUm03
EpOwSSqLIdK8QSVhyTnbWGeTbAIvTYBGXZ2QjGXlr6KqBeZIH4LgzP8toXs4Lr7UxdT0EpOcFKzG
OpzIGnMzPteXWJy3N2P5PEKhkzE9X4cVJIkcHGStRmLncJqF5j/FT3RTLVP0epy+MjZFzTKemk/d
rkHHBQ0+nieYtiDgheZCbfYsb3iKLcLIdykO0VUqMa7fNRx1lwQBf3YOrITbiX5+QNJci+s01DaS
vZVrak1dTFgUSVSFflaZzCiVbK1bc01GEz4YNLPkGdFOF4sSuOOz0ZfjBJffeopxPLIjdEfFNjeR
2EROmCt2UgudIc91Y+LEOPZ1m4O1OznrG4rDemHLjcRZ7b/6VSJN5veOHB/MqzLntNo7L84vOHvJ
6ZHn2V00wSTwt5uNVbdQI8Nj+8cwf6LcwqOAQgioN1Vy2ShdyI+lmyFtxmC4EV4XVxCi1fkfQcb+
8UZj72ZIXqllDHG58nMltVp808c9Tt4WA1Ss82QDqAbT/cO5EFeMJmM3UeBmhFYosZnZCbesWwrd
kM617P8b2QmdwGicKHvE5LXhY85v9l7Uakk2UovMfKpEnoJnBBSMX5OX9sC2SakYrg57/J0ktD+b
B2lTBNVKVn7L+DF/fFxUJbYGzCkt4iVGVBygQBoUEYUaDcLSD8+6hETZYl71FZDtUugzNQuiVPaN
qIgk9BJORc6VZPJrWDqR5yIAvmGSzrp0dBvDN9pL4Yq6vl+BVJLszrSSWo6VJRBkFVO0o15yiRLD
3yqNtYVZOAmECthYk8doPFozBlCgznHrb8bTcUJTkXRKW94t7vedMzgkVZvlDvetAZ0Nkmc5tdhM
IgJu0aw/ci2hUYVAoS+R4Y1YOkufVLMzchd727r3mYAS7Y+shIlys+gH5yQ1w9neD6S4/5XoQYMk
zr7lwBvSJy4VYGJQYEgl3hRu4fG4rkMXaLNj05HCfhtY4uePkjSOyFbY0bGLdgpWR0+YI3ANgW1e
PXZBlK4m3kp6jVLY2uBku/F6bY2ftlvOKEF/WuNQWbrak/VTGrtmbzE8sS/Jcz1tMOLr97DrG9mI
m0LlCG/isGZEJzPVv2wTYpi7060mw+WaDUl0McpypB6RZlBAU30GbQe1WqlUvtB3ZBSeGpxt/yRC
srvu4XaEDOVHvoZlFqlj0gjbPhP/6Un5KZxfqbZDIa1iRlUdg1UuQ/MzHUeZAqqBnF+lHFvbMReE
IrsIUNRX96YYoOtNzv1d0tnIOWVAuEwIvmZDyVtGCej3LjCGSCfrsgKcNPuY8KG65roG30nj8167
wKMkZ5hPIOnkDE/UsbMmkIeXYguXDuVMxUbBtAMJbzUmE6TU3bQWwLzXKrnam8POMD5eEhwk+s3x
KfRFlOlzvu1VeGaog9bdXFD+w7yCgzbevBNb4ziPAgF5ecl6dgbLLVIweKCAWgXKC6zQHvotr26I
UErHrT+TSlzSO8ZjkZwUsdv7SnlEOLT5XvGQB/DvhcS4+Y4yI16TuoXYTEtzn3FR4mfRHqAXlGtK
HhjoEfZJZdzwTMJb5VRITAsE3SNEtvIJRhxRB6QINIenvd9cMswuShc7gR9D4FMsZ3Y7eXzneisB
VI7cTnBirztf+rGtfGgmQ06W75+cgg4D5/VtrBV256XyzDou9qgBKrmNP5SwWh72ZzvlTp5hnbYz
HsJUJdmqfYggRBSaZqxThZvqynAYmB1X09e48pAEAcpLZwxwrP8MWzDXxqevLp7qyXAynXMG6vpn
vHUpqDb4kaV52Uz7HCikA+r39ByOzB9TYVSc1UYaxKIKzx8yAkgXEC87668kSmuz4+fqdld6PoIO
vpF/Ud+H2REg1KjpBpVAJLyvBcc0uHRAnNspCaZPG9uRjv4P450iMwXBgUBQDqs/C4pBpljyhyRN
i6xpwN3BBx6L1Aro5zC6gt7fEh8+1nEGKAkPFfNo+oA/Miyui2n6032VeMlgC1F6W38beyDFS3Z4
MbWNDXPsjoEij9PL4mwV6ugf+HZLQ1rkq4WlHGsb6tvYVjSG94Dn7Vjq58AXuvVMynbsnQlBRneq
rdIqGhjZ89wtqwOvYCcylGzo8iPhaAAHf+9QHBmlSB9JQw1dNBeZ1ebeHBLmwzgEJVN8fGoKZZwH
/kAICP7f7iNNpvcdBgvHfQbB80qlE8nFdopJ48VkAILX4eLb5NZq4kwxVwgGM2yM/c8fGLHD+N8J
CmodxC1a+ekeVMCp0t9WeZS6QkM2spewOG+2AfHok1DImgWW4f3bc13pIX2WqXoOdfT51yZRx0jf
QgXuuulB/n36RozMED0IiyR8wDWlVONQIBX0+LI7f6ezYt0fS4Cy45+abaP8+wtrl2y9mJASSQKl
V2PXDnoWqEcvmI98htDhAXadq4Dy9+xuYeqlpVDVJhsqF+qYRIgy7Lnt5wZJktA0q6Lc9vqH9nSs
AcEE+mZ5BZQ5z45MnQxcaKIpaBX6EoJ4a4OL+JzWfM8xRHkPIWGhenb85O2AKLoH9cQiXyDOU3Rx
KE+BX04OLvyHNaQM8r8XwOzsdQubWd1ZiCsetHnUlyhNIF42PEvC57aH+KFyuM1CYmt9a6TSsb4i
7Yo138Sj+c3doS5xtJjAcllKsRfdyprjvfIf2Z38srjCGtKFIiwjJiUQG/sjivj3FUl2GBmMyQW3
opsef1fY35OcLqzH3F3ltWaQBAHdWPjmpj5Khm8uJ0hfj6gPNCNbfp+GDuNQ4nzxKJEpWOkDMQ3i
4gcVn+sE5LU4cSkoGDArEZf+6qPxBcqCphUZrICy+XN49D3CD0/3/LwLM5m1iYSV3DN9S9riMNMa
f9MkJbuBGT0rNmqFbXUSTR6pFbL3702/bfkhtJbvDDpz+DIGkZpk0hmJ2K4xEkWLYRZKoELWqhva
9NguptFPW/3xmI1SYEh5praaVndlnVg26S/2KrwTIIClj8SHFPcP83q+AXWk2mOdiPIxftrIXgsn
zn02gywCr3K6lGeka29iyaFII6E1OY8eBab0i76GBDrsGTQZNy65LLV2KT5tKH7R9lmRMyMolnJ5
6ho8ABO1+3hysWQasp8dpYbhY7GGHBI67KAQbAapSoYUQ83MtuQJDN6c5sqJbpgv55HeNEzRuHNO
5lAS9566R9Pih4jCJFLa92C8ZTzNIdMPtS6v0yNCGiCuXZSPidFXCRi1fMnK4YGLUUIAtCtXrghJ
bcyglh7fYvdgzs4X6jvFAaoyKPmvfUYAp19fZ1nIrIIriaRN7ooWT4bw1bElUOWDBpBTjQ07jprU
pDrtn5c7DGdQBBwuQEeGUoP3PsO7/iFw9ykk3IK+oBIhF4UZMcGuGMSBmTCmFqZYls22+Ejy9cUm
4pja4JPXdrRceOpXDjQIrmJjJTQtJuGjiuJRtevWwPXGzVVi/fG/XKtujojTl4Rl8SWXE+UzmdbP
TUr+fz8rUNLnW/v+tIA46afqTQky+BdnaQvmOIRMh4o9Z1qnD+dVEUocriidbgcgXH+WWB1Rvddt
OGCz/KOzCSa22z8kqvOXOYhjn9th7TdJjsePNqRKLsSQK6+jcyghEkK1fKeCIkCQUPVFuXQY9umx
cVBKvRA5UhpStNTuWcoLL4MnIIhy09zdtstgudiNDD4x0IBuf0a44LETyMeW3XGgj1T4JUgNbShJ
AaF5ZWMI9+/MzATd3/O9RwOPfu8lYld6LSvqVNw0Mqg7kO4m6Klv/ZBM4Ar9lM7McSzooCTuJeLZ
y0WoF+k9STZBJ3dGVd8yq1VN5ObzXLK8HbGP1XNJ/dd7ODQ1JYGaYlXFeftosxiCcfHslc11fZzE
z8xtkLXV3/K0w6d2IsKykXep2+Xd4+42ZE+KGt3UleRbyM1fPHQw1zkOoYchz6ydHewGnSJZtMxE
vv0hcV506KpXUvCcv0Q4RSi98xzay7JGFxT7MjixLyr2y7/bP61MPuOKBRT8+LoNOzUCK6vFFFtF
Xu91EA14QpOhoDVU8m7GMGAPX2VuJOz9lD2I9IiwVhV+RKbv+nZk2reYcLMT7ja4PR3P0WH6h4d9
Zj/vMvZSN12ml510s87OzmaqFOs/kLPQBuwEf3wRgKfMmgZiQ4Uic/3P4SxRNrTniI8FI4A/jkkW
IPCRrCqScYTLYx0HbQKDEAQavU6KDyFqFpdirMFIJ/RA0yWoO2q9dtNWmhZwO6iI+f7Ost1yjWto
VlFR/4Ff0ObCAEhVOPastNv/PQxusyDjwePMz9VhhkvmGIJdhrqn6cTCLeK0ZMp68XqZMu7Fg9nA
xARVguJVD2PDX5WKQxgzjjiyaa6hi3Brmn9ErAxGFiBAC8HTCTJoOoTA2WPvJAItB25ApEF3oHPE
S537unATMxzp+zAXxkzQZdDZRXpukPH81hPaJgtNJwTfwqbSICfBOtwTfI6zUJSpQ2SAANNKpWPk
DKE5c7V9VrPBqqncZZr0cqH2dOI/QyDsamlag7Ofl2YBqqAB2Z61L+XjHyCx+3k8f4YFG+RqUymw
JhSFmUvJSZYgDO7cnJTbgB5CPChnEVCDAQpqit5ZlLBmancX8msNKAIRQKhhdX3Xr9wgUOY7515M
319O9HzMWkv0G4Jq/viwG9PS6WrbSZFS6JLRCDhGxECB1+IvQjFhOJ8R6GNH2WyyYCtG3zHotsXW
hF4Cf4OX2D0GgbRQKL6hntrLyGnZVHxhekhCH+pDhdwxmURBjd6IxaHA1Od8o1MQ4D2Cb6RrucCo
82vABfFyTMvnrE1eZVLcb0ryN8fCYpvRfIxcHosjeiJTGv5oVc5NIrRlFw36mDoAikCUpXUfCgzG
YA6it86OWY5tah5s4W+QS4XItnWneR1LVveQmfPpDkwTOgOJhJbBsusdggnpsa9LlpfkyApYXH5F
uTc+oRpZ+TciRUHWTzbTTaCyIeRYrDijTetcHdcdNJyRSGoTKRoL1am83kk2OiiS34wFycecZkUc
I1/x5wBElQ9wwfw55mLFz4h0PBfgDT9hfGLfjzZ9kPCbCt9e+e7rdxXNX6uUKIsavvDDn3G2xSpR
LhGGdtv/rEem1eY43QXlexOqNhtNMa+WaExdkAoW6jGlzdFaLLUyV6YIjti3uXKxdoRHswrMBUuR
l4hSZSSstzPVKMPKdgIzBji03ojqGJobpEARL4aKl3DwlgX/Uc0LUFJFp37ecIlSqxu8rfFFYaXs
BRYUbvtrK+TMiL97LNcNK/MpKblPUBvST61A4CbV0Ibts7Nr6dOa2QDVCo4Ck68IUR4oZ+Xu+a+O
ai1n+UTSDkVXVBYf2LGN7wuDl6z9tu9mutGqnIChdYyPzK38hc3A6cohwtcmHSgTMe5L8FEJj1zR
BFgRiGuCBmWpunFYWf6386bOkvn8/bQLs89+CQT1MVjHz8Y5Ek5IytXkA1JTe8LwxXGPMLd9rPMn
YQz74H/iwF+lvaWCOB+bec+hy7YmfPIZhOVdju9J21r8CkSMq6YoV2yvNZ70k9yFwR2AVQ7MM+rL
iO3QMMFQjqCqQOYRWDALaIyExDKEZ5pjevfvvNckP2OUdM/6svGoD1ikVLTL+EyxhxKbj+Nt3ayF
lk+2GDOE3CuQ/WyL+6Dt8CG86QdPnpPkSwJ+v3/zuyMpL/WKlIE6+0fMsva78k6zsPgto+ueYZnC
pPEPfLVEpvvnE067jGJLSDJzKhVHplU=
`protect end_protected
