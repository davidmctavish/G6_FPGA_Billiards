`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qXwUbNWAqYbdpqBgu5V2Irr0yIHokdWq4yIsYatvbtHKhU5sTXcicxiWkZwMlmh7JxJXXORLT+ZU
v/PLV06P9w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
INsIPl3meZGaPEpm/0hY6qn6pNkmquxWy2FiThgvPkXiH85UtEqY8o5v8IRoHwlNbiFMfARYDbEO
+OZA2Z89jPi7vSGZam1nQVpdb9tTe8gy3sT0W8L8+/zNcgLhbWP9KgDZMNF+3YJnaj0hueORxLD7
CetUAimRvUF+Ldr4nyU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gJNTE+b/peQ4Oto07xlVbEfbFZ6nMfBGBuiUK4g+q+PLYtJWQI7QotLPwqtbFK07bXzvTJuyp/V5
wl4PKEJefSdYOEbPh6MIoiuvoQGJTFadYzFpMqBoF16yqhXJkL2oVtmXvJfQIITgSFazvP3qKZh3
NjuPtF1edJvfzpI7PLpFpZGoayowx6z/jtYsnIk2GP0W7YdZ9cOlkiSH2S1km12oKXLOaR0rDUTJ
ebEra0Bgy/Z3Q2E/7BECOXrujkXocR8xNi5Eaeaa53/ccDlgYYbn9NCrztVKJ5qtFbzqTQTW0d9a
mJndrp56FTBESQa//wxKfj8ZblMcoVBhTmzhNQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xGHFc5dhsERwTBJ6HzSxtgI4YwpmHAsH9SafoAvaDa+cI2KAeGL0jrTiG3tkhsE6iSwJrqEOYnBt
n+EBnh1QW0+XSDRvU22yYrXld4AFAowoDmmRvGl8seLeA88PptewzCsn0OcE/MP4++TlNv7LK5dv
mheDDGnWdYqkYHdJIIs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jbuyhmw//VZkr7Ws9+6WrN6Lj7dPBf/FX+UDLxKbBrhbv56fo3Y5D7icn71R0xbIApuFFtR8Iwcm
uySbAa59erYexsrtv2JwyehWzp7rsT+wE9FVJrZ76BH99VmVzK8R26yYJmnQOxniTZ9Bpt/l1Hgp
bqR9KddxVv7YR/TVF4FIjFACcu1LMYgxNBjvUjYUdYT1kFzIT54fa5kEBMPS2KGJrfY9RdbMnuHO
JIGhONlUF43KljQ2n+XLyCeaL8y6a2Zgqg+6lrVG6Ztpt3ZM95CTfiRQvsefR4QauRmUQSbN7I6O
wmyxcB0504V7UGeVSRNaInvWNlHwpFrgxy052A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19488)
`protect data_block
ZOdI0iP37J9pIcofeEB28BfxN2U3/rji4ipjw5lr6o3x4jhbCjwb7Ztbz/CLVL8St7mYcvoL/dYq
5+gWUzsl7Ydljsakd2HM7+lvdUDYlMDu1ak7l4pPaH7afx0UDQEPoC7zbAM7mpb1xLfrpqGnpVW2
JbrdFDxT9mszhfrRlEm26YIfkwPke8Y1y7yypDB6JxxAn1+nYfiPM1gklBA/wAmNFZ/fUDPztbOx
fr+b3oAiKEicuQhOXDU2b2grmWbhknxewEgKnKv+W2/jdejqfVh7P4/yV3VnVWs4fWuMZRv91LRr
Fm3vspLbkewYDRcreiIAMYIyc7Rt6gqq5p5+awdEBeWb14JtRbIG5FGJRFY6yuZDzFP7Mt9HWu8v
GpOIzL522uTZg9CYRRXFlBitsgVKBZiJy0ni8tiLM51tYJMvrl9gigTn9+YckK1bLrNGcxIrwzjt
nHffYtRVHgweShPwnVv/aUkIiUM2O5lqvxwKvs7dzXxv2Q2adgle1XLlAH67+p1MgkWk+mbXVU6H
wJUheYWopF/lhgFE61ivB1qTJyd6j1lMaPiKTsAAtEuxaBfbCEXNH1T3wPlCYZxUtB+okycwL9oC
coCvP2Geu8Y0Z1mNKu7u0R8xw9OB1EJ6GRlt3Aj7C0Xguq6pyRnZrSTNGRaZDZe6PLh3Dx2Xdqa8
Um7mAdWU6wYY0qMQxPOmrYxh2n1XILRKUR+dNrHLwP0+8SUdSN0cMr5S5UuoX5Ob1ppAwFqm9KEk
6ifP2WRzfl0YqeUpeDOGXruOl2JKkdlldvfm2LgjUXgm/Ei22Bc2gPEmFoRTYyr0QKH9vH2DaJDW
Bxr27qjuywr6ffYod05Czc6HCqt2BmVJbhic5tbUV1TJs7vYHLBZI/LmngPRp090E12m2t8MpsaQ
iOfQQO5U4wLXFut3X12TKMAHeP7k2TBQwGDj8J+4qe5FuoExKXd+WGpIA5rWm83BPjZb6k4s5aUj
nH+x8zoZet6NMQcvzm3mHy7vvXnqbtFBC39UEXGqqO1XNNaeNZIgigmeCaA/C30Zp9v8TRgXqiWi
g9NM40arYrmkXiDwNOUx9Pk81z7g7JAGAtzIdlYeCt7a+vbbhkpWODL21g4pWMDJ8hepuU/Ji6CY
2VAtCQtkpi5p+tunmxw3aRdrqSNoPfi8B9Y3SgSgfvBGzOPonbaDIdGJJEuxcb29Hxu6f2FLVA+O
KpKRALtdUC/kLjpzkkJ1eAvNARPe0fccPhw9fweR+kIaAncKZuymXizBwJ+IVqoR+rE6v5PtloS8
Y+9zQQ6zStv/79cXQQ1H7dmZBpqdeyQj1Lyv2lRAcC+y8t5Tjv+rcg1JLydWS9coiEt3mLsLhuS7
mteHH+MtWou51Ez4DLMgXkanfxi2BQXV8dJrV2tNEwySHkKmER9y44AVhUqEQj40EMGUWxTxInDA
ESfN+BZgU+1qhi6yXqdSHiDd2J5mfapKajD4w28dQwZ1hEMfSWqRyPObgUHIzd85zk5cToJP2g8i
TOJHuiObOhXQWiBtYIUms9teUuGI1+mZIy74ikDrmh9KcMXZuV54+jEfJG/F63QPQPwPlbomNbTb
t/QEWX0gkdwe/ZHejgg9lO5KtVVeY2W71CPPS7pBYs55eQFlDv7Y8tsi9buPuoF01KN/4cyGFtzJ
FDWRo0prEZVw7QN1HyyoGO+OgCWSJ9+J6cgQ1pFodl9NB1TphCx7mWg2t8aVFfTkQnaFcfvcpusY
6Yn53kU9irRsop0uTzTea1wKd01tWzA52vKPnFE1SLb+Q5xwGLFAI+xej7gm2ooEwlb2a6mSYxlT
YxZtrtZwBN5i7j7UO7FYj7rNr1E8Jn6gSErhxJcgO2hPdsx0RsuSCvWGtefN/GSkrXQesBzAdu2Y
mhgFEEk8LmYSlwQj1rDpWCCr07lzqs3R0y13S64VG+aYH4l8gIyd7vL9LURq5kOyAo0Hxhp9uvdP
JihCbqqBK11Sr1kXE3cL7l2m7U7a11LRcNLMFJDrTzezn3/7INa8q36MwZ1eh0SHcyQaKutkRd50
h9UEA+lnVTIzi9VjSwe5J06ax+ANn55f9UtPIRGqQQOuRkrm95mU86dcNeoqKAOQ0VEcQUR2wwLv
xO28IqToexdE3JBJbOIE/Acrz+opvMl3gE3T1t1CeVw//jc1Wg22ZfVG3niStXvLtetMtZA1qgdK
Hk93Hk2AsTdMP4EJK8O5uqpGNGrYV2dD0YpmxSfDUcHapV0gXDkLdn02Veqq60L+VM8yAs+8ZgDB
AalwWM/OOsLPi1kNzjfoy1rgD9mbQIPMx79nfBn0ZYOldkgUm+4pc7ch9ASgS/UOoaQobUfGfTxh
DrqkbkoJY8DWgvSD3LgwlZ+dfTqLueqxJaGEf2j3CPrTWN53pjW5GmsjM7kmwd49yWJ3Y9gIDacW
854gKsux7xL1kQ1EvEbIpzynvVW8FwUSKaQIXv3QXQehbvBNe2+NFrG42fm6Bt1Jnn2EpTZPmmMJ
BAM8y7hqIqJAEJttbS+eO6WqJHTXs3Uj9EfGLVVQM3mk7osvQtCw0+6qgal2X/MGFRFc8Jebq6n0
L0aAFwCmGk1QX6Ohr2nM6o3xqF+a7E3y+WFlKuvrDsLQzHEJY3duKaR+E4vONhvRJfqUgvFZewMs
0cD0nWCm5Ka/yfI90gTofvZi4Fgk24utJcaOqVqBCPGcu9MaPidFKgKGFnyr6M6mqyKQuEXbY54g
ifbECttY050nG9H9z/k9mdEuEHLhrMQ0kLmY5SAR3JiFIms8dtKPIDChKlPIRgI5ynAyoa9HiAmA
IWmQTzK9dkUvKE7S3+mo5SoulQ3B+qkEfaitytlI13392Drr7F09ThJgADrcTyMsN8oF32+AXh70
rpc6mltRk269YM05X+jXsfTNb0bO6Mc5eAesoLYSwqm1CGCb/HY5RME2TlqNUZQZPHZI+7Jo1wwf
FZ2e/pehzqf16buKyw6zBCoDvSJX09g7wnzGn9aLKIuRKmRE+3TgvvHQMLK2WzYKKVthAW5A5pPe
rRZ7RqJ7eAKRNf27mgY3XnVA6D+tK8+N97w+zQKprfVjpTrZ3qwpfhHEuzv2o26vH7ExL9HxN2+L
cLxy5aArT6gdlf9cyhHLLUh8XicnuHHDW8BsKRtq5JhAg5zTf6KJRN0uhArS1djeg4MgOr+2G+8K
4gapi6CGS0I8j65GpZCo8ZW6Bcgc3i0BRKVprsXfScxkip29co0K96l/tGe6hc+SVuzX2pM2mabv
KiolZIb5BUaHKV66YIoDnQtgg/dJeCPkKt1F8a5FfkF37NKOfsYsxG49crqXmFnW7t+OFJarMj71
ZvwVNmILzHLaNJrT/JOOnsVBqxvOhqWB93VDTcDFqz3eooibgxeBW07NBVLwzjqNK6BdFzbaN2zn
mTTnx2iq3oLwKdblWBqJtUF3EbYDtodJ52Lq0x0g88JuSDa9TjhY9PRog+dv9KcjX14bMsKTwxLH
7kvjetk2XsiMJPW1z+Rn/7Qpn2fFsjh2SO6yiUj3lwxIlj91uK299l0yyu90Xud+qlvA5OqPm17c
wliUBU/xZso/v2DmL24cP+KGT1LjyylAkqnFx4LKM1ZGmlG7pPNW1MlXVmQ2Ix1Y5vIbQO/ck67/
1DkqUFNDzljtYy/UVtBSJptSsr/EQkcx40pNjmOO1AFtca8Y7rsc9a4ilBz2sqfQbcQvY1oEgLzw
xHnX+6HLkz9u9F01n8Pu8to8TTYoF88QkE2xrpE/s1nh7eeTcUydzoSz50VNK2Dp+sELeYyMLbPr
quzG/O3SBcG84HmftvcopYAiCkvKoH8gTwdWNbP+VeTr3gu/se5YPo4Eh64kGMwD4s2pHI3C7WjP
OHMe8FfgFBSP/00ItXE5PAgWP46iviqBvNLeXChWU+oTNyXnIuAAXEE17vYDCvusRbCk16RXP3To
v/LDgUlNiQiFZ3MzaFFoE0cwNy3GshCm8sNTGQaXOybw5lCJIsHhFRLvhh6yp4Ejy4+Xf4sODqC6
VybJlZkv7jT+sG+GgUyIG8hHGSpM997CqYi/pKtbrK6AfXU0tlL+fDDdxFjv88D2ymeVIN2JREmy
0m0kOdP2fYA7p20Nct6hi3VYi26+g3nAFgWOS9p/uCt28qYHtuMUqd4BH+WHeBDwzgGpjFslB1vy
d1JtXXHmiFz5fUv+vCXFPGNesDgbSOwXh032Pkv09zTgXwIL2pcF43Uc57ISMKf01sBAw7gRDGFp
yDH+0KdhHWURhzKBmgm94cifysCskBxhQtiQiFznh2Kn/Qr2hdHqIHVBFr0/oCL3WfLjhztQgpeH
/XBEFo71zvd1nbpq5mCaEJuR3napCAaaht1bmTRGt+QGlZysLO0js8V8N8Y8vFVsA1+muSmyhZ4U
NeOxfxrBZ4FGHv/neKktZyNX4qKBBjJJyCHGKU/tLmdB29Jk1Nn2JBmaI4+GNcM97t6EBaSDoFWi
O9Ww+w/13btpNXWBrFLJgPSdN7YDRhczAsFIhwTfUDmEdfSeFLf1XkbbRDgpHOdyLfAyTWSWs8bX
Mg+XifY7MTVYCw0IFNWj2w8CpW2VIFVKaAxwpHoCS1aUSMYN34zkkCUB6leskZ4s13wSex+BHur9
qfdwvHGk40WRwa6xStvNoLfcN2PMiv0z13UvsyFLv9PsdA4lrzfMVH3HRlIz1c9+6o01uPuGQJyb
/5jIMkJz2IbWV3WjW7HZDM0et+LpVmwRKvobZ6NTAyXOSAJQTOKqZwOo0En+FStcHJyqysjhoJhQ
XN4q7KLrCbrv+t2MmUIDHrlXbMi0EhI6tF+Yl+X5wxB7w1PnABLrOU6hqOgBVhYDVGjnSEd4vnhe
mg77HyXxiL8VfKFFmblCGsv6XNHfvbe2apWbaJLouWczLl/LeyrZF0TqvLjleHJCmCysLVgE9gQl
fv0yqg7nr3f5pA4bPyZIe/Cqb2LyWv4nems9/2B2BLZQMTj6ExmqOPnd/URjkNGQ1tl6UBYDvjU+
SmE+uYVPPmrw1wMN1B0VeAlAGLSlHq6A/kSumhbQ4Ozmbv6Jb5WPZfb900wbF3vMkGRVun+zjy22
NH+4MaE7E6kLEyu0Gz9X9F9EvMkjMeLoB1BrW9lgMcS2MaQC6ycK6bjuI3xZwAADZrC07Gfv/R4k
hD4C+jFX/I+l49sSOZ+I4Va7WvOoqBv/vFdon6jAfQZUWHTEZbIAc8CR1owkpMK0ruKEny+MGM7q
bA/EeItFHMnZ+8l1bWGHngzZH/X7BgmPhtDFU8OaZouYQzJ1gxLFkW9ylUBJmXZNS9X9PfTQx4RH
2DuWIoWf2XZdlOXgOeZolu8v741TXGSdjV3W20X2NLD7Es4on7oHPJ3WdwfpL+kvFqm2vjQwYeys
Gjz+o0A0uMDjCLnK3ubECYI1aaNcOKJRxML+0lD8nFaSHz5InhhkZ8AQesugPedEsDMkXJL1ODY3
04gEn1/p/j+zB6Oa49ti+5Z7IhXB2jAAcnJzDfiwSIwHPzOJkAvbAwgqKM4k0VIq/mhaWBmC+z8O
ZIzpotsf4G/GSlcSPG3nKrDJQpYaSH7WxZ6P/lj/eDFq8Kcbqv56PdGJWZmALsL9xXTTLH5rRN6V
kmaBHX7zGgUlr8iSqwaD+8uUL4Nl3QKj1EHmDoxpFtkzgoqqyRz5f9ttxWJ4Fh99q8DsbcXyUFzB
Apf567qAGFb5gFjKlOEWCLQAv4tWjONBwZROOHN3MEBYZi0zI+0NSpHGcIzzIKIz/FLBqG/qlMne
7upS1NnlCSBvoHFxzPxEYW0UJSn59C1EpC2Xcpo/ZDegNfmB4Q5Y1RtwJN1H3BZFtGcc+pBu0gaR
8ueMPiIIUMrbly1C8DFn2wGpwFGsIdgaCDPKAcHYQu+56gKAmNFXHntiMyzJ5ZMQPEKe81SEJbyP
pZBUKiJtcacOhGCRtEraA0b4dZpNv5avVlbJ71S8o/W5w0XrS59r6RS2H5C1jNQr+SyiLavq0nR+
L0Z8jvFzWbZeTpNWmtBKiQJ9C4y14hyPqpBzGYZXYPyDT9PF+P/6JLG+nWBmphjAeKYIskHdar9t
WFCHvpssSnGuNM3IKMWdpHij3uH7EBSO7k4PQFN5Sg1bg62JHbx64ByZZdl8mdeCVMDBH0BbcfJO
ZgJnRQGkY0AK11jtz2QAYUd572RYvLf79P7X6y3IWcKOELGKfoJgf2nzoZXve1zrbXnKZ5I57B1j
KuTBbm4ohJnTxKTBhJxBRrABE2XBmRrHrq4ZSVXlOiJ3jicxVR3IsIb0Qi9tLMZ0xZ/ox0ZTv65c
Os0VOgThk7tJ7SSYdkXCZUusgEezAv1HcaO8qXQgqYo5jrwVJrg3fFLOEKiB1WCddKthrwh7ucoj
CRgQ64q+jfpC4UlpEG4Y3iFHg0oiwVQuXfyOqrXOe3LYFcE0OjZu6bTUc79lvgVMmSaBduPOeY8W
ACKO9IG5MtEGNOXxVAEivJcLPs2FYO6NvohsA19nJFw42p0sWFyO/cX/ziW+iQanfx8pmE50j/Lj
HDX9D7GT+V0fXaV2OPECFtOK98gYHuTFjg8G6Vg6GYA/LcJoO8xTCpeH0hxALcKMC+sUfkKv47L7
I6MZs71b729VW16ietYBR2xr45jKWxmP90n3F7073OuxhK8XDEl25LMNdWljP99CP0T+8W+F2t9M
COpLJt/2vf/AFsHPD7+zpqmLnuKhJdaJt4Xv4irm558MLxmgVcYult4szCO6epTqi8xBO4lgViOJ
L1AQ34yGCDsdWqmlrHU5R52tgWjWR0VU6+M7DBLkr9detKgC0iUBPHrIQ2xE/jHlqjVJ1K1zpXNd
AnXJHPSA53dE98SmHldQA0XqC3gnDjYrdfP7m5CssIRDusCQ6fIzhnYIhdvCh5yvnRx56LUo5kqq
jGzTxfX/7lXKl6joSGrxYafMf82zWpGmkZBP7HMIaJOaiAbqEqtp8FA+gX+4ixw4RXkTKIyOgKqC
s6t+GorHun2o0zjflqUl+dkoBTpEaHGbgLWnGBNtsI6sPvgJNebKV1JLH5p2xNZboBO/vQ5eP+PT
/pPKE2ddDZ4xKOcJmd8l43ztFtAq/+z1OIRdxAvseuHcTtKqo8+S4MoC8A8JBNEA0nDFzQfTgz0G
430uXYaVmT3OHlBYclptDMuAFqx6ZxovFs6UEa4kHc0mLNhWZdhjmo8Aoo1Q6tVr5fJWOJYuTXSK
og8w/n91yf5U97nHbr4LRVe3tg0GV+UTPnMkGHzDiqY9RMdG+jy5koiCaY8jm+loir5BZQmyrBmW
65eDja2+p8o81LSAaKntGuHfNvxJ+nna7lpJrIJm5dCwKs9oQ58htKhUQ0WepBnaOQtZHl8V+wMk
t5NyunSHq6QZQyCwQ0LOyLlYvLhCpz87qjH6QKc+5APE8G8RJbVpX1IQ01MBn96f6s3SlKlRXjZR
kEUyX8p9mWKPqXhQj4ewGMHrlGr44ZFAZYvVr6Lz0lkK9c1d5HayuqPwhxFlIDus8oUh6xpPBj6s
1EgaS9FXkkLASMBsjLbWb+zODzGi1UI35pyKgxsQ3UnUfUWOkg8ui0hxlsWuYXKuEl938GklrUF0
V7wGhzbZPSQ+LduiPiUZjBv5HuyHzHx6WvwIWa44CntdL93hmPW3c65OMP/CRE53kzuFrjxzVSmc
xUq8+H1FYD4Lzwd7TzIqPxNRNYZ/WCsyXw00XGDVfAI6m/48XEYF4NeyH+Cc4szS4gilQbiSn2p8
/XS2J1BeltZwDzkVOCOSydzJuuy/HU8mG/wfTED1PbJo8klxkiA973QJ0/YJyAJLZen8BiQRgVWE
oZOM6nQlH5qRpBIDob4O40KaFnvvRMQlrwgrDmMAzsO9jQSW7lCjQ0AAVfzmKQYswGrugd2g7r8h
nnMEOroFe5e7AjJ5wRbAmalENw9dShGaHlMfuTZ2uX29Axr7U3TQjSo8gkaNnfSyPlXg0kU4UT5n
RhiE7yi2Eg0wjjWBe4gmaDIR6okrQPCGiToeHkQbBMBin89XWsyKa4lL5WT3vOqybyK2HxC6iUYD
Q6jGsUaHT4wWkxqQP6I6LdwgmvbwXXqSpJtb1uTAehRtFg8DkNifsn1PcyfP8g71PZBor5BPcvm7
VG6eF00tBsxZXlR8OcGdZia2NOUG5WLKA0s43u3B6TrLWeqLCYyH+je/y4wS94ej3tutFHKWFoux
VSXzgZNpzIvuDuYEAvcISLuM+Zd4cMAztnGYnSd+uRo026E4MgjlU6R4V+/R3UypOrzL8ZNgGoxC
16F4pQMhQ3duPwW1GqLqNhl8D/GVA1CtBbuVi0ypa7vkp0l2Gphai7KRkUbMXhiB8Wivy/yD+sFc
9xh/L6WInlTgGYJX5zYywiq3zEi9UzpxDfMos40iVDirLEuaQoOpePqp31hMdUjP0+z0TCfK7Urm
57MhQkhVqzUGETerpsEEa5BrJ5wBXzc85hNnfLkow4HljHEQgPDiG+IES8TTjf7P1l5rn9a985Zx
wBWwj3MvlQ62+0zqXuewp/5D8S5Dij1AdZ8Xt1lTvGeTOWmavqT48i13AcK7TUvH6L1jGau07pU9
yqFoz7D1MwYcSQbD3I/Wjqfe91HvMQ7Brkn/5FM/WIa5d+uat3WBf8fkIEwmJM3ENDekN+NEZ4ZY
QLzuxEgU3KkE/woVVA7siUEvnZHGBl8SJbJRoEyRiVFyecbcXeqX1B2X8ALSWJfDQg+p0pZSUczD
14hLfBmgqiVG7KrUeFm4O/FcLXBxSbxaFt7zesVQt5YSf3s7jWRhsMhmSuRsdOF6Rihe9+v0mFGb
yC9Um42IfHYWn57Q9T+nUTa6bIVg+PRnvukAKBQJNGQ2bWNJdfm2Q14PPg8KZjyjQaeLZmEw27vG
elXzxBY/uTKIV1N5H7B2vhyIQXikKCAErO+PlmGhKoGQTiIi/6c49q5c+GSjOe2uCOcUIhr57Iv4
0LO4ZUBobtD6gQlshJqtYL53YNZWnKWJKQUigaASj7xbFXm5hsoLLMm9dJHL4VjcNFxjwkGLV1Uj
CDWuM+vuDTi8ZdMCywHxmsX/eDEKthG7fEsqfIc7PRtYXILMw3LHRfx6B4I5jzhHOTX+6nc5yXrz
QtVmvcCxkW9PYg3IQTdJqKFOPOlRJAkDNTZqp3J/zwLpHvTLBI465TQwSuudQn9TpW1vJOZivfRc
EI7qtVcvVuangZczeqozQMk55FjovFRAwb0EG0f+GBZAqVRikwMrHn0my/sahmY2gF3dYC9aadPp
CDDb4DVCHkRc7gG8Vm3/R6O03bZoSK34U+RaZZSz+8yAG8gZq7ju47Kc4f+bGoe3Gg57z6jf5sWk
orfEilazEbr5JglorSuGC4JR5SVHvXgjXmuaEkQ/KcnH2IFS1XAX1Wqy1Zes18OA92gQLeFYTKQr
C+Nh9BjqF60bG/R0UGRYrfku9slEx4DtdaE7rDMeTKaYXL7HUD2Vsb+F50IDvTGSi/NHW+gP3f1A
Tntt7UG4hG3ZD8MeiquXQBPnrFdS+9cRMhrDaF341Pig5IM2pCbCHdByLn66Z5DuXyVrdmgJuTEF
PdMWNuVft7XZZd5rL50fsYFP5cymcutTtTQE1HjO89/otsz68b79N6Bo/fVI4LhS722PM41ziTqJ
j+kAnzXOof4Cm2ReYmZs5wI2dVRjNE4R9jwhoy8997sUpqIWgLDdgE4EOjK4tGOo1zEShO8jN/61
+PQcsRdn4pmrd9/CBiJA65t9iZk1CZ7wP/7yCFX3AZsUGuEpLYTuO4ihhcfBav59iYQ4bq9OTaA5
SUZEmlFvfeEiBAXMguraIWgZQC4Hgcz3hXWC6vxzNxy+Lygia+Zkg4/lWKENEDmw0mmnelBIPjcG
K1JkXaNkwM2+ZFsXy6nbhQrXqzPBGZIuyZQez1vjehRNvo6z2wg1x1k8ID544Ny0Pd6efVT06cVo
EDf89EuQV7K0cYianx5272OXQOiGwOFVsTLgxmiV/pQunpt2bkccDyH+mWo+kPWY+KeuAN7CbolU
scATD4td3C8sZMzVuelvzRiiCoDVD5M3glOiQmFkAB3ltseppJtvo5npKFKkiWItWboh9DMTjq0u
78HJp1uDpD486MfP9Iu7DHLNonjcE3eo6eU1xe2T5nprH+K85t+ZFSfTlRuZPFItLh/PmrO7zk6L
QK5VzkobTpC550XrT1GXQ51w0hTdXOblpXewLQKhbsP66lSlxFNfr102C0DD+SmMZY2pjs5adlCI
eG8hOTnnSa4ePwzMGQLmlVSi3n/H7QUYu2ZdP02JLCGY95ODI6GQFcsFNhN7ls0Qe+20T70+pjWl
c6V9/Hw9zHH47RAbjxvC/uqNmS24qlaUAHHgeo/FlHh+9Elri8ulMtHME/j8wugCm8y/nsSA+Osv
/zUx83XHyRzxoQA8U+xLKx7WPAdL6K7E9kndfFMPieKaCuqGi1pKVOwAAjd/8DeoNLtLpyJ8tO5Q
o9yhp4oBzo0o8f+Yfh0ME1moCvQfh+eAVwHirX6M0s2AAB1mKJ6ysWEPNuNae5HIbntrtQprc/Rr
cKRA/T9eT/5wsw03kxwCfN6NF8N0JrNfAt+YJE1oDgsniOQUKRCgxVTR/IChSz8Im36opU+6mPyF
ROgk83e6AlTSldEBpgpvRNkdM/pTwrcujr1hFmu9Kbv7gT3Cztynx9Q6Mm2Gh2nUgrLYBi4QNFY1
ZG1pAQxz2RBkEFZbQyBBSXSrmUmt04pkD68dr9Yblh0Xx9Px1yN0K5nQ+ot/XjFhgsNAuUAvL4F5
Rt/DagoRxUnaA8kvBsKsS7Al2Cr/+/H2bcDqW5OM8s7soFA20umhBHYgTPx8FQjJxTEnruTS0hIA
OVjyIC4hE+phkDW6eM3sYtfnTyBPZplKM6uCnMxSQy1bjF7I8I8Z0uydWQsGcmovcltxr9Kmkal4
ok79yKWvgyBOqmxPSYZslrWWqVQwWUEV1xNHCSuGZeUaZN1bnbzoqYU5+Gmi3PVSDQmvZ7se/S6C
pQ1moDWW/Jd2ucZJSaH/0+IR9o7U5hnlR03DmTdh7W3lXpgcQxEm9HP6tj6x31WhgA6qk4gepEQH
9MNHAdbfJ8O9WiBKHWkPD4QWA9VEYcSUpjlXVvB2n0CoB2Fg6rtWaZA0O5xDRl2edLOBeOT1PTW3
VtFcANlvNv1rKaXbMkVcCZOEBgt7mElBey/aHJj+Cf1jY79r166vJ2bltKppZO+MRKTtGYPabNXw
8K1jKOH2t955EjQn/Q2mIBUwW4zbI3fvgb8FdefF4zhk5LmyftMwYKC3e6QO42NzDDHHhpJAm4Yp
wmZpXCp/7cEIDTGc0s8CFVIkBihKIkix7NjwiSBdlrJqYOjSeCk7CMg9iBnTI3eaTXpk4zGzJ3xj
Q2z5G7+n7oZRauxksfbK7uD9XzSa1noiYCMDpex4A/GV9OgxSNiSIZiYejXVYyPVdcaNKm6bRtGs
DfFOM/v5FYr6GwjsmCuNFDzB9ble4pO6FHu5f7WaRKgTT50M419wqccbNQxgTVJ18MrOWDAtPEnU
zizTKTly9WCj03A1QU2chy4caSCdY4Dan4jruKnEBcG9an3z+8bVd0W92vpWrgVpwEzgiMKrZ9LV
bRz3hgSY7ducWWVVSp83NtnGmzUrknVo2zBk2ljyq5vduUHUi+vlIMJllc1AeWVjEuV4QoDRg1Sd
TDaLtmxeTNkRhflWmxRNzvknKbEYkTA78UZjzHGOe77VZq746wPsunGVeXwsUuDBupXJEO2/bb6L
lBvsHfl96lL/2ssXHpZG04FefSuMvBanmw3Nq+aHyxAnZE9Hid45tiSHkrnFgHz1YcljADC71HBF
bB9XvDfuMjknPWEB5A8MGT88XpXwCIrj4dYWoeaBJ7HNCirwoi6UBEihUMkaHf7xHLXn6oQcwPWR
KQO9QS0rfZ7LNvRWU+kLnHhah58DZmBiyQxVU+Er6XsSCspcKv+Of5p+zYkVi5ZxZ0CDi8B41/i0
9t7znMKYkYuP+XkYlIox2fc/7LudYWh1HT1GLKQHIMnbBaa/DllzNeL2FlXMa4BLVfp5nSddVtC7
gQnwLyjqtgqCa5gC333efhBWK/mD308DHTnrL9FeWQNjY9zu9nE5yzrKxX7KKsGIjts0iiW9MOL7
UF/1CZYyyGivDOJvs0TuYfzE5p8h7cLx6v1MLXNxfZNWKDAIyoGvkjJJP5bu1m9s48wS6X4IC0fE
o2OHyRifCCmuXL3rZ6qMDU7c3R+sq/bUS0obCbQqQ5ACvo4eEgnLV+8DhmYOGBs3t8sdoEMPPA5H
G06/GlYsTMWsdQTXMs9M+6mprdSLafqB1ljpYqi4I9lax3NCCpQC3VBPmmfhadn4dgW1ectldcUb
SMj+X5a9Jjejvd4WI7whQtCsBhl/1pRPRd6XhFFfot12PN0YI61ZcyYMvhkUAUkB8UJjdm3t04UI
Q6L43uCsc07a9NzLp5k9SdnLU1eChbaun3hlkvmLJdH6j3QRbig3icPL/UrsBMfXIBy4SIYSwk1M
3Gsyh8k5tqEyqIiCeGUifEnjh6GJ/TecFMU7f9XN3hjuGWOtvjEcuH0lCGX5qflStQmSv+gSZy1r
+zaAgBqKVNKPHI+NZVjqaFN3JwPXczXJB5LZDd7kyIELjMd7O91j17cdDcH26KX1mbu8UQPYhKZ5
nJGYx00MGTAi8kLGQogofKvqe9aCoIHF9hZlH9dwnC+4QwepTuERjGEnJAIMul+OT8WGZNXE/3vS
N4gZm5lC3WKlN20xOMzlGYXKlXgoIvfzn12NYE0sPR6Qyxd6fA0j+xBhhmwjS1GxYzqrTuFapicx
suu9jvhHhn6MNYit2B4p9ITIgUdsVdlzSYNjfQzb/aV68+frEMap3ro09ee/CzuqgQnl0XmE3JfG
h6lPdiVlUMFLIoIGBFJhCh3uMLiE1OIgJJWe79Ko8MPK2AqNhh1QMz9veFn6BIzjAEb33ge9Ha3z
wKKrgsvx1/yK6RlQ56nQUcGYfLNrHaoI/h6EyOy3o404WvJvsGMWN7kB2BOnvtCwxErwvMDqhZkO
HtJyZqlUhhiGrv/4JJ8sC4s73OCBqvAPNSYYGrwBN/T6n7FB0k9xU1BFq6rsRwjE4f3uSbIzeFiA
RV5iIYsLuBJRPDxFeOUlpEnVPK1F2hyj0gRCfk8XIrIv+xg7tSHY3+L47y1wY68vVSYPjNbBaLmN
bKrftWmKfOd8LzcEBF6x5UZp4NBgn4rkxuHCxPxFi8gWPWPhNPvN0kv4RuqwCM0G5IPqcbOh6EPR
jJcL7wZ1L+hZ1ewFkgD0Sq8JcYKNPM7oqaEu+ksFJi5lj6zyggc04pGiC7M2HqKMmMTaK0xYct8l
9j51jPJWBcYqwlz/1MU2BDtagClFz/kyfWkx0CRzV6D6I+Jpfrek1sa8VRqL/fNdavEfwlS/JpvC
ToGWBXEgJVvw+TKO0w3z6vO2w1Yi7grCOV/vjgQU1VrMyJGfjVsvVMO9VPJO6omjfq7tg0Yh9WHN
Gt294DFtRPhQVF3hmkpYb8r9ACTpbsTQ9yh3PYTjMIe84GcFNItCVU5+D+O4m6U4qHKse5yvyYML
nYh63MO4MQnAuNffrr+Z6sBOOXTL1pBa70y48XWSXxGAzImmrFCb68S5hR51wh4YqHS3C2veAtYQ
zqlTKcBVVZQ0JljYrnnsmgQBlLRiqNT00BMZTxYQyjKoeanfCOogKstRGShVPdF+we4+dd3gd73g
5nvDRTECRXFDKm1vi88YnHXqdw25zbwyjk0m0V3mbpEMEwiIV1PalDkb19Y+YHUR31K9/UsOx7ij
3Eh8pMNowZaRPhtXv13GYO5ZBJnlZmjUVCiXSsa/a65bG9i3Hvsw/4knTOeiqoxVLhS4008Wz2ul
j4mo68lfyzIsCtlPer5ktt5aiPOZEL1138tTGgPSV/M1GK7PFl2kWoyDpOYtiB0pGmGwJecqnvc8
7kdDPeF8mBQbe3arEM+j8zPR4mFp+IdlpDL2VZaVI0gNwny3zQjRJoKd4IYrKwK9tiyt7v5Pi1h7
OslZd6jhfnnbb2+5YLisYP3QLPMad6k2rr36mNc+hXaLp1NTdYXXKJBmujpzfueN7kJeJG92RzgA
BQGh/GemHF/dxf86KVdJMbj4zFn1+ZDnALLRzp2jg2oyoxgif5SLKF4eEI7qNOO+9TbGReUjjG96
8vDnL4wsWCKvz9p2LacSzQZ+/lBet2wM94jK8ceCdWmD0ELbvY/eU3MFyecVPbNprYS7anWM7QqI
H1G3QmTXb+xNtIcSPpvUisdDSfLTSpwxXxSOk1KPZqQtHXIusfAW0sRWUklURbOJ+zywP/h0oAJI
6D4Zg1q2asvJzkMVGXMKd33mXJSZmk5Q+2YU69TPoyYhqAiebDmJqfj791U89zaHJ4UfiuxFfWjx
ADjsSgS3FztSNpq0AakILVEglIng8VtDKNpFYb1R2QO39r2/uasuycRZHznbCB1AyzmYAel0EWKl
AOzqy4v8DLQ0MyDQYDPNBv9NPsymXNZkyfODrfprOEl9uuZdIaMBE6mO78L9VBU6AIdwU0GFD1oS
kq/3kUNpS97FKOnE5pDsz5h3QpywzRYwGBelUtZQeo7n1eS1NuzHKcjIh66Ps2SBHQa7WZtT3ngg
tXVI4ObH7xowh3BFU8ZY+LbHvfH8246xA8bNdQN15rIMRwZvnbXLKKAunF9YNYB53tjPXzhYMCpH
oZnmALAqU/VkMJLd3BsNTbszTNgsFobR44oNLTQRaNZ6NDkaJ8YvbdyYp14+vKv2neeollbMWjQa
3iYIwrVzEBESRHkdqgk6g+C74ZJJqjf2nmMcqwhRjyyGJxREiQ+krJfVBYGDkbTuCYQH8wu/AkmR
aJJjR5ZwKkkj1/Ol43aA8qh4wVqArqu72kAoHMiCE8y2Yvxp/kfz5nXTToDfTeA7pkRGyj81S97L
WDJ+mAmaFbC8/5dJwiUgeIpLbMRvpetQoelicvJRPgF9j3nTNWhaqI/JVVoPvhty2568j4ptv+ch
+KGZu6x4HShhnRPrKRKSuph7AXDkoQjVEE/GaiCBlucTCUyfySrMf9dTi+rEcWhot4OhKKvBuybK
qvmpBCG0uXnXvg0IPg1cxyWZWPWZ9xTBgKOYe97JBtCFFCO2uq2b2EAryG9eXxzRkQVNmMul2VSh
pPGpUWf3AwoefWpnrVofFdezR2wFY0ItdYxzSOPgXEC/er0Oz+9DikwFtE6sjmQK/e3t4lw5JIJA
icw/AFEnT1dVRSDDhMB5xSlTzhZ/0y69NYEPWJ1ucUA3APD/78tqEf44N6G7fcaSfb7vhvU2BfKM
2XqDMwewiefFPYld9wu7WDDLzoDCcRCFaDpbo296a0cDoTAbRJIqumrMAU/N8q0o4IuuRfI9NRTO
pAmjPMHH5A2sMZn1VfkR9fcroTtMBCZodf17robntScYst+eEezFt2oLFWvt/RGmXktF8g/+j/0e
qqeEPnUkgzq9gZVpY9PLC/RdAne9LxpXxza+sL3BbyBSNSuzPdodxfhov896WNlo/EYCGDddMfDr
w41x583iv0CFpxW+l1XuLHlqXLJhzvXnsrsFPQ66alGC79XKo3S+Oml+Hxl4gwrWaGJJ/lAJbFXa
YmYX3zGMcucWi9nMUqheZ1zCq6jE5Q66559+ZM+wlgIps7xtO+MCtz/Mv9aaXvkzyjezZqUz0Pou
FdyXhjjFzADhsUWTYBRO6cyX3ui/II7CtA21jYJAx3HniDgQeVj415Z0mA9Vip3xKT4cs2pt6Hwl
8NhG1ob4rrGdyyJuq3znjFScYDx9tqYn156Kka7G/yR99+7VpolDqfEzmyNz9fh0u25MwWXyEZ91
5gHYmWsCFZnJ9GKoXXmhPV+w6nGb3tBdjybta4SG3uI3gm9umNxV3cE3MM3ZF8KQH0y2auLnEWCY
wXM3n5S/ZMI3gV4Wcv0NPCMQo+9f1Dhazh1T5NxwcBTJ5BS2vFZw9sMO72TZMSJizfOHSCR5v4ra
Bwepv0lMdtZvG7YWdUWiYhIR2FmSnMP0BE/Locptinqnf/LMGiGv0frSnnD8KpReBVFvBc/Z11YL
YjZntdNhkrrKR004cIOiAW1H/eoN0ypLGaE6wDnMrIs5E9emuFzP0vkBfrfrZ8iSo2U7uJoAhTZ4
FT/bwDsyUj+2WxF8jfliczSAvw0KA7cPqc19+DXpkyJpHKQuSxIb0TF/Q9nH22i/Dk8jZRT3FdnA
ss0XHeX+I8SyVOYpjH4FeWaSdhz0pj5ICyb2H+g8KUqOohZq/XLG2P8GtU9ctoHET/+Z3AoE4VK6
2sgfTtKnnNV0PpjKt3LrhoVB7R9gFp4igZj1Jjt7/5gNnq3cjIU6Z7GJQGW6INAbBxFDiIZ05V0r
l8wxCeDr4QGhU96osl820FbDEZ9GJ9fcsMqUIlHA+fZpFZ2q2J6XsGQYKLIM2Zgi8+REF++YXVrw
3jkws3HW4wW3FEMXtZddrtSjbh5lOg2Kn1vIWiKWvVm09eSzqDUzxDHy2fcDgyvxA5hgbpMmR7FM
t66ELVZmUoBG7lgzqV10BN9pqj2TpghhBCqNmNhJhPTTx18RXm9VNQVw49iM4yqMYb6PbkVfFwxL
XOTYymQ0woqVheT6fgWy9mpvuXrPh7aXfeoBRC5o/AVS9mmbeHJoRThzVrWJ9q6HW3s/xhfdZ7/u
stsMnKrRK+KfmANE40pVNGMppr+YxxatTHj6VhsCy6/iQV/mxGAitcngqvPMgdASreskAHJIJEEJ
L5Ck2Ikw+3kswdXjz77DqCXO81Tjv5DKZN596CCW/FInU9ivZxmB4rL8Hdfhu7gjijvA2yBjCHRn
+xZuz51z28hyLlWKlmeDAmdGQGLOC4r7+Z1efxrgzAOuhQtmIGdUgB7IMi0F1twVaPHvoXtK74hV
vAFS2fk8CWm6M4rRC+HULQgc3TbYqJ7Oc1w2zhAyQxYHUyQDs9X+Zl9QCyY2aj0cQuXFFgDxCu1u
CMVVzbDcmDxWc13cGi5kHU3fTeevk4/1mQ2QFM1eTu/Ymp9wSH+X3lRsgoZrTkZ59bXzgD10XTwI
7YpLw8/VNynn/G9o/Q0DDSzlkn3dNEHh77H6h6UPhj7qJWK1XOZHw/dlfxr2jKG7Aw7FlPZIIlki
wtEmp98EHkwtbEhl3c7EAbhZ0BHVGt3LRS15OcyM5q0aToxBYEc/H9bA6vltNMKgWup7GFoyWzzS
PrQsed7SVdojLwSjm7fShsQtn6iRYr/HF721uPTyJVxr2rVQkkBPjxztsjIOJbrDjFXtA73As39/
SsajCPElnI3xi0vqyzMqRNox8YjTX5OFXKf4N5lXLeB8zBBM6tfafHAl9XoEomiNrqz7SRro1pm/
AN5irpgT9MagZ4GxJBIuMH6DjH5LFri5BfYiSSPgoonrhRtkjQ0lpuDwVg1ISdmidDHQs2fKaUg0
F84bjODLCLLTcOIa6yYbpKrYhGGAMNBR2uqV1cf8dorx9WXBK7dIfV7ZrSMs8u3L34MGDanAwCGE
Oa2Qofx3hBfjTxKI79vSt/yE3fcvOJjlsgBTect617eEi65JxFIT8vob6NpawJxzA1Ba1SbvKFdN
UtbEgbtqV+HFAR3lzzApMZ63feuScpmxArM/1a4CvSZdhqKdM7kOMzOymt02G4QkqtAvJTa7jfGo
8Gg7NdSAln8fEgc39C/oXTMO1V8yy7IJBUuTnFymU6Js976h7veI9V27QsM3vLJTA9nat6SjJrbX
AW6eGw3fqklYB8J+TO8anxWd8WRs6L9/EaRCYIdExXa+ggeHWCcwnrJd3ooAT7Qu6Y7Z8ZiTFwpQ
XWLFUpAudgN8BM8iQMxnaKig0zf0yzDTVtjUNMGews0OXXTlfpQfRF6IbQ2O759fi+wcAycyTL4p
sFoWnCUAjCrdPVCW5QFsYkkQB1IVxcTSN2YLQlI1jB6ebRW8T8uRoTBFM46e/UiofESlku5RXt3R
RuZKA2kNXCnwEEi9WsWlPnqUkTk/a1mr5HYzvQn5Z7wD1mjI3LJXzn3ZXggyJn0/7Z8N5+D2Wj5C
Etc0RLE1VCidAgbuCZXOPI7nmD876eL/tL2Mb9mgeuUGF6hhmopl3ldHGIaC02IvDr3C8qyWPA11
ntJORuBtzSyip1mRXxSX1oqW3ttVk1fxE73bXQRKyBYZZLYLvFbJ7QUKYcjKgiYj9houLyATyQUA
FTrUvtfyn90gumSw0gU6oKEnpuj5Pum5VGH+RrJYyCL0+Rr+0Wc0lv8bvsY4P9M5WnNuQO4QwMGM
SskrJbXpQQfSGEb8CiLpKxZnOcNPq/zx1uP767azQxnGhNQT1wCVPn2I1JgOs58RhU2+m31BE6n0
NjwE0WhUV42ovkDYmP5Y9+2sjZnKcWI1lwVFnxtOCkHW/lau9vYugOjvylRwYbEa5VMO6p+e2UPz
aYjpb0N7WH3L9kVdYwycoSpGsalq3he9pi2v/N0xWZeIbCh7kSuqlyfc2aBh5gdwe88e63y+LNNI
Q+cv4XtxApBYxEacJSeAdMkZxxpWipFPuZZrBqrFIiu+H2XpFzIXhdI2msL0a7Ya/299xdI7yV8m
lafqp9Kr4E5a2mEQvqf931l3hRpnTtDRhRkyHmVYNwCJmTqTPfijzEZddiHulzW3DkY0I45WYzh1
cOMg7CFPruB1xl3sFwCF3X0AC8ZtGM2+2keo1+bAFXy7Uv6Zs6Mg8Na5AKmB99z9re/n2y1yULwg
1CQCcfB0dixNs4sa4X+RoClWqSKjG3A2YfCd5oVnEigdeHh8snESMoU/gFdxA2NwVXjys6LasXAf
Z/I2n8kkkObF0bDpPyqk3BdKdgZ5cC3TtvWJJzGYLvCybE8nffUuxddFuXHiH20dufRso9N/UeQv
ImcxMGuZMmoJzWbre2g1tyRT2HyQcALC3KzNjN/kQVamUrIzLWnuyfvnk1UslfNjV5Oa6M0cg+Ul
hhar8m4jAlo6nFr91maBQyGR0IY1aqMIp2Gx5M4kqHoKPB+9LLGbF7MHf8y11QG+a82k76s+WyV6
DDxWXD0Y+y7QljEZd4ePpZpRUZdBUu/EAEdprLG6xIdRjub0j4w/JBb+I8ifAmuH0ShqX5XadNPm
b/8GQYy937ZMLL4h8gfSD0T9GV9cG82C0Mii6iZUm+yN5v19mgt3YoYA0vrH2ggIfTX/SVqsI7Ty
geHGCEkx1SLfsJDSGZlxm/vEKiCuQevsr86HnQhtojVDkh5jzVm2M98UnjSym4upA5ykcomvrOLP
vKODalzuAqaBHVSVWWNRbANtxvtKmW+e1L7tOY/N443Y2te2CJMbSDFGQNaICSV/5XovuKRbB8kg
eCT+d4NWMaHzqwDELBbga2TW974YieKMVaDuEtxEmUwZV5zkh+2KAVdWmDXINfyCkiLdq+VHRo36
7JnAEsa/A8cLhoOk7ybGqRHqLXv0cVQSn5MROmAn+GNRV192FoReEVqBeHgAvnF3BwICG/JafxM9
lvgI4eB4icenASQ213UMa1hq9+pFKXQaXUgmEj0c+xfXxMxiwY/z6Q+pcKVY4CS5dQuZidOzMoeo
/EMAJjBVTDm1tYyndt9QoyQxdFlxixRe2fibzBLeMrDdEjFbBmkpNRqxJ06eIXpx7y5/8ikrjQKk
pmIU8nTb7p/BrPf0dfOURlbxCTJDEtPrOFgtYer/VT78cZdyrtFpZJrBeOokMwcL+JYLKW294ENt
F+SxARXUAVMukKQgwpkIYpnVWDfLkkUOfB/an05veHeFQhLFv3IVfjTiUqERktn4+ECNzfqeJJXw
n+3OSYU5bSBRC1IdTg6miHAQo4Z4f2B41m9/nImK304bqiyZixgVHuQxl4rBNXBB/JNYmjoJIQoB
gAFTNSrq1JzqtjJbZV56DRMWxwKySe+bDVbC4lJ6SJjXiLgEI0GSW6w8M+hAGD5rWlsJIl1g2hz0
z2DsOnShdsdJINW9cUqWGCIkc0zVggFSBa/0UrRK3xcDvlFe0l03hoIFtd+KZx2EUb5URB5VwHi7
z7WlNUrprlD4LJ1ED23wVJaQ6VXGqze0QLKCkA1DNEfBgxFhuoIiXZJzk/2u7MhcjRlKO6uuO/44
8hfr7Oqt9zCgW2EUADjI7Ba+yXeNvqxY6Ao4rO8hBrV3z4draARgiXrmW5PKv7KCGRa1OKRw54Gw
uqBkh8vi2WdRv17uhVlnoVJdDH8Y4J+wb0UXfuFDyhx2UqSfc0ruVqjIl8PuicuGGW/44SWcrWtX
xE1sXyX3OMpIX2FrBQUCu6flh+cc60WPR9+vTFUGSwIDFyjPLQgGjnY++MMRoS6T3NS/EathTi7y
R2CYqquXR4TIyLJ7ziqz2AMNroyAzF8PUE9hObmzF0xUdMZiAnnAIn6lb90R5QC/eGQptEQs/qCJ
Zfs63s51JSmVg/ADR3E+jB4Lnv7Fsxd7+mRr3VyuASp8aGW6nROMxmtZ/SmHRoIpNP5TOEYuRTCm
hCjREBzknilmWOkMH2A1bvoEHA7GQLhQ1fBcY0MhRvcNPrJrwsMlzYAOCGUkP6/NaRf/t8wkfwHl
YHUDsXJVGmUTX5AQoTcNbUBh/MhO5nSnLTh93mzYGAQ8GD8v1x5KyKq/r5ZKXv7i9F2TcMKguSUv
CGss7zEMHJxAdgx6kKvQSwwwM99VOZDjNgqCt2KuesnE9yarhj8ZBd60M0v+9Scuo92XIxRU6QtX
aNt0GjQ0iVfmyHR8JbKjgg97AbusfS6ni8IsKaxfkpuC/tuagvACU/evu21Du0mDZ9L/JaX2e4Ml
IX+VA3Xa5bmd5Hd3xpJYsVRzeuGr99thqGy3nxcSmmWanxv5wirTuBvOIvaZ1kGJuZmgMkTU4glC
eFe2Z82q7I5HEeH5fQXJ7y1ksNsMqWPOkcfmiMBtPZp1OGMRPKcj76MIElqGtkuxWeXB1Hzl8uk3
49ObO0c/ggdHszqUhTKPDZ57HVyLG2y9/wa96OMwqmmWc+arffjUDSHlbPF2wTzj4YMEUWhLIPm/
5sNDwkD844om/S4ptW4pzcYbziCJaMYlZrSV8UJVj63eX43WTNoNDlw1rzGUtDRxZxftGaHoTnz9
4JbV4o+XQ7X2dnJps/5cCWED3uc1wa2ZpqO+D8ZyfAwh/lNHEhwJNgwDWkRoL0ke8QUu4VX+G01c
EDiXFW3jzpocsTbKWiNpkEQ/N5TihZBSFnL3kSVyWXBvVl0JqYv+0yUzjHct6yWYVTj3s8uHcC5B
TxBiMdXaj3SIMN4L75WUWl8RbIS1MOT68BeCFV47jyb9OevGA/y2l/1JLOQPx2b70FTntqfxExVv
Y9e3KuCWc5gYV0wPtruXKyblVTrb6N8nrg1y69Nyi3JHXEJsXfZearWax3mAlebgpGC7xspiIHUs
0c3S5rZf0zPHGsmE4Vh0sSss/afKep+eQwv/fI5pEWfYBv7x+tJFERGQsnmpkLf/h55ELbETr+7A
57LSy8LEyns5m6XeegaGwne6CLGUm9A95IKEEQNRVeTcO7TlA0HpiKnttyqBkTpqB+a2VZSuTR5+
sNHqf+UVVQSDEn/EDrToC3rA5NzUjn8JJuqp1/kMztO13ukT73fguQIUj11jMb8Gh8/3C8e1fxGs
IodSNyyQq+0ex7gUcyMQHgmgwQ9WTAFhketK/9DYZ9l5+EAI94xgGvY3AYF88l5AI9Wr+y6TzhHY
vbMZ3NhU71LHgl3WQMKefqLMc9wfFVWsMKYCsDV/+yUYBuLhcS3JPJjP0KEMW+wdPHPSStRipOqZ
hcT1jKRV1SM8bH/Sa6w/+3tOq/dwErKjEsRFntaM64TDNvydf1u4qHpuMXN17BEg5ZDCM53T+C8d
djZR4cgT46+dPcPsyGIC3kKTQsr6EGjVnRIrYVW38+ECnUoP6B9mwnCEtgqZOryVNIRP4rlwrOTP
Jd0+pIfxgqbnCG7UIB99iBuIOppnEKrqYj5wJlI6Shef2Uj2MK60XFkJus9Gfch7nOX3i8dZMGha
n70CM/htNZHriwrT5xxfGyci5Jr87upRRypqUMo7pARA9/53ZsTmttzAmV0Z7KBkyxcNPNLnOOAT
KZLm7XmqT7Bh41VPzQvAahNuyhjaj0kMWWWoMjzfUVwq+7Hz7o3bd2cRTFwryKE5NuMkYsDSwD/T
lVHtoRd3Lu0vN/NLktoLTHmrAF6WqD85IYO7bykQi5R1gvwuS8sNGensOJ00NrzwJWgJcKX/kxZt
ev4dFQzB6BzXppC/YAUiB6aAzVhPL9t23KCrer4loKJZyv+Qv4DF5z5JVCBVI/UoOQKjA41UZ8Q8
H7WZnOhY0iDMrZ1quP0Au5h+0JXz9BXjAxyD6IDGF+rOBo8x1ep1UfmjZDcivJ00iBkUvOAgcraa
e5xtGFq/+DTej6dq1tQI9AFFYUBL0Oh3BaZtnuJOUCq2uY29RKqCGGMq1JU3phGpsEJP38Zcn+Gg
XnEwD0SQup1vdL8SWAaOZ1NPWlyaQAbKeRwp0FtKne3NQ59HATniwotFrx31L1OEKdGUultcA3J7
l1se67mwDb1FdNbLR3LyWgWABXYgbLfjn0RPAhKFxW6TvLTudg6sY8/MZLlwfLzTRBYPftv5xX1U
xOHTwCdo6cQZvhpp481kmq8R9CaMEfMFBrZl7VidCZM8yEtsAW1deYenF5XDzYso/0IdQMeFYiRl
3yM3vkhthhEpq6agRoVs3ySN5MHKJb62TKGOV3b5135JHQcJ597+bxVpJFMkIVpy+qEUDZ2pc2iN
gAPBomntZIVFOQDuEDIGHDiXSQUKCrMGP2KyY6aTd9FM4aVINAnqQmQICEy6oIsj7/iBLXMfv5Jc
YvOIMnEdXZ1DF/gov+hE8HKuHEfi/IEFrX2j2NFHrIJOBsXQJk8uHB0STG7eVZ+9OpjQUfeDJDmc
7TuAcs6St4Vzynd+/ggNtAYf8A3IUHRSLFLwu+2DsDioRsb1gKf1hDwmiaO73uuhmTkseqs1AQvl
4ccuQnVAUGYur2Bly9TG342jNS0LZgxv0N+c3sUvnMUbzllAoCe4VcWj7203vJ3wM8r1I06uJhiJ
iYY+EjQDaDDVcIlFSgtOhvhtywfNXHyfNjRD42tPV69+B0StoBtivTIEkuD1kllcwrz9tvSlfO7u
CVuK5nV/qL1vKSvDL1L6vJ9CnKZwtWKl8hb/XBpDLtMaBVL+izdhsGBzJnLK8gtu8fHc48KyrP5Z
5+8s289bCOA210dBVEiz48sje66Prlwf1oxCD3WOr8DqMsqk/RJbHxVr/bGMUxw5n6uNMJN1U31t
+QhIfCV7pJBpjHbZQg2V092jeKsENGQPR3fE32vwTfvM1urHFmjR+iKtN1FXIxXEWIrAVCZeDj/4
DN5Ta5WvpOguJcVkyfbT6PALIeJoSS+ixBfz82o7ZvcAHnUq2clXr+wLytVToQ5XB1mFsmDk6+ni
uY/6HX1NVg9KaCaij+oQeaUVFHqKoDXjYcu5va0LgWyMnso9tFCcjcO+duqMJnKP4rlLO7r6fDy4
FyYpToEtal59IewWItYeKpicyodgZgYH8/INu6wW8dWBQ2oZAr+IfO3UwSxuovhIZonWjCtDg2gQ
IIOKkbOPiyIwo2/iluG0K5tr05R/wdCsObJz/SKiPvorUoIwVRtYjPQ/mCNCZ0xr/vUFBQ3m0arK
7Hzr7P0RObYMl1zpd7MuttYLQHrKnEwdxoXT1VLWKfsc6X57B6yG1g/wl3YMvD+DMFb0OxTGpn34
eYR7PbfW1hCNpCFYjahmQ+HyYNkPm23FrPMPY5g2BBpr6NLxJOAIb9NGOq2cBlCH0p1E6t4FOHQu
V9BQdmcaRYaMjk2s8BO6QA5W8NFMCrZBDPT0BL3UxR7RZ5JcYxyQeE+YwSeYvwjmiMYICC3GbmW5
OCVFs6oUHvXqpGqS+PomMjd6A9gDjzws9r65tv55UQa3ZFLBhUJH77YP4AwTohQfQSCiZnexYtG1
Az3IF8oHv3pYxRRmGnhVSjeNYNlEmXT+Tu5EIqslKza3d14S3rhBPF9k5GnUvDlzwsc7H/bH7+87
SNA0+sty35tFalhWo2jwKgFGegW/yQ8cVAP8eqn5yek0CI490so/Uyr5KX1D3USP7tEfI3OJsVyP
rlo5yxaq2DpA2+Iful0AnGWq9XzcexGUNFl6EpsOhiWqt4fdSjIdHlLuG0kid3HDEENjW4qO/WO8
ar5bastP0n5LwvpMG7k9KDLqedJpO0mencyrpX/vrE1BWXRKKOl/HqgxbnkqR7S8wY+0FgAdqmlR
BmFWAv8hEQj7DwvXj/6aN0FPa9todqul0igmaGz/zD9no/IhpYk/tEoEBLp/MHu3c8Bj+J3JOpqd
ztOSwSav34Q7yjh8wAKw4WMNqfARbKSXBq6nZgA7srpxb4wPLRrkWQ1YcX9GT1zmg4AfIJPuUozW
v1/lY8bo0NXjHI0i1kiqTPvRO2PhhNU5qcC25Xnww90VmLBIzSm/KaEkrEldiBtgaMClMdBpClv8
GTFg8xMk+GfL6lPQPF4i3dkSaaVTF9/Sswqx8X+5oiWh5wjtotAsIG/IDEMpN7q/rh65x+9aAneO
XjnmsxjC2X6LS77qCgFkIghk9c8QyObdM308aoBE48molDaajypVp4tQkOf0bU9Wy4xVNVul/6Ls
Lny1/myGqI9k8PG+t1twLgsbFfBFXXkDldpG1YiPQ1oxV44f1xwMrPX8qdkbPq9QHElnSpRdsF7k
GIXSzczqTSHDlhY2NpiCNgZcZMh5S+iIhEVBHRj6sUudkbpA29p8sVhglBKTFKyE0ulb4UnAivNW
SPgrjzQvYGVRrMgfFfq4/wFlO7MEBlQ6Kqs3nJ7usbWCLnxO2MrZThbjDN0hQZjmat/img2tUFD+
JgzM9+JWgp/GFs09DZUxKlv/5lLyWhSPwdBftSjmZjUad/USMj9pD7j1diZC9Mj8ABdV6cJ2ScDn
AacZC4f4ikQ74cbjF2F/+A7HPopL2IuUpivg3dgaP9rS6GEf5j8tBHeAwCCmqODFxStKdIur1bdN
7FNufbqr6c0GrNQYygGuF6+lRC1VY3wXn4kCbcviYBKDdcsNzhOx6xxIPhIMnOVKcEZVlnGFmSiv
0a2XwVyi9BzXTCYSXfhJZQa10QvhA31UqROzffr/LnaqgT8cCqf8ZKemXMTNtBj1lFzEMFIvLPih
UlIae00z1enfMvhuXE2aJjTZy3ZMXPQn46K9E9CK1iw9nP+GgQng4bmT5QTmsX/fRToQerpAGzpB
bJrCR/v9qKPjXa1s/zECJ3RuAA/Oe+BKBUVixuLEzVzHqHNveNQ9lfcm1bcRnLJX5MWt5vOBvS/j
eFit44556ZhhZgB0E88YE3upTaqrnRtg91LuHmaPumkhFyMBFUBSReebCNKv0IIcwqNKaVMlKO4u
nXBz4rxmiloAO9GyDrzNiCLAZXImQo+jwS76r/QAyDzGClBX7ttXnPjFFZ04VofQyxMgt8c13VNY
AURx0gBSIHy3kAf+QumcbZUjmthr4fwGFaHCdnlBQPhVPmHGaygyF7uBBT3LmDOagcYqBG+lSN4j
bq+D+UXZ93x8LYiKyWnnHR+rbjNxGTHlsqO7We/lYrZDPUSlzgwxY+XZu6Gx5h3sTpoFBxc1gnCc
DelspIu9+J1IOO4/CX11UTeT6F61jkEDCKMpaEHLILfG5F10dhiyKmBqPXUSKSlq7mnXvg9m2eK/
owWpjEl0KoGy34XW2aSyu8cVwYakgD0P8pxqfiEK9kzhRleVyVF+HhDUJY4T51GwmpERDzDYayA8
1sZa6VyW6mdCT9HBHcl+0OPn7DG/ook75wSmReX8JjokJGpId7/kS25aY6YKRXBCejhRXriCVBuf
x3s6rDYgmK6z9kqDqmKuibMqxUDPruZDkVBxYb3mR82HEkiQJf2RLRzylCcZQKNEwn7I
`protect end_protected
