`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kOs6tXJzQbaly6q1YmMa5yYN9ESbbI4TG7psRElo+D3cUANPdAkUaP11Rtv6aQHEb2T1YtO9U+cF
QayzFykWaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kpFYo8t+C5u1/YR4XqHEKItFVPkWlU8IwR+gPeKPSzKkec37IKe9K18s1a5/cEFm7diJTPXL7HF0
VohSaTQD/umF1kygcF2dRUpCZFxiW+tRJV/6A5p15sfIau6KYPTJ99Qood+MhSdY8SDBgJltxPv+
mPAUHnNV6iJTo40YZTA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nuHtvxJNEzsHpCj0HTDVYIIPhkVs3FpqR86RYOR+Lgls4vDSETQdcjLkJffsedVITnrjzagoC6OU
ZYtqIhFE+nAuFdTu+Nfeq0/XsIyypKDERqipYVA5oKT4O6e0B5f7WDKVLUdIXmxqGlNYI3n7xunu
KlmuCo/9Vx1SdRi2srcsPh7NAch5XDhhsoudnD3wThbSF8G6K9fDtg4OHGtZ1p0A9+kCEFOp6J3j
SDkl9VMjNadLGP8mDeN3Fxx3Q4QwBQclUhLnMg0EtEcKXjDtNvVjIRk9z41mT0ZkvwYpgMo0iEvl
2bB9KT6yQTFz8UeN2E2CGOaQRVi37eKhp+oVbA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BU698lf6zciIHkn7xp8lnUJyUCWQ0HaTNdk1/2z1r0hZZ2nF2bvMM7ti+v39w6AcGQwSTYVLbJgJ
MTQ3HSB+aKIwEwGoSPoWpUt78ixT6W8zYoLF9wlMTaeLUNOZ3MOViMI4RSZfgmfGn1xP8cG6lJWc
Ss0/U0d6OievndqJWLQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LIY0j2vauyVeQj3uiBvFvvm8E16QcWzsNq85IRlylxI6WJVeAqbjJ5OQYvJCBd0ynHfPWSkWL8Pu
cLuATqKC5J618+iWZIZpqlH3QDcCQT/k6zYzz0TWv7i0LLV+EftpiWlSVXka5RewWs0n5z0s0vmT
PPVkUjb1doz4k/HgJ1s81qAUT3zd+t38rGj7pUDz7LL8tzGsO2VhuAcS4TTIjIiRLaPZlyIBSrNU
RRDEgRXOXwNJqdKCAQ4/By1550ciPmC71ZUGFRTVnx2IqYfaKhJjEoNX+pHMIsNx034TrzeTz78k
EDcVF3CuWM+LXcdtLj3VkbgGr8yVX5oMz2u+aA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
JOBK7m0ZMyJmKPrn+jaU4o17VLkIHF87XExBPEfB83cxsfmR+9gq/XFR/tPz265SULCoSChqXHgA
DXcJdA5Pgn9ora7IswIK+s/ZTpZc++NAEPcKxo5J9QC/0ihqzakOUvfTMctV9YPEyX9LfV2OOHY3
Lqoh4nPdnxLJBD8Dvbob+zUFGVqqyikCablzsZXF0Z6rlH9V5slFeJSnEAGd1LEKQMA3bYm0Pqlt
w8Hj1IvG21ijlsyFFqcdi8knnCKhnBRqIob4bsNNTzeiXB0fmVS4m3rg+MKw6nS9Q3lRiI0iujAJ
yd4S0KsnRBAV2GxNOq91Yr5xTSEXx1iffvN6wYXmbtZ5BSSk94vX7V1UoQkN8PRhdjTDPqmFrOxb
Sy4Ufj852WGbYgeWz6nj/6702yZrY5DRBUkYaimi0p8/zn3ihNbmY4aTDFemYVl9gviyqM4cvCUX
XgonO7aN2Y0ZQ39JsqmKUI5HGBaMA1LlGULif461pEZuJBLsoUPjmy418LIccwa00KHxMJ7IcetV
SF9mNPVIiC8twZUHtDCWe84k39mdYoVD8ddhgDN9UYTgdlCTS83e7LYtC9cUz65qV3WoUf9sbHbf
wrsTO1pDRTLfAGxLAtLg3leUDqRxceEtCWg2dfMMXOB72AHYDv98XT+Yll3b3KmOTIEsezpu8Dl6
U/TK4IpzeD1Zlum6GaEx+wh4jBVvcv5ojo0fuvr6LuQ5udgSAqmZzgJQZvC887V/inzEsDT270rb
Qgqypl+PXfY+rya/AaKuz/pQDQRKgXla6fp1bQAbECBBXPJx1RmrikLFqgpw6VrSXSP/BZPB9MLi
LAY+bpegmr0BHmtRRuRfXxY55YA247ALcZtO5fWZLEcmXfIuAeYuWQnwbN44+ZKLn54zj6U3B0DP
njoxc1wdpHOpfs4UWUNV0h15XY8r7pJ1+/NTn0ve7Zn4GxmSMq6q+y8GHSDYn8M3qPZuDSMcqbUj
08sreI8NdEKsBGY+9UgZJEQbvmFq2h6BIVTPLWwsA2wYcaNhdLwjG0ruVROXkZZHr2dEe2MOdDXm
Vl3bVXgaahNVJV2yR6IwEkQeX6v4yClKea3NHkq+DPJCRzN5inqk8b+Q/ggULOplIcxDiYnPq8B7
o6eVO10LsCPGuCkAuDEdTRS0cK3fuBquRHbNboSZxDGb9l+Ps4acrxPzZoRkbrxfT8iSC7gbVZkb
oO9VQohnY9UHDPHIe03UkKb4oU1kuDLI46SrzLIcRztLMHyG28cJy1tCQP59OKoO631VPASx8hGp
G4ieRgEs69w4GUyHADEt7RWYTBRKVIWzx2v+UHcH5yE72qevxjOtGcJsKAbqIbV3o623znrq+CGL
cf4kutlVJytqnOGEcYpLjgvH6XWJ2Oa74K2mA7ew1UZy8NtXDYcpbm5N76pAWIE92cSGyaK6DVbw
Y8BHxtS9jQmmOMCTMGaEnz+wVtp7hO6TWTA/v05siEK2sFKpyV6NiklwLko343x6AFMWD7pT4hV3
18HMWRN6/lDUVnLtS/72PNZ9ABIiqbXJ7dNWxneqkDHaBYBnznqQvjfw6Q/CgZzzY2+Ww4fdmF6C
yKHFw90aRAQLYe5deq2ukiptLFbsJtswC900+gHVDdNf7AHmqk/ZfZsN2kTk1N8o42qQ7dIgP4Lp
EJ2A+nEmQbLHR1c49gtYNAK92bmMcqRkmGtQ4CAh2pyCGWPXabT+Bas1zwiFtRJzgNo2+lLSfj0D
3h9ABFt4rQGuNqBhAHwP3U9IdQAsjahjmpOMgfjwNc/afIJ7nNXhhkuIDYRoca638711p09i3SYq
DJmVuJQhHanEWlfES1I4znawVGaZQcF3W8XLpllwfBAeoNbT1cF6M9KiJCDXXfLJ8SZMM3467qpP
CeSqaY/I2GNKQZQQNqEnKblWFHHZbrSQimJJZh59lCpo3iiTgBLTziH13nHXT+nxwLezxauGB8zi
wM0Gea2FZdwUiVjtKCmsGkGsNMN7biSiaKd6GcpWnWkH/LlXNtAhnFIVFDEfOZFrnZ33oT5qu2va
Ww5BlfKlqdxV0uQ4SvFMYGHVQjTZnxmgxHaFRGsBCVmdbZJlLS5TJdC/YbvdxIOE338BhXniBxrq
VkVFZTU+n/pXBgiCEt09VsCzlzScmTR7wu5cc/VMVEd6XeKHUoURMbULPh5l8q7qekHDmKkC8IJ4
lGPNI2DT3GOvE/gHcZIcJZUTvE8FFRqb1rS3Hbdw/m3eQZgDEl1zNckxY+aR4J3udpoU8wE+X/+T
FvXNC3nluq1/qPmpshVizSua8LnK33lraVGI4BrVQpZZb2W0DK/iMcLV9GXce7kB78vYoqcYdrSv
9AzdGaG15ii5ri86Z/21Xz5T+3mzQZVvQ5fd42bnhIO8LFWEkJVgnRNmym7SRIHGNciaEF6U3Ymt
bdo9C+q0iSLD2UE6wiEk4+ClK6uibGKZC+usuZ7hJQUqByWgOB9IZ6zG2GdcheYOp8Iaz2iN8UNG
H4rKCFbKO0AsAY3n3jjU93+3airEAONkwT1HhXc0WXKzZPabikR890xwV6uI1Q0zzYeDFDhYxLut
bndk0aQFfz7EKTHF2YbxszuVE0LLUWtzNmSfRo8b/Q0aymW5jzmB6opZ2WV2NsI1yPQD0gQgjlIo
zVbPkMy3UstslI3xa8InyeQFoCV+U9p9Jy8d/KNwalWJORskCkx4YkrJYZdFkMQd7l7mvos3o7i1
ADKzwiaC837tPbyDDr6nAL+gjwfgfmz/z+kJMpRZoreXdghhgpuPs0poqXS6ByD2Q7ESDNK9nLmw
BMw2ojA0suEJlaahSOjm6YcWWGFvnRZ2sMajDUtlOAl7O6f/qHY98Ga2RoL7w8AROoJUXFGcJdQV
ryDILoRxtTup2GIGamtKN31QAJqzZkgumHEszF/XnqvK7tRW711BrL0cMc5jPXJtXuAajClY86kH
Tg9RpbF9WsVtt9ojuVUu8oXMD1XIVja1n5tcmdieFonmHjrw+VZoxNaAtZm0Zaa8mIj8D4WytMNi
hFpJn26D/TMp2NQIwwoFJq13xLJQM0PNHuwhcl0Z/YoEZTOxFznxMbexTKqf+jG9PZpSn7cX7pxu
I0OiDaneAeR5k4tprNSc3zTYsRHUEFshHt8UJ3ZjJPv5GGk9UH4YPRFXcHSyrPOCUy8d2VMkfr/m
CnykqB97h2OIQje79Ivghv1L4verQqWaSN1qjJ3VJpijTqsraEiZ8AvDzkL8qeBMHrPHnsJLF85U
ejjp6PkwnziSzKU7LYggjrtO8WJzx17hj1qUI/sojRhZ7JsQ2nq36oshsrMoX9dKJx7++jjaYZQR
W0aH24uocxjz2mWs25X4k1pfUfVOkavrVVJE5CQerkexvoUjlsEQCkCP4g3uAV1r7F0kYIqoufmc
4QfOUjTPKfwLde1o0sUvAouaDF/rsxTEsqoB6ZBdrUsXELTd6LH2olGrRvPID6shkYAaLa2zK1yB
vnbhKTKzYp0GjFcodnXS3UGrk6RoFMdJkNQtvPztr5xpxVZANAKEZHrJd1ysbDtRb7FViwnz9zm6
t7aG1t9M/3XeRcwOsi7MG6qEtaS4YYVEyAWzTcdREcy6Xh//hDi4sNe46R796TqhgdNs8cTnDnB9
lttG9rwkgpLF1tNz7PZCyQDcTlrpHRWXFb2KuePG9jZln2QTm59jkH4cNfExRIKXrNKPs10GoILu
Zhsv3pH2ZNdOzNPGFW7/n1/chAciYWuom4b8/PLSwrCtF2+AhDrbjM6wffxeUH1LxuOYppxBnMFS
phHF9xF+jf0bjapBAksyAziycsV4IxtmDy4L3sYkKvVoOk8YDWfGYm+FNtNgqICdvK6L+kXn36u7
5jhHG5yCIf4OcBuG3bMq9G3WmgpFsmtQ5eX65d39jNTsk1puU7wpZ3bAw8dhpX9H3pSP7JT7ndZA
c6Q6Sy094Abk9GtwQc6+JbhorM9hSyEhu6uffg0oXcJare+ub9YOsMPcaqJcuNPbPfHo4AjSTJrr
zvBHwBr2DJOS91fqRN3NnYlAVzI7gvvdroLUWYbEtGTncCUQucbR/nH8zmCiRz9Naqx2XUgRJka4
bjxlCFK/x6JnzhSBPPgF3Q7gXulmsgAbOTK3N+8ofvw1QHaEjJ2CfeKLNx7e+xu36Oj5SZoevqC2
KMdAcu92xix79O1veZLA1jXus1HhMjG3LWGSQCPsFM8BqVR1kFVg1HcejoI1m1girO4UtN8A16PO
usa1TqDtfU3zNlyeCgPGcLQvyLse6kdKJqfDMM2K8UiyGUJ7GvSyNjYR02R3Q6XPKHTdjgO58Eja
3GF2N78t2WsU4pSgSFZQ+varhGlb0pLHRdFGERvSqPs4sM9ds9WBkXuWPUH4mBE00mpnV7B2VlLU
53o0ZZMQs+clV5SLZC65PF9mcpBD932smZ6x37DkBkEcX2Jdm0TJGCWVIWV6bdbFYnc1H9JyOlrD
o746ei4GTqtP1L1Co07F0zD3PPB9nSPIpogwgNq8vijcB0eiEh2Tw3taZxy7o8GGFb3bh/jm3TQh
C00rFYQoZFNug+vvnQs466avCQFkxuzxD2CpPaY3atny55eIEsbuv8Ga+bmEAC4BxtM7OetRvCuT
PPgycXtaMcsDbZ8PK4FdcI2Js5uV54GJhcICbGRsXd8PBSCWvMZSrWZkywql04Wb71LrpUZoRLVi
l7Jeemm/AObsci2Ki/9lO0CGfNR+qEN8/IXyUe585XhxKrkOBQPchhPEWNGJDk+XRbSKQA7v5FdU
NGczWGeSjZAP3yfRaOKa3MrFMxjiUg+AFnmNes4gB7DtLDccp2qX/edSDIxT+28FHFME6dqroXLi
pbrO/WFlyowooEE2luYeAf7TpiX8m7YcXdf5eZlc85wSHxAaLquObf+bQ1azTJ/LGjSzX773eUay
rAq1ug1QYXo3uBWuV2nXDVfEnbqiwoGJwIvPq2YC0IhlQfXopwy6MftAP6Vckk8RUEtFRye9Jrpe
DYJP32OEikKv3inXOhXQ3hNHK1dQvtR+4dwsT8j1eNwLp4BxMKas4Ix1q9Zo1oQbtN4rsSG8JE9H
atnB1fYhk3rEYsi2G0rm8CeUyARtS0fxmOgn4/EF7p+XEE+lvb6tiNlyiaQWSn5Vfx5dEJmUNzke
K3ahg1oqPl4NWs6IYX0nUm0014jc1KPveu5oSnFf88LrkTX1DyDO7lCR7E+aPDVa46eTtrRydMyX
qrKE+QoGTDXIWSKXozVKOlZJmFGFcr9oMbT3S5famoRaTfpFXV2CmGSFpxHR7VmrJc9aqJcmL2e4
c0NIAFcgUQL90B9LLxMV9kmNZ2jq7/wL3f8qATi9lrvn+hCcH6xCdENfiZD9J5Ev0rEZHENX37j+
VGpTRQkmwLDkZwsAADyS+YFTqrfL/QLoQmtq5ixCNMdzYgfxEgkFISqk7q61e14TwuE2Mb3GXr7C
LxH25ocL6mZEpFL65fXGz5J9jdiw997rFJFZMXx3LKeFFGoWkbcbfji/Um4Jsr3sqUErFrYlz1iW
GEXzipmGBmQ/Rb0WbrxKgg47kxQBAtu1YZ2Ch2UOjB+qalxGcAY7eBC83c7HWPw1FHunakxjb1MN
X1qLP+a1IAZfJonx/p7MpPzb1cl7nG7WWwLmUAKNf8nsH1umyDM=
`protect end_protected
