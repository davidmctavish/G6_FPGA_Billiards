`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LGjg5Z0niYiPQov/sZ8VzReH/zxXabKdsZ+0uw6HN9LQQoRofH/3Tjnkm8Fg0Q8DQxl2mUGCpfnS
4TeMFabfSw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A9Ju626SJ0dJbCkZA+fMWl/An98X+j0zRNbChgaHotd1SbYSn9cogqLRewLNtMz9rd7V5Y927+6O
Yn3BK73P7H5IG1R9XgewL4WuOH0cjcMl/+WnQsykU39o+idh35cRQFzLhWAAgGXIU1CkUKZj7VRd
Yb4V0/deAvI4y8Oyblk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JBNYHaRgM6pJodpGK1yNswZoP1lN9C0P80MsqZ/R5AaAVXauuTF+PnoxEm/vV2pe5CI+43+ChwsI
OgVN9FWS0jRL6SN+wyaK1w81P7wmNPLZMV84Acmo1B2neze+TBJJxFzeD7YOVshJmxRSUPEeQLcD
tMMxahWnm2+mNQ7cMpin0oxwpDJQtrqx2iCnUSV7g/i96u+y+ZUj70jsmKyYuI4CQMhfum2h3s2z
FVC9UjQQUaLSkmImRTyNjceV+Miq+yHEE3rr9q4RPCV1w8ofq/dBbnw4h5ZqgJyb17FsK2bf0wPR
Lqmdi8vTIKokMxb9uzX+N4Wia3jq7JfQS4UVQg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DUg4hze5lHoRkqBO2aABu+BVS/bhHlMets8Gj0c0Cwko+nlrbmrXmW0+1a2Nj1ox1lzE+O3hlZj3
rOAQURNlKnXHIGYd7JrS4csvCICLWLBzQySpWdbuc52I1J7rg8RCOuSG854Ej3zm+o1vnv2EGtIu
CJQKsOQcLwmqfL24uHk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RoRO+UqATC5A1R67ifWnVp2zzscILREvCjkcVyQmhFkBsqBm1Dd0WBVkrR/sFQN3B9XtIIrHRsN4
dJ0x7ejdOhaoKkDLmLWUuXeT8zCIvykNIEURs4Lpuaw2JsX7KnywQlhe8qKYzbXkTS4rljUihp1s
2ywd4GIUzhsgJSxWX4IzulMZm5UgFLogFfhxdK/WgRIysiB04IcVa21ktSFOuIzRjb213Y81CEc/
nR5VH+J3ZtDD9c0tG60Qb8WQLQ9WtKD6aoHnAs7FXBOcKqjTOvJcyTUQtglZoMhRSWeiJHKrbNkp
gOYW+TMFBCtKxZGpv8mH+WyXIPlRwnd59zQ0kA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25312)
`protect data_block
YUCvoiKDAMI23pwpChmz5eT2FUwwC6pRAHOL+mgH6bRPw4e/Yy89QxRnNLEyHVPCI8PouiBiLKnU
JyMCOmgBKF8Y1ogE53g48oUPhsfzERRkWZgkm+I7yQqEFb2UW7R/hQHeCRdHKorResDU9Zy/Qzeg
x/GNxgBbnZ2QpT1FrD1pKmzspJ//PyFP9201X3zseOer/lkInBRJ21udSLcPRlbnrI62O1bm1T0G
w3PWBpSnJpRWPetD3riMMCYQFvm2l+G4TG/zl5OvOETtpkt4yw8E67h//DaaQ5ZUPIpCq9eMON3/
y3GNCvYDakoVvzl/Enk6zCQASIbpmnop8rymI4xqKv4IH0kv5S1x8sabIXk21oQS8JaPhAIhusx6
Wj4dwkftiteVXP8yj80PcdwJb/LBAL6omdsKUqF6ZxkJXTrHvQXDNsqVVDZ9Xmbw8z/fReOMjX3U
XuUPpXqN7suASRzI76+q87wmlTShtYSdx1d7kWzr0kgj+nlJh0KLNqVCPK4e5CRdfjBuSRW45PKj
VErMnAz0NPIhwHLTLrjzDFMBKUDY16Y7H9etAEFzaXBMOG1uONV57oeCbGs43qCGdHY7A5ux2+U9
W2Tr2xlvraRbxUy2irKrxvd64G5v/hbesD0jszFqmb3qDCr6TV4M9SNEePUB5EqIcOvdiDSxIc19
XX1WIXGu72Hg8XFrH1In4GxaSbyZ3E3zAKLTob5Un3RWTvSg3iI1UtWyWtXABnoNTOixJklo7F+z
qxWqcVuB3dljYTgZmx6+cEul2zLHCZK3AJbpJGl3BTtzNjpe4ujGTyEW9IdEr+E07dmbHvxllTAe
v7LXVHW9pUBJm/gq0oNvdjXVSTghVQ2C4KvdW3zgftlnjuTIfCfTxSlvowFp3Z58NalBWP8UeKGK
82xZv+blQFJQQeFUwe1fQRVLI+ok3fb9jnYGrWe8PImYJYBQvgs0dfLVvHTktyMKlXup6XvUQF5I
TthbgtG329AA4z2dQ8FJVLh+w22UekqnSEekX7lA21SCUzDbF3iEI1CtDsaiYaYBMDwkqEWSq4FY
kuzh1bbl18R6uZqA1T+ISxrwas7RjlMeie4gMbJ37YGDDoAMbJdRp1nJfxgCJH05oLu6xKjpMWlc
AID4+2r5rmNHFw53erhGGbCoFC+7MfTeW4SUNs64ZwlPNgMmehRUALeGcS3aePxf41Lw4WCMc/NO
yKzaond896cMpAGbY+2fYvVZyeAwAf6yJN7cqQWuwCVsPrdD054Ct/K/d70hclUaOoZXYJHPTGE6
00RcbUf35hxXp4T+WpQh0xb7by8zs52voyYEthDhssfGdFbjaIx5jkT/1oK7nv7jB5GSbtJSlmdr
/9ZcomUzRQVKfrVdH/tTCIEaBHNwuYNswvyfI9nKblYGasDEDMI2Xpy946EkeFeF4z73TJlAlbKF
unzWRsBeWkDoz37ORdwluc+ZLT7vIuWGk+zImR/C5X5G+rJBl8opPG2ePtPWsJsTKbg9t6j6Y7+d
5JKUpPD/zdpoCfkQ42If49/DUzNzbciE+m/+yENPHr13YKdTumNLpp4RywVrz8A4tIrhNDrqUVHU
VOjTAXK7YZ0YvJdcxrTro1UikF37szd7iOwC359qIZbLj2c9KtoOx9yaTDMDSohzBatve/2nl4VU
Q01XxDswPOvUz48c0Gqh6l/tthFiCNYK2yo4lmnSSwrrrsVyBqhUIpXf3RMWF5HtazrGn5sXz/0g
Jt24C8LEhxjgdx3fn+fZc/GO3zY6qMh4a2mf3wiuqDryScP+09AEp136/eklASL0/qZTsvtE10M9
UgufEOBDtwZf3uTnT5ObLMoNZsD+QwhSt9CI4bnUml2nV354RgajBNA+2ozuUJWSHEnc+bX+pkv4
Zw8eouYDbej8HBTSRJy8XC9nWgp98xVHcbU+xUKepmEd9WT+zVSBk8onm41kZgUCDAQLy8eQ8KA9
xIfGNB9wwJBwb0kzF4lc2IxHilHHORWsvynA8p2BjVPuLbf9g9qgo4saBsyH78/VESP1O1YMRSlh
32tCb7YBD1qKZOmAdJ9pQPN17ODZGTd2hKU960mqbrWUz3NwnXe7mFpNnqqrxI0XTFKjyFZZce42
gEkHs27Q4DKP5tliTimzGmEBgBS3B/NxvQwLYOAxH8wkEZ4IN8agLBBaotZ5vV1Fmu4HgDIvu25U
VnR/4radYYVh0xo/rBz29dFwhQdZkB4cIoYA2DOtMaKRIEC/vISS7f8/QL3yOO5PKo2OxgDwU2ly
uRGTNBX3pidgaIok4/p6umaD4Ym4O0cFgjXIEBCVucRNyPVJysO+tvQuNax0yUs7kT5gqklr7vhV
08KOCgzLBixHzMzglaFeXwygpH9s9dr0fFaqYO34SUsRsaG/UmEgGySAakzhHUFha/15uZViWWEP
2ErK/PKyX8a2unY7Oi+epMC0QnFL9HP5xYjnv2NV8KYC5r24HqarrQ2nUp3fGihzIe/e43+35ZNV
Xw2yDvn96XHZif3rHWSrVUHGBo1ewxOqIf/4ilr2zjLSRp1ECiONx0UGFAl4CY60A52vzqZ4TZrz
f5AHz88WOJdQ9dymw0KUVGdocI+7ddJemW/UugxWuF69hrHEH0GDqHO55fvHHfoQ8PlgDpS/exfq
nFP/Ts/pZa5QCEQwhFsM1ujq32mIpew4XXFLE57FzQlEcLEBamXVUlCJNcsGJn2KMhXOvYRe9RSa
AXIIOznXsEnYb6715a9K8Ua9uXNynFSKj/hp/rzq30nqHEaEo00UCZSTUdKns5clTYMDGK7uwO4p
U7X/NGfj8XGkuzEfJWIffIQ4CPOkLteLpUvcVwcrdcu4qYzazH1NLMhJSGb98z2LcrfcNXJEAfFR
xGTl2r9vbNfA/XZCqDp1r2YtjDXle+16bFCZECZ32V3mV6vZwc9s8VHa7ZRaReAEWWnIfB7SJCuL
nt8xKJcOg3vLgVFne2sFoU1eKxCC2hkiS/ZOdqdAVPesVB1fMEskbai8cbwgTE7abLEynwFYtCrM
+0/6BlzKmgxQ3ngkmG3Y1uF5za5RbhfnX6nyL70rOWEEpWzs0gGMG8k15mpDcw015JWCScU63vdf
/ZPmJzPBB9fSK/jfcTiRJKnik3OEBXY72Jp7Xc7eytzxpOmAtPwHVDNOXhS8LVDmlLnv3fPFMvn8
v+AEgk+quj2Sm1TLb4ULMM3tTinqLYB/ihLCB2NwCAGxrcPAzQLhxGELXE2IMWrDEwtVoCQEy7pO
pjXnyfAGLpEaZf7rHJy8+26ICEh7zSTfdVBB/Vd4D7eEgeDjwYlTZugSMC5d1CAxzl710fZkAsw9
U8UuMpAWVYhaOFUWEp5zJ1jPNM+7mWERhXGH8Uk3C4GuIdI9SHmlFlptLalAZuztIuhv4KbIhcpg
olUue/9aK5MNhe9/H6rdtIKxstp9eSR/jwDOaZLW0QxKCvb3XvpR6lFhlkb9LdCIdqZs2VmuRe96
r7SxydXJCCkosLzKRn1bQ4UnsocxjFPeuy6wsvWkhHDCBPjG30wV+MMeAJoQwOIj86bkcso2JgdP
0j6L1tr9wf7L+oYBxOcUGjvaeFzYfNkozjlY33vUk1Cr4oIG4sDZ1TAZS4X0lPVBsYRVI2tuKxun
F9s41/nJ9Ux28YyexjJB19OvH/2lUf1P+ySocIUa/oiOsTwDDsv1yqJ+IaIito+7QSDajuqCvqLq
O0N/laXoBnpfKLWYzBTXm7xA3ZVMO8xJpscc8A+xETfTUCmqrUtzGWcjohcfmPT9iaZTVQwOA901
3LpkLl7u5e/U1oHhHEEXA7FXnrB8PF5gED9bjqtfRfswHsMnWJZjQxFG5mWuQ0/pFWL/39t03dQc
rVtMKPdFkc2//pVsLOV4SCXj+hqle5knSNmCZqs+9EMMEle9xnkpgU8zBzRks2mNJ/BX1581hqHI
MUbsgDOYF9dWBQG2Fgyq25MDFdBOexHZH5HA9CN/89019V3JiB+ImNqW/wB8gkrKsjyiWs18sEw3
g3pnnxSXx/1eaOwIsFaIaCPhfM+b+kLCNScM7eIe7aNJRfEo+ootIkcamQ2A9f+XmwNgfTOdwGIE
BxDHylUoh3PhSncBWLwSmiiHcxmJ60tcuOAXGH/Hpe6zZZV8/b6pXgOA7Uf3geb1ObsSemeKiCFt
cdXlpUkqiRgkcS6f4I6i2ONWZvM2N9i0XAwJl4a/F+XuEIIxZfdwFZfkhhz0Ik780dk2QIdESSbX
Mu0xJbh+rjVGW+hQ5/w/RVR6WN+1800YFIXskPGaZ1hya5x88ydwmx3ZejSGBKhS/gLLjwJRPt9k
WFpIFpA6mAlgb1QO+fEIfhgmWAIUgEf+wfFpcFUDKrsbVkuhLYKBY6BilFOu0gGI8PCXHdleLpnz
OgQHe+NzaLlqnQYZNbasmcJvZked0A9KXWl1Dv/41VwZ7mx/qz9pIvl12kLgDLsmuG0Vq0siFVVs
Pd7R22aTBLZmCNi5s5LtXPobiZjmPeAnbTgBQ1TWAGP3WEoIUDJEQqGEv2mhEwBTH8k8wa8J7MAw
asUeJwW9ohgVoPMvZB5r+lhqd3RfEKKUnBM71ZvLqo073KmCUJvf6zRXLHAuLpPsAbBuReKomIhF
3UDc/yxduyM6bTZiMKN7TnuG6q4TA/o8NaoJYQrxiGQwyCR23jnBidcBZAbK8UXB7kN2vjvUHoJz
m2jOkViheqL2HA4Ri8Yj05ia2hghoNrDfF+NSKuMhFglebpv5ZaNzNcmHntItsY5sS59wA7sScYz
jHxcc1miv4sloirBxVYEWpUxzxnX63Ud59tV8qEWjRUw+JmAXU9Z86bHMjfJpus+LFQOmVlRYZ3s
Juc0KIW5wZisL2RqHZ6Ml2n0mJWcSjdq7PK0IdLexXoYqUvHLGdwQe3kxpPFU34HIXFqn+JDvElV
WWScekfTxuLn2V9kBbwfZOVwrSEby4++XQZhilbYUQGilcCzOqlHEjSTdxduue3Oi0v8CeGwDFVA
Ti25thq9WvtmKexv4IBMt+Ks+eGMvuuKEOvTQrwzQ+V41oqQr3pU0QaDQBWEmK2LMcqE/aIuYB5x
fsf05lqOCWbHFLX7KAsQLmtMi5QS1TNlJaWpbIxGuTr0kF8AC8CaPjhWFtSfOAANcYZkLqbm4jwg
uLhEVh3KVorYRJ8d/im+0/pabdXVxM4Bi55/4YGYn15E/YMBxy+OHWS5BTsSlQE0l0DACs07wj3S
doZMRipzZSIZm2gVrFp1lMDO+woFfZpNvA5qQTfNOPxLqQq//AaQt8LX91kdCGh/onC+NI1cVjO7
49dHJ9sBVXi6pc1PRdhNaXGmZQbzNUa2i39NosAvw7S5AHbZoIvJowxjMxBv17nOR+DPqXOYYJ1h
qEGvYlia/UxNcKvIIHySRZn43beP7ouwbSMIA45derTZMDKlkbQ0Dy037Fg4wVc+hNDYK/SykJvt
cIQ8PR71huTufWBwqjs5wzqCe7zC6x9PmDZbxhGGFeckJ6AQRkl5rho5KdMlUS3NRjLt+rbOnDfT
6XCP5RaNFs4Ruy5k2xGaytwTIMLBsRgtAxmTnOeB0ydAK45OWRe9m7Q+r/1klE0ePcD7Brpf5H3f
ybxaIJol/Wn6nzhFwuXa83H8GDhqH1GxvJPzhM7BIbalE8cOVIPypNR3gW6QhHDs/MbQq5KwyNQ9
Kj1NyXRG59yZpohaeP/jLLwz16OYbn4pD9UbQzKKA/tY6mw67GcX431VVkWVijbY7QE4nT7NxL2s
5/VDi3K2OCpSHuQi1li/IietbwAkqLRGPE8qPPOvFH4wnrc9KqWR8MC1rMYr8LWgiJCa7B+Zr5Bf
+A7xkFb3AIS1uVuhvsWDcA4T/DaZaMKVidexxihXQqwM57NZeb8Z5MAkU7eKk/Y6WqdLbg6Naf/F
jolkjQ4DVJpQjYQufLz6z0hqaKcMVO6bixxjEdrLpIgW7SypW/JHjdICAYk6tywHfoeEXqpRWYwE
eyI+33ERxQSNqNLY3nDQPvWcZdXinhHqTW/2it+a92FvqSBTQOK4ICIJdwLAiHC1KqPW/TmflgO3
ZTcaR2G/shr65hmBL4xH+Il+9NxkLiU0r4rbvAVB8B8SF0TsEVAIc7K8vnGnMaqLi5nKsEvrfm0L
AHgS3fydcZ6AoE5ob40uAyqaGF+3jgQGOmG/DNfCxdtLsAqMiSdNprhn+JVgUB1M/4gX1t9tkQEz
eXh6Whr8yJSu+/OaiRdhvQQhajMHsoKVvZ7srW39zOFRg+6gY2i3jW+zbLo/NLJstvALuKA6+03B
OBU4Ld7lWC4/VoSPSCfgNCx52c3HNyTyqcLL1qpyemCsAxbvFax1z1PdquiID030ROhPsoU1DhRr
twwBK7p1l66hXtMhV4Ed/1nsnW8M2yEdRajS9Qjr3l7yNXxg9qA7pe8UL0VqK3u2qN/OP1Qhn76g
ktZV2P+H5RdAnlNcI8eGTWNalbcAB39CbgsEvlvtntaeyr7G0VwFJBwOXqhd7AdG1jFvYIXkfxBW
asY9bPF275mJSO+Vw7/6ZLHAoyez51X6UulLBjd+ovbmmCoe9b9kmP9bs2zgBL58U0BRKR6twysp
+waqeoOElyH2dZ9yg0JxYiZTIbxiZ9tRCyJWgXXr1dHBffnUb0Eafcus8vII9jQhJg3Bi8B87nCK
xhyzNk+HtptT7UJIpJazAOColXat6zEmLXMcm8H4hdh6Akvuoj4dzMeLHCfIOqu88sGGGDnTenXH
OWll9Ae8HgVv2L4xiQO8cZFpRpqIEgVN2s7dwjmRHpe35YgTD+3X0IOAnNpEJVv6N0Kfrqc3Hnc9
n5YsT+ivJ+300FN1+lc35E/pL+uNp7pD5lxtqXY3AHkOo/B/BeEIa1qYdJw/3Dui5+dpDaCtKtGv
eBgX1moyhmg5WwY54ZQBnhMBQ8tQMqm3YCxSsQ55v676WFl/77UR/XYXZQlRNU9pPFDpMWGvu+fX
aIPhUiQoUuYTXPVWycjDBWBG6nMlYBQy6+iv0lzKc1X8XIG5DEJ1rJ2kj6KeKQr8FxrvSL66/4C+
aXCPcxrBEh3arXehO/JlxWe8YlC27w45eNsPHiHjWVSBoR95YMO0fOstCRsh+gUDB48HPe2GTQPn
QTUpVXdF14KijD8k7YBdaMBdlhv4m9WEx4ml+Xmj02efZq7oqLHoyIe2YTGKhoyFHvYJklfPpKrd
FUYXHZfn9t+CJ9+3+6xL4yixlqxLDM3AZG6Gq8+T63Ij/97Ruq7z8g35MTjFY9T92/73pxTw2R9W
HLgxszy1ni5Go+e2T5Q6hr1G9CB3rU0EJ9w8QIN5dAl8rriwjyoQxJT5pVjkdgFxauuYVuRu2euH
C6tnW04YcGpL2TxSePqIqfyA2k2JkoUcLZrc/tXHhn6l3USbU8fJK13UR7G/ZGUKE81lY8/aghuf
IXG9pbmiocFbn2XqJK+A51htSDMRHeHJKMGB+gH/DelEKi4aOr3gJl2bFmW+kJG5siI8Khc6+Hsb
r/jR7dEykZn4JcsFMhCPN4hRyIjVlrIZJHVSVm6gloloc/DF0kLKI2774vsjXDycVONjhL6RRXQG
hLVtepRo6h6WakTw3XOMU1sNPZAYcRuLUIG1P5RbIxVX0fVAkLsA7kESE/kSNVw92FyvYBC2+VYI
0ML2CGp0T2UNhUaCJHvhTW7ZM1XZAxV0e4fv/ZkY3QoneWZp8i6CRmlLz71p88AaJb//hEQLFAH/
v5/h5RVcdBiZEUZG7bbi2p4ECXv6SAWDr+b7MZe5UGyrKmD+Uf7hLTVwMKXnR4ZpWFvV5ioVAgPm
0vCGbpVBdHbRiNnD/oiMsjFcdKex7zJ5ssXBlln9h549yLNnIuPAZu8frTKE64d55gd09WS84UJ+
k/vSbMA+L2E8vsRY4FOAeGyTZZIn9yH+RZ35gvsIAu+rUmv3stVCf84BQpP8EM/bZgUHOsswc0Fk
VCSSNe1tFWwa2u5EKAE6fgkghAkULp+o+eGIOnMDAk/Nu5/16UZJL+pwpyeAFxqHyBdyrrxMgt2a
+l1Q9CMnC0oh3UDqELzJV7Vze6OPyLXN7j7Fv8Pz+auOfF10cfCwp/kNM6A5qTFEN+t1TZGyDvXx
TNTP0Ax3OySbXg5RcmuURk2FsqkOikWZLN9gWfubxiqBM4R8YIJpF9D4L9RWCfo4zqe/vAPO79rx
RuAWNsxOyV0aRH1uUJYUTObcdIa59C7z37DOfi5CksS3cYezPzMdBFyD0IooS0bdUTXgMRoNS9lk
/Hh1000BTS6cUzRemEVr1io1v56wlvTU3U4bstLTal9ZB+tAz/g9eDUl7NhaitmTa35nBe5MBsnh
Zq23D4ulaxe4af2zd+0NcwAuuYxZLQhlL8n/DWXXhlLxBw4Nrr+3ju6gUQAGn0iCwHw21Iv5tVKJ
HFBs08K/KmJksBaaE2yJmYT1O+KwxJfZoaFTuV1QolLciyWAFzQnNdZkrOa594mK52fpnt3+BJpm
08PHLAiYVC6yJjzOR+81UrOi2SpvIGTXi84SW5Ox96dunL1tUMSayXrUXDcUJXKfXf02G8IwaUqn
Bwwxx0mVld796nICNkWZROPll0UVFlOm0JqP0FeQhlsL3Z/C200GeaEsfFqzYodj0FdSnsEQab0X
1zdVhfb0xlSOhqllQxyQxfhWtklDt8i1C7zJH5XeJAe2kA78r1IriWBqIIJNxLfzVk3bGRCNUGHY
dvfV+SLp05wLI0omayIynSr1tDhAVSqIbKmZQ/CptqEkdMDVrqDiFktMKFGZI0EqSh7VDvAgr5oU
ELqzy/f+7OhZDWO3pSlNRCv2RH3yffvsb8+09KwVFqZf2LUG8ffd6KyRB5aAilRz86uub98NtaPE
HRXoyxjopgTz0WAWIhqdhJx3eGSpOlrsbVYMVaWta9xlC/M/BF0J+2vhfmL+8FMPmXWbgnH8e6q7
MbZTOb9Cc14INa6bIVXJIvItgzx88wLXerFLTs7cGMMOKo/EGpAk/ykGGFXhE9JEV2wrqGcUG7Al
Fn291lvsAv2nQ+Q2aJuqXz8FhRJ1jHz25TLjP+/vbdfU81WeWoq6wzF4efC+xHzYlnTKb31YCUE0
nfJqmxng0Qbi4VRLwxxanLlupher3g/eaZp+CBF0k8nynYK779FWzsryo7EWUa+Vg1EuEwJ01ld+
l1hqrjD7gAhKFSUYR31ws3qZuyqyv+rBKrhAYLCbyNRTeVX+ToS6E93YmIvrnUNUmCKzdW/+lsnm
xcwOWU3X/Q0VD7MBhk9BX92hSxNIn7qmh+p+HOwyA8Irlv/MwToQbSp7SaSY5i7Q1+Qhi18R2MFP
xivvP+KQBek54aPMVq8ANqDrTkE8uPoXMigWvdQI2Y6dbRvrLge9sFXKGmUniC7CZ3NIV1Xv+cFb
jJy5FoiN+NioIsL/P/JrMo5/PrHhXgLYwWkt68qmzrqmbmEVl7tE1j4GbxpXJkWNLb2p+GnxrJ7i
FiPFexOJ4axFWBg52w/Frh01Y1QS9UJgV3sOPLYVnQnjcMETIDIKT6N25uIzhIwlNB1nPHBwTz8D
ctDIP+Mat8O4RvYdi1pnr5AMufpivL6zDYMRYfna17yIZpfzuQ2JL2t/02zWU9Nx34BuPh4DX/96
GzCkGcbXpWeBo4aeAxaVU+v9jmVpK79+AFV2vJU5j8K/9WBa03l3s0qfPd+sQ0buIBdftTBp79a9
6v5xg2NslY/KWDIK8tjS1Lrt0u+ZVKlGe7tFn7C7VthykWqgW+ujLpQ6BmtqJ042BhoCpUBrTFtO
iKWwUeY0j1x5aDJQu7CqL/Ur2sS+hB+S24RL5gsSkxkcsqrUzLxsu0wFLMVsi65X84CKgvRx2WlB
xb9lviS762kuShQmAiuNVDs/Cqri73Dw5fm2s+d0hxXGR/mo/bNjP2D4W/Z46cZ7jhyNY8kchvcG
sDL+GIYmYW+1o/57XhY+HtDwSyZsp/WJVcNNiKaW9iGizz0Sfr+K+QXn8O7FG5erCEvwurK0pefL
OFLDRMAQrSvP4b+6iBK76xatjMGiYafLzy3EHw+sjpvgH+CE+UJis4Cm5HcCQixdEAQzY0aySmUi
GItIkGUj/cjC8MzUw8kP97oZw5nBj31bMluCq3HB5UHtUO0lOI4OMelvCXaTggmSMLvu0VDeW24c
YXImeOGnayx6ObmQFHtJTbKD6s/ktdxaULjGojHoOP8lafO0oVcfOaaZucGVQCx/dmPtItjghy8y
fL33Hh564yjFFvRChtOgcY3Veq/ZusUW7V9SJcYqRLMQXvw6vSq5aZAp/v8ZhcY0jBFiGS1mMag9
56+wf+uWolq00l5KcW/Th4BSZ577M/C0OCSJe5GlK7edIpO156GJ0IBu/PtILhjYOT4ieCCWa7Gj
VUlsIACSjkmaInb8WrZRVPcfvVPicLos4oBRPKZjL47zmvTF5Xl0Kyf5HBCR9wvlpy9C95LIRvXd
aBZrgiXjGCV+qOcC3HPvvZVB1sOjlMUHkJwmjGXfHzkf0w/Kmv26ADsXWBJl4zihWV0t0rs/GDCW
2YihrB5lQHbrDxKbH3Q8MnqeyLdcDHXHmlkztLm97mD094Ao5PjrP+8ejlBin8XtNn+hbublbyd4
K11CM8bMDT6x140A2feoYR6KANSkgtghDoBdDthCagyQfw1neSD+MeMhr9C3Bm6PqmztX9cpooqO
CQUnNDJDAvAcd69CjF7sGy91R6u0aDu4sfgdAQs7wWCdhgxQdYgKC+frSOI3jPnLeCXl8MrJmgYE
mgMM94qS/sxTKt00kGmVriey+I2qK/YPbTxOZEcZVErhwiHeDaqNY6k3d92gf26/5dxYvCDSIgdj
zjm8Us6j/ZYUXsY6uBXGUZH2POiKyxHZZ91pUIUTnfJIoC7+wPUaDka291mMqdYxL/bQe3oykUst
YO0DGFsGBLvyOEHCpxJ3PLuauTT0CcsuoAalymALBbEil08IfqpAF+UcmcijLu843eOrOhOPBP8j
d6Kc9w0Wll/FNMHQGTduohS7AklDD1lhYP2w7lMxITr5NLw8dGqJVO8BzQg6NNf1nqXX7Jae/m1O
azx0snmXzXVClPhjfh1XllxGTtN6bIGQak197YSjBRqFx/ZQRD1iOvqGofWXV5RyUJNqVgLLO7pb
f/hmdlSveCvee1ju8BN0dt1Y76udIdKE53qfe7eVEp+bYZyD4rCHtOel25wXd6N25ImdvDny3pcU
nULyGg83DafSOKukHQJwszUuHu19cd66ysx9TkcJY0G2LHofYIa6yos+Hqc8QZqfUms9zMeCmyXy
uGbvA7Gx2shSoNm3tmlTryeEMngmFtXDLJqzybLWz5+T6zlPI87k/qpJyKv9IBN3s3XSzohqgA+9
wSOBJN/v8PSVakt6ugyIA6G59q3LEbIqt6xMoY5kM/SylUeRed5QZOm4ouUiKPgd1L3i8K5qX9dQ
oULD7d+f56MRGo532ktttMctOORJwhPQ9sKud/fxpetSdxVLoyBpaI6MWlTmR9LwMjJiJiTKL2+m
fKtMFP5x+4SpQEvErE2iInsnj/hJs9nVfJHuOd24WIuN7JR5SfsX58sLsHH7weWgLo1E7XNASJ0V
m9bRDqKHwuCiJ9J0soF8HQTqdpQpyH3VTHz/Ev4sxWUh4EnUgmiByukWWEhIosjFYSGRMVSgFCV4
Im7P262fAxONkmc23HCKZUKlR3b94/N3hT7nnm4SujcFrP/En+cO9GifDFGhl88Pn2VxGV/nrpGK
sYx0x9XXy7zAddjoM1qsv01f2lXLK73KZ9hdv3/vBmbTlfsTVA/fCUioIY5yWRdLcZisuGglqKp8
Cb8alqvqZrJpTso0BT7ZoXF8jPNpS4iRFGuXbpfFCZoF/6FI2qIbjywxWr81heQvxLjnC92wNUGd
uGhQ72XeVDu7OXwLruLZrpUqwae9aani1hDwcq9TQuIH3ERvwz/7Y2L1zowOlY8mTd2c+q7noe0m
GIBTkp7M9c/pa5fu/jgsmN+GHFBtg5/tl3e4TGfKaKs4dLPiu0Si3X/toGN4yqRpiTENV8XgTeeP
2VOKdeLNkDY2zFtqyOgNl+OMQBHKNFLHAoau7mvbVXqCFkkGMovjWPDwZ8cx5vtVh+ywcu2MOUtC
lPD8trT5kNgTTLhjhhQkznf/9yDzCmnUObFUzWdQTTT1UW6ryL/Hmb142JyJO+7ubLd6TxLPC1HE
5+qxOG2zbEWI1RCW1tR1zHc5AILO4oHZeNxn4MYlQFhwtfX0Xzd4r4nCrFhMxIswdGH0QHdUl+T1
YPeZvw2Eq9geTNcc3DD0pJ0UlcEkxkHIyRilVnixn8+WX97W1xbKoJEF107qlxzCA4ZKwp/J8zaj
GI9QYmvSV7MBDchmfMr8QmL7acgN2l5+12UTIbAcg8y7jlj0jax0arRmI/K1rHnvocgaiGdVt/kS
YLXF7ottxGJi0F95H8HYJLq1tTlxWqtKM4EhP6z37zBOCC4vprKshi/nomlTLEa89Cyz7re34Oh4
PlIIE4OVK1JEnN9h+z/lkuNsSnxmZbOeUjxgEhenO5lZOfu3uBU66U1Nfk9zuV55/Ag0SoEjK7qp
4QDYxZ835/EiavKUlnGlMjC1KnIDgJMCGk0hZhi8F5EQon05twxdd426gWKuKlAENKjRhyo3br63
BOCGRCNffa4WXkdAZLIHh/t3ntxiFbab/6jjdl61sxQzYFR+IyC3uco7h+gRZiFEZgasGqkjk5KM
NU0da++4uVrfqTOI8kO8z3GfSLTIqEmI+skoJOIn+hTH2PhKAdRRwSAyUhiobwpXieFGFuKXuZS7
MPp3UP6iS/5gcdoxNrdePj6GqTIbYjstbu/wcrbE4/+6et+P+88fOJ6qGifWebvuoZCwxKoNe83P
IT9QLwbqwryzd0sFvHbOubkFy7eg42EYj1uxyXjnmFM48R0+zw892v2o1dRQkhI8xsUspK+CkDSE
EJrzbGr/ChPgGTA7U7kLlUVjiJpoMdmdx0dkPFoji2M06NvApghm9VIudXqnXIMnjuGropQfZrNo
GrNYaIotYAwk6jV9aflFKrmmMvhSfKd7QcVeAcebpQHX36HwYxn4J8C8vaY1Xww+5YcPuGgLVmix
xHi3PQXfx5pi7Efol6cTMkk/sxasGPXBkesJohJHPdNshDgZk07xvh+4V66fuWD/CZU4cxK89btL
UNHE+vlpPzkR84+NKOJCV8x2p1l8CRJCOUFJTbuIKQSuEzonRXV/mqor9XTJmyO/pA9VtWKqP0PB
p8e8tRTZ0NvqCKqkmpl3prrx+ksWKUP+AoJlgBIgR+kQ08qaKzGiyoqs/n4tg8ZoDKXih84ChqPb
dVTsEM7qn9KuZl8LsqMUPkcMDhvh59KdlzGMP0a5uJCO2L1l2Ag0r9sQknrq6Utyc2yexmfp9PPP
pEuEsh2LRlceMmUBqgjYcdZCqVo2Vk0Wd9EYyoD22TNGYrEAP0Mta4lsj52A+r079SFytsgV/JfR
wJwnRjBJwXfW7V2+0xIRnEYpaRWNqIJ8E0y2JCQ42ItdAkGMHiKXObT4vD3hxVUpJ6D/5aL9cA+2
weSCArZMHAjK2VUnMEn/+STadb7lYUKOYFd+dx6l1yZFtxUugV1CVCioW5FG4OMwKQxGbOf7KKzE
hba339tJnkueN3W5E6ZeyidqWnb+8dDn8JgzF4dVFgQk2PHLIcCUzsQFmooIdcY2OpA97rccGHs2
/6FQ723iL25yNFcTOjmsZ251rweT4zq6H3n2SFvZc3d6KxKKbAABLZGiI0pVx9UukVYNsqKt9eCp
HAGRZ6yOFtr7/HaTK0FyapPdqVCJGKQ5x2vpnKtJA/37t0tStlRBSiWwuSxOagmzb/rJuYGCwgAM
ecXQJSFCaW6Vhbu4I2SPt2wYM15FY2Ttg3TxW1B+jyK9PFyv+HYNW7p6wBzd+KXRQzPSHjqwNk7M
4nRjXuiEZiax4h63qRyqZdg0c0Il6p+vUbXhXdJqPdI0IgBiqQbz5uupW679sAzWAJcqo5Lr6bOT
PhrPsjP9mamDkibTc8k8efx6d8oit9yD4ucBQICfPn2Y/ddJ4yc1WHKgRppffNco/BC/AQOp+0QJ
r6fnCDG3K7OkPGvO0C890EWAuxOy8R+O3TJsfuZGA6SBpi8DzuAKDzlwv9fjYBVn6nXOUzdmUN9S
Di6jZkR009pSDjPEXWUh09HBlYYqb05xT6T79KjB66wCPn/V04JbBO5Vw6SxCTHJLZd+W9BQDRtY
U3win7tt4Je5b2nRqdi/duL6mccJ+g08e6zS8j/qLzoUKYET/Lpi1Z0h6XVUfoNEYH03X5jLiOlm
3Vc2R29Ck/OOVJt5GIQsofBqntMeGCLia5Z+N52IUjMEJom1BOa950RmdBu3ZPPVxElmm7fL0chg
D8Wtf8DqiieSOvgPQDrwkngMHJkkOYp9Vr2gjPiXsMhwRZYDowb0fUw8efG8XFVKv/m07MXO9zIL
3N3peVlOh7QsYHZAT1e/LkWGo60hPhTSADMVRWGM9BKXwyAsBsJz7ApQhJn3mvLIsvpQVGFpL/TG
7pLxbYhQ/qbfG3Ww5dj6JISL6mB5IyJPxjdjOAkKr57FOPxCh+CFkMRGoPM+6n4gYFgXw78GgNU4
UD4I6IN+up/MM+rsjsOncgN/OuX/x8U6se5g2MfCIs16zh/2qmKaUoZ40hoBL6CXuS9GvEC0LJwY
C0kBP2T3O+B7KayBVWfS4LG8bVWglnRLUzTmIid/EIph105uAgmy8o3PjeUVxWF9JKDFIPEqc5Uj
HdTZj1nK1ddjCbT+k56kIfQKuIWiHC4YjbWlLgRo6ECfxDR6fWT4aTie/fR6FzYKjU3d1Iq6m96r
VSTjd7lFQDFC825uVMehsIIlW0kqjKGvMaV8/eZ+IupaT2OuTDBhJbv1DrJOS0OLkASyfbWKuBuL
nJ8pkc7eSN6xYENqMgDxHoUdZPG+fRKidJmC5YlOEdkOZa/qojdk+qf1ITro3e8/eYzBnNwyvA7z
MawTDKjkPHZEGIR9cL1zm9+bpPKHMfwHgbThwUARrNjYAhMfFHIjnM7M4ksaRjAavwDhaERB3GCF
AewpXKOM92SATvEeaNujn7lhA9E86sjOBNbweHxc/LE17KBwPwdTvim9XfbgWNrR5cxbNDXhD/N/
7gkbNAroGrlj0xBleKHDqet9R/ELxY671THEFZq30J0YeWgRsRwJjiWyiXVs2h5C2yOILGGLvcHA
Rn5jUDfc9qTsbX3Th2PHcWbvSxDKsGya19Y67YTVlRNf6LSwoE7VyLCn9JAPqfkwP/9rbD00b/xp
6pjVTHzvwbD5W8SldkzF2s6EPcn7YAE4PQvCxl6BS0q4Vu5f1cbg+kWJgzxySi8EoFwwnHXlti9w
DQgVPXAhlzS166g5fC1+5rX8BaPbNMrk80sJ+wJiVV+tvtH2An8STAA1OuPIpgyVbFoA5OHx1Tz+
Xjjy17iIstdfs/sjEb095UESj0dKk9XoaP/LwI2CpuY02MqAtsPJbKlzGveSK5Fq4VIHtToBmgPG
3wVHJW2dt01VxSWQGendBugXUpJ4zDEEa+2/8S5/NtVvrxggRjfR3Up1qSY7kFOWYC/5i5oE8oU+
HR4v3tzw5ZOzLmEf6ycU0AemKlzjMEAq8SXNMW1xHzjlucFShDNCEUw52WAKPdZGFtRnMU2UgxuX
iAZLMwLL7HYWaUGJ2Bzu5/ZyasrUDYk6jZoDMp0mxRLSZXvzha+9+vgJtohrt1DEfVocCwzY4ecb
+RPVP8ipqouZUWfs7xwwJY+SxhNsmSG75G8KxwRmUnMIbkn/I8F0rqdWbbBdEFN4+PRmVd0ft5c3
c2C1DPx6TjYhgzRxrcRpc30iWXCEGeXOH1ZVuzJ08MZY59cohpYp/JoBhgwYY1EjphYNVqZ80E6D
0+KXAYKBGFRdbY5i6aBHs7uCJn8SuDBIwWXVp3hkKlA7owDWOl1pixbt541x2FnFS9XLsxdwIS6S
RhmbgYW0ZBY5EjbGACXPt1PprijipLCFc1wbT1O5h748SMnEx1QtwG+IyYlnFe8VDnJJUy7Fu0YG
gSRdKT9l399L5YbHKMlLR1vWI35D5NvRIxgvoE1fwECeWh0ig3W645XkPHgtdEwDu/D5SJ6+4o21
HfoqPkuUczjYx4B7x1tDRv6Z5ewe5QqUqbL3cL4uq569iZDWAI/uxNHP0csNiNxh99zHwO544Dxo
DwtSJku6AKxcUy4GL0KNOH2KcoK59zCkKJ/JUQFOFQSvacIZ24H7kvTkxIEqgXXybw/fNyM5BL1a
cH9bN7OKDjp10gdT5YtDIVSEgVSPJ+MRcWmy9h84yaeNKttiHP2bG7nozBHZWza3wrPdaJYjvv2q
a9YEWjCbY0nvN232e4fw1FI2FWgy+bEWPRTlif/jZtAW7sz109YqaIhj9Xm69G+EmPyq9WrMxRDa
lp8UKh5i0XE0nkrcRTvY+lctGV04T/Iq/96zUf6v+F+Q6MaDRjsqn5wkAZIrCfnkdRVkYvziiPTn
Z02Yrt6W8O4XlFWBeICC74aTOTKryMBrYuBD8oLM0ZUWoi8+aMDaIwyjBAvPNX43s4ocsWsWrpD+
Eo8LaMyI1eq8CDluQKBiIaa0i1bkLPs4T8ZgIbjr5JpfRKHuZWELJz+WG8Wg7IPfx26dpkGvvCf/
P1yHDXSdnYmXXCCaJgC00o0cnkcDiqRsATw7hS7nHoA62Jjpaj73GPmiQaI79GmoZZUIlHdWkUPl
fn2kXfc51Q2V3QGEB6+jGjS1oBnIyDCLWPEKBWTus8wlnz4clEKyrRW5hCLTLAvN3CnCFvjwb9PN
ATRrH9YpMN8y06v1gNrvckQBuNKh++ko7REowgm+AKV+rwI9d15N2K35PK/s+XC0GpjbOPQeHNfM
FBpj9wuu27cQUm75tidXGoa8mcZlEk1tiS4Ha0dqo2qCHVi2RWp3+RhnbEd9Bc7yx/1VHqutJ1WS
CZWUYrpMF2MHvRLvwDRSKX9+O4HC239jKa9ymPCu1Ipn6898eNiRGt9aK8955JxwwXLJq37QuFs7
LSJXTUB878vW0LETz8V64Hxz+xsX2O+f/3lBVIh6xJd9lZThMDhlcJC/0JFgC/zCM3RQ5FlOt8p2
gCboAfjO/9pL81sqeOLLcitAsuZXZbbhE2h1cXPoLZoGN+hXMrvvyDJ+BYky6BROlelMzFcS6n3y
Py0e8HGqYpwAXyht1dKlljYicIU+P8csZeSZchl8wA9pDnsYmtlqIZfueqE7E4b5Ke2G1uWai+g7
ZwcjwWgwY5uSWGYP4Wc+OvgZuUW+cdC9e0qA52te05RWikIHNOmGAUA6pF1gyHkBJDUEm4Rk0nmP
2qHYRJF1ZRsfvfRPBwcXrgz9IkLNj6gqUAykcqCVWwdp++JPub3BB8XY1GHjoEie1R7soJ87wwCD
/6Asj7VjVIRoNx9uX+l3/c+K/62xqi1JZ48Q4Yi6RQ8bGtwWiFmcOkMR8FCZxd1u4xGZTzan5l96
Gz5D2waEWxO8sNLJF1HPS7WymNQdGOZA3wbsCFu0WR+WTffcJgdYphQ9UvM0TboQHGTK762GbF3B
/Z7rPLoQQHpkb4xargAHjKKnBceKc6pUiszSKbvLHYwurJoQ5aDIcGo8X7Jg/bKVvPE9LFeDf0qu
QV7h1GZJRMIGyy7Kb5A9YSOPOivwGHUbyfEGxqhNCmAJmf0hHOqXYiNWi1ejIaW+XO7cgyGzgDEa
u+3bX5QPsxFbNMc/EyqJpIKaR2ic+wwPYt/6RBJ1Dfj7GQV8ZntlJa91lC4zBxgqLv1d26HxOe4O
BZV4Zmb1jdOVvCDc3fw7lLV1sHGbrlJUd8CEXsKZRQZTOsKBzAWKfKMyjEBYxP9nU7ByggRVhj2I
KtuMl6Rlu8XZsVzKjjNKiWbVbo7PB4Ql/qBys96zPlg2y+ONUOOe6D5t+JBoXpR8VqHw9ZhhKgMk
+i+2qaDJ7OIXPX1gzK1klFivO1vDxgWnY8gRsf55jxUHSYoZvKyFV3CJQaAc+eqPGxVaB124kHp8
vl1inRTgevtGBYc6i1d9b1nnCLTJmr155r21FF+Mbph1DQ3q1Xft5plQLCPN2v2Uox+vDtytUgtx
WvIHDx12O+nBW41T5jAzjBu/th49fwJKOFhWdD207Y6QpE6+8rJsnUz53K5EOq5vQaHxZAoviNT6
RBhdEzUVYha7iS+ZoPjAAolCxf14TkytXXbJ/0iJMR66xbs8xyU1kzjmY98ANg6EnDECqC3DdQxu
kA+tkY5V2DY7bNn6/VDrNyHKy01lVgrDuYRs345dEpPCqx1+6/7LYABoCelPxIh72f4f7ILABrqz
oeYtQzidY5vlHBe8MPeuaiUEocA2zNU8vr9flNauOvW9zIy0ugYuYLnJVqF3yoVVVj2FLYahe5nX
wxVA2m5er5K66pPH6w1/gVYV3sbcfEtBefpHZLF69BCZypvXDyS8OCoDPHwpbcyKIoFv7x123pr3
/hngYGxsjU7jET+X6iCniJGxWRz+1dBbH3+rv/1CvseLghXHtrovC2gsj11nDZss6A9O1pnHJqUU
0TmA502jNdGCAL8F/KFljRyWZSkVRHtMqh5fDrUQi7MLc3aeviM70JyFtLqbqh6OjmJgYcwQztx1
/g/jJJX8tTH1nGVdVhlWGeuLcpbSLsiy3HnAWOta70fUO6GfJ9+iAjgD1EbO2DQbn/HG+OwDb6SD
EMr4Wux23cLXvvl5XxWTv+2enDrRVK5pEWCuiCS4ykIBqQD1nVOOcdAXP+10mMUraXpuIjA/cDze
fEKTkyfYJAi8vX6Yja3O1JIZFNyPsZ89L5kppqTdJwIJLCyCAN+w1Sm+ILoTG16s6ZPsy59+l14Q
0c7ik61UIa4gdU3/+LR2fxl9v/VwSd0Ox/rpEp5oGLs7jdxRYwJVGUpbsjKHMaxqYPnFqquPUseQ
ba4K9+LJnrF1SFMKdmXV3LxhOW9Q6OUAwB8D15AZ4qJNOJ6JL8j3g4rF8iHWyyQOYASb8gQIkrV+
oAri2XTfe485M5atFDQvc1sQ96STpg0oR/2KB+cNu/6wnZJXDAADI1+b65NgG7BIDPgTt4ogIwpq
R1G0tLqB6FINcg+kCZQtvJgL7R/4UXxMuO60fWJ5FbRNppmJdGcaC6vygVL+1kIdusYI//dVzJer
zeFiBzKD1BGfNsvfB6co132GgOMWDD2ARA3U8HrQ8XEl7tdjqMhmg/atwJamfRUre4KR7LK1NoYf
exd6AI6dpR79NPgBjWVuBQ1Wshc8ARAKZ8nEDoMuAftd3th+kX0uFH6i3t11J4yiVqz9yomXnhQW
InG6HRGGJPqSMFVKQbGpjhCdWJQOUz9LkedjDmhUQp0UChPDtIgDzMmYwmSgFPs5Jjgl8NHz6Q/e
ZT3aIR2C3tCI+WZ5V2PcXY1eVYDrcO/arWa8WB0Hr0AmvFLrhViVA0qbUJFA87j4OZ8B/IcRJwwM
jRJwKUsRYTx0JsQJn/KyKTAUHnM7MKy1joz0ChnEak5kVD0aHfAWkN3dQWe2F+r0xdEwKpM52kPu
Ly6plPDQPZ8rzWDHb8OHzYWBf/cs9U10CV4loEWqcjDuJwunIyTioPtmhRgPNUAs2ymyW32Vu4Dv
CnK12q5yF1E1u+h/hsfmOXEImKu/bzWrMfPRseqKj2GLMQyPeAC+/rhaGHuOpAyaz/eeoBVDdiT1
Y96/HqX8oJPgXK/XYvzElNfF7aYOLkqPQ+Yvmp0OKyItMd5hN691UuWV7/WBVwr51HHERDD0RQC2
8yPqBnI9QD5DemryQv4dhSQRT9yfg4fAC4CYcVKzqp7yOr2P/dxjKUVTR/jxA50+xA3gzL8pJgnQ
CkevmLixqvhXwhve3wqpkhe6eQ2lonh6fYf3Ee+kWyNFG8Zdhn8YKp6hAVlq5jwOZGU0C3XsTVOn
BdHXuhpMu1AjvHBjrjCkogqI+t3DvaYgFSOZHre1f7Be4v/rcsm7yx6OFMV9fyMKFSMOH9jGGwxL
XCLB3YqItv5WSqA6fnjtq5cK982KLcTv9dWnrND3IyfoDYg8pUCbXJhSA/BCLB0bxg/Yc2V/qrOy
ymGLmw67XMpuvQ2lmhPdyUDHRvVYniOb0LQSQCimkS3VLR7rDiz7CB9PIKw4jV7V7HK0kpYnU0cv
e7rS9PT5si+E+5RQOZiFT6w5AeRG5GURbVotcV9uv6HsJOn0ytmUADhFgjf/xh9c1X1E0RRHDJ+f
TJrzseCddyJCZPv+CjBUwSYZ4MOEAB0UiKd52mu9ByRvzkDvpHkBLmFCWykSXOKDvNB4w1+JgTFe
zUrPeO4nGsymDPkPJp+qSa3TstdpcNoy4v3BusX0meK4jx0/AFmgyADMXBleiJ3YQ+IP5n3DOh48
Pwv+RDVdP/ZhkAN0kaNERNTuluAzkrJIkkdsmrRfILPw40bOEXKl9W+74Of6dq62yAkTYdSETaZs
Q2mpBguGSjzQXBXT9AcQl7T6zchCYPTcaq0ta0UhuoJzqtAplvy7hjGPFUyLy2PlLyLUs89TRF7d
CDwwTYzQIO5Fr8gDCXxIZaBi7PN0QfWTN6VkmrqXuoF/gpMf+sAxrFJZg+9bxO8eLvphquE+hKZr
UKucZwgNHoVArMj9AxwMcS/c3OeLhMtJC2SpFuKb+aA9pKutRTXh5Dmx4SLmpKvMSUxzxuf224HA
zCprcOS/AinajpfP4ZQ8z2W0SXIsWIo1xm2+hcYSLylT+bm8O+lU894yjtlDIupXwCaDUEGiaprs
i3rmWwbRUrTbZahSTbWC9n5I0ed75PPXtzlNqLiQodqCuzRDlcT0FQsvHWMUFU3x3LsxLa9PzLVy
53iyY/NSsJXRicAJqS3IIrUnnYUatQFE03hEcaMGQLjogQlNvG7PANJNjjXF/c8OVPUy9LGDjDt+
rnaVfUcNSAbbAd9xMCUBQIMkxjjvZT6uFBZpMB5h3OevEWiXb8URlcTD57qEvTVnfBWr+wUyWrl6
HA5vO1WqaTxw5thV9eK4jDGprl3LSmZzHBPrMT+WRjo+7Yyagarka9MEsaBUU+g6sqil+Co2U3Ie
RaQL7YNfx1BWuPjfreq1pLbtmhepeR67Nh5GJ6DwQLfXrnAmvqB6WijjCCjSfcoDOymmYz5cwHOv
RwO02Ytsm3KaxsElpsi3czF2HHPnF/m3gDcKUyz00+P5wHxQBbOstIULCOgdqUfyq6/BeJECHXrE
43I7NAc6cV8a1z8Oj6N6oZYFjHYoEyXPUDSnGuZXhlgLbRj4HZvVfck4u1CSnTDLrOzshD2q6ufS
KohXK12Dc90bKw7DWHvCYtfLENTy+nt9/ZD93CElneGjo9GaqMtY7FcMge4xJukB342m/7JWpWw4
DyPdnaLy8ACuI2wgIwNPIJXPHVqF56kK1kR+J1bnUT1k1dAZxZysoTfJQAPpsV8AJn+cIvLox4v/
wXu0xSfaPNv+nYbe4BcIonj76OpBS3tu08Af3riclwNbbbWMz7wV3OfwBDHatzjD6/n4boPswijg
Cnn0W5hqx9E6FaWDKqP7r6BWw1Xw3XFjXMLsXfOwOcrWumoLSUbYrsSRrt8gyjnUa08C04D8wp4T
Gre/Kfel+I7M/Q86ODzTw7GQVc/08ahvSZ3d5LuARcSkWZkucnqhqTvxDsFo0hODA5qPNfWjdlwe
wUtxOJnIkDerg49H4x0gmqmX0iVfvbZDDeYGiVzMkzzd/aFTJX9Nzxb55aFqcFcNNkkkLWPYDyyD
n15+PatsaVyEs7Lb2C0X40G9SKA9C5sCfyx/ViWb+sVaibFjLtDTmWfTX89D7G7s1gjh6ZUpgBFT
8jy2jAK7fcCOcPG9q1X+oOqtBAMa+ZxpJQVv7EVPwoNncZQf1chT4l+VxdsW8Bbp3/kDiFdYIMu3
QI4dN9KRTgTPj0XTlBIR6bNY/UgBvEaBZwWw+s5rUUp6Y2/Vk9P6kkSkS9LtYmIaNf951ncIG6Gh
TgeKl+qJNIf1An1EMLdrgT2CONnxM07N+KHOnbl0MxL9sSoTtbzfVkfpJDtRPehZwyvU77gqYQX/
6LcGc4/oywmYU5M7HzLL04j+tPcP5ndyfZnQU63LN6vYOrPvJgJEcGCXTNABrqvH2I8lUqFJjybS
2zaopZpbFXufje8yd011P39c/ZpFDdovhl3Dvuwh7c8WEcUCV43w0oCQcMvZav87kCb542nuu8bT
QCuOGlV2aoznPhZAyeV/1UExliYbPQqflEG0W4PGoJ+RbjYJR56jEkyAPF+E7kTn1wZIqjxshY21
ptyRrN2WehYhMT28H+/KAeDYPKBZVpGPxOwcM+RU32LaYdewACdHxxPPhHQyPDcAzk/S/1M0xuS/
bzhUlMZjGMkmzSBCLd9LUT9Z0WO+eZhALnS0Co8kn9CXJvO6HwYX1mZR7bZ4YYsQmqxrIO8b+ows
5rGKcKqMGMoR7L+CzD93dF8aDEeWRwPIs3HcGL4kzwj+gzOh9yoH1WlB9aSkVTX8LH+4j0Lc8qg3
JRnmaVsN30i8VUW2rq++gfv69u2EzbYvhmpbOnUXyCfkAsttSVxU9bdcPQZNu5b0H3qBMKFpZhz7
HiU5XttItlbqaGRLRcUv9tk2cEdnTuadIfOzm0/Vz+MVOuSjG6tN7GY68AEfd7c0UkE2lisXgl3i
1EfsbgetA+AEgPP1q3OU5RcjtgKBzyDkFFx8ij/0dWIliYrtb49uyg4eIVDHde8lhXsJvj0umS/i
e9HtXoAUQhQG6j5HfhzE0enY9MUnPBQa4hMW+yRSedkBTXpsVfykeE0YSNxdUvwcA7cntx1rMcZz
Ig8ufwCXxq0gaduTXpxjmhfouL/Hm//BUmtzrQ9BFYBvg7Iyo9ISHWeVN7QIXoZg/aKbGD+ckaQH
lc4xI1meX2vZv55+dq/Uuk5QM38LLOe5oN8F/JyggcQWnp/mSU015DcdGxbXgEyXyRZseW3A66yz
QmQ2+ZyvdflS6DPUPtvgdWxpwXAOyBSq+0LAJHWQL6X8jt++SLFRHgVoyMrFtfHF5exd/7fFumt3
AJno+q9z86r2rvuVDLjKBVdY3I0YCuMIC8cGZGYuwE+TdpgQqkzv1qHvLHxY1hmk15mwdcN18k8I
0wM94vbg4MBTkRbj0u4ath7zaSlLZC32V3SRluYDyvHl+2pNC1JU63/oBEk4Y8GmqQEretpEyogY
i22fIvUerY1RuOBWBX96VB64XLgD5XcJcOHBMYgsvy0M+S1/8wYDqPJqnqso1CAGoHXaBnbjLO2J
i1a955ZjAcIDEuJcWZ93wY5HRAAtN1KiwGYoAV8HMIf0UcKVE6SvAAd7Re8r+bvNHjYxt4yMMIXz
OeDPz2+1k4ylvWRZhQLEgynoPnnO3Xq4hv/KW0zaNN+bDHhFyfch6bojTgNLtHC+EXACcTAaE4jm
gHdOziKgrJISsnjKBEUU/mT4CHXL9gK1F/en0DBc+94jU1bbJzGAyLXUOIMm5d3auPMuPsHZ6qDw
Cp9M2gUxqwnvJcOrwj0bPH0BPAcopFyHpPoRv98BPW02PHRtMGApXPLXKRYenTBKUB6EoouD7b4d
n77zUyPGzCYp8nzuDOoRpHT13GnLAMtDCUsF/ANtyRPozkuvLQFOVaPsSwJR9IVPoIxHx+kXY2nt
iE6exRjZVl8ajcYiOO5v5SQema2ip0USsXXFNCgceWMuZXcGAUdf/HQMn85hQMAil7yEBvn1IT5M
ohb5UhJSMKxzXPZT5uapwHPuFmkfBl/az3K0zSJbvp+tvZIkIuIay78fr3UOc2iNy8gFIzDOIy25
/8Ipx0LRtRcWSUvLQGV6+MNGGaPYC50nDKiJdX6dKxMDG2d/zFVAsRIFC0lfDQty476PLpjzhmzY
8buvZo+rDb3+hAxcXO0RsLxjbRb/nHgeeo1e4MJQTgEw8ZxKxQGgWac0clASd3WBaiIbL+6mfMIM
hufTpqBpkYgB/g8t2b6MSslKGc61S0X0C+Nvo65HvRT/rDhdbmIIjVZv9vSP2n5ndejRb9cKqiEF
twX3Tcv08mx4y8GJxdXnQ0epBDKVxybnUEtt1AkIsFMqGhlAJrdEcDKYYTVAIXEzZ8XUkU96wBVq
SNSF+V1eciCGWJ8bgAz3wrnitBIF6oQwNJ5MsKBbBWvvQrCJIbRXbIdAWeG9DMZpEHLnSrTuEke+
TgabzsNJEhTSTPnRhMHg5kD32HvxueP8v0rBm91vcAJXimoEDPxx7oduV1qLdkWl58NkXTK70M0e
AOIO2tTZtrtFdwh4U+EpX2JU3EogI6/VAFtT5vThw/+JMtO49DaCQBzX5V7BhvPyqBLDj1CcODZn
vj0cW3QHIbQczc/OCpqjW3HTLObJGdA/OIjv+ifWMCyQqSoxmFRIEdg3VEBHLL8HYZaS4TJCUB33
1Gbr1H74M0wGDTEFwPn8FbzIPxY0mNzt6/r6TUyEn5+WfWfMu90eJMvFG+4pbfxV6xxkACy56yxh
iWFkYC4o3zbmL1emIRS1WVRcGzAXKfJm8w445mxeX3qsuSTlf/gZOwGYyA6fnnpsDuJDbY51s2Op
HQr+nd64u/nwhWlPDarc9095J59w9aZ7PU170ZO8EXWX1euSQqi8i+rFPSXIcFzLNLivdgNYUmkp
ij4+a2K4Q+KY6HhusrjbOZMP/IroXEwHtLv4I4DPU+/O/Z+I99tsuhRBoFC5tr37xEDxJ5rzFjFN
yv7FPd4NAC3/bnT333TCz2VMV6QlTXfWdpUJWccqJ2q8jPyWlr93w/8Dg/6e0JK+iA9ke2g+Htu0
jO34letAwotCwUQei7AOJmfalBIhxTmIAD8fX+i4tHbTXwH0T/jxj38s9W5MOm7XnnKRNNmY8eoy
HAq5AZeC3fCgp6TaeAWb1VMBjctdzI+YFLAC903bngFdh1Sxd82DPrSlCzpBEYUTORePJZu6HMMa
PWwQ9K7gT0tS2f4jaGA1lp500av7S8XqA66MVGkw591l4k12TvSS7szAphLEo6Dqfq5aYL5WHBw1
F14RLuEtHuw55y8NVFvWqlmcodrXAlWFRaL8OboKSZCar3Ua1slxDr2vbZOsRcGgkEUUfZFgDUrH
sk64yfQtmZPKQk3nchxCsnggMFSyLXidKwuVMUlqApQnItV64lVmhjGr5TRH0ixGrMhie7OpUITp
FrXiSdX8UIRTRQkpcVmRjdRBTznmfD1OGCDf+eryi2LkFSFE/JcCNxV39i6KZ2OjU5RwR4SI3fhy
UFF/4WalILTgkSdbvJbBuUet0sJxuv0+eHZ+pzmZY20BTYxT2pOiSWpmJSafNCxm5Tw3mxC5K4DV
UZk/BmpecI/Dae+x/USGUQMoONuCSOxduPQydauTlROkX4bldiQpPRLBv2d39i4EQV2xVYpm6LPA
gKudoEWV6aupBGBgd4E2rSUCaNHpT128Hz9FljMyz107Not3FySpAJPT4GOhh/tNwek9W/o/XxMp
QH7KvQ5FpGUY5ldDiMLfJQC5A5gDFz+imbr138CiFRTle7REAgd0X/YOQ0kg9JVHNwBsT7NZJE//
jwaQxdSI6ax4W63Dp8d6KNLnLsyG8zxYWgCLhBKe2VqB+2/7iOlm33XZQo6H6nbliLOUr5aApkUa
iAaWmZoI/Gv9dkTtGQsNyo4wwL9ly01UIy426ILQiRiFpx/ttBos3WoAAAHz04f2PzKXlR2FVsC+
e+x/MRa9Id9iePhNRAgnIX/Oo+PSEiBrCpI2MSZo6jq6QEJNn4R/7NjhX34MBkR8QHxnQ/iNyHcw
b/vm0IHiKURabTVp9mQPF8e5iDltEoqY7IozfvB7JO5pc2zEAzgYAPAvHYaASZgxVQHPaRyPYTYo
x/2IayudgAzZfn1eM6gdIuXgMr5cZkQddfxFa0dpgTwb4823C0FUO8w1aul8U9+dr54SblWk7Bdz
17BeKZVb6zTNXwN4dKyY+0CkRxp+qGUmTiTO7b7HM2UZGiGhDCHmbzZ34eNPWws4DMF4tovPIqvj
/bTtaRn71sXEKaA+q8jADGacOyBIH9rO3geGYd0j7nNaQmw0hueWrD3J8U3n6tIIVnBw4gSOLgFQ
4jAz/PecEVORQR/GPlEvlvIMcppItrCPgTCW1CeNxxh3/gMhrJnvfrjlYwiU2BOzeneX92mApB/M
uk0ar6/15xDM+bG+sHsIe04CSMTGPzMHzC/ZgY/vo5bF6kcqDxHcPbiXKr3rPMqqTAj5fh/J1YIQ
DdAYgstRNeqXanpOr41OqzQOmKEdJ4nHxja3yeed3pMkwDaimNz5CZkmKOJTKI3/ACRuIqCc8S3k
0aHYkcVAvfUPlV2Abn0jBJZqJ7JLyOIM3ZKFMa50EY6U5mGQ+cXr1Iez2sNHHhh11bjdjhFsrTAW
l2urLMXgB6RRc7rM+ltiKMHTlCB0GMZiHoYBt9eDvtbsAYJGo2iM6yVM2uTxhnjXuRa1Ph1OMUx7
GQCx0ApzPBZQM43ycGbb+bKIq63WIMnNRhFFsKZRNVstKpNwQYEvbA+q6hK8Uxhhsq4Hi1U6/Iog
EXds9Kbqh3SgJv2G5TP0w33H2tCCoaBr5ls3Xfwt83pVv9fvZq4wT5dc7d2C1DX/i8ZEaTTFPi0t
KJMnddZr6X3dodH12OWNx4ayLx7+gufN1F3JLXJjt10+b+FKw1/v24VIXC/Gj62csQfEcm8uUuDd
eUa5J6viA6HUlw3z7syboGeetNQuX9aNHTvr63gSAnkwhm/yNOloqK+CfmymLUWwJd9qWYdjYfEo
HSUW+4G2ylQWu3fIdjEr0Vo+6fkXQRARAGybGy++aFwKF8QG9AB69IdMNdR3WFsGXCmWGNI1uwgH
85tS+0C6VcCvYRm/qWKwoq20XiTH2Ug1xU9Ml0FX7CsU+7+1hNyLE8GUIZRnMpiC8zGTS0EDxsxy
Kf5xjBQRcKDvX71aivnFNvGSkrhnNYaicneoEDXUKT9Gk9mAkITH1Q+2rnuubTF/MAwR2VBvXqrv
zTCNsqxdWIt1eWlDzFoCwB7xs+e+duGLNi0vpFlwuq+gvPuFTT7bpvYb3A7PXAr/jirgMPGBtpIe
AJOkDxjfUriqYJ75IR/qNoFk89s4QKRhNwahKpYTfAyGfSC/PH5NcSItTCcrnmWhOEkJoIsN/fea
GLu66O7dHMNVVBzIEY1hnj4f4RZhUkAZe2njjR4j4h8lD79vJQ3bDk3ubY6bElsfwT7Nkjpv2bEo
BqVHE2Jl4ILEJx5bRgPVI0iviPZoeSQLAIgAxQtoWGuP7Nh8DyEbdHMp2b35ZHak0jz49F7jNqPH
KUwza7xAAzlEWMpvMjT9T/0RMlzzSMLMjwlU6kvvJ7LkKRwLba4SILkvo74IxK9ikshvkSDbA4Ay
UiguimX/FHiovV5+WilnEwFdvun+5E5njAxFWBaL3MBSFACj4BrKEtMNE5yp38+i08j93QC1Lugg
GRMSOejuMXa7IXyCu2PENyxiTYS+gqScZ089pt1zuC7GD586cpJn0lw7AnY/toiybq0WiXIskn69
u7jBZC9/CXhJa1oWQTyBFc3HnWoytmAat/PnujY6ilcaC5yTiHqOV4jxdUPawIqf/j10I5z/YNbx
SOZ1LVXGgjo7snlxEy8Rma1NtzhgBLz5gbMxnk5iGMJ8Ibmdjpj0xAQ42ZIxNPAgG4sPSvgXX1tX
QN7nyuPS7V9Q2xgQJExEg+Hi5WGbnk32RdZZdiWVZHwIuvL2gz3Uc1wj7bdYSoA/32sduSpzeAEv
XnqlNYvALmywVJ9qivP5io50tXmY+9DtqVcduyLVeulUqhuTc2iFB/DAjgtMi9WKsWHAam2k2GbX
CfX//mU6yz8gP4aKCQQjXXGkVaHPzdofK50fpzYOHOqbWcTqEq4mBpj/7sk38kEHnZAN9chNIRM0
MVbprKPA7MNHyNiIBo7aVhviFDRgR6uWqx/0rFjHUh9eGiZWG1ExRECcK6hjFph1Q01fG4E0NxJN
9IOaeyowuQ1JykG0fNNQBxZuibVHmdYvroz4rv+QOq3cQPzZuZdTPdW73tCFuir3Icz5rBhylkAY
GEyef+fS0ff2NQOI4iNhe1UwRbFvIIxdg7fRJuOFWpuMbxC7QJiikoj0jML/2z/fF2qd1ANy0gVv
u/RhYmQDY9h9QlT0y5fYKHUkLMdjfmmf1IBZESzHAB9ewT6a5/2PtHBZJ6WyiV0F939AeGnFeEj/
p/PIhuVKBUw/ibN+QzfeCn2AjmQ+v53xt9Y1qRN+Od5mT/qsdjj7NQg++SM1ZCK2bz19xxn+ntq7
1AusV8Bd2laUk7LbXogPl0JUwdS+uk/ge7Ai026IlT3r9Epvc8F49QUAzl3H1sQguED9yXUtKnBG
5J2NrBvW5anJ0xVFIqWwkD+ivTbxjFG+v0EKd/tpUVRI1FwNTkmcbcuhLEe2crpbXnS8FBaSmGIc
HP7WEtXvC0WZJaKCtXWO/r3FR7jK6fryZ57/mRlRRXdruTYWyppRMsSrxDR1pZ2ChzxSHtGkqRkd
W2fU6/4mrcjB0OPQfrWYtsCqxxa+efVtajP14tFYcZxS/Dn6L9LAJLYlkucMvoQ9FK+1v97ZupAA
TfGEVNEhb72o4WcwugxEzhVTmoZlPFoJ4g8NJOw2dmjhZ5fVGNcdp+6ADDh8urStFJX3AS+8YPv2
KzSwQwiELUqokLKwnO1/dMadtbBbmzSHNP31wp1WhcmlyU/6grqhy3kwEm3tyKapNR99agoZQDW7
XJQ+P/Lg++EA/24BOhbswarnkgl3u1LAVsPUMesYby0+NKcZypKoAL3ZHjq1IHV8E7R/fGPwbgrq
Nxbv1zWJ2PBI3SFCN7CjQhQR6qXuwYCyPcvNlkG7K7AwEi86hqS0goLwSSeI9JmXYv4zlSISoRqS
cstKSS+pqqmPgmq3Rp0o+FKfCodjsPzWhk6APoxU8MTsR7Dg/xuGPknKkKvOvEmb3QZKaq4I7YtH
LWOWG1H6GzhwdO1p3NRGyH3zzgYKSA7Czepo6mJEOtJw4yV91W/ozusIwrs+KJLOZzXxrbF+gEG6
zKiuT+doVckFo6pqM3lhamEXKsRCDkpFdBdLor7hilScpanG8Tq7/9TSdhjmOQ5VaJywVlc1pCUC
dwAcWJZkMBkgu8OdAKpmp/4I0Z7J9cN/26gwTa0/qD9pUrYgHcGWievMs4orKj6w8gmTIKHRNBK7
huJVKLwGjGUa4+fztE5FCXGewpAJzGcbTpXCT6zFb7BqXakM28JXqrJA6bt/o/Iu6fcToIaCYRB8
HAsuF6r+qLw7Y5vab2v0qMtOleDAPcWWEe68Eex3GPNgMSO4WIi/eMprWH6A1uAYCigftCDc+Ii6
ekYmdd4u5b5b8Idkm9Qc6g7of2BQCHUqZbAIZ4QWmUIQBGuXkIxwqfIqKE84TFeBBmk/s+rQHNb1
D5tEr1KFy8u6YTj5sjdPLYoBB+s6tFnhUarByD9urBoEYjGotEM74FrGP9nPEIa1b8v44p90cUdu
pR27Gl+ITCotTNYKg+dsyrGFrGKjDEWvK0fL9q1OECUtKMXpjNoaZmcemeNS8uOVzk+vKIOvHy5h
9uztwCjUZusHA5R+GNwSwnWLbDI5EqWnrYlUxB7rLh6HL/8bk0SeJIZa9PqI7YsJn2xi+jSjPiPQ
7FWAuEwYKP8Q6rfRkfXozIzgp1WyeUg/jIWgF6rsp4khKXqfrfZmo64GoTgSlIiKYqHeIKYgEYjy
srvEudAxeKvuZKzP6+M+SOm0NzLfohlwMEzRz1zca2xnsM0HzqJcELjMUzPIdc4RcAMRC/q7px+v
U2KjC1fRhb7JmqTlITFmAERPgno75Z/tZNiEXrviYVLCvG3d84Cr20O1jGYdlkSWpnTtupxVb16B
ch9c6x60Ovm/iuOQVj90OYGmqHNV2Lzb61i5l4aVnCTnrh6WMR3+BpRDO+v//6GSJPSvBUquFMu6
2kT1Kk/BCBhbqWelyk0vcg2RpMIJ7eCOo/utE0jjl7mQwXrRXiQ8GxSwD2LdI24YGepin+jjhBSk
RTaiXDSSzWnlLTdSg/7Z4WN9MQ+pnmPK10P/gKJPeBdJDbZUsyV5R174Y0qxaUqkFqDu6rsqRtT9
bv2Jh/UGLQdmuVENFEBn8YwTt8vG6GT6DcsAlnrp1c1XxIVKIXJpTF0wX2fH9lWXVBn1c8Xzw0y9
MP6Nw7FBFcvUBZi10SYdRTptiQU8wbbhFkUDuXmzt0frYSwA/EUDRriyEfw/wuMTXL6iIifgksT4
LfrSbOGI5UAbIf66kVt2+qroobKPlOztXxiCA59ofearYrXjMYmcwVej/JV1uf5sDnwcuoiSzVue
edD8A95tNaDC378nBVBoixg812z+JKaRlgaFhSDjCP20vkiSBZdjqwD8uARc1MnMiJ6jBllg8TZr
XNMqDr2HZGozSvHKpFhxYkq4DJo1Ad7NOdlxy2Q4J3/aHJ+hg6Y8Jymsa88YogtSE+MwuaIsQk2C
+2T6Bl759ZJNPl7J3sxVZdNzFcaMlU55n0ZpCJyV3GouXcfQhb4zDRTW4kzXKA2HjwIdfnUIaLLe
eHpqEMc0Da3NplCV6yUZid0wNLXWYBGctrkJFCgjNkCysD8eReDABjZRGetAb9cTmNWNvzUvaw4g
IwjbookdiMswUEuEF9YuJ+fh7c57t/U9hVUbbEf0aFnF3sCt7dKlGWN8nZOwD8j18ueXMH3yJKrY
LJXLss36Ii9t3g/UQxODXlgTiOCucOUqjn0mGA72/EXx8I0TVUIbTqRy5ms7LbjR575VvZeyE4F5
VCS7O/QdgDO2AV91HGAyE5aVr8IpN/e5dVJy3CZt9Q6FTQ+6ZtSCwG922fsSRhq0x9V/SN210gtY
2BJJQu3K3jb3BYhT1JX4zSgTG1LYbIM3Wpn7yTqJYTL+9/MQLNiBZpwF0fSX9x1WbwNUVxqG8o6j
PPqLCwhcqDk5Gv4Zt9mDN/tEdcMdQa0t+ys513vuelF2KdLRfIg5ytKVIkM72Sq72s+C9Xjyeq3y
mVNiMew25lKnfh1P0kLplNOB2Oea0mUHzTiArRlJZ4AfaNzgmmHOOawLtR7v3c1SQ4SpLYr/LRyh
9B/0up3Qrdb/bfRdDNtOFkPB3IsLj6OYGKz5cijmA6qPvPeiguVbUdx1B96GgEme55Q8w8a31C+F
ZQ8kHjcTBkMi+qCCz7JL3iIIBIAOomhelddOSF544u02lPt0I2knHNNW91D8PPrIZFupzAqJFVwE
46YlQ8iuQQKd6sPGqjTN1aQSUCxNtsF4HJwshnM/AN77b346oa87RELHCCyTXqfC8/lDExWl1XUS
UrDH3JuK+IdtgXQoOzrUPqhSuWOccTSNRxxr9BaezedM/iTnBHbSMLFyDJOBDLFCF7Mjgi5notCW
F9EZsQIJ/qffaOJkXcuCZZ+wZJphUl1t7DF5CgWaZaLb9QI4QzfyP5wvYFT7hEelQ/Mq4LLbM6CF
I4VDs0sG4HirVlcIHE3LmBQJVVkAbPZkT5qvsZjyQcVotvI1QKbyripCzoRgH9zSXcFdKZLakeV4
TJc024ha2RxODV5XkVKmxiBtx+yJQZhe7mJoUBp1TeJfH7XiYGanrNodjlRXPi05IVfVLZwDGfqN
6hDYLcV/pZK+erGq9JVAFGyB8YiMjKoVRNugVOtnuojnHlCTuDl2YU40gr68YIrgkPiajiY44QWJ
tlGd2GlmbxDzrXlTaUuq2eLlSa/Gm7LY1PGwVeioTgpX4flj6OEcr8zwEC+PWWZLZHXeeJOk70Tv
cW42/Cikl/BKlGh8JVBDC2G0P5g/a0UoMcKznIh3oIE6kZFsYBJCtwz+KngoXuhvVyvSyZKhxMyH
5UWcE1EmTisi2ZiMUCC41taFdZA1LvFUw1dhxUSQkLb2CzY2tAxuL7ukQKZCae4EjsUirRyyf3qp
rRMUDWMjEbJFDLnwTfHdojiLnHLN4Ruhe0QsAeymxXZe6TuzYww173yd/9mrNdoRLeibbMq4UwAY
4mX9eUvxEkmyNxQrRgF+ESP2pX16GpgU9i8iY863jyzZP6SukvZUlMHppvKXyezxomJvxu5EYLGI
Si6+hJ3JpcsMBVhxIpwIO+Aik+JuSH6nZ0YelHnrjBWYB0gpbE+RK9Cj1QTM0z7MTeIFQBvfNHkw
pM7JSdxVmN3EV1/A6v7btemOg2x1bGY4X6HqRFAGgdIaObVu912cxI8ta8m9CBL7KEbMW1woXuzg
XhjQeGKfKK6ZUj8XzxbSgIi65V3E3d7R06Oj+jLW6TmwNvkSYEtMr9zkuCcp67FracLwbtXkAALA
KGxrldSn7ulDvaqrAYoGTfjm3BwbuiONpRoj/Jg56aEC0OLJuWj0hfEeko7AYBMsPv461aYCgPHW
7TRg/JX0RO1ZPOIVXpE9F6JBdWf4SXw/0KnMEHSLeDblupwjwxRZMTk1lMH6na5meUsuSDYnDVP7
rnLXzuaaM1dvp/dfgfM8HcjKH9v78tupkEHSZZGPKMR+5t1r6sqx6dlGPG/se61v4bSi5RZYh3/Z
p5f66f9d/vLBIlX+JzKk0ww4n5V/BZOphIVHWdHmGNTcQype3GcnL/FsnCN8U516OQPxQL741xF8
WBM4hwAK8erBp5L+OECtbKqPIBRF4MUtWXTA12kPwhfrT8iL3pT4Tk7wvlPgSh3yT2P59LnhhzOH
0q6U+UXfhM9cESQOk6564FFqfXTCTL2Q1dRptSr1K8V+dbdyJUZjban1RoiADB51P+AhVposjsKQ
dwdmxLTH5PYi1Sc12nhVO/Z6RuFbaLAfNzZOG+WZH+dHIW/iSroXSV2CrASwsmV+LsjsluT2KiWZ
eKD6CON/qoM7/Besl53wXGZFYSW+cvXZ0CbVcoeuvJUFf2cGdcLPFJREbIhBxA9oZTp9Ch0x6vJY
RKquugs+OW9uMdYhlVtbYhxBfQGPrRl283eCrdo1wiWf0VPJeKdYp+i/uDX3AqdHzIoktAqAfrzQ
vno2xC2H2/CMg3u2Ixk+QcNrd6DLu/ipioTyLDJ02GlyG5iKCu6pZJKJsz+6/ZSLfFXD2QC037Pu
qDL/aFQs8zDxTSwmDoC25GqbhLTVHuSDVVeLxeE4MpyZGobewp+4mI4zHg/2Uuz/T7JVlaI/mZjr
ZWhD6K83wEJxZeWCckw9ObedYWCW2YXRQVPme3ojtllt46a45bT4wHKw6HjReYG5v0E6gMcMbqm3
sx+2XDva/LjGeLilDXIMw43QAB+wi3zAF+mTWFc9ox2eLcCwgmCvcXM90YhoR8wolwLp7Z/j8yuz
JnJvZmWDmUyNAvB5TWoSDHLs+JOMoF3FMuxVgHZeMNd/V+kLpLmMSQLPCkrLZScMX24Tu6Um8sPf
WZR+Y683gD6xiV3m4EkvreTHnEOP5faYs/45XmdGhqVUwGt0iJLsGHplvCmNj+90uyE0XsizIq1f
hdAfHIe08c/3dUjImlJTjOboQiPcBlfoLusJteJXQoh9tMAtN/ljesrEDzoW22FtqH+9dcFAvo3M
bHOFaK/It2097eEMp99LfMpvOX2xxOeTAleP97lKnYcOXfQAVV6ThgkCDBNTD8O1aW1d0GxcxEzD
hce11k/k2x5t7XV31mXiDb90u6AmOSTOSojQHqVQFPCKXkSa5WJiMt5KFZWAcxXHc2TmWJtUz5j3
YIuvaA==
`protect end_protected
