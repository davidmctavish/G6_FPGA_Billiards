`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ql0Ey3vkfkQja7unzC2x8goyLZRmr5kNKdo/Pds8njR6urujoaAruCnKQRX0hOWwwWpQyh7LGcbk
cBL3Y8e7iA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c49Bl2DfcpF4ruKL1EAM8GrfrsZIyB89jJi8otP3SoLZ24pZgCQxApfea5aD7kfLPBVnjK/ZT9nd
DwsphTCtnxt6lWZKj+1j8mf004hc+gvTddMvZxbavl9iXCfbkqaF5kyxR0XQtBh+ps2HmuEyXrvr
jPjk92E2C1PpbQ1hP9Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WsV2Bfn4pvJXcR7vtWn3MWw2FdTHAZp7nid7u2RKDzXewosVY8HqxZTHP7+IqLtG8FLlXZoIrpco
3lMZm2scKLnTQGDru92yKl7S8gQP+i9XvkiUGwf+2CdEvkkDvMtvdvR5Acd0jZP+4wHRojoXRDte
u6FjEI4Yj1OTzZfgYBrLVAk60ibuZo3vjToT7zFprXpdPffMO3dKcVCHgD0j2wxAU1KKil0saXlq
Y7Gf2uKtGuWJX1jEIN+VYjf9lhK19J6khnHxwcJC66/xLsLrXC6xpCQGpnqExJDjWgsIvvZTGPyL
Qx/CF4aVIHamMvzeOPFcVFKlcJyJemowWEK1Rw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZQO9nV/LSel2c6ZKcXCMN+zCvoXbe6NCTqbBoX56VKzlAFqpiSpZQH9SX89BacuZhOG2fhhdrkWo
xdWuTH3KmgFeohXf7+jneoj0VjgkE6XRJxAUM1zCFhDPk3RDU46PTTG4MKqSl8W+0B1eVt/r8ibu
VJ38y2m1MOTyUBrEG1w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
he7DVBr3s+y9UDHdMaYoty7quvHMvbrOXKy0WBeGrQyjvkKYgYIDaMrdIZnhi3cho/UrUFaZt2Qc
oA6SKsQ9uuQ6EFAG1Ji/jzo5g9qjju/0zdImzV8ITjF7qBId/vleGpM9RghCNlBHbOz7/0DDM6Wo
ZoBe6uw9rcn7kMV94yb4CRCcFxkoErnWo1dBBAtfBIrwUed4scS5cbMCVhLCmETe5RBhrH400OU+
2/jBC82zpwlMrLFSaK2u9nc0aeQbte+A4we0Dk3NNiP+mTWhEiPt/1RBz809EFSzTXiuc3yU+Cwt
G4Buq4zxDgWdEuJDvzYqUrQwU7R6Cf+U7ay9Iw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9744)
`protect data_block
H/xArCsppJD2TkHjW3ivjAK6o3q/vl86gb1P7fU9wpof0QaZ6eGBX/VBRfQlh36RhcHj4EDMdzSv
IXwRhuIFnjUdPgg/4Dm0h6RisQ8fXhB/eBpkk08lIRzI3cgK0l5Apw01BEMYQn6YiFZShNdcslOR
ZLjcX+9TuieIj8vui+/8kChUzWcitzpCpX7xduRekAYnQ6FLNwLr/tRjZpTMluaczswTBhFBzCJ6
wb4KI54eCzzMouWbUgUiaixkkGRmHVB5hqRmkwctILDXcVAnPpeK82AiibQyWRo8SCxV4We6m/WQ
TUpzZkGMO/eA5XIGPrEfMBZuZLQtDqAR7wG5DT/WX3BOS+jhrd1+m0Xm2PsrissFvlZCI3KgfDhP
B8nS/BRUG+eRxiKDVSB4/lYMjjIXmd4W+ZaiRHdv81mtpeUFQzJX21dKKLvEi0y5Ov/RHjnNyQNS
Yj4JM8XxZ+InawMgmIS1y+kZk6kE5aRDl/g+O69uA+XCsQFWy49QreamyBy8iv5oDS3WGHn3TVHn
AGkJsOIfLneeSMA+MRni/Kh/URvvwGbfKTg17Yt5hi125ZCmD1YIZThQw6mBGpVFTupgNT7mgE4R
n0qTe7QFiLRIcEgouBeEBvZzTf8ofwqK1eEL12GUIC+fhIG4oqXIFQtDy8dx9cL8BESNGxMvXOnN
Fi7dM5qEfdNnFQonhDaeeSmm03xqz9/t/FMNWhWoWwHryNc+ADWQbYGCdVgjrA27SgF2HPzt/pLi
uXDbONhp36rR+P0zekHyoh6HpknHTtBZhn42TIlhEgFyGPCgcGq3bV2g++mFYg+8FPiJ2mI7Lvrg
o7nCk79hUFyfw9b1wvAxp2WXLVfmXcx9g7Rha0fCnisIRXDTspy3o8breRRv1nKG9JHKWmHUuHXG
RkWMZzAj2UrzBATYZPWVyEZKCPyYlly3/hD0rAdWi6dDI2zRsiu+iG5CbCiVf9MJ1lA9OpLbAU58
PpVFzsZvhVBv+GOoV2SqR8RYwBx5WKVZkcIwPGUQN1M+XcA+Xc3omwKi6PIELxpQsZhYRRswGGq3
fzuWsb1olwj5/pTzQja6Hwu5Wk9+Vmd5gnzrW6/wlbmym6rYU5NM5ERdZL0snSJne90a+5xqKx4U
rTRYXKZptihCOGJrHcgK3vU8g9VCdJofTUvqSCdxVWqSVf+tCnSHVqzzQy+Ztag8JFgygwlWg3fs
QjqQMjgVBa53OFRqpDVzabgZPImKIwsg/PKU49z51/hibvTFVrDHsdsaR3Xrmq4Q3MOhc/hnId05
pp6aAYtGZwt7OnYQZn9caPvkw/O42D4Ayr0/qRbafb9VC3thIEcPZxklvXPcRxCWhLybd/Uei6TQ
FTX9O8KMk0OVyPlJR/2laWnOPHevO0/aCoevGBelm2b6oqxWY++bsooee0XfFKoHUgrjB+kILvI7
1KNsBTagZ1IYAiZgCC8hMaXrUDVFaLbFqUHMb/P7pYLMlP75yAgXELbF5LlS0fY1ELC121/24qO8
ZJILLdzGDHV2ILQ63TQkgoRirIUo2rXVPr7Rcg5EsvW/S1BbgfvURc4w3je9XT6YQlafixYMnAhY
syFCaeEPDXwgAOAUnReKM3Ut1ruz54JwEfTtDnq4loXKR+2cKUwm9BwpXI7VMHaS97OfHJnDegMc
EsxNhJcqfAuwC69IzqpsU8APaHxnKomEAFUkYXWd6Rss4tkeZSVHkmMFgkNAevomnJM/SG5BESvd
s/PMbcdVeeFel5LrFVNOCmd42G3Wzbga7nroG8XDbLvkYMy5bJfpcPEUayTdwQBBIGnk3qR2c5oW
yU3+QnReF8gUyw1vajrFJb+NWiJw3Ucq+gsjanfof7uaSfeqWUfN8DqrAR1f6slEqprONbh4VQvR
ZMaqemqg1ZaqTkQeNh+XcNwrPrcjTi1ZSlGAZUFv1IFa6AijYFHZdCIobdAqp+nw8FX/h5zIFWA7
i4GXX//wd8dnVQhvPgGeZbRFFOsZhDUgXSF+XIrkvu5k75YoCtcHpooCD8A+67mrSP/Pof2CnbCx
1PirPMOoHjvnnK5XQt+s/LtEpnENZfKlTIIEgf7gXtc8vUrIwCkb4My/OejvF6Q2Zu3DICTAhA4y
l5RODTN2uee2xnYApGlHz2aFIfSEJhAYq2i8cdfXM6ZSvN9Zn/TbK8byWLs6t4mh5SnoHpZ9aKw5
BXEwvdB3EVNMMPBp8wRb9K++PQ7ie+BBqG5H0IZTnDJqPYUYqxOJOE1akItGlGDBa9wM9X/POCkB
twIJqfZjKvrOMBpUloZ4xNpZ3+0O/dUBew+b20UpjFNLu1cM8swSh3Wla5SD09PKyY0/Ry7S7caS
QIEPIpEG/6CN5rWfYz2BywrVaUWvJxfoM2Srn6tN8vYHN9dbknTcZs+n1y//aGtRe/bjMel3eLn6
iTrBaaL9T0n/GY54wsjsWo1crTssCcyh1agK6TPh9WbfIf2ItLgaxAF6gz7oQcS8dx35BhDP9nKP
Ht3OLnzFHwfVPSJuVeC2vAK1JtPXVYCzG7vnrTjpdfYeVoPCCAJmxbxI0NCvvUeyrraXHIbNrlE7
1/tOMgn2GPriXK+qMrUc2tzcr/sBTOOKHN4Bs7jaR8g2m2yR/nMdxrVKhTdxHpgIvweRRL2BTUS4
xkXR/aBvtpiujG+cky6xr1QHrE+bWXvR8wIsWhNsA8c0cOAleoTP/YATs4C2FVBojt6ZiljlsfNq
RvEMfmGmHZLFmm8j9HOoObywVCkek1VIB5bznea4jVvQI+2dm2mbvlVfbfZwx50GMY/u7YT4XBIl
29Ly65Ir6zcVF7SFdhUMuNSUvxgGSrU5sKqGW7qpsD9g5DSO5ZNZjwo81iNaeqqBD9rjoZJXmLlE
Iu9NK2fgllCuNnWW2ZO66t+QI8c9VGeUN2okUcfwfXr2j+5GF4I/4xvzS+gnONvqlD5ceVmIkc1v
Eps0LQ00Nj262GVZXkC98MJRlT915nv4n7oONV5qHilvdBu38/Z0hP8Paz1yrBEZfWDMM88HFt7X
mb6mrPMwV2+HpMQ7luP6BFo3VPiWBQOLJ8Kzg3GJw0ZfnMXeZFbcRkbQU6v6KkuaEHytvjPql7/g
XIYHdSDdpoZW/kxFjwLFecHA58g9rr1/Q2NGAjg6Gc8k3xnuD6lj/XzzgzNG1N/GMD6bgrzUcWhm
ATPCNMTIw5AdwW4jE3gOvu3hcYzCbTeY+Xhk+bkqy1uS75e6w3VtTb3dnq/D+oWu3XVLAM3fSxk0
hxcx9SsT9cj/J+6kIw7zCpxLiWcG19GW+PzoXYvPuVKR4R97fxubD23ADzUgILgYmTQYmTEPaOv8
NnRihcAQvUaU/8ZuK0IItyh0hdrZ2hCYTtDS+AezrtrwOClsqTcfIvf92a4agLyrG8Mjra5sHQEn
xWJLlAfIXsdpsHPAl2kvFZnwIoarRDDHiBcDIXDRKONZAuAuYoo/MJlB3eWYiavP3On4zPfJcUE9
2xR0p9nXPf7XocZHOYXEnH88ZJPnuXmwcZU+UsfpixgOQgz+7ZuLySjXZLz12sj4yveCXZjt309d
S0Fbfded6H4wmkfpMM8OOfZ26F5FInRNJIP9v08kvVl4OXinTqy0XNlU/vLJvxca9C1ppeWcL1XI
P5JlBdNDXLCJyUqIXQMuAncanqp8rBqnd79TN3snlR2JbOrtoNk07dP/qljzFXhufPZtfPGVtxhy
ZU4dB86wmYRBOcz3wO3DPP3w3thCzt2NchlO8zQ6jzdJ/qZvXGr5iPGzqwNM+IbbsoBGwczLUmky
WIBMJ5dve0gOAU3x5kbOjbmh+o7QyDaaQxP0FrwF0nQ2rjWrGLTIxz3cEoY8v2CExDeTJpm+2uUC
oNB2TOuCDMVfmqIqVpvI268f7N2LBMBP7STfOS3BEdKIJH0bGoDd0ZiSB9WIWliURroaJCoJh5Cf
Tadq3/ia3mB7pP/thH1PuSFgSNUKdoqRnEC345vekPOvAvxMareey45z/8jKRkN65lEU+N2vFEqX
nBrQWd7qTdqyHHiwX4CO3x4VMH67RxCrif1la/HObNZEj/sB1sHSIKxcKz5CWiPxtdsNEiNiU89U
BIXVOGzQJxlEHvpXwxSnPdpaXTa5lNJxohS1G7heFqB3UqLu471PT3hJ++0PfW63mCh2vmx0lZbi
tM0UvEUIjNp6gCm/H++VDOZF4W3uHRZnllEUZwySf6Q1450k5ivqUnbPwWqKKw/2Ir8G+gu9SpY1
2Z+80iM+7urdyzDA4l84GMBa2xCvjwZNtOu5Ky1h2TegurRf6AjKuKaItCDOrJUYUXVrn1wO5CpD
3w80FmgcqTzl5+wVHsZHw7nOwvyKwgQFMI945k4D+budZqkSPf2gxsa/yEogYrPdZt/hUlJQClo4
t2yYAgrqgV/NFZag9Rb/84mjQvVX8I/bEYCON45aNevBZR+Sb09MiBq0yPXPGD7gFq+f0nY9Rn27
HDCJCICE+H1alLzg/lMaxhzy64OkH7/xHev4R4t8QfQP3o+5TU5v6D3TUSVbESnTSy/KjcMDifg5
Q9l6W5XMjrLkKiagD98ruN4TGull/KOd0Y0y65w50KlawfabBwV5PhRtcZj65wHnNVIsQCaBNDtc
IYO0BepEEd6+Huajv1XzpkPKmQpoOlJavLnYIjqoK09CgYY1T7ndqhldc55UYZy5WygPBOiGRGor
d3swACcWtQelXDXy0bndnjqTDQCoSOZKBt6iG6l/ZzxwTNemr/mFkagwkQ6yywPsuMp7ptVAu/Iz
pg7RSzYOKJpz7rCE2B4YQo3SAJeoL9dXFpfzulwwkJIjf5p4ftPGQz/rLcDbV1b/ZLh7+raTJP2B
w73/aILZrvmf3K8v00bWyvOm74R6ZKK7Nrsy1SGgKGguX68DL/pRtBV6VAMF6ADTzuhaiGP6zbiV
5Sa7t7XuKcVNs/V0k2i0/p6czadkFKwL5FasA4q5Y8+z0MiV4/p53PEnEb7N5R2JWLMjEa/wGCMs
w4pMvBtyjpMyi0j7NGDV/6KS8mc8NEs5LV8QkZYWIa/nYCMntHOlmXw2uHxfnDm+aMx6dCLbm46m
89jeMpjjnYhlQf92taZL2B1biTbrSbzAqIl7dksxcWS+dIxs6OYQZB4/sNqvqgrF8cM2Big+8aNZ
JVAHbJyUMEGYcS5zPIhJ0XLTOZZ2vHMn7wRd2VKpAbTIXeM/clonyGe+j6YSX8TGVmqh9DOZXVda
Uogq3nl4rWyxpZ1fVPL9pIM+lCtR9lQIAInPlMkIJaSURLgcLE1HOdKoB7LNKWPrZy62xzt7EW8/
dm9+KUXCKNTeOdnZDOONt3WB61NL+Ibp9ErR3dOdI3Zd3QA35FEskDTm2McMLfRGqDl1nhLn1/Ae
88dKwLtIiTUx2MRj+rUu/pawp/5+DD+CNPcWtRpk/hnbSodWKj3yunjW+UUD4P0t7mxyqdAIO21M
U9ltIgjWV34PFwmKsSN5a98Nf2s4atNN4rF5fFPdHyRiCD5klw1FJkWuMUPznTfkjS2L/TnAc2KV
tmold1J1VnopcN0ORMBY7oHt3t9e6qiPjCNWbiN4j6w3koEZMtmFvIWObw0nSPn1WXTiuFZAyPSd
pCPymlCE0fOn9tBMhdOuy9CmQtTC9Yoret5NMX2NycMQyxG2oQL2/e7bI+Nk9Xf4S8aZkTSe0ou3
xCYMok0QKDXz3eNgxHSBo71/tsiFsjjA2tw3g95Bou8qm/HwylQJUY3gfIHdNUiv+4sRvNqy3KIB
+EWCJEQvMLOVpVM/vgBkipRU5XGm3OqZMMfmkEM/+OeoN+QbFefvJaG6QQW6ElkdFkH+0ZdDBmhR
uJ0Mw2Dkjcr7+loebvF10+GU5wtDs8sFJQncJPHTKOWXL47M/OwS0GHmcX4PnGxb21TYfXN+tjZs
JlA+WVVf9V7wUA8qMSXByK7Jy43SXzwOVtwmKkm8LS9PaaNceXFVqDLYiMlcT8jgU1Dxh4bDCprN
1lm4YB5SI9K1eNthen3+tm2JE4txzN7exUbCDBw2ngojAgzmlRqLbn+rL2wFAkckHkpF1pueiNsy
0wD7tN5zeYaSS9Vc7Ne9u41CBvJgOYAmgI4ZPOZf7f6Vf8cd/lAuivIJKGMzYtg+nAje9IaNEJHJ
gu28GDyht2dtLVRI17HQRXbcZraJumYq+h/S8nnGdq45xt6EqNmfl1lGpvkPZ/5Go12wJB/3xxst
sb68MYNTqgiox6il/IQE1AD5Msq+PAgsIOV3xtaE2HFN9/IN1E3e7Y6C9oWIST5uRLFy+Ith8z01
jk1MKOlA3BLadbx+RDRdMB6WM6Hr4Mymr7eQMGfJnuplPTNQ9FnkI8vTHMyg2/1eyi4mK+l0F5xM
GRmBBtw4BpEZkTufvc104k7FH0y5naoZQsUkDcGUZI6JQ55KMcHhLOFqIDvZA0Uz6EwLnUZ8AG+I
pynec3WS8Q9ypDjKBBu/W4lEfnTz8aZ2WEp8tQxLZIsufFoFFU0qk0Ks56e0Z4TzmWnCNvvgxDM4
LmcTICeeXAikJZVc9BVew+IiMikql5ljJjXqrBI4AuJdHpNpCZm3VllijN9qKi/7W65llKBsj6wS
roLijWgpNcbuh8Os9NUiBB2Sx20rCLzaS0BS43BJKf6G4V2BtaMU6Yv1AVGHMuhScceuqCDYub7U
fjeWYMRUqLfnhEcx7uXADew0DbI2BspFYjginVywne9XEckyrUyYsWjeWxXMhcujDfKrF01YeLTo
5cjJU7iuoo+m/RcKn9In0U6MjFVgEUiWsodP5lv8yc3IjPb8+7Em0leh6ZQ1ZbEGzlcwSUP+JrWD
CdsVA0m3SHoXFO1n8a/xU3XDzTcSEMkBuFFOs33ffvP53fbTIVQP3mCzypCLm9CbkAL6aJzat0XO
JNaksgsESayHE2ynWXEAAbA5ct7yyjN5V1JKUglqCUlHlOqm8mAUvizltQINvfPk+xsdeE281gg0
TrQo8szjj/lLyAahWO6ZXigXS0TKbG25cYSqnSBBZiS1sb3IwuLzOKXjdGwuVafmLq1P8awWIeBy
g7pOhGPqnqY9mmyfJjHh15NApYeMBW203f+5nC5hHhoLrbCt8CFrC6qJsUikDNMaQmkMDqYdLCCU
I8HSEG2NGqQZfKBLtnHGuX2MrVFhxpQOpVrXuo2peGrxAoBV2E5mc/otkxh06xJFwQEymOrlLA7V
VDMriKU9KX4pWqjpBgCqWHnQDBwgSzZl+6JberSF5LS0FI//f6hfKOymmymHMKnorEnlp+Kr90nl
kwaKT6aCs7Dr9Yme9vUEh6fsCZPIvO20+7BEoPsYoakdxx8fvkHVSgx7BQCFNDs2t2YkSEo1tcp3
i/3FWab4Ur9Bioq9HSUdC+/JGiMCnvVHnpcY3OtVDxn1OIDWfPNjQSavAWUCdPdWuvK63xKicOhv
QkbPdSkj+LW0nWS8EMTPCe6f4uAlKMmasVFOXfWpoScgxWvFk4T+Dszo2xGcwxlVe7+8BzQUwzYs
JpXKlsCVPbzMsSdwWBaijabul+3o07mcxmUyqWpHSiZUBuaaVUOUzIzFS+tcvZpGvB2XZjZ+Dfjh
kiRUocA/maHopBedzTuSyYBmuly0lf0m/3Y36+V0keMAPUUPg3B1aDGcqKeSTre3loS3rk9kDQVY
j7Ydu91/cj13Cuk/UAmRmfMrFXuRGvxvJ/7TvYG4/hNG5uFDDgsYEDpDh2Tk2iyNjjmNamtmVkye
xxE5M7p8tM4k7Z36cHk9rO5jieLS0NwOSJOcK414yH5jgNNgUHJvf2Ty8MlMjrehDKn5ML29habY
zY/4lR/PuXA4e+/SAtTNkxqiMbdpnkREXHdp5/T2rqrZYfVq4A7SqMpYpOVzDS2tpdnuN5sYuEs1
yUu/bVzdhn+/LSBY5SbleWGFNBrtVcSgI8OEMODIE9FRD7rAWcOYBE1XFLFVwcw/liWUaCi+4mKd
e0WJi4xWlvl2pADaG2zmEZRkbXvsi+2EZKmB/GKeUrXYB8x9Tg933LEw1IIwMn7cTqKBJjSD6SBk
wfCSENH4Uh/ekKF/7g3/AKkUCn32EAjnqnh5N1eC1g6AXJlsy3SYSIL2YrZxmRoq6011Nnvjxsyc
E9jvtqw/Y/3nrrl81mhClmvM6kg7dMBlznPB1mhdN3DdVTPCqd7aW5B2owxo7vAj+R5qT7olqb56
LqtOEY6F0c+nCqs9d/GhieJkDFgyz8NL33dK+tOxXJ3rM5sa9EbdQ8V0BWRs9/vTMPdM4wHM9C54
rSUwdmNu/oTrvN7lHDE1oQaFoYPwXiBox4xwD38iKr909thNiPj9it+5p/raSfQdk+cyIbeXV+xi
yCBnjHONWHx0IOooyLXBG2H0PHrNCzHTfurQDK/V7ygdZPN3hKPObfEmfZZLhDWpjwxS/qllFKCZ
2UaXwN3ok1zE/J4BJtH+Cd1dZfmyN+LE6Jk9ck/E48OhX4ub3qmRZZzlHjg0WsUe5+B2dkLhXP+o
bNTgANFb+MTyw6k+5LJ/3hWxhZWsysT4ZTAmGxNFewdo5ALz9TKBQCQpGS1Dwk6sXgjd0/5ZrVeT
YZRXR4JzpL/+wHqQNV7iE9spVTRnP0Qm3ImBWI7jRnwBaMrI4KclSBo4Oexn2ypLtIjk6C4NkPWB
xquvfxCEWq1ywVnRdUxXllwOXFsGl9jBNbEn5phZTqzqbW8f/gg0OgWX8K31pi4fAVQ3vyKQz2+p
WngE42LTLbLft0WEDlvLOvEc/+qF6ta7O5kpeyU+/fiPjWFlcZD9QZJEH33mlYA0UK/cWVzwcm4b
ZYlQBAQ4HmLh3jU8FiyxGdfS3OiRFBneFjwJWr3a3NQJ1EMVc8RbNW1Ix7DQfWL1RUNq+VO//DQQ
wOEb8WGbp/g4u+dHYn+C8ZvILFKkLkKevDlf2Oe2e1RyDYrcnwMp1prjpe9WXbYjg0M/ZF43wgd8
yoKhbo7UPgfR/ml1do30zb44CP2x0kSt83AHSyVZUyd2g+9CGUbITxN7mxJW98KptXijJYDGTSe3
JrRpw3OhN/SfFDg0gVSOfVL5f9SW3nJrIF6dAXmlnpFb4MEZjMZ1Hv6xzfV5iqyhgS5APEH5lbuL
ryZ3sik5A30wUmxRUh3AiH9f1FTTz2Jc2HOyRws/KWD121crBTASKDlOib32ulzknC63RTJD78m0
bsoe4qLz9P5N8LyK8rUj8GbY4eBlbUJCARuo8XzMmvmA2xPof4L/1t0nutcB7XDTXiPld7Ivk6sZ
PEeBHGpcKqrALVea5coGHlQlJIO/gRwWbE0SaUUphCEKe6IPDcvIcvGK40Lkff1/tPa/sMNkw9qz
yskvJ93cVQXpScQNn46fOk5MeLuwlHVYBKc2K4Wd+GmGE+7jQaP6bB62rbGA6pkATWjBS30nT6lV
f7aRZfCPnaATOJ4jxAH7h9pDTPPBybCgIhdY8ykoKiY+67z6209SBrUfWBNWXy48N/3tSB/R/XcB
53FzypPvnvfbWtxLGOMMjbMq+bttl3w0EHcUKGc81jtZLFvw/Pyt4Kz2g/nmTbkhGHDX2o32J0Q6
hnkADuOBU9TXXxnfAxkDqj6LewajLMSsJVvyoq3md0SQZrqPBG77w1gUYANOt9SNPp47Bq5gujNx
8deFqPxoeq7kJe8kAAw3tooqUCvA6vP9FM9W6Uk3Y432S3qza/fTT41sk7nF3qgNCNuOvlml0oH0
HlpTw/3POyDWAMBHaxq9DnwXsNaJ0SOmqyX2cCtw+opkvxCleYoZf8OiCVdVIOlxExnoUOycTqhw
9zR0sBP92D7Jawg9wIIx6ta0+63D4sC213R2wYlD9k6ESQmYL/32Ng43eOOP6JKL0H4wKHgSX+Wa
vxRaevXzbpQdL+AOTWEjrOW3oO8m99k/CWYHlfogFiX0bTui1jsWHa2gP1zqnJb/kQyBF4p6hSOK
u+5iULp5SN3LCiX+dHDeW0N+mPFNipw2DTm6Trn5+XHzwFp3r1lPd4j4cxAKUqgXBCW5Keb30yxL
lJHW4yxwxWsOmP0ojGj1PEib9BLWbBnH0Kk1nBaFyyOVJpZ+05NnU8ICPewZHQdPRI8pOWiFq9Yd
acIjVLt3BiCta6LnWyUuugDZEnhn61lb/tkTClmREb7xYG6BmNx0EBh/HDJIN5LkKo77NRq4ELOi
HJShA05q6/emP3r4+5rCmz2L6viJg9kNB+7c2gWARGwgLgLqq3IXB2hJ37ANCsaJgkboRJ8+Qzev
ZxKh+JXC4X/wlfr0qP95FJ8ISh0u8ovq+2wws5afYGZKzgyImCwW96hNO5HO1w/AtviZdkiyM8y9
GNJFRdx2+1phcvuRf3EYClNgkMmOyzxh803g+pGANxmpHDj6rD0K1VxxbR+SN1or35/ipvSgIsLx
/j3KrebJauxfc34EzrH94OgzTJUM7CQrAOyN/uhVWEEnub6Ve6dhX9+CPYy6JtmcvM5KbHqvwwnZ
EbdkpNn5CpAAX+Af8k/7KWuNI1LvwiFRduL+tGYrYRCy+fqy5AAmswwrE/rMdlBgduFSWo72OYoD
B35jw0ZTZnLnwFCriEZWNmTPOxuego/5/vOd0XdtimOjI8sRij3y3KoRWJE9KcQ6pxmbHMTwgYuz
tbJcNnteyGhjYKKcB6QpkDSlnjtie6Ni+XWHLN8QjwDwyG0V7hyNvxvrJ2ViNXip/riAITrVr/mB
cp3LO6hPT8B6wobAVzEkPlzJMJqEOiZRs1bkmzfBDvHfTzWqIA0IG848pnWHAYcdb++UEzac6MAW
41qvjC5WX/i4m7Mlt2ZkOK46mAKonLznuHjy67/TVcmYGjIlZqUujp6wkgWufxBG3u7wKoKGlODk
RokFtgCG8AT9S1v9OiGY+mcjJiPtHOTaoXYWBuYVyQI113DG3IzGCbB07KnzHLT49cljYMfbWiYk
bXSGrMYvbRxHuNXJ0DLgEPmNRnMedSIGoRnJg18giVLAg7Mol43NVosMheI+ZQRBSpqFEL85WyZB
DtIwswYmY1bQcxwb4F0hEWoE/OTIujRkJEE+GeNsewqyul0D7DOzhBDbC2W49+eDtrPp7miIsYSM
ysJF2na4tgAmm8JIN4qdI0wfHe4sqfb6OyMgvK6UVjibwPw9EpTecxnnlq/jla2kdUU0KX8m1Ksk
nNqKHorrQ5Np6g3YrosFwQd3qTIufjxkxZa16eqdBULdoizGbXW1e/B6YoX7YeLQ+KC6Emw64Cin
PWdgbIh42mVI6LpdMmQwNegq521rggjzcQTgnjeJGVx9oHBIonyV0uUWpuYc1Vt6AJUO3pugmqoU
uWzP95cCKCAUfZzqpSpL2rjl9o0mhp/S5yn4lnON1IfpzHDjx7F6OiQFOwSSoNkdSDmEX89T+YfX
r7SXjaZ2MOn4p3dbNEXuE+YHPRmykovaDYA2ZV1ZqfqZP6ZBiUHehgLg5GBZrmRBL/6OzXz1ctsw
j13uOG44Ph1A+acs8QVMYUDVGZTEpPIaQUkdIDNQXCcNr34LkNomdWQoxDkEBqFBQKsGowcBNX/g
NkBkZizcX8cK40icOeGxaFDRqD1gwSCVe/qGDNemErVFzrwu433QPR43YqCzVDnOXYh/sYOXRsiU
UzUwJ6SfOZKP8t8voIG1E9U/luWnUKosdLBpULVKmM5hO9EHLVkdVhJCIg64JEeKFvubBWYH9NNp
78OVQcuEQDMBV4NXCIwDbMA740H/fJkN6Z0ecKfoFUyIYG9dodzSva7h2ucCiSdJ0ubyKrWo1eJI
EvbkiUsPSE2Qv/eXsT6/B6TuaY/0WgW8nd/7toJmP2xW3oFYCkMuoB3KBxfZ7JaPUEnfWTHPOk7q
e2qLMWp6z0gtdG+6m58YYusieuN4G9Iw2zTvbIfQHf6f1G5roDEThT1WFltORTTsJR5SQDb6fNWS
hkKthfIJYXsmXCrq2oYTM9aDXfjO+8f1C0Hm3QhLjet/ATVttvAiXI8qDvEuT55OoOB32/8c6FjQ
Z+OLcZLOZA/ORReB8/Zub4X0aVurBeMFMNFj0PyLAQvlf9UgLb3xX9WPZ0N+Hhh5vfp3Mmv9vjAd
aOv+64V2cKgBqi/7qVzMfH34ghfwpi/kAke39wO0DntRAaEIcDILMtOBK0j1k3YCaBpSeMKOWPuU
UblRLeToGIZmPawiEHxfXhXawMGwDsEA/Ti8PPtzEuUa4QX1ue7GC5xfqEPn/ERY3joNjVcuVW1R
+ZyUirNVn3nRNKsvWTW8alTinTZQ0diz9nsOBZZfepr4KXrM3eePHyT9FTzaLOU8fwjA4eDUcnDd
fueOXjEFNL2ZrCn+xc+K5BIMb+EoRpgDaxa8VNUpHibaZOnZUjgyZ5OV68EHLQPeRAG3EgT8cQDm
JGcbloMmTnILmoNtpKi29PBoldQ0g4DYRS8XQHsDiWF0s6E8C+z5DCDScSAOvFuclejkfYvYOnFQ
lTm83hhdRHm7U//YDlmpM5s15gu9T0uHC8Tj+VG/5D1Qdxie9qsBrZMCjcwE2SYFdZ1qO0uUBFuO
0PPrZbnzQKl+3em4+vHH8sOK+m52s6KL+y/3M46uSXJJvrsPdzj0gkrrX/YN90ZRzq0dsLF0I4mo
pxQsXz4XpZrr0cM9jgiBy3sP3poieJGTTFE/Ynr8tMIpLhcdbL5IpVNTP+sQwalrWMEnDT+Dbask
iJfm1RVVxalLq0wFovOZaoCMnvMAUSvDP2CdCx6yk5iznwQvqzzG0ZawlfNqUd0UiA6uo1z7Brhj
/4ouHYapuWc8eaAm2P+OU4eGGhho6qsclXYaq7yumSYZZOAk15J146/jiNyj8nIJ80zrmX1RPbxs
1JaP2vIQjHTZSOyj9PDYfbbYXEdjcfBOspJpR21BFG2HLFJO1DPln4UxEKVSzE+A1KIBLukQ1wL8
h04SRenWhtGXz3ZCkxyoZsr1Zw6fV3du+pXyCS+iiDa6yiiif9MtAiWaMcjYfCEa2BYEY5Rd
`protect end_protected
