`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPzY5ac7rof36eiw7l7r+1HWVeIK/1fzWUcnTHfyYKdIFR/7huevmE7BHkaBLWn0CPsDJvANqpaA
XYUzNauhxQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pl14fIKDmlbQFDvmAOmDwtv/KnPM4ihgExETaozxmJVBnKvnBfZ5kkiCmiTUpMo+e8NUO2tWzzRV
rszGcacUmAQX5LZCTIHebG28KD4369LpXFeR2EGKOkacdUqlLAiuVPVROiWQF93imoi8nA9vJVHZ
F133EfDPApQ3PHquz4g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QBM1cDfnoAz0yxKVSO0jYLV7Q/jjDHZLi8N9f1kjEEuos4wAjo7CG4u/xkfi0JyPN+pMasE49oP+
XwEE4bqFtXpTn8g98qj2Z8oOaHQNm5PPbGaTsqkJQCRl9P2uPoTc0IN4qWQU1PfQH+hRzKkO6KXw
LcDbtA0+ThKqEMr5Lm/8THMMZbKFbrvpBJFQGy72YVgbxojHwblM4eL3LY/1dEvLyb5reWB0COI9
EI9hkeZIbdESuDBrDLt1Pg4CtlbXXIPodh1Ev0Nroo3aANcr3WCLQvIehTTTU6iVBvpQm4TFeg8v
DEBTS212sYZTl7glvSZgj3WoJpP2jDROkQbyGQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K4v8WGTkIn5id9/fEEE3JiW6VjLfxF3CvdYmiBs+95yyBvZwz3WcP/uUGBwX9YzSrPS7VEo7zqis
ZLrxCVp/gjEHeKg88O49UL9B5/1zsrPBnzDgOBdd1zLV5HqfNWCniZtLJqzlp359ROsEnhtNo2V4
1GAhGNbb2qWnpNiMWpk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nQo7UQyeOXWCKffMAM5rRDWnCuhOrUYrqVoKMBh6D/7EYgLAhK/dGXkQ3/T6gljWwQ4c26m6mOPd
ENqr6dQ/Xq9QIi+vBR4rJvW1Pf5I2oPF0QUqBetnWGvswB1pzJxMXj718blSUZUiI2UzOhbnO9Fi
4aUWzpo8mQqZk2RzxzQBchm9xJdh0QlY1XcxARvLpdUbNVypHd70mW/FqVuHSzTxpyeyxB8E9qN7
s3xsiTZ/kVAym/92FxhQ9LAi8kHEEQg13uwCWKUml/Xgm/tP8pjxW3m/LKhqCXFPSnXfofqfTpMc
bssK/0Af27JsqNDgvjH7G9TbQlEhv3xPD2iRhA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37088)
`protect data_block
dGX5+p4KiIcQxZG2dEloUOeOs03K1ZPKvVAVZi/FEIAh/y1WxbWObWXo1y4BtYZAdJ/PRZ8b+Zl+
uz7anEmGRTayTcNBd/3s+F+SNok8anQFSfIIUyk61Dylf7xWIZlSCmYKgx+sZ3lrOU/IJRkUJ4DV
tf5MmGAe7vY6xdxLHoYJBSyEzC06HHYh1LRlReHYKkbwqEuaVt2Jpqov0srlvo2IYclgpZYR01+v
YKI7VJtD4fwBQw9Ou1NIEvGXNoZcrtj6HRdtc930qXSURp/HG0yj9k12VEkRTB1xJsx+lzGtm4nh
HegeFTMv0nq1lUOKWOcQod1VZJTX9AOBdO7VQ1N7yXdrZM0kk8QEQ88drIkDfNJIg1ko1HUqeZc2
hDPnyJgA13qpmRswcl5lJPPbP27q3Dgzx4bK2Lu8ljVctTErXveAY8ZAR+reXc6ULVvfH93cnd1/
fuzNGnPrznXFgKMc3hR9dsL1QKkKKY+TL4DdAyVWLkkzQNmmR0qD2PCvy7+7xdiwmmcy6O60jZ0X
JZI6w2ZLXSZBdGEcPbelpFguSR86eDhJ85GX3eFKz8HzCgxDriramStM+voEMGo5cZKxqTzvVOHL
Tp8F19UfIZtjsAHFAWYCJoHoLEAnCL/EsmvEPRX8i4teI3SgUpbrhmzZVRKhpumq4dzx4wss/jXa
oA7SpYrGdmotfeVDM27fYRLSaSLoZpBKZ5nEUQHU4OxYE6KZTv6w+1xVtBd7JwnRfB8u5adOaB1g
fioBcvpW0VDC+cDnYITgBhP5QnccIC2AIAUDPtNQXrDggcv9bsjMnyAW13bC8WgRYdl6XbuWjR53
3RpwAppvr/nLEEN3muNp3Ff5b/TldlKCXl8oi+HkkSQxoDqaHMb6MkyID3NeXuyBmdeGBygoGp+z
0yhmoM97yepS7Z8NkoLfwn5M8Vq4zhsw9jvtGLWd0RoikkZVVmAunGDwISToVuPM5i+TUUDQEJoT
lgtFRouOL1eZjAzlhjxmiyFPGw3AVVPT4/XeEJosYvK+2uc1gYEDpqdFlFG3kWjma1OUgqM4Dyqk
lNmwOUKXm9CJo9Njqlb9s3607HjN9+5ocXCxdz/hMEZO6SuNu9qkbU0S6YzFE7dfEet+WQ27Jdoe
peJxRSF669zZyCwHgJlB+06Syu+HLiaC/gZHxlBCzldfG3aCoypzl2lGO+EJUN/mT4Z57pMWsJ7Y
ThFw01Ln9/qZTJJ/FRRqBBBVfkPjRKvGr6AVStYVHFoWm1ccrCD9jH2lNhBTXQlOp2u2rjAqyjSr
lsb35xZeTobvs/PaJwfqlaOCDNmvM0L32pt64kyTVgtJAQrxAOQzc0imI0WtaDWQePoTjxa+54hF
gZwwPoSmTol9PCMF2ypsNnY5rZBnYrFy6W0X4hJOz8vrkD7gHN7ycaKyDwLJCPWYTq7nxNO8RYwg
vgP9d6NeLoGHzPip/BtXw1jK3oPvr3NNXhciv4e3zLnJnt7PjxDAqbg1zcvhkN1uVHQPOBt35TLm
X0PxVrDSMZMDgSdDOjYeIwEZLCdGpZ9kH/snMpKiTZhbphkX3ytsb6bR0rI707FdOZlhDxRvZcod
6fQ+ccdQJ0QnngHeVpG3MP++UKO66p/wTk8QLxDLg+pi6icxtsXlCLUxnz/OXrfWdJTDOzyvnEED
Vk8XZJOg8xc6ZOz4TeZ8YyRL3NXk80NJP7j/V+MoBBcWVQBpgCZWCdHZS/bvti/HLKJSqVqLDG5t
pA5XYGMQt2iZ+HBcf1dh0oc992DlN6f15QRojbKje2CmQ5mhHRw6J0DP0GLVLq5ZQQqsnFxcnZHU
G93rKPwYDG6bzk1KzvQh0VyrKrf6/6IZzoUon3Ap/ohE09yMe45UudMzKVM3DN62MScpOWlMSh8o
Q+RG6Zi/mOMmEVUJTJ4tyJEEM+CkWR5uSpRq4+pVcbnrFQk6bbnHmPxEhKY0y57Dtk5Nkztcaltp
K8r9ZJkUIKnUa7rHFk4PiMUg3o4qE5yGo3HKkY7LZeBozK658SvrwtTvNaTdT3v7sFr41CBYhbiH
MWloqm3dxCUA6bDssG7zZyBYZVRsw2hSVyf1+u9tvkAvWmBeoLPlKg82c6lNlERfAfnlImyj1gRM
R8kobgN/3UpOiXV297Hjy6isPgSQSJxx/qfttAa1OfPx46qC7ezP9g63U+edIXofPZwhBCcbvbER
j6cv4EusTstg2UDvv5dzL1NSdYbg6ZjIAv4Zi6I1kOI3xdcOM8HFWyR8ZA5bZ1hJgLYpm28PgY8k
qXVSf2Grv2E1Nt2n3gwaSRzWm3EY6RrqNGAX7S6tfJXM6TZtyvALLVWwWUCynuiEim4rlHc8sgub
x/rr0dM6Z4kdtozOeqbI7v51qBnidxhWYy2lMT5k2bzTAK/Rt6chAzaKHxL6rPWy/CegkBIk9MSo
L/87xk5yr2K+JVI0t4NBIVUsLzeHaClMMH1fmeKGthAwbD0Ucy/xXKUzq2AWq8LNT/PhpFp+6p/Y
NE5rUrwDMRmBS6YVdUmjF5D+nziBHEjerNDfeL4Nko9/XpFsCgFtARelUIzTlSPGBz7Aj1BE6R6Q
Saayh0g5HH8owWc04qUq4zqUgLRCIL2sDQQKlhlABWSH34OI4bk5zAp6ip8IPAkf4Jlxilskzzcy
J6tulZeX/5bdemGwel9tyr5crpQjc+FZ86iZNneQvBPnf94iXuBGhyH6YzyD2w3zgyTJaMbx8wH3
uLq+7IECDI9Sf7jZQFDT20PrVLpoFhZiBBx34bG82RiAJiUfQyftIvOvJR4dkqAN1yyd4OagoSLY
lEIkbYCF2nQg8PwYMy1x9p71ZaJdvYLmlnDNfT2qWno2ibIB2+kr3j4oKmRAjbejILMgzCPUec/B
x4bkovmr64b3+ZwwDEqMLmpli10RHN8s2eiAGqKpVoqJ9aT3qYYHn0aowhHXU2TgEnLC1s7xgT2B
pQjHn39nlYgjjuiI73OCrXpNrw63WaIjseNrif1y9QE2VSAxib7MiPtCUFjVv0OmkDB+J2H5sSFy
BN3gpmzjl9zC0ChVTL8QL/QyQ6cUiELKvagqpxItF3zjUJTnH9f56SCy7GUzfHQIA7fYz5DRPHvi
037ftlYGgtl9qPwM6FK76emeyB5Yv6pzwHhWmWSjtWOPfgR6LgG9FKsOwol+Xz7ERrw8sO2gPdib
Cx+a2ZsDr2DoyrodwkEWUkqfKRzVB3y1h9AvKDiEw3SunS7FfOjRDwVzPERpUMkowEf18z9HD0Wg
s3wqbq175k/TT3iy0QoakOpYioXPBgmbh7YeDxI9pXdIUx0mSxv4c9FaV+JqrviWyfxp2vtPeXFP
MRNYta/RWVpEOtUUAeKUwUE+MDu2fEFILO4tYexKdo6U0MXDYjeR3GynyvWdMn485BbZMBOd4A1K
2Ubo42C+kKLmD0/4f0QEdo0iTU5ZnkIWgB4gsZcf0UtWtEt3oDn85cgcYtVRmjKZXU/jMtZsRuzM
A9pguXYd5MYeYQlnDkZtw3mKPggXthPjcNsoK3DJ4S3BDtPHoTrTH7jkHAIhuc7qyr+6hU/0TMtG
qon9gg1O+/xJ+60mhLbV+EDHBf1jtxrcsrji9q5OTXIfc8n29KgEg0cq9D5cue5BOrhfKgvL1neV
rcWqkvSFs4oBlduuldO5gs6fbnzWWX1HhTPLpHNaP3WbGAlneRa0dfCQvQifWxd7E68tQ2wHIqgL
GyNa61E0fnVB3hFRR+VqrGC8LQ7SAROwgBGFG+n3uXDdEPMWVpBb6lynjYUnrf4TBXAVXNa3OtNK
7KCB6G7Y5hBkeGqnlRhymWrR3wHzlPcPqOq3bduxHsqFNBLcFF0u5GPXLO1PxOPGfsTDqTWr2Li3
vmo4HdmBjMvUaIrW6NZeaHOcAiPU25TWgr6tAEyil0t7O1qXoV1eNIg0QRYhF1Te5swUx5H1u85J
wzVyKLP289qFX4Hw4ns/xX1WtS1wHyUnerJATsmq3cusY0m9wZu6mxpvKR06sh+or4y7kqRFv6c1
S8R6FDvi/niYdKOdJgO4hJsmmmolUm4AQyi/+0ueLo+Zx4NWgXHMRkeyyjt34kSKE7Ijmm1N8JYd
L20JYE9FW9vuIYzZYA897ASS3/ynTNHrLng2TA206RZKAPca0rGkxDHjURqGrEmogLg9Bra78/Ke
75TLhbarDv1KLLYqf6Sa/qpJkUgin+53Edg25e6PKENSC8QDzYmEZlPlA8xcZKT0SsMh2cbZB2ox
BzecfYAquZAvFBVY632lSToq2pZOyCEo5sKXX9MojPVYxs5yXuKPdMKsN/UjC+UoY2nyL8V20G0f
kbvqJHYnXLWvRbNcReMrNO7ltYnTkpsKbe70xHli3zb5ASibQ39BUP7WtM0h8XPOQdXl30H0ukg6
6p7h3zxWe3lldjgtw7yxyTvs+gee3yULWKMBV3Tv3yr8Jscw5Yl6P8/AgvOs2AuxRiWkmg+xhlv3
O3rOTuuoRzNXXvadR7XT68IbgxpvYUe3eL6apSTRvfoxZz3ZzQBVSrTLdYbWThn470p1fHH+B6yc
zVfQGuFf9+QJfQ2DT30N+wugr9Da9ey2hyfcMMKG9i3O6XH9job6jSZoId6DZ46peXWwzDSCJ92k
RcTPpZAf88n26PX7Jn4HKFJOc9qdvdmiszkYdy/XY5944ctheOWGKPA44BvdKcUEITQT7RT9IbcL
X6Cpt5liryJogSR9YLKJ6u7xh2J45RzTBFkKnmaaOxd0xDjOhkIRj7AtrrjJr89XShwFK9B60UoO
CGogDDpHOnp3MDATzxT8MMElT9C91X4pUgTsXeeNPXK5gHX+uxjXYCzRyudYWMtRei9MQN/qLaaV
yWTHh/TLlZBLXB/FEh20de7RSY1gZvB5FaxC/e4PeTIZ1AkpfMHbi38OdSEfC4YwFPnWphsz37PN
l/pR7RKlFoqx1wzvQuleHjExPCLoHOTq3PJS/G2M/LkRZJF3CUn1bRYyoDo20Kh8KD0KiCF5Woda
szsWqtu8szyPO9CVBlzsk575ClSLqFPiRIyg7U1HJrd5hxI+pQ/uvDJ1kjvrBhW0VTiRVTJDNbHn
0q4SqsHq75/+9tW93IGYw9y1pjgr3d2P8ribR2voRHcaAOpmdbwM+D+oRWYRqCu14zv3EeCvZUuy
hpGDE0XigbrY7Ed71Kxta5NUaGc9KXpKgevWNnZAk2b/q1dfhkNhQM1IgNZGUdat7gu4r46mZMKi
tBo7AWfhKzsShcT8sTk6IXH9YBntXGyF7chz8RlA8fykQcLnS5Ipx9EiRKbD4JXOb/TeypauBgm9
fyzGgOszW4O2JIbp7zDroHWBqU9m67DpKA11RlyBf4L4Yz+eat14p+v8yxnjphQkPTZE9ubMgFAt
XX6TgTBiCRfz2vdFc6Vi2T6CQWySzwMF01kXQyXewQR6C2zIyff1Erk/5uQIiiu/ObKJS9oDNsaw
bNHKl9N6BXySy0gMm/rcSx6S9Reqhbbr+6+hTuUCIznW69asExLNy9p1go/O3PQ6+lM0EtSvxlyp
IIGTNlGc4tveG4MqTFhCHnHm14NVZqzenkNdGJhnXka4+mAhIBDQIFsodYIqBcIaXUes14sohTYF
hGTc90JGkOqLWXX9J9/V0cZVopNWD+1yep9TJlxdCrbii4MBzORTVpf2uCYUt2UjdgjSHpgJiiKS
jgNdjUH2kdf+4KdNhmcxH7zXshVDXBncu9TIPNBEECG3e0joYJTp4wNFD8RpqRW114bfPsoBi8zr
wiPrUmR1/YPY2rYL48zQ9GwDxrl4HjMSWE1BdilXfAJuXGKoRg87BUZDQfJhhx9EPrb2dsMFlMl1
jPNfwP+JqEri2cFf6Ak/0TJ3g+rZ+El8GtSrVEZMJqQNlHSaX5ifXVkJVliJanMUmjeVxhJwhUDc
jQoWgZkaUn4fG07WqauDqxC+mQXLw4MIw5L2BktFJ3u8qNlo3TZimqNd8GwAKs9tYw2xFi2MAsgL
YemEQ0RAzrEHJWdPH16oW/+J2CeyIyO9iSHxc+e6QuGECDRfqa/nbVfxUmI3CTmODT0Vmo3Af1p6
xuEw0RYt7PfNyihF5dgb2VNHifHkvzrm+Re/eyldnA1wgEs1zcF+P8MI3SQCahsxb6hC6//8rm2f
yL1/9j/yjSS9e72XFs7EO/BknAXutYCN/2f5/HIDqPhLasALvxH4xIkfPk7tPPIQfc51/ZK4cy3l
3lJN3kOvZpj3uN4LPBQlwkBjEIcln20RHZCM9HPAChmSTZ+Zv66Gfh0FJAFJFS1GcdTlX9hQIGUc
g2VZ+kFummgPpmUJ5vkY4rJmze67AtKu54V15smJ8Iufd7z1sA5ikCy4lfpU2+WKDYiK0QocONUi
jzStAsbJ+iUnVn3UV8NpWKkvL9iKHtBX5/GpZFQ2UQz+r+wsyHBmWooKUe1ZO1Zpl9VB62mNcu+Q
TH/Rla+uuLfO3DfsHAM7P2dR+uj7+DHNa3HEOCnchEVcdc6kAsYLvI/b0tASIGpdcUuMimoUF0iG
GP/fxlykURMxT6mxQkkUdxfcnSOpKINAFXWQfqQ8mVccGpsjQ6+c+XPHTC1TmoZ+ht6KDvMt5nll
jB13mJeebpl8bZoBnxtXJRxZGsK28PnLJIV6odW+aRLv7F63AtSQK68gubsccOS2q5WQwGqzymJI
WqVkzVDNXg1eitgWs75nteVSpgJpOMLDqcV49pGRLn7KNvKGnjIJRITa1IDyhhu178c5dR6Ncd6e
NsKvxffq8ZZVNIoHQGFOVnKHzmDB4OsuENJtm84y8p2FxqkYq0SLO/RJUDubxR8th+w3AjaKWM4+
kzVPO4O96g9KmMuOwOJN2S3+ZzwIvSq/Bk8o/AbAoLi2swFc+cHSjOGHQoYwXcen1wtbxvjz9CL4
Ql93O13iggWpS6pXOuQTUNEZ4Ne3wzqE+Qg3scA5EKCnrdXBL+hL0Ash7sqZdMwV9pv/7HMG1f2o
rlwgynMbLt+5JONgidZuHQ40AFenq5fna7VQYSbzkEbGNKXhlPvtSDbMJun1SvUfha64rX/UHhst
2bilQG7+YfB5w/YntqjZqkOlnd5b3PGuo/pg5S88X1A2S009w9H2KD9KKHyjjn+pcwm7OIzCFc6a
0Dlrj4jIygxyIMT/iBt7tcglfpSh/L6tYuCLfbSq+glULbJ10/I12X4ZazMLuTCFeDFO2lFc4304
1+lYhcrhqcfKrxqm+BbcYzMteARwx6lfUCcjrPsd3WYVuLVS7/ccFD2SJ2Gifcjhj/wkxiu+b0Er
UxUPPhEQGH7DFOiw0DzcgwAf/f4wKRvr2tWSDuKSYIgGBhI+FugCx31uRfZZM2ZLjzHJWa//YcH+
YQQ8lfjpDMU8XyNsin9sr63RhiO/sdPH+MbC1NqRS+p5P3yV4WySufiH7gJFaaJN/IeiKTf2+q3A
XTBZJlzb675D65YVrpOEukhYhPqtYmRnVTWw6Lkcvc1jK2YmFirZmSGOJorlIcVQgD3h1cG8PMW5
4FhxaK5CMDED+CJZCg7QaJj8eAHwteWmxAPuU8+Lpr+GFI66BKjbKAB+98CXRBKHBIOQTV8hHZlD
b1rzIeZBpX5o8ptLdrfcQ7u4SrRJw8nPXcOSMpMy89aGOEWLgVjFcrDtDdX/uGcLWWjtCwjED/DN
7DqYIW/MrWlbksD3h7cGfsBVRvwGnDhANaescQ+58xzfEdyeRFWxrEJUgTsNRzteUFlFma2j49Th
Ka4DLql+589tKuuROeTBvrNBGNVDgTD6gR3KV25kuhvtnX8wb7rRyCC6flI+stecieIELsR+eZhf
SHM6JqlpzUNDX8r0nUkALMBzHKVu0byM5A95mZPxw1idVkphkajgNxDOMghdKr7ThENg+5/zN/bt
Nie4TMlx+5OksMDEmETbPTdpNfU4o0sDrM3dm1Z232E9hG7TRmcymwHUWxZcoKqP1/G++H4w2Xzc
1JQ9Tbes08TThDAmdq2srhP4day+WNcL5wawH/5QefNT1/UpViGQC4GyqKG9VoTrKjffKm4IEoRT
CAOXD8ImxzMYkPC/XEw06oWHAHMMo/6RazTgCckhg5kkIPAabl8kfRptPuv05VQB/DIb25cz4AG3
DtGDtg7L5idRPjdN0uWEGLOvisUKv6WAws2j3Hzfxs/WFnSsqb9zBoOo3ia+lq5sYFAuiE6jg5Oa
l4iRH5LM/doCLuo/Z6OI0qXl3y0TCognijpYV3Y2psjvIpSF4GRPCD/Hp/t+TfSfpH3vfJC99bij
0THMsRDkxlDcw93ckRdNIllggIPCnIFXW/QNHj2kmM23aahgkXvfGal+HvvlR4pe4HfNpuyycvFX
rtdM7cdqFil3X8RR1fneacr7PI2Cv60yJHSBuuUEQjrVRFtj6BBp/N/0Swg3HIb/qSKUPy3+VIHw
Y9Qww0ZHn7h1gHHHWWwWOGGwkg6PBhKM4nPwGcfPQixiBT/fK6nYh47oGp3hqrJqee5Qhuu7RoqW
5qNHAVTX53xTLSQT1vrg63W3AHWvlLerfvQxqxIZ9Br1XNFIDD5K0o4J6GpletVbEDdP6nEfam79
iog+iww7rGVzgMMMgCfJa0wbbaDDNXf82luFqbo/hxz3xuDQEPGI02aiCUo+DQE75CIZz/iBZV2w
g3cvpqW+l10sxdTQMfiTvIdJ/46UpjeiTj1GGvBgrkeyT/5miC3VvfklrbAT8pdsbk9GoVUuhAFV
JzK090ox+GUpdGHgNBkacmtoBR3KVLKTHAfhtno2chdFeF8EGC4ObyDhFZaL3OAuu0XaNcljDfuL
s6Vbn/wJH8b5pjeXpUq1V3HD2uSbQzZ9aB8WUk0HqsDm8LwEEjp+ChAo3lOwIc2u9D1R6edomQvg
jMYlIV4cWbCnRAERffNtNkHSZYuXqnpvKcVaga9rqv4LDvzYZU1Az2eC0F8vhN4xOViD8ezpM8k5
vA76Ko4znlwrdpBkqohqcIR93HP5nh9PX1Q1hBXwZByamaK+dKsIqK2Uwm9wxxsRU28a+GW6Pd90
gJpXSp8gDYQzNAFCfaoGbRVF/+aC8u3Ap6N+0L50HnepEbmF8K0IdyHscbDesSpDvS1/DW8Lw05B
29F4mOHaDP7kTH2blUPLQeD6yVHRJY1T1SEOBTib6oy6Fs68YxYIfTtWxvBptPBoGLVdS102iwO6
NkppeW3CdrGTFfGG67g+4DxQRgwmgKTsn5pIqECsQbYc9zO7W1/1qvBAPu0gpphbet3shixpKXzw
8a/+twGdJV91Lqsi4VtEQFaU0Ds1CeuBoTXO89U/8/vt3n95RvRG19DfqnFpeUB3pTI0yStC6Tzn
tgQhjVdz5maG/YOyYAjNr03B2Vr8hmJgAMdNhsLZvk8QC2FOVs/6WRUO2M69WOHjxzmchaiykw11
ZOY7MnVeJAJooCM5JWfKqxjl34UcEoVmZ9o29mI7aBDVGIxbvvAPIEaaFfeTrva/SYg8haYHU3uI
7oT01E/BzS9gBrfGCuVPjg6jXChqcqr/OVTSxgPEoXh+StaTykl69588p22KJ58BujuDwZgCvu4a
GiugAsa372YcFbYcRSmLExNGxIgtrH/xv4Fo/69XwUnObkIN5gHtF2SqXIzPA7llCnnpnty7aTxa
uzB4VwJfhXEc99PLR5XumZ9dGhFAUBG9La/E8RT4gm4xJ0dp4B6FMb/xcLbIcsuouxqAPO/uk4C5
3V6RGnKZ9luOZTcCdMs79ZBxuJMRynxvKpNvqa3FECFpog5vtLsjV+VeccKfEDRzsMZloKHgE0fw
Z/AZeIUfO/TPwMZT5suIvw3BFOh8TSivWHKWJE9hw5MYj8airiK5tRKFw42E3NtvSW/FujoDkJS/
DRFJRYjMXLh2y/L0JXJt/dz4tQXi4pZ0qMD3GUa5+xQr6Vo206AfZl0rSJfOSvGQSxWArJkllSil
nKuQlq41EdByZGVC1ZxnCnxQOKJyupfichySiQjclOmgcbI/CF4z6kdXLEvitKHQsX0ctYPjMN5b
H5V0lvO/atwzcEwNntb5MOCXZiS8bAqPco8FBMYB6F5IIZqJ0g2blhWx8X+oGkv6e1l3aegnWPVp
RYeMMZ1qkRyNRsvfws8Z3rGreSfpMLOju+ssSYU/hgMbJtrfbBYERXT0YpRI404JK547U5mniWxj
o70ClIi+PZCZZcKV1HO8CQkbbZUit9XfIuUEuCLcwshmS37EJ2D8rJnUfe0HgmOv/y9I2YHewjeh
BiKDHOj3yQzpUN8UKHU9UC5FeGCCpsvHV0/VFCKgoaiR2jMAO9SfEeYvvkx1PHBeUXIIOQJ+v4KV
UsJZZFMUgfIRzUt54cGVIS6RypgIkd+I/EC5C+BQNIvGKGl28yXoRf/rwJBb7JKSwhIk2kJrca5v
UkKNkUNABXJo5iuDyhCXPNFsaH46mIHDTepN+zq0u9aOh9u/4VI+Azv/B/aZpNM/pq27VWCmL7dd
ODhoQ97LyIiZhP460v2k3JRWoLUg+A0b/9ZnpwpwRu3AERnA2XIXQsDLJS//hF8xWbDE22VBfsOX
0pBgAOTXv/iSI220zn9TRI4WMWOBm47knBDSME3rst/GyDKwDaR/Go0Es+jeEMHzCMixAKDgvIJP
dSU/h3eAqbMdrB5ToILEME3WsBjUGknZ8XUb1jPnCKaCsi4B5Z9/94VYNTbZ8FHDJDB5IfPvTiKA
zoz3LtfMUu+r3McOOYlNQIfGdo+MNuaAf5L+ARwSWK0l95u3eXUkp5vjPw4Vu32nxQd4nKuh2oyB
1h8z1K7Lg5irciijjIRzLofg4rYH1JodZwGmEA99AZyQmepeC5yW2UH38gZVY4o2V/NtJ7C+1/h9
kJTqW9pU7P9Mx1iGmPtuZUFwiJ2yQpS7NDbNi6v9YINGwMAmR6qAvddZzX0zIBNjzWYUjL2OZl8Z
eabsON5kSTfCRboxvqRLu2WrHZrEQus+YfoTsJCu/h9ljCUexs9FvAMhckEKeiM8oflnCsyufasm
TM+U3nSF6Xj4gjLq0r03VLD29NZGomz2ikh5Prn3jbHdjBdU+793GGcV0keYvNlTLjs2UUhEnOMK
ewg3WE1ysQ2eMycS40q9hm1Oqt1J0m/0uUPRB774+nEC4ijFmeG2Dejnudv3eIrAmabnWURodZOt
r/ry7yvsQ80lBmEnC9a2clYPpqbtLKJoIBnOT4AgCOCSmoGXAGBRGZm/ruYUlXa+87KAsgYyRnIL
vrpAeBzj88rCh6DYEXuz2HrJCeV1KMpfpf/20ApZwrptYd6e50Y3zkD7wK1cx2GUs/K2t2mf9dfH
AqRttmRkGQtpckgpc3G+AO8LqFDRNxnYDy1fkusDxNINREr+Q6a3mmT2wHmRtk1w8ilWpMWlnfkS
3I1X7k3ZH0ctHPDV4CC7f8sbAkmCdArBYl03aQuDrjWlBIBURF3U1wOes2sQtfg69zp8x502qu+J
jKwD1uKaASO2sfYjL0tVKZY7mInSGdyN2ep4Zloc2aW3/htFolyPCy+hXSiuumTVT3P/h+SGLb3R
5U3fAiltZ/ayUCPjv87UguhUlAmWquiIGonC3ldxmwaDknQzHznqSADpmUKvzGA6JAP5DeO5LTPS
TkV7M8+DBPosKEPwAjjkqkIDSmzBk6g2JyXKZ9DuNX07p38R4RYjhwPTQ0VEFcz9rHHZdfUQF0Wa
GTQ035bKWGIr3aB6ST7AHI2dNRm9ynDpIu6RbzlXc68TdIelHBIKjviNL+Xvx1qHh7x06jfJTpOb
mmGynpn+Qh0Ux0vtBkuWjOgbyGwrIAMGZie0vZ61MS4eAuCSKFzO+QM6wMhz3ePOi73QTVqViJ25
D5QAuleLJ56P/9w4kACxmsW00c3j5N9wHP4f1+c0Z6xaANj1+i/MqYL/Koz/ZWDmTeDO+acvWstz
V4KYXjQPbSk62jH0bOwaA8e++sV/lr1uRDdqgEdhYtUPU7VcCpL13q6NX6x3nTTvlyOVCnjqrmVx
qy0ZORw9uPbhEZY2p9f1kYYAR1NT/Lm461MM/yq8VNfv4gmNqBl54Q2Bq7+UYSk/Dgxp2XHoKrfY
M8EJ9N85DAEuhOJho3O2Nu6E5U3DDCxu1wd8QzCXp+tJx9pZm4xT0gRQwgaRD9p++2EtAuIq8Pcz
uO0zWGw1Q5IjLte6gUmkUTySZJ0Wfz5/7YaNmdR94uJi95fPD+TL2q8oNqxwKVvfIfl1toTJhez8
5s1wGjP22nIZMLrAUx4qlBkzE51vAd51lqHM6NlIgxer0MIHMopr7BotYMOihUdJpHmQVuqhru9v
3TjV8yRmhVv0H1LQ8lUGSnoujJMPj/LxYFF6UKeW7nCzpWH2zW8upJUwg12jsNymCShgimbXM2LN
VbMI6HiMNNcuFTQ8nn07Q+xZjOwdZgBbOoQm2EkpXa36R72ZIkvtvNxmmwUcpvmpPC6KYZyu/p+V
T/9V3G1LXjgRA9ALr1ynT7AVaoVRwdFWTKDas9p8m8q1t55iaTof4TY+Al6OiDVQF7hB9TbcEw2h
bRQo+E64NRgp3r4w6yXM45BkDS/k+O1Yr4sb8ycC1ZPtk9ajrmN/uh/9oJAiI0kg/tpKD8ubp5rW
tzKV+lTQ5puCc78Vp+nCUgfwo9NLovzWTWCVk01gF7hXbeHGX7ABlctrGP7zXO/e4loFhnqdBZo0
zNJXEh/bI/t3kOm/H21N9+KWp0TayNUgBk8/hznb0zsn8k/GLMgzjFSyosV2q3TDNQ4pC7Q6MlF9
9Dg8e+tLjBZhjIVpShi+ypCPtQnoaWvHg0j8HL0Sip3gl/+G8rSmDhZ/7Qw6BzgXepAqOvO+PuRz
/+nqYdldThiitriZ+eA6N02UkAeyTv3TTaGdrn4IY0vgVHebC+dkzo8p/BrtJBygAnpIMIkkSD/x
cuMh4bzj5aS93QcmxlpIu2nI4z0ktt5fEFQLtG9rwPeu9bRjBA2LgLiZ5QpE8wdJecPkOvyp+Thm
Op+rKdwC6PpTEleonGSa4a18ZOK1hg+fyjfsKf0NVRhWrRmsP220TESsWnKrTIUJsFIvLTcJ10RI
qlvwRcyD+Wd1yVgAvONDctJfkXA4dcyDRn2GjxJahzZaQwMCIyUgsrf+AsZL2H9KKr+GpjL/4eeh
+A8YzbXKWhQiH0GkcHdTDXh+uCfhsendO40LyY+eov/F7uvKwCGENspBV95/S0Uf/4GYCp8DeEX2
NDtspr//jlrMFQU6uVS/S2IxtEXOrlW9ZhUsQ332mUqBrQuFv5P8m35ZKRtCVHGGmxXivggcLwRl
7H1N+ur/yVIXY2KlIApiylhJ/WdjasvGV45YWrSyXqtDrZ+PZQTN05wulykBIIS+hZcpkcHXNbv4
jxnRqeIuqgwHcZzE9ArHTuJgC0PYRxW7IIzL43IhI6Ztr8+nGA7pIYvBf6h0oJ1SHFbdZgRAXbfO
iGY9RYaou2Auj2aBQ6b88bq/ZAyFs1drxi1jWNyUaGIqM2H2rjnzXg/yGdIidh/yudBPYc/v5YLN
kfxMIVSAAMPb6bcMn8yMuNniFPnsypewvuj3pPU8U/e67g6ZHKbvBlyUXkAsUdlDSoISxXo8vwYl
PKwxM4s4RTbH0b8ShUAlVn+Idp8KFKgyLWohUiSm3BdVnvx/pqAped1NR4h8IMQnyfcSwLCvQXmm
g9uwheDv3HPHteUNq36CWOrRq2jeI6PyZhAe7QyWwKmDncWBw8bw7DAHYD3XxCFncxyET8ZPImlr
FNMNTkjMoAeDPDbOpCtbIkRfvED3gQd0y4NmBi0YEQc3YW13saHIJMWynko0FI/EA/JfJz+h42T+
jXfhRQgZzWA9nEy0/302dOoM0dL3TCm5PRu5DAvd52sa8OMmJ2j70MUpuO8bc+TaGSIWdOmRAQML
RpMhqkxrQCAXmlE2osVDM+/YmIrJA55J2l+pIkwdVOHseHEngHR9St9QjQA/y5cg4A9OYu31KE20
kx2CU9jsb6TeAEADTvot9F3nNibyX92rQvqxdMyp/lWdmDjnvnsTRoAcbLZRMY5vmqKGkKCxTNCc
dpJ2SgqDHzK1j7bG9+4nEwduV3YQSm9sl+2xx03Lr597rD6YORl4ikwbM3x64hGLxXegHPaZfLjh
Sq9WC6iJ+2fkLEzbd6WsIRAahSvaxNOsWkLry303zQPaOKCS63UtkpVDAIS1Cvm83PvZnOnjJvNi
H4gLxfF+m0my+JCwWThE33z05ZgAblfBkIZi9ZnYX2Mnj8beqwX9XMw3+sBDp6/9EDNnipjv47Gi
ML2yxjo5ZCg16iMkuzFmbXAuaG2HWtbZnhy83XfEUlwPfThHVFaIgfUjMPVKWh3No7eeDHyOl+ls
lskGabZSRlQhpZYDMGfiYl78CbW8ynlOHv6zIgIm865KcqMryXTIVrs6CoXccJoQHmhrqZsuE155
mqfOaOX1UyY5EAE0f/PDqKiGb+zFuMEZpzqQnw11R8MCktz2jNgqLGoKRRysO6KK+69x+AdrbN9y
mUnPas8AbPgkluZ8plrdWVyAfhWwFYfjff1zg1P7VA9qLKab1viz3on4t8Ivs+wcEVNxocN/36xY
2/EsrGyM9i6LabmU7uy5pIT6z2CwnNkbudWp37xjE67lqMZPOHPpLOI5t4Wxjnzy/8zPkkXjZvqm
QkQFkSSgYrtO+ER9Sg7QoRA2lSi1XIhZXusMXMW8POreN5wMX0qKR3hILfWvnXndBKwgzi+g6Wyc
a8Z4B9tvMQ4pMzK4qC5aiD9i+NkUBE+aUXPseqo5IQ01ktHXoBmq/hHDa/7/edjNgidMj2QyTcn2
jtxzMqG9TCtKiEbzMQ5mEwDVzoFnjfTW8XDuvtRU2I0vpX2ogxypGvhg4XKxaCl3cwM2VBaXIcfK
CHCga2IigzZdXGM0YsX7wHkR9cfPcYfsvZnJ9veCTW5taCPLXqPEQZdn+4qCqzU7A0cNR3EwUak/
y+YTNvHMa9cLBMRe/grSuAEBuTgBUZHTI9QU/odPKjHbhf4peeFMmFQfldXGAHWHd3rJVMgWaYkZ
JDMoTxjVX2cxVLzMTaDjriyAiVty4/EBWjrQzb9sI1QAw51JP5yHIRo6I4S6fb5i8bH9WFuOektK
NGRQNn2fGRpaDKR1FpDOq5NBLOS4x6uhWEdQOjsFyJ6NCuRBrrfgQ9hlBSAkVZPbUCojOdUOL6/N
eanx32gZIu82fMIwp2A53a+gZx3QnWl0MihMDUVFFMAFVOHDBl92orBxUrlNlvZVaBzXq7u5hTgh
Gp3kg+w8iMrz2t/Iw67u7tAmSMh0fiOW34XLkUtVzNW9MrXKqTZHQdrphaWEaaXu7py3e+ToU/KH
G64dMyIaYISt9/5KqDsJYXvZETHXL2DDbAJwy1RzPO65T7BFraorcKXWMcZwoTKYC4s+VWVYXZEh
RAjh9BUeiZ9ZMQ54N9kaMDvhjD76ZcFPtYm0POGdbIOgqQa4OKHZJ3OXYo7jJoB61GJSFtQ8m+ec
IvW+QRa7LfE85cR+WoCccu913RmYaUkKu9WcdzN8GikiqIe1jYYGmWyMFlzayMcvet6k7Rxwjh2A
hgM0X8l3nCF84Qxh1dKdsvOMJpOQG+g3kUxyBa1u1VnwaVrGosDXQ2/1lt/cFGKya/bJ/nHxWg9Y
7VbGthBBXY18j5jMUPtmZfmtBiguQ8yAbSBNPAe3aUAdVZuuJ6/JojcYMmkLtTfpwVtbzqnpCPCF
3Y+14uTMRGXVKh3rPgLemPKGl6Hlv9C6trVEMuIqlbYLuCBFZsNu63D11huVwSz9uPtK2D83ljnj
rzUAnl9Okt2ZETs+2SiJ3y6wlHDSDWWK92HHeuT3XpXdQJ/jFbVIPGzaa6t4i6TFgquCIXAOHyEg
Dm0RUV/mUtvBFKxmsuqoVEUFCfIwvjAjupr32d4f145wHJPFSIIB4QDBz8kAqCbScjVJh98mN+cW
KUjousCE7r5R7/vOOMlBNzJbOIfOgQWUmnJ3b0bqo+aAFNjSX/wztChqzL3QNUVL4/07CopmGX7+
QsJb9pgJ7CSKevIcRi8CeRmvfDuuVlKir03qnWGrZZUtspN7++iRDU8xAEgqMEAcy0eW6Qh6bZAp
XWygI4+nS7oTv+ztb3b0BQHyclddcSlB8AQtyWoRbSSZxsdNCTPR1PFGy4B5Ju50gRjEVDhBz0mG
J7tdoid+dI4drgYS301jusUvK5FYCqhzmia+pDOmVdes0Pr5vMfjxdYVmMxvHxDl0CirDSA+BUvW
G7BZkCmuWAEkYPhriz7u21zk3JLpmaXECr/tOvFVNHzESM3nyZneTHdbTVLWtin5muEyMv8OXECl
Z01MlWA15erYmsgAEDMZLbw5XIBOCHlsWEEZUfmmFnncxuYbRzegCb1T8xIZ+/8zPwcNIjATC3zY
M+3SoRYmCYsoVmjYf+kRTEnxDU3MlGwCnabh3IQFnxmjuYp0wgussZL+5si7lMpzWLbcrlcPRCGL
AKGNVtG0dTt6U+E6MyPTAYHWSrRH4+NqRD05pWdWtWWxXJ/8UYSFasopQxVHX4IuFPGgNhStOh6r
0xbNmMzZsvDeO8edA0jzdchCJPnYiBKzwzTlvFazGzt4OYj8SGDLKA1RM2MhVatxSmvb5Kes5Dm0
p37iAZTy7UEik5qqosiUU+oNwMBfYq4R228lXXWtjc3Rgx3qN3PPVxJdDCCvy5U6FyPKJfEWqHMA
Vo5JhRPh0L/FhjokcDFEpuoEUZZyLGWSimdbE+vASKyKoSulBGnT0KX1CNJPy3iKtBCDn+de+Y40
TP+iPN6gyqO0d1POkNx6W1UTW/PlJ6IInSSAh7B/ad0UEC+1Cd6UUNUK/UHBhMQRHzfuH0d3JXh4
lzTHSfg/ODbtJRVPaIzUcAL2EvMjKAxzqrHUH00o78QTkjYezDd1Bu9vNoEDPO90q4Xf95oVysFZ
x5UDnxGZ5A1SOU/B8VJ6no/o9XwUBgI91ZAxm3AJfXBTNuQaaETVL2Xgy9Ew5hTZV85GvYopZMwX
KGDjVi0AJXPlPUNQ8cCRsJtWGJTOSDhi6kfUCGSq+g1/gwQgq8XGozNaJxMefWvrr89/HfDK9HdR
AwUeR0qjLKTF5lZjG4cCU1CuNHCloNHD4Wo1snSzX0zLr+ntdvbvzUvhFBr14TpQdcknAqOV2ECp
qFCNNVp22WRVfVrjMHyfpJ4tUY6gWLmWSBZKAj6y8z5w5PDUjIBSyQaZofHokdF8wlDkkYHF7EcB
Gj6MG2lYNQt1Nw17DHPqUTV85CsLbebNPRNCAeErBWRd8keij5jevQmuwAxOm/LQRPg8Q2UXDOmX
3OHu+RB5r3osTFyGi59iVzhVrWhJPOUIGmYv3eygFK/NxQ3VUkSWVbcOn2DtAAhUH0ndXNHtsoqF
o9hxCIN7OYKUsPmRh0sAF3orNtkt7pylExS7sKFB79uTQfv4EVYux4Mmc7FiduqI+BIc3IEmZjIP
2Z5uDuBga8sH+Rsmh+QDlA87lsBwzbrBD/cYAzVwlj4cRbHT9pjjb132w7xzVTo5HI7iiIoPEU8K
f3oTM2H17Um/OI590jw5Z6ivewQq9Xew8DStC1TrcNXy46msIiKs9D2S/fQCJD5IciAGvoBIoxEr
XNTfHrZ1xCvy0V6302jpzte4WpPkD8SumfAL8YZwArPUwnIg/aWtwv0tYIRdK3JudS3vVsBXm7cA
PAnvzvtP2wIi70MnbOTm1DxnSaBfAfq3+NuTvlIcWd8RoKFrYT+7WjLeR7vwJ6w6QQUJMRX9B6e2
iiGZ0rCuOUHVvhVm4Vlai2uRNpCnMcKpRlNA8JjGGAZDqwXewlNvbgSTiegqpfLVKL+3g2c1Y1na
zIojnTc9fkAz9uviDe5/iBIxf3Ngm43T8bPgrA/R8FoU7wE1zvC2dmc8zChmyMDcuJ/IavLYJakO
NeVeiaYY8BE0D8Uup5LG6lNyRxNd4MW97HLBpxqU9WVz7tYguFAdENatvpM5WYk1VOLj90eiyuMM
rr3z5o05Qf3217hKx76mVnzHxtKWXp08I64fBNedJDmN5orjyNbEym+UiluInpGz3N7UKEl2f+Kh
rnEagLrISJRyGbrIOzYjwC/z8aoRW4p3n4af/Zl17jC4aVDBjX4Eln2Fm7XkVNv++HBnsuoiQCCX
kijwVf637MyuheOn4PxH6oTn/VM51KYvgbCiiwYVk+C6WHXWAJHrKyYPc3lprbeB39OPO6MPZ7Be
DmD83YYu7XMxDQYtJadogP+qRMJxg0ri0LjQE++0q10nb7pNECYZ3/7cIcCDGJtxvitjKOvk12zo
ecCSLkXVWP9jnlnCMfeBdxthwTj4thThMEMqYn0jAxXmpWY9MjCJPa/kPk1Z2ziYL4/+pufNvzzY
To2N9yewgBz1D78f3weQwIi8xuuzhvLawtTDXyJNUO07CtwJ7EUGUofrSx7qLQ3+R0KEYK46FAY4
WyQW058iXyWEOS6P++Yaeku41F/vGiNI3Zy6RtkutCqta0mXlo6GcHOFHRwn5jMAHfMFpA06Oumz
m5ftpGWsBiLwXe/eq6vGwI95f4mrNrb+FjNZnnDtmph51ogMg5GKG+HiKtqzDKJ7tXyGCV+maOcm
m5wD+o12219+jwgOUhybcQt9JpBRwxqM6jsjuRTgtqdM9Nf2PMx9v1iZfD0i5TcSfd4b6pQJthoO
kEPRDLgEbCp0qDhcU9m76G/VChsXUXfSH32IXdItRKjGf9GHNhOZfKBbUwNENwnw7b4q368od+gB
uD8zGibVF8bxLHPxUR2MbX7gEmadOQbPdl0zsNa9rWGUptPCkkj56B2XrsPwZNOympqhDeuUVD21
sbWRJn+pNXwMCXDz9612+Vyhj5NSbnPDoYiRXlBcIBRKMWy7WbRdxwifNqUTGV7hsN10/pZFh5ac
MQt6KTCFyORHO7dhWxk78Hibhe6r9dYazIjX6iz/3HXdBy0lrPeE8aSJJTZ5C2XLO6tiyd3dm7Bn
QIXjii0AufIkPA6uGYIjLoIBLGNMCSO6e+2aqCe8w+UATkH7shyMt3QfM3ksx1oVfQK48Xb4kAwQ
pCQEfO/FNYOqFSDWzRW+gglrt5FVST8M1ZErB51wUWg6k6dRu9UKHHAnZGZzx5U5pgqTIBfKD8Gx
O5FfBbSxZkzQVf8AQ8Jb8Q0xexAO+mMxzn9KnJ+/9JMnqggTbp/ANMMfJh5JudavkvGocrtLTx2r
qcVRiA5hHsyqU1EuvGCq6F9BdgTCxMu3E8nCAMVdHBGxZjQtEI/18Z6cpngyORRE60D63Rbgufbn
E3nZi73652mAt7ul3vCsjmLL/lpdclQY15IVpUkDu1G96ZdgFKS/jGlKKwkGUmtk6yhOvZu2rAIv
2yXQNIU36DRNDhIXtemEtZkU8qPUt0B/t38l0VbOtfCV90QI7aAHgcBKllMaJMlXn4IKMX8WEm+p
Yj8c059l3z9MuzFHkCLJLDBHx5CC8hLOzbnmg+zEhfUwvlBjB/eABNdEdGAnQXhyDhvXIMep0T89
ujvXFmpjOufeILm7ZkEmAKcEf8gdgvE33f+Kd3vYNqittxA2ELEi3DMZrp5HSWtxo1pmk7Qerwsb
bVdfJTIXgTpj1RAHlq5UcK9Xo/N1VRzjOzqw2yu0i8CaAZJJJg9fF1v7lV6zramI/liI311gHGns
bwGNft/YJExRKi1F3nFRkhA9AtK0mBBgpLIBNNM626lbjMSPY62iQoUUx2ZLI9Sp9Ri/1fE/hJn4
2OudSwRdh1qEGKwYPYm3phbBxz0Pw20HWezDGMIYXX0Wa57y/zLwf3Fxmfpy37QQInMeryBO8Sda
zZ4H7IE4zviSVKS+dtVJRLVwVkQa59JxW6PdVXQGMtWGw7O5G+nsZBJdNBHvrvujMG99Q/40azUB
E/6FyhF3M/CvFmpjl1YgjIE9UHCkOuZySfDhzp1Zn/UncS0cg5Uoy+8n9wbszn71ZwS6/H0Mb+cT
ZYdKt7LlFLSBbTN7vkfINf5OBbzPmEOjfmRoz+xUZqhjd+w+YFMFYkloE81GBIaKNhJl/JwDBJ2y
0e0rtvYnHNixgamqzPYIIi8Bpd5/rLEoAU8eJNwgG4PQDi2udJKLtwAYEO/SAC1cWqYEE4fmmp+o
SX5pm7mqgXqDnP60Ifp9W8ZD3AyxBwalVxR+n4rw/XrPkB7Oyj7SKB601jnXZjTGL0u641rFauQJ
qDz6AK7LujhyV2I1xmL5XnynXUz/ZAkuyQBWTGr7i4209eWKVLy1rYuX+QvfpBAxX8roaTIJ68kb
I1FaTtBuRNsA188gd/OG3pSi6DGcR1gip4nKc+wd6Ira/RtjZXwZ7oZ4LQU0GFsVDmChKCdWnPoy
vUmbaSYxlWhF1ppdKjY2aoe5P1oSmVfkzzdbBFW4D7FTEY12kXNkrglrWX72tg6vkq4zRWetGJPc
XGiaX+HVPPVIe5teajd67YkfPshSE5BXgtEiFd34hZTeVLDtpBCY9fneyaTvU/Q5B9YQHZ3k2Bj6
nXpNN/pX4SvDuVnyr15eGAYQmNUK4A4TC0wJ+OIYrHkijgmiRzolcvIg2MxN3oj546BgvYlMHJFL
XqZ2LzQ0gIKfwtXWgB73TnPMP7OkuQP97yakLFHEDW6WoWtFJy2zOikEsdN4jJbo5xZnHf8nIbuu
Q1erbywTCoGOuIT+LGo0eDl9es6+uqRLL7nnuzrF/c0TeBLGwk2VQU9DyVdPynSNVVLTMBwbxi9Q
K0Sab0mC1nXhufLfahg0yYe4bOm7aUZHoBSp0K1T970BtUNo8V43QQuPQ0sWm0E1IMlFyrN0yP60
TtUuuXxslcIz03/+Z0Wvfs6P4VR02AsovE3rqzNW6xV0DZyLpeLbBEaQQ1EdFzAQk93m4MJ6ga7V
SO2YAn+iXW1HTz+d3FVUeTv+jKA9Qge8vyQu6ZT9o/tuqB1MJI5oLQUsuzTpcMNHN0JUTEHxiRc6
E7DiyO0+UYZN5EhZ1B6hHYTuMF8c0Yq8+CXvVT/j1vP/GgehoSXnXcIfh3H8pO4J3c4X2P0K7qMq
Y4QnVI57lL4SHv7KWbCjyQ7GgYk75eHn1m9RJrDiJe1c79Q1wFIJNx3aTyT62kYs9RgH7yZulg3U
565crkh1eg0A4ploArg4ZRHflv3KKeQgBLIrEI5wnCjMWx9AbV6ZPkYc5SPhQfHZrx3Zxa7lekvp
aObbbDArZ8f2/h6muRSeTrCaRXdTJuREaIpO5Xibd/fFfOyegDvQ34r/rXfjhROMERT6zwpJW7/j
hD+Cd+Zvu5BQ8l/scFL2QX637NxFRU20usMePWSQo/XK74pQx/pyTfzmOzb26MlvVAx9OZlUmNLL
d02IyHE98Sd4b6bKPks/r8aAdNZYRH8yRSQT6I9/1j8hUvWSbb1VEP8Dq765isX80DI3Rau6X5PK
W4H43uoP/Ua3wWXV3xCebnh6cUj7esIrIS3x78Y7iiUvcakPz+8egN1esZavTtJzPehw1KbBxUSZ
IfHecxVxCDfqtPoWGh2ykzEHkL08gK3wxCxWjS1CA2njjaY8728Ri/CGH7elJeWenyB6O63e0+jJ
C87SZxdkqbBYEbK0Xae8ItNCvtDKvd+A+rdDtB56RgsqkwRdf8GTQSjjbwAtXxnYgzL/QWqObYRZ
P/BGto6SnufnfNj3KsmlYeelVjJBqDp3od0TWpwUvZ4HjRlzIPfLXCKSDEZU8nEoD3bhVK14qX5Z
e4oI9eZrPmZCdTV6SL2TLiA0qrVH5ogdTdqOh3tDkPRUqyI7Loa+MZkP1PkjC/J11ozloQz5ysG8
51zO4ctwcIoT9idIInk+3edEHoPVDIlXmnZVM1GvM2DFYXyX3q3YqaeqAv8wn+m/nKM9xTvTnv7a
hdxJM24ZiavTbdT0RZhAe5tNE8S39BjcGZp+6B9aRgRNCQzLpCVYc2NeCL+DtKb3wjeaQe2bqmDp
lK0SYAmciuYrJGpPtugtkzx1JhXUUMToP3DIr3NAReSY5pEEeguppM0cqSSC1uZcETe0kN8vpDTN
GBfQzSAytONBIqAtzprkKtM80fx9nL0oBvsiUOW/DV9+xZCbSrbcANcyjPbXEU574O4IkgWfbI0/
is2+pUxBmQBDGih3o6MWO+mVeMv4R2bZUpmAq3zD7R3l4+cylZ4T1rUqdK0aY6UmLhrTPBV1LVmg
uBPzLEjuzYcAnGKW246N+HYE3AHf4LBptfS7dfWjNOP0NeIb90bDIi1isBi1T6UiOuVh2P98hYhV
F4Bm7Y+1Hr4zAR2LXfA0n2PL5BlYZaisbNnLSkX8/Nxq89BlGd+syhxPCb8d9WGv7bzHJyku1/hz
eEQY9cX6PJqNuVGXhS5fQLqZpBLfV5l8POTBdTQSBhRKD/gNeYsHSB/quJoeZ0mZYbMgthkkXJPU
4xRdp9RcjRudy9ybWkuHMvut0nNABfBUrl9tSHVbvN+iThBe0bdPcEW8txuALaAxKl5m5R6dgvKp
hljJLo7GIWEdjkJ1KA6zAjqBLO4S/PsSI728oz1L6pbfBV2VGToXgTj6G2/R9Zvc7TT8z4vMek6M
UzvuYR5buIec2caLCE7l6hWYPpRVb25kNmMN/elo7aT0cjO2ylTSr1HOoPkfc55FrCI36iUAsOzL
dxh3WZEZdvk8ulfh7RkwLWHdvyFZuUYl3hpovcBfoUIwUzf88fCBwGMpViREtjKIHPpmR0SFdH/s
N0pLLxfSWoBnLpUBpqsZCjDNp+PaEaCJWujnCCg3i6v3I+YfirvSA+dXbpAzwgVAQFtB4zOI8NIR
/qCXswA+YFlwxj06kGbJtou8SkntvT/u6NyJCsgPStpqjdYr0CKYjEpeYkLzLHuj1Q3FRmLtTiMg
MXK6d8Nrj2Y/10KuWpYwRRByTm6ion0MQ2aEYnRWFLc9ylQYMp+vsTGCV5AkkqeXjNJ8NDZmf8HE
vTtyjqh0G98XB+IpY9u/n4JheszySu9lHqM5jvn+cCYaM7+uS4h4aIaBY3uSfphLBgtglU/7DWzx
l9SU3QgOpLD7TO2uLa8LDmrsXse4D59MgKChu+dT+CuceCOmb/NpCjS7P81yU0trRdSPG3tzvbpT
Pr/EN+OfWNrxP+HsvdAPOTeU+d+D+G2j+Tfbh0KRGENlPXi1osmHF38Hw/xbwFeh0WZrMO+b21LA
Wg1UrM1kVCwlmKE58nVlYzVNeK0ytm129n5FC/ieDRig/r+sNcNuyorWoEaV7EKAuZ0fFOQFqeKz
fTC2ff2HZZ4Jo+Amrwl7SVFw8FKb/d/JxCWc3liN2cDRlO0UuGBk68ukecHCc7MlFdMprsVIrOwn
TUjZWgy37adi242WOiDrLC5tC6qYmTtGWyx6PJrXhlBRon9Hw/VFktSE2y3/23CU5D8Rty+jxiDW
XKDOLGy/IzHapu4gra6sfCpC1NuQK6Rorzaw6SFrq1Wstjl2kZp9wjOtMRGdH2yvREfIfmimTqPO
W2AWXEm2LBRbG5mq2EVQ+JkwlXQG4rKhVZ1dqT6AKx2cE+j5W3rwdGnRWcoWP/p9jjkX+8gfPKqo
h2a30JFYXGlc8Ac5kQGGaeHnUKMR1yUTpm5wTuy+c8hUSNxe0/GBYoOBQufJ3oFrqc0mcW2M0oK3
ING03UayX7k5uGtNOFMxLFNuv+nH0HI/0EVMdsXZaxBON0ImNn4Mq2dJU0v28t4nZydi1TnRXa9D
V5OKNMeAwirV6+EJvHb56GFgQ1ojrw99Cr0h7rQLTsDU+u4tZepkUUPI1ZFQZKUWhSaqrZKeg/ql
uEpqyUUPxO+g011xSiH8HdagGy8iU7sBQ7ixNLa7RL5IBxzshCi7EDK6MkYDNNm+n6uCqbwFmXjW
5QthGyNyKf1+1m1adJWXhGKT34IDiG3NppwcvqHjKXYboDRAVYYweo4DFiTRzZUuCLbVdFAi4Mzq
nS76IS3lgCdNhgmtdFvZJMa5QoIkNuEOPMEk33SCSn0P8w4Zaztfk+UStKfjSzJqK4p9CaQonYmh
3gmZZjz3H3ANjhFxuS7Msdtl544Y6KG0O+Ai3H6AioqxbwDq9qWCnyxCN+TmnmopCRGn7wPWXfZl
0j8MnviRC3ssUC/pCDpRFmPvfQEstd33d7Hm6fN6/hB0+hbPv/lOlPo/jY9f5KY47m/7CAY0Y3Ef
U+gRPEqXD6+RCon9LBCWtIPAIjJeGuegtnvh3JH1oGs90qOAFuwDA9H6UEUM3J7FQgcRsbkvujNR
C2QydSxTHibKdOM8NSoFnVvk29a95BPJDsCdzGw50Rk4G0aeEx9AiT7LZQoolkNdWAv1L9xiKsqb
8J8FH6LKZoQJ1xGSM+lOynkCeJSSeEGOxuAttgp5bYrMPW74wvEu/FAgZMUbh6G/Uv69sg7XEU85
um0eeiGk58Z7z3//fytbUc1/E/RHtOFbpds6AYrnZoAhTw8eRI2QeaVoH47aIKixRzWYyrzfWNvS
A71M2yBwhnx1bLXlRD9t7bn4XOAg8nwEnpn9vpnjFYOYkU7y6pmyTY76RCvf/c5m5dGsm70sJbsC
UPXsrA+ak1GnGudBMmmhsvTm40B5MU9ToBnkjDcK95XqA77bAe/v4PqiOA0mwrdLnVfrCV6+3fdS
tF07roTat6CA6zNLkMK2FPlmS84gQRDejYKXMjZylXefXuxb8m9MRezwOfhEIS2eKgOXG0j4qWQr
mswkDeQHtkjcvUUa8dzFDUSh44MDDuH/XkwvDT860257mxQ1RI//bQCqtPAT5wVNlS3ZepF2CYiH
MEDjMh5ZNBHyx44dF2SPeLyGDW0VPFUmqatU6FBcbwT2Ud/Aq8Na3MZzDUWBoWfxTpWzC9Gs38PK
AQN0yIwcIwOLv625ZSddV+5rs0AvIBtBfX0lyO3O+2Tz5U507Ovxw1ETLDFMF348hlab2UGSocq/
bnZoQCluuNT6WyrKLswc3+orCU0ncuMGpYsjVlzRzXvzgTErkIWdFiBGgQYInsnOkBnurksecYfe
FH3hddE1EXd35P5gtzFONQDtb5QrLSyHjinxA6Wp2+30Itnm4XdT7TTyog8Foh3lMXePpQYL/dMa
JMCAI4gnZs5Wu7stUwRc8OJrxiXQ0MBynS4o5cWzHq4gvErm5C5FeQm7xPW4Ds4YR1SDzSi37hyp
aykRgeAZn+pVjjechvETXfuXwDORZLyGVpcuvlSuuKtJgdENFtlYIWxP0NF24utPwpUJG72gaJoI
8PQ3TdKbjE9T56uI95y2rwdb3RjQE1tYXDrajrZuxIWsjvsImUTGPeerXatRW47qqAzbv3PznWAK
79tWxjjnFFDkgJskSwQ0sdJHBhJCdpvWveFITVit4Wm5BzPbjCdvZ5phgmXqmqWzSJJNGWg60IDE
Ri1xODj8YT0D6tviLxSCuxRg5ZvNyYEP6n4YaXz/P9z1dyRBUZM2VuAxDmOzDYzBDclu+jLpp7x/
PaKFC3NryzokPRcCA6Q74yIOBtNbK28JBsio93pUXeSESGAKPWsz7F9YtHtxw3P7B1mKYo1PbG0F
+BAppLK7l8NDSAhMlRkjSeOq3fpk+dApQ6od0k3DIWYLWg8K1UI4vkoyLu47u4I0kMyJpYc8a/7V
k40myIjCQCpcHMpj3V71oJ+dcXho+pjdXhQGdfdp+UFxmOs4Mafhp9DwyF+6F9WTSypHIoCLXmub
N1s9Vnt4Bx6+m8CfdBC65mwOdppNyOtMYOtsw/YM/JTEdPg9k1zIVrzculv8EPukv0Jd1SpQFtzC
ZUhPR0UT6zVcbVxgL1xlCEvuaaJNCbNi+V/CQzeyVsl0cfmYJpMpto3/YF0D8JU5HNM/56pupAZq
zkvYRdeUKH8mYHmd2RJJgl2nuyeUa60NVVqvExzgzWV53GN/26PwyMQKxBgc6ievSZI9UefWrGTn
2I4Ff9TBQmwn0BvCtIocY35i3ZUvNJ6hgbl30QzU7A6f1RMGxs0l358V/9qN0kEJt/TbD+fSPJ67
3ZZqUBZoYG9BjBsHE2FHMYoV1znBF2dtmgFurGo6iH9i7ghVbKkSsJcPnOhW+YKGIrjm1q4V8vVy
4FzuJ6hfYjv9TWZUWN1Rl7HZ/qVZp6JGttUJqAr0tCOfJS1UYZpAzk8LnbegMWA4KBicsXusAK01
Z8nAPqWamJxZyKennsx2xSuaJ/3HiWQJ8bE7jjGUcH21IL5niexVQjKTZRw0LMk1/lZHmT4PQ1GW
pcGB5p4j38JsJWKwrLyH+jJ45TgINShbepHu0fM42K4i1ivygy75cnPeK9tTUA5LuxIUwP49sODG
ErwATF/cEmZPl5HiiikJOBxnQA7TJysT3VxMvTTTQezkQebnasj+Uvue2Zzb2/p1rdhent4ZDsD+
zaFCCMWkpjOSQQMq66cZUuNXNNJ7chTK0QziKzSM7LWfCQLFrFitK1k3XJ60+BAiAglsyD2CGTfE
JpBsu0xZiVPjD3JHHMnyb3lLN3zCEWm1btlymQ78fCFRwF0qngXLhmH0XkLOwXJKiJwEPSwCn0XE
vJweiogIw3tJWX8ffUFn+9I1JxlHsDgd1YEdHbojh0QtQclxVgTFTgK+ZbFn9U2rd3IIvx/JcRsW
VIOvPKvtJ2rG/d6Wg8KUdttJQXJ2UsGgXxRCSN+dMUDnsG+icTbZGwQ+RMYsUeJ1YDn9aSSVsetX
m4ATUWrwy3MW3tM3qpEgh9o900fihRWX4QyIP6P53fbc524/2mtDAzqbA9b32hWz4YgmqvzLjtdb
mRQ2y4KC1xazyCD4Q23bXUg4AEspfesKt+i7POmZICImvz63HbRFe243fRDs+MKgqAXrPSogbtMW
4/qALRzm9J7q1lWyelbvcxzADOo0TBVB5CCdaIEP69iHarT7G0DOUOLWa1NR7CRFruCk84PLipE4
XZ7SIrlQZh48ycae7+Y92ExnrHFjedHijpmdI7l3HRoGWtQ/wOYW8zHLOgbPGCqb5LgcPEvChMH6
17LQSrqnCGyhZt+dyqy3/rzdtRxgecOdq4aX8GJ2QTa8h0KCrKGZXJE9NJct7cmVu3/GHC41gki7
WlHolXQJafUN4khx/YdrJ3EuDjs8bU3Ps5zHLqDi/REvjM6eLZxXReIVvtrO3RNmkqaQB/PmpBH4
5aolvHmg9Vtv8YvguiEC7Da5vg+ep5Vw/4ixRrReOIPUUwc7zd8SZqjUgDQo0WNao25hV1l223MF
LznISJKuOiNuygIl2npaSMcwtEIrTYZ45upHzVk+4MS6DZhuaSYKOgcI38959rnSu/sGzMfryJNB
2Hl2voLuYnZz/diMFWlf5be3Rys5Tto97kG8j2uqFuez54Yzd52mFvSP1xs5SXJSrP9POeH1l1tr
283SUoPUmRrMulUacx1NmxilsDp+iJ/dLD8TkO8Fr/s++1qCV/FXS6dcCptCvkas1gBqZRsdPt12
e0VWiozSUR9G4EyjAhQc0BmVktXPwz/DeYOogiAWuXAvTaiUZGvcYheMcYl7XYYyw8pJaB9jdZGV
Ptv0Ci+BqxKtHHFhi5VsHpl0R7R6cwX6ogKjt+sU9X2/YOSLfKBjgG2uajq+CExgdmdAUutri3FP
eP4NkZOEbbbD4PBk0mWC0+Hw2m5xTqpS8MRsCqPWterRYYU9zCwr0vcrLHIGUKRAaRbpTdWmooVo
G3UmYVYp1Rz/5B0anwIWfqndco8uC4M8spIgEuKMYn5bGHCVagNbU7xJDEoqThY5a+FyIPh7QuFJ
Fskj+AAnYhj3Sa82kGoSDcySv51fqzxV+FJmwV5ckMNNVGnxcv48CHKQvvSv4589uxceQUE1VCe/
lHzKwOJVoiRWpFLc8v5Ok1qI9357mpJ6adSHljqXxNl90qn+Ty44vA9rUwmky7oqyDSlFUkSBi2+
WuaGKQ7b/xoCP1qZUTtKNO1xfD03Sf4f7G7UWYEJCBx8OTOyDoRwhQY2vI+gHOiwZXWBkmPJ84ar
iebzFCBJp64UVx8t3Ue6GPby8SVjgdT3X+dHmUJ9k/BhrkLHbwe8WNjKaHuAulqZu97sR8Ev7nRA
4iw5AsGcu7GAkzaHIL2zLC/1hUVtBWjuweJF9g3z9lICuPXMosYYmvrmjgBX+FAbqDkqRYVDbTL6
b3CzGh2pw8vqRzrA3Hkyf9m9NfU9fGVkjy3NEXoVebNkGXP+/qZ4CeYvOx4526HC2PXaR9hlvm9D
PQdJWL7b/ybVE9fIesREECX994pjByz9kD1xNKf2gMyGW6TUdaCn4jbIkQOjj9x26oeqkd0aZM75
+W9b6gsPhUwm9mtrCJx+lImMySd2QLapbf8ZxnZ0ANXTgYBA7OteTLhRpqJkJ2TgYtMPUKz3LdTP
XLP5TldmVOcN2CY6thBUU9SKMUbs2Epz6PqbTlzf9dlbIwxmYy/qBozm8RHpkNqfGLpfUxzy0Q+I
/lUmrFPOk9WL/PjepQm4ITR3I7AYHyj09QIry2fIfaai2TRZRdRoKTJC9cpzZs4AMINifd7E+rT2
qI4oPI/w7511q8CMQ/NFMutGjJPmwi6afdPDJ8HOdgYA27LGeuFqV93phcoGUZ3uwIuSSdE7HL/7
hah/H1oeNWnUdrod7ax5bnUUnvudiUXCjbEvYixUSCJsrpRUOUTlPKuhOnjV9CLS86YRA00Eag14
r+xKvFFgEXyo1aFAHixXomuGqd3dGCY9C/xcvKxZlNuUTvlrvDdOkkY7ue2MWst8PCqEkereAasQ
9NIsoaJneW1zgde8iDZ2139hwZ/zMCYUiMEYQ6fgxfrGUKUUXiXzVnNbtZz699NkoM26MCEQTqdg
OWMYrrFAwywkXxSrZCcfpEzv20C719AAScdSQpiQSaPjFcS0hcsRXLm6sy2w6SzD0VXUzCWcQSUK
EJjUPq6r5GIPPqSoLe7SN+axyGGqFl5OIgTVoAqoVrB/qa8ClckzRbI34b+PMsMN/V6BTVZtrb4r
SXfVpIZ769/OPIW34UFjbxhXmEiSR9ACEcqnr1oHGKHLlAjPmOkGkFFs/vdq7cRGwx8j64lY8z/n
xGF3ifdZxTGNpv5Fdzj0k+GZ3Qzo+xqwGHP8xqXhAKyHlkHdnNu/666fskoJZvWfF8illN27pNb1
oC2yT6H6koZnySyhMyaI/+kknxZZtdkUxxT9zHQtshOMatSuF6aHAEc2uMB0MlbY+++tgPizH2EA
XOsfGx7SkbKcU1hpK5R6Q3XgR+EEfPgjmzpwbhEemsuvNQc0lecXFTxiAMNGVXRnMLMbWPcqniT0
MNlMaAIEq8bOSomMXSNgAjnAggIfgUfZ/obzQXdAdKkysJs+w3H2iS7kYOE7UCFtIrM/OcZi+6uw
ydN8+LG4IGjNUnlXT/5BijisIKAqjpDZAQShyofxUJyo8b7aRSfi8YkIZVnAu/4lnThMcO1Ax1vF
tH52w+fnxPtD4G/P6++emRQ+Rm0pk+cu/BjthDsWhGLJ9KOw82taAu2gINqWi5eAxtYNLBhByS0Y
jXSiiYpNJqsF3tbnZLmc8vxRzM91OHnHH2Cj/T7Zn4UeaWKxzJbiNAXNtgtwHrb9gNBLP1sFV5fu
zzAvj+PViqKVLk3/1HlJJAy2Su8hoWKeWvNirGMXJOSPmpzrKV05qyoNgDIz/5h92U9o1u8BNurF
wvFZf+OVGsiWIZ1fYAUlKhZ1LQGUaGXAqT9xapdpf90/5OX/y/pgtWFcMQM7maevwUvRmZu7lV6j
0KVKmH47absFhYJ5gzvxcDfRCooYMbBb65mLlIY8XDtl49XgUbeyVeH2c8aO3Hj7eUqzpNsEyGxm
/vw/6iFsDAw5KP28Q8N1kOsqjUqv3gW6SBRK55nkeH8hfzv6deptvov7+8o21h7hGQwkaHVXc2V3
bPzEgJyornJU87sgiKddYMUPfcq5SB9bl0xzd7C5zH/bYXXTNMz648fOrKByz+2FCrfuCNX+aaYI
UQQFOQtfnVw1DDD3TeGZSC+LV6+os2udeyoUar+TmBOnSdOnyIJ76paG93InYl1djlVrN07GnCPy
6TBmX+hqLr3IlYsW+xbTFjQLTyBQfxEa09d4nUp2JqJNbi/irBzQHs6d47UvWsj5/79oEKwvw4g+
OllMH3v9OMh/7ibjMGMdKh61FaIBKumaL/XmNukMDVL2BaSS6jR9Ylszv0286KCy82DMgMREH3yW
9toZZQZcLgBOHDaYjP3SRRa045ma9zZZypold7BZD+tADRkFkR1MxSb91G1hiot3G1qQrOxR0sAU
QekdEskxZg5l3yeKKqCMXTufFLX/Rjy+6mpcnaqXj972VgoVIx4EBJiEflOa61PgNjQHZSFtBNdk
OV6jLKZ3KZsiaxC3Zayy0DpD4IVvukCVa1ZlCzEFsjkMAX84R01RII236y1rupk3PSaBMtVQudG0
S3uGS0YTZnSoinWDUGfdhj7ibnMTUZ1u5ITUYnenwPqm/Ynv2IY6CvHysIKz2Z/HNlIMSsCnGIoU
+hQsbjf+zLGFvr+YoMPfCzYT27dBIwpHVL8DPxqHnLN2OYGeTb1xlqF9R42xSVyGOJjlv1mhjlZd
TBugBxllOgH6QBR1H3Y0JtRjfnpXgRWpePOVPem6CGvslNhtXT9x/LKyLmole7HdwekBG7hd8V0E
ZRyVW5McrLO1K8B0KV4cbdqE++0Hod5G2RFRHegaEaC7/+kDwMERFXX9Bhlrk7jBSUny2aEtunnT
xALjTj/ex++LCZUEA81iSAk2W7jXBdjyRkQ30MdIlFUGv58xVW8e6ObD/PfQcIMPs2YCviqBChWl
v05oe3CLw58mNF42vfccx1mkdIvej9m97GYgFgYifeHXYFr1yP8ilRTQRdGbxghWMkQzfAba2uhF
/wIWWhaql3Uq7JJ8Kg7vNSY8/zX/nWCdDdnpBd0i/rkdL0XF3b5LzA4oI3Ncd+iZGBOdLTLmc7eb
vsylEufJBhz2ZiDvzJeBQqgSzpVamhnSmePldQvMfB+Qw7NVNTSV0bSHeGO4MgVbwS3a+ScR7ST3
xRB68Y0DGFHApFoh89LJpCPGFo9lVRFdYDboWzig/VmnzWoVHMvbjLQPvv2pOcVbaXKym+n9YBVJ
RHQg0c/hL/QI0hZbqgG/0cDD4zAbvZnfOZcoNZDUrBs6y7+zjxlE9TBNXICkO4m5V4MuB8etFg2B
E1eoYOU6Pbqf8SzLpGJX1wg2H6lnMf9OT7Ux8taVAptujXimu6pENwnPCjHtyEmUgvHGfPe549SC
dYa6Gygh03WwcEcgDtKkIf/oP/Hl1AEkW16vj/84ZKk62okTRYZzBPPOt9uEk7kYmfu6c7MHxRhk
Opq1WTKK/jMV6mCWcJCDh0N8QKr7VluFeo0/RhG4hvkXNLi5PBRNo/N7hF0bfTM2tq5FFz6pj8vX
xor9Er1dhBweB2nCapNuZUl93x4I7HRyXIBVLY9BVPKnhCMTqc5RyVycdjltlLkTKiew4ZlIVqJk
2X6vsPyobB1A3hxs3wkicRQFzayjE2APblgooTpTyv64Xv4uXdzhFdQjyhpXibQkwPFDBfFAla4p
h7gLRL21G6TO0c1w7Qe8ZZpRiE2t1yY6NWTz42GrLPeLxJfcDzC69kOJNsDzQyxybFfqc6JeS0+G
pccfzml91YBqCjxeWL/ZMlUH4voduoYPgkmrfzbezQz8nVkO4sK/Jz8Elgdo/nTJsbWvELE3OKs7
fjlH6VVw8k7pd/Nm7pvqe+6RigSv1doH1cvVmAAZUiTp6oR/I6fiQSOOY4/ThGTmQNmk06ELVjVf
wxCbRwjslXkBVkGa5zdYheIqbkG9qmc0UXHQWDRNYgjJBlPQv1EcvS0gn9PBHqwqyXy38xtLDRcg
sooECutWlvrnXmJU4vf3I5ViU+4J6h/JvfwGsSs2zDyOB0znAb0UI1/PjDJwkkCwhtJ1wWh3D6Z/
xpPvXYUg+QJVaQ7H1b3hGlGdBWTWhVrgo1nK/Ho8aLgHxt5DaJwcGu6ZhPzGDnjuKpurlnE7Otcr
2it93nFEDY/w+nCMC0BFombO4opk89DrPise27fSu1nZtUNzjOs4ePa9NHrPmiqU0NPuNKl6T4t+
pwCtmPP2IuwmFOJLcOkfuw6HWqnGaFXtVnb27miSO/n0OPkUCVCpUTu4F5WgKjdQBZm0GCeU3BYP
iccP3Hj3BE/5xKBFe8sQ3l4ccARvqLYBgICc8Jgv2eBDy/vgPg03cp482pLmp+73BhU8hwW3TUmu
P5Tsy7qLc35EHWt8dRx0LbX1flo5YYhoiTy0HEjWtKFK8tfx4kAnravMCOKtAbO3f+Lk/SMwuE4L
0IDAXoE/jePJ0Ck5NuIXJYkkflSqhqicbs4vjH9iL0kS84tlusCa9oLdC0HJYfdZ8osOYsIDTD1W
+I7Lfgg/7cgihQkRQs8zNejSGUsC9rLKqswT3KIAJxDzupof1DcqlPIG9+ntA0QOjsK+2qGNcal2
DvqkJC6oAiv+vRANME8WO3k/ab0zQsXFGEnbG+hpxLuuVyhifkwW+ZQKGrPe39gmXg7SmNXNF7g8
TFkM02HC8N+65qtf5YBMJPAwqqfnP5MS1SSvnR7RUC6TaGNr5insuBhJJ28+CS5QlVe0J/WNxUsp
bAHl7y6mdd549VRtOb3yVFIyAp5+2l8UN9ZI7FsodrKu+fhr5XfIvepvLUz7CPFHHP9DSwlmNIHb
xlgALwzB8Ahf30upDXp2Eo1Nwidm6Z8eLm5ZzbgQ+sk8l2fRTKUHVfZ6cMQyHKyZRnGbTOhqgDk5
ullShYyV6MDULybmz/qWOM7NiIry780Z4O0H6vTqOfHz3op+/73sLDZJ0oqhnwuW+Nk6bP8MNWqB
n/Roj112uOKT5n4x5WO1e/Re+v1QIm9qMVMivBTgIw91wYon+Sm0+3izf6opy1QXry8y4q7Q3Rva
6X2QJ9UksyladMz16GGibquejoB5TZDPkePKn9goE/pRCHXZ9xRXFaR88lhwQ5NsSfUQP5Ag5uIe
UPvl8e6SO/fxQfkgf7z9Zony8vxQYxRint9iu8P8V7gjyNUN3zHIk49jZwwPDJZsQWjmuw23RS34
AYBNwN+4j9iJ0d4hqxgwvCEljGHkKcp4kjCNiscnLq5d7f2oorOORBz0kEM64hKA8NNFZChlHlcG
7w2DRMtzDIZ9jjbksKxeA9FhpLjjJaqIloK++ElYQrLR1Je0yEbGmzrVDQGtLgJUJCNnBorbWjjU
puLO6EoI8+Pb8ZweOOt41QOSBC5vn7tiKdnjog7CfCK8ZGzMq5ZPswDd+xKwN0rxne/dz3lZs7tT
+U9Am7Vcc2XZ2Xtd2t0wnJzXMIfdn8fQhf8H3TRWEOyVg1g5RLYceSC1qEGWOhdbhWjk/utIWTbA
RzfPGZi4s3TMXrkzk8+EZhytQK+v5eRHeym/JNr+cS1W7m+MkGnMENww4j9MqmLUrbepDaDWfs91
Pn105sKXziWtkxbmk3wr7hvr1ueim6bNZ7NHIvjk6cH/KbH0wXXHVcx+SG/Qekf9MsHVF7itnvYp
3PUW2KWlQrSuwa6Fu2HwFOhSpyYBcnXkPhPT0gJRGPDkaXV5KVhpMAkGZvnb9BgbM1TsXO2uVf1Z
5Ge/vK2W5dIVz7FrGBqln1F50NmkLOJ9MY/BlejmU2d1+yJGxfmoGjuduMFWGOKiLpkuIaauFK0g
EmwECd+FtmoSdIO50suI63DZstGBSMXKYcW9cBkKD9yrM9F2L+OsB8+bEcwlMA62OzO5236taWOm
vi9X1sMeHpXrII6zjpT8uaHHuzjQJcnqbwFQzSX6rRZWXsPjVp/zCePrCPwZ3RrxQ3hGDduIedJv
yQqWv4riU3pc49suTY7gwPcE1GTVp7MC9b9SxlO2dWtclvZ0JPeIWxqVCHUyke/O0vw0dqtNRLwm
NATNbZxuPmCCU/DuH5oXdDaf7KE/4O0Wl9d8Q7Cbbkj/Zq6Xm168dMUcAgVHHgNtYiKlmXn2lE5F
26G1okp68P3AZOMutLMrLwuBcCzfMjfgACYQDxxotGnXTxCoCwZSRrB/un5DvCbWY8jQeVj8N1hn
Kq0+uikR4A7y+240RfpMlRpUsXHoAHKGj78oo412g5qZAbHxHNHAp9vm6jPo57HESUB5BNLKZ+jZ
CA4wC4vUmekdm4MVnspOXfqveEqWJWktyzfqKBBzfvnrG2I/ccrA2khQLDRhlL1jMoPAverxzq9V
8pgkQ7do9s1MN8CQZxPjsOfJ4d0gbZ6fQci5/wA2yEQ0hm0MmrNWOslyR1etC+IMN4SiVWn/Qmm6
RDhnFp78VeMDju/cXuHUgd7beQ4ip/ZacGwhemb6c8KGlyXXkonOE6Q3GbKDfkASiiRBBS8gLwlK
NPzJhzF9YXRnhHKdkCX2BMsMFfpQtv/eh/yqtiRWouRouL/+F3dxprVLrOaelj/EFNNBor2jUZpp
AzyQiJG4sldw6zaNEVgpkruiESTm/8jfHoz1uHUfoWZF2bJEKRTOD/1Bpwwsh5lMmUYT/HXrqfs2
h/92paDKkBzPMTdQ17Cj95k9iIjgVg6TqjmbHq2ujSsWJmrwVwhLOlOMqqktgTrD6XIAk5XtXWiS
EhVHh77lHB/8zH8Ip3MHPg5cXbtrTQi9QB2cSZEt4RYgqCbXtaxEWwLlGVJa25A2kgfRjxSAVbiy
YV9idn19js/P9Yli8ZRH3zfgJQbDTeqk5hwkYJy/xDl55/M8QEiKXFiDMopebSd0SeDiPeYikSTN
voJnVl6CR8qvZrVC2zJWUH5v0Z9gmAXt3efdzkk2L1c+nDBvXh6+tO1R/wAGyn9829k1Hu0a8dkQ
k8Yq0v5pILXMLKxMZPN8cmUT36xqyhZabWk6vWzQLy5LRn6GOZJNS3VA0lklYG5+lCbdyZCZu0Qz
fBSpY67StUR+XoteUHQix2RjUaZgTUlrOtYOGR0wcLRwvsdcNxly8UPQNHl7vZyknomYjjFKsxaF
QOwnSRuOEhKwRd+B1oD6FOCg2I64HhnR8HW8axHxCnWvjWrUaWmTQxJgRIr126GGm6i+EkMeSG1c
YtEvs+g/XwSlhSnqsmVm3YI1ck3wd+BYhD/hzIdUQAumFLn8APi07ctD8WCPch1Xlp677Hqf+08n
Z9QjASBCWw3BEY4WsdY+jT42e87UgC2IV79Ah6d4KCiFJH04V5tx+7wIIjNMd7vQFGSevMPtYm4s
PKl+l81yhKH9oNwaUI7MLTulGuQfUvyEHZkyCVU9sYuYG2Fag9S9ZgXiaXEUKqopBo4gYXHi2zT2
8jw06EC/ERJfkhdmsqgnx94RFpv1n8bDeQlrA/GcjogmaIiRY0Ft15yK7ECrMQAXYsxbtvaUl53P
S29xeMHxEH+O3FadZR2WsDEahWS5GAsDDlucPLx7/9wfL9TRV4hFypt/hyRVhIGxl2il/gn7FjcE
Ss7wQPX3+c4aM1QQW2/2lRSoDBjTnbzeCwCqvyXqnw1faeoV3qDmvitAR1HaUjrmEyTqFHW38wdJ
umBABG+svpFb6GwG9rxQW0FrqIM0jmuLEESBFUxzBwjjbgt7FUwDq9W1OWlllEtZg8RBlfJSgG3K
hf90xcsJptdAZUPrOiPMJKiO3D3Nih6hrJRHx5dyrfeAEdOFwwY1686ofCh/OzPnHnB17Au7VeSY
fPQYW5M0uJ+vBS+9XFdMiu9R44rQyqbfso8Iwu2F8LyUhlx19Wo+sEuZRuqlAsnT3RKHSlKzltvs
ynfqEJ+gy2Tvf/n9lG25kibagNkNjrpwakvbg0/wdGVTJzgi8ipP5pKiSV/iuIwtdD1fbizTo4Iu
RC0lgZTxmonbB6il5F/MvqvZJQwUIFZ+Klwn83FkDqVs8NbTkYKNdNWJYHWcBUMt1E1rDVaj25XM
jFbBZJCvGS9Jh7pvlpg8fKz43PZ55n8h2rtxkOBj2sYKoC+sx2AU+ArKW5Ds5qx6wMOW9ZbhRl+L
FmRygiCKwlVCLvvPT2uwZldVRj8oUjCvX4aJQ89X7WmcRrk8vzj8yT1E3sm0O1uCmWjTGMZb5z20
UcZp1aDF0OmLTpX0B0k7FHIMANs1yctgSDd9iavHXQRurOZldLkNvE35/sl9fu+JxtGVazEFyVeT
rj85mTqfKI6LcbVh4qV2UyU0iiHmCAzq15fpwNnyJaNJMNYSFdY+4WMZv4qkzHwjCo0K4C1CFfUX
wpng8ySxDfYfisWirf7Fksl5wemzvCuHY5LR96G30Y3pBi4GMcyX6v0JL30m35NIGlMTsOZRT1WR
/E6e/gc2agi6EVzf6uzgemMYq+sIgA4GqPiEQlFQ68Uirdvpn2gpvc8BL4DGEoNIZQQksjOhHqgw
5ZFuZhwNkdIfmMp0RdRdmI6i/WqymzWlxznGxdIe+Z7s0vpgwFexAAAR0lOubEGpRqtLXAu9/Fgl
su57eB+agYE31rzaqp+/AYb5htV5Juh8+zrIjvH4UBaXntiYlS+FVUDRX2U2SS0qRjtjj9C7Pv/a
RlSlyK18kLxL8p2x5W+pQblIj6f5/Xoxp70uL3nbG0JZ+hKPHRcBaqq/9I07j9GeOfbp+q70l0jH
vkYxf4UGyzNOiblq77bGbL2WKYWlobgsHtvZBwUz+Y6h8wIhmsuvlSq1JBVdZWBWxVk4NH1ypwER
DD8iDQFJlT8eHkutJACsbQsnT9EY0//mB8FZpseA/YppzBpqmf7J9gcwVl+wys0/onwBa+m/2dH5
DPnofh54ufy62vy+oT3bVlAKNbqPT+KRbPYiIF6PuUreUxM2ZElr6keEilPhEMTs4a1rVZmTVwaR
6iTHYs12YwKPcXvskK1VnL92iVfhpS4kQF4dTynhpl9xVhyuI7Lkxap3JnPK/PZExDCC60RXdTI/
2LMj217i9yta0FFmtKgK+c9VSC0Dlq0Jfns9ChaYiieRM1maPtoAXi892YxsNdirHv2R7YM21aOS
JZ/wYgSo9f72mpvTrY4bV85KqpXY1RqmrFwPVi7HaSP+Pm4rfOmX6o3hjl/YydfPFeIZjSZHckF6
tjRd9o02WnshFmmHft7sWw+1vVNJWan8ZEbpzkcyEq3wjVsCmqAyDNaNtRKVxnBrWD9DiXF/hKZp
miEW7pfH052ncLnLA9dcy61Kb00qf2+yNJ7J2mDzGqIz0R6Xgy0H9rjRfc2Vwt0jX5A4vaidgqYS
GlJduLxyJ/EAhPbz1DieBXdz6DNWZMz9Ij0GAGN15UU1qaUBFcWCW93FjBiGeYHbohqsPtYD0Bvc
VXvKez5zxcJAzmgXRy7XjhoMcDqBcNX/dBXij1Qa+wxz2BT6x7Vmsmj/tT9CNoPjwS0U+Q2W9SgI
WNrnUU3TpkuuT4bcemttEwOYN+u64m7pjagURfvkElkfB8CVkk8cr6Q2r6PjIavhb1/BbiXv8C5Z
MdDBjqQ1vYlkMRrrY4xI7lXNbXRKorrJuKXrNtDO9l7PGLSw8VlFPPz9qBX2zJqCMLSlVaAhuMrt
LE06asS/Sh6Fkafeha3pgNFRHqUwuNoe1SmAoMfBghjDBggwtKt4d00oUtAFsFP+bQX7vAm18h/9
Ce8OkS8eIFt/tVwWfMwSF4H3m72ubHaH/pI2qwC0eYB7tWkYrRKAYO6UMRqv7P6EBXX4qZabwoj8
RwcqxXiuqGiH9+HGVnjke84jyxVeuE9tS2YXsgkNIUfwzdUKrQjOrqIXXnHMeTr7ZqpZgRmIF/qN
Leh49nvW/bTPw4Z0jwf5qqphMQvXddomUeDPiaFQpPkvO/K6XWSMPX7DOJtNmciNplCF14qKh3ZC
uE2ECIByTe+Doy0XYjLfvC/UlKD9KQwPFgmrqkbXZkSUwm0SRK1HQQWPYjYIn9KF+GeGcz4cBHf0
fD188dKAEfT3UISyLZR+utHKO2DEQ+OQC9HnQ4vSwttju7tl4tL5kSFUH8gPrwLGHh5jAP+VRd5G
SMUP1zftjSaiYQL/Bq81goAD8qG5IsUv1Bb+7oO9NfLB7otimvl7h4rkNMrEegDxblsFloSDj5HN
Zgr12Ma/4xBHh1HXZDVfki47XciKTyDgP5wFmzJhEZM4mC3uXjHQl8E2yz+dCpMkgA07rGnLBtM3
4JiAvp8choICMenlIM9Uq6U8KWlydTiCxb9/YxSMw5XAefloUUR9eETI4gkTAljLa9oTtUHVf3mw
YpwI90qscJe+iw4SL3PuWq+pwjPl1aMgubwYrXOjPikkJRN8VNiwgsGjxghb0EGGIU7hKeAomvJG
REn0Aonsv7Z7eCjDofjoiqGjCPhfzFLyacLsxWRM3McLW3u1s+aWPXSA7xzeLaZlVLYMczG6hG6E
DsT97EOSmkSf9XVH54dRo/63AJhIvnNsMqJl0JnmkOneiF7vqc0GqGfgiM8TeFU1yD3oLfK7VcPd
Fk5vqwIDOVousTeuFl9vcS6BaiKFx1/vGSywNPE/ipRf+GoHQT8gzNkNE8bxJW5xLWW2SLudYTuu
xe+296X2ztP0YM+xllvym6gcB801LH8bRlREZzVJOHsQuphWRuBoPYkM6c7naN2+3D/aipBAp1qj
9gYnY4Ej9S02jiFVW4GROqL1w6RTM0c73qM47dHaErgKV8O7UAK4iJtdgZywknUuVeb//PxkXg4X
P72qdUhfB5CipxECJg5oLctUQQpFmtZpIRCe6ZG69622dtc+GuLCD9EH3JXCC8/7pF3Ce6uYdL4Q
qj4ms6o2f7ffdSc0lMsqSAhfzexmX2TRhMTTlS9N1iYDnIWFTT7CAC5PvpNhUG8gRKpf94NfiDJN
kwFAhdtXHrotsyd8RtsPtzM88Xlpc4zZWkr0Lq6H2KPEZvz11r3yO8DiKBmo4Sxi61nmdhz40Pjr
95oMH6fdQ9W/ciorNDx+KBfrzNASRX/cxXZeyflEH03Tf+i5VNd5S+RFHuQJ8pQlfQxvs10leA8D
iwUh3sVto2wVpobJF2wRCcTUKShbwbXyZn7vf3O565nmGuSIdQNUddjIshcTJi9ocsMM0CzbweHk
E+uBGOtvMcANS+Z3U/9ySo2h4j50qXXjQEYqZF7mmY407ICnO95TCLZzpGv6XPsnh/gIEYQu98nj
gixE7dkOFEURzyJ2GT5vSB7251pw5c0CzfZkdRRpWzDDmKLw+19kRIbD2r8Py6nwkFJZzjmSJWtu
D/WlZBteRUFPWgEwe4COUano1v9WoAA8u+glmw1Q0hifgWMj/4TVQlXvDIzUfZs0cKu2JEVOj+k8
X9/s/jtHdByF3TpQTmtUJc/RSGxoQcrNzlRGpOKXvt8GkByWuk2kh6ner8yXjB6M8RWTD5iX7D2N
JjkLP/n3zVpm/F4fFrIfGq1pQGU9Pr4Brlzt5jK0jG1zfVM/PysAh/1Lvu2ArERhRBk5bWqkirmJ
/CaKpaTpYQR1qBiJi45Q8n2gc9WHud9dZa48KOXMEv5npkjujH71o7P2p5CumBNJakIY+cgFz0BP
AhJVrbydjZLOI2cmueEVI5MU8D1sAwCP5wfq2uVqC7KIFW51OOi49Jw+MYYutfq5KRt3R6l+/Tui
7Y7JhDcJFWOWnACyA3ahN8K8w0BuL9wt9HslivhYsDEbgRTE3ulArzNIkoETY9ruuwxp6A2cMNxJ
mfxP5FyLlk5EcpFUURbVugAslORZYHX86Z2ELoGqGdANRbmOOf7OC8QF2u1UQVcDLNg9R+N/rytT
FA7JlQA0/A9+aw34lk5q27sje6Wjex9WVFZkeKGPy2lLRp59uUW8sCAQIw8VtPhN+Tty3GZ91aSY
p6T2+/oshTlFHV+GgRlIXR4WgtGOjYDeMynG+B7S49GS7cXUtf3k0cqO+Aqz32C2LtrIkrFkcS20
H69qs9IU647Yim9bus2B+PXqAU1TbMWAgAd7E/KIcNN1T1QDCxbilUswEAs88f3i49mqYFa9ZWRz
mnf031xZ7pA+xQWGhIvjqqNBee9aLoPNPFT1yZyq/+JfugnT8vB/9XHLmum/fqC6yfKSvvialvE5
SpMGaqKscLJb3ZPXw5waWM/Cky56h4NCPGU4EkJvqSKUugEZnHRLzqANIx9urzFoHPVBlKsJYSfF
0ZdDpC27tIJoyGXKl50bej2pdz0V8kshbm2ngCjBE9w+nTUjPf2fs3aWe2QjCFQTO0NlW1OOOfXY
YaMltI8qNdm+kArYzprR4sVwEjdNsyJXZ0GG+i2JaLQU+m7BgG/uUEjQ7WHAWdjkTg7kC6CFLMuc
Ahn9q35+F1JVHYEY1J4v3JsFb41a/Qj7d37ZZrwX7YEvAk5LleUwGvQPCOMf17x00o9uoZXyeOzR
fHQ1vim4zYjyQKPaSqDj952i04n8cInusQjHlt9xamFlHTRUOzg+cqOIizHHOgEbNu2bJ3LBa0IH
kZ5WyT2pgeX48VCPcXWnbEwZmBDnM1X3gmH0vWKx36bsFM8NWHfZQTMFjc0EX0AXdKYMKA8zaS9o
gVx8crNcNV0npnsk/HPpIOj2d7BOV0tVosCor6KcRH/glW8BrNuoMLYM5NF5aDqaZtqUok3rFzIM
AVQq5Fn3iRpbr/TV1PxCNcYlGuT34GM6xDIgnmH+T/cJKV5z6GaBN1H92ZV3FI5UZAcuDbT6kwM8
DCf476QZb8T8AAQ9CGQOFCpnvP225HUO5UsXI9mQsPUQjXm9npFHvrvTjZ7P9zCdYYpnD6QNyTDb
gZxRzk0QXmWbMR+T62WWV3fY3aYDtG3A9ocNIXH+h/Mau4Qbvx/WYt3Gy1MMXdxI3t6LzPiQCyx6
IanVEIntfL55Tjf6JpX2E5vY0DJ0AFmiCBxMJcKByYsWUoieAOVGxwi3/4dHaQtqeVnL1nCJ1FBi
XZ4T7KhpMqHv13zM0lbPIzHU7D+6znvnVtsBuJcBryrb5mUPYXaN/Mici2bLNaB8otCYkk3Bd3GA
sN3l0RwJ8dznegVBrErcyW70S6ckj4J0/o1ODGFVyJ91augfiQI9a6FEN6xKYAaLayJoM6sCoa7g
ZueJUxQrKbWh+9gM70paytA14ZQKaxbxs6YclpqrFlxxd60QduLzJy8LVsbHLGrRXNzs1YAIMPvS
EVtxa27/2HpfwlcfX/BfN4BpL3fHcFWMm47JTs4Crg7IV56Xl0QxMiaQlwg2AWMUygkSGcqi4oel
1FSxpjIhAvfK/uDUIpnHa4eKFSed3P+l1h4v0rZAIZeBjD80F3sVXgSKCUKVfTebLuhXn7DBx93e
H5CwhFrKYmLzv/gRq9/6fm7Buv0YCD/uoDRW6lYq6nhdyb0/1bFP38JKm1TsNs0S7eGQcoiXYu8d
Rnafsj4sRZyyrRxU3CH8Cp/B3+vHalDa63ip+YHnRS+nKiocU3o1VMHv/CwoN4ZxaPlXNwngKt5h
3xFwr3j1W1rD2eGy6XdGfqC2Daae6pk0lgGLg4Opw9ziiX8I7GIzm4tgpTlmSlBIUGFdxhBW3u5J
WziMal6u8NKpDyI9bgDus3jvGgcdZPEhFMA8RROarYm0Q0PCauljWPfdHDxh3aV7cu44SgvSUQUh
hiuUSRCgkrdPE9aas9uSdUeHRhTpzXPDkcmAtoT8lyLSFi60k8AjFKP3MjGQoNfYAPhkps5wcDJn
EonVd0DL4AZRBZkqk/7nxA9sHGSB9L/OaRC0qwEzf//Wati2ozGddDBc3RLBLlOOBQoQP2+CKVc/
dk3R1TPnkSsLwZCp7XKWovGB4QqvGiOURXe3rpozTA25ZUjLdBWI2+1Sx4VtoxVHAZjhb3sb0mUS
jK4+255Pm7q9hPF+IvUbp2GBOzQ6LiFvEkD4h6unqdQ9ynp7IjNvuP5p39zL1bojN+mqoUzB6fZs
L7CVfh9EUyQ3BLsEaxLiiO9gQkIPZFV5eb92bbA8RvzRfm0JTKlpA92yEpJekYZoOmost3+MzX7W
7ZwP8MChGdZMh/O/oev/+d56qtvpSZMDrPoruLmkgu/TPrQA+97HBaibJ7b3vKUcL7uuqSIiDPMK
ZZGiBOGiy7zjGRSZQNe4/MH5B857Dk72BRDQDnDQSkaUD6t0198mCXS5dbqceTRGBeHppswj/a32
NkuihuA/9UMKb+5hllaLu+3ZxybAobiz8BP1WOxs2Spj28s5usAC/zc8/jVfsyOzIepFfxMwsWYv
3qz+6s0rEp/7HQqSXQ/5m9+N4ezgNW6qhWnOzgsVKtsJ7AQ4Too6fSTax15LfY0hKSSc6heTrMxq
laBvq5WyVVo6r3r9ptox0TET74rTNV9l6dhomDRitQMStztS8JUk+2fJa6JoT+vfbuRSVf+rgpae
sKz+MwKK6yuKVVW+0kKMFoxc0KF5yAUTBucXtGMK3a5ws8Jd3DyNYE9ltW+3JGgoujPEqko8asIE
csPAmNaI7wy6OnTYW827gKc5LFsGul/f+hlR2vRRW4FEu4dfOY+/tVaB1cEcii+CVwPg7sYpD9t8
8kfff4ufT2dfs5GdGXcM90TrFY34di4Rvk17uTMv4GxOtUx3LzvquVd6n+/uDcg80K52D7LHBTmB
uUgVpK7M2PRAE+9Mb9muw1LnJ6GQGUcN0qj6w1ecfVoDReyCuTc0x5KhQSrMShPIBvd7yxk8eBm0
YshKKRuehxJ51ruti2eLrtPTp6pxE4yO2fmmvMwWleCDrM47zLNGeMgm0tmD/G+tB0/wgm9xrrxC
Cp0sU4d+ZDLJT3cifnCEEdfqCIpJYsy+xfKf4shVlG7x7KlyS7sC9Pkxm6Impxb0AUSerhIFNDKG
zduCOGg1gUi+XjxzZgU7MeMLdQjRPE2dUeI2P3v0fbAG2UhKwdk/1m/ZORXWhFyD/+546qmkeGj8
7NvEwvLd8mOrlamvTLEt/BSHz9BlaitiwFdeKKku+eCuE2MuEAmDGZn297JZCiw679txittZmE2h
vR1vpCpHweKwMdPjRC6ckXemQfi4Onb+gl8Tiq0C8MGYLGcuVw/RwOGYlD+n+wQbboUKf3g2CF85
gMHlQcetqnC+jR4PjD9PwvtPhTEON71MXRRabrsRKuC0nFqqns0Av98yegkgkNceUEzjOPafcGr/
R7098ZGLIXN3Cjv5m74mcJfG3OYcWUpJwGj7C3oH6hsYutAuSFqBJ7DOGmRmekHyVqZrPrUzdKsx
BPd32/RE2QcToZO/g95YpvdWVoGi9Nj5n3+T0M1DlX5bsW1a9AZFrltbiaTmjQRM5XXtWfnQN+Q3
xdr454HinaCYCaguTkUtCblzCfIz46O+V/2gUS804gM6mTpWwmyTAxNAtbEFJBQWVbNIO4nbGBSo
rlE8NstRPMSwvLSK1fiDe1PYBxborncjeneFFGtR0SsV4Wiq9CLZr4Hd2h6KYAJM6sy7r6qtoIZz
tXqCZbr2UTm0tl6K9ypRj4UnmnlT+ihtOJvcMclxdgduanP1y8PTasI/y/csZ7qtU/RrSfm86Bb7
cHMifLtoO54X1FWt0Q7LGL+jj+aDnE4fedOVXD5WLy/5kRvg+FLQaya7NuusI9N09M4awgkRRyov
QGfUD8bGRfbMO+I3NGt8mOTn3SvNFhnId2txPQlt9mPR6m1fVoxx/ncyJPhHp8BDiP/X29ke/h43
YeO2rpLUGxKKz/yQtOOz5/DC6VY03vp63BYXD55UKGdRpm2uWdBCuYAbI2cnSrwU1fECM/aJ6au5
bQBc31/caRq6jDyvycv8MiPe4t0NqJeLsoPHPsWRbq/VK26hYSCl7eU0A/1IFAQp2v9YnTWNIk3/
Uilpx4RML8GDHWKLTbJAfxKAJ4nFocD7d3vPgvWwx34hX5DQJHyXWxQ9K5axyejCTFl04JUmdtUL
r8WHLYnuheX6O2UodEqTOMkEWjqaA0NDi/YoOJ28HtZdAzUVYDo49TGgzGXZZZ+WKw9YU+0hjvbg
tLVAea3p6XrtCECAiPPuJlgI9HXdzQS13I4/NBKvEt08ujEspJZg7uazAdsx6Y3xQku4ib4X07q0
iILovygauNqBlp5MwauGpN+P+IYkhj1hcCe93RyKgsrjHOwY7Ze8SPr3Pz5rUleEZZ6KPO902wJt
LacO9aNNL6YNn6IWxgTJYRRv2CcrWoSFpjxVtuhuJ3px95TzKrlaAFyAfgdLo90O5U5za52pxbzw
YHYSp1YOzchSCw6lxJ1mSpz+YJFdy55Zrd8qbVcxdWhf4KKHolIiabiNucm7Yt6WPTI3wrZPRXRK
BseN59KyEYhyKPbUBrB1en9BuY5Or59faVpC0o3MgGKJnL9Ch74Mj452T4EYDIMWiuiml/qsp/9G
ujsAkQzD8fX36ylwb/xph7vOHiWgI18sr7TaF+Ycvxy5194wjV5KrRvmWaBUNFG0emm8PSAnb8g3
beKVRiAkSUg4RKc3uckagXI4Ddp21AMTKsjgFA2TVk/YH9CDESCqEznkwm5VGDnG2FrMVtLo5hg7
VPNVT5vojudOOo/9m6tEbFuUa1DlxCpqg+AL6yfaoqDbzbRQTlLaI3TO93tboOQDAv9CsJtgQmNY
lfG4Jjc1stWk2xUrXDSc60JW+mt9Hd6NN5Vt2Q5QbS+Fm0+Z0SJXaHBsGQWiSIg8DVBrR0bTLltS
/YAprKLBqbnoos4u3OjQetyKdnFVstVDhb83rBbX8FTMYI8YiTaVzpV/vJlkHBmF4RlBZ+qyfdbp
XeDLbGE91c69h3DYfJX2z4jtzGsPgyW7Wqug2VnY4h2+sWsTocb9cuqhYHzX5XY6ZD7P1PKgSRcK
Z/k1ptj8BicSgChaBNxitmkBhYIhCVZc1vTm7R86QL7gb/zigfOtGnmPZ79x/TizaYmPMigow+nw
ZM92gTjSILa1JtgB1VjqKJknvVBVrdG0cIOpRpnDv0baE1MYwTui9AL2aVKCiollSbN/YLoCDpZE
e1F6meWYXaKhWz/Aig0SQdJ2Lc3pnOx5XbAfp1mY2gBPIthoLCOm4TUbceh8PyWjPuY1QumOc3CI
eQPTuGIx3RFc54glZpZoWV5/CSUec8k93lg6SVv3CO/NUoFOLuAREPxlXYSCxVk6Qvp4hjkMxPJi
7itnE0pinBlSUmaK4m7YsnjA0T13aPRUFvXfyUJlJZknvXFDc5tPGXpbCi3aK6enpWxlH3YBV7RR
eT3jBzuBiZ3fIbDWnT70w1G+A/yirPaUKBW4qMbZCimR7ApsYs1qtZDMOo6qwXYLCuhQctYW3ccH
t0Y7IjPC/H+l7rURqI/DzwwpVB1M2xtQlznqK5ammbMYbpNLwqwfo433ERDhFVgywJJR4ShbGVVy
2zlE2UUIq+EgbS3T8Fom3PDhYo92HUPx3pr/EgADO5/Hy4rip9Q68QQpU5itDhHU6k1KHvExYpLr
WgZ3Ldfu+huGmTi/hONhfYGA2uFc29YTzTsJyNc3tCv6u/sS4q2Gy2mjpdaOrs7ITRj4/H8Xwxbz
+w9apWpQczWUHHVO36/EBy1hYjyTHXiC7kuguQmSdT8cxa08l2Ykot1v/UFd0vBSMC6howo2Waqp
Hj2JikAnx2mmuIWGOPrumd0VB+NORG416wmLtQ6Jm/9M0XhxklEo80vfBYPbnHuQtUbh0bO5f3D9
FDVKZeXyZo3BGN/Hb9/Z6ohu+O3u+VusrnXH2FNddx1XSxCDfPrzuRIJ0C3FBt7dWCXVpjRUhzpI
FNSUOiVnI+qjN3cp5hj9hhu67aGJ3zRaM7ujAKwxESkl8NfEL9fw6JKwlwNwS2rPqxxzHNr2Qwp5
cSP4om9qBeBGpbK3ReGqSD1n+OGGNqJm7qFlGYfhPqL7QOQewK0/bKLlA9D7CGQpIra27yjuzimX
AUAR1njmrBRQAVa5k9OHou/raRqSGADpZzhIUxs8TtNedOOwRn/1ci+QirxZvEkN6gXwo++Rw10W
VuCdNyfhaTltVmi4afl1C6w6cwkyAf28LAt1a7DOx4C13jUGBEipLIJrvgH4ILeYJq7ZL+XAU3XG
1DiNRgqNWtNOOS22yqVmwC1GSRwogtA1dyERZWzl6TqAyY0YIDgj15mQ4OMrDyCJThD7Bd/TKB0m
WWjHGp9l46XYDS90NFtQFYu+a6/HpN/MS63ZlliHw8pPQeFtSb93yIkStEix4UduhDVXa1Lq3Tk6
ETrx7TCi7MdmSSG9U2Ru/4HyG/WWQH3IdyjsrpWXhZMwcTGynic0axqt0dTfZuS388PjRR/4zlJ8
tWKOtukA8B4vKtkx65URKvQSFSMKdMhqdz8b3bJGYz52g12blqkLwPcJY2K0Jj4dgsxv7qhQPKr9
mf8vxZwTfxG/pWqOY1deruIzi9gxZEiMWnvC3bwAD5SFoSfGb4KS19LauKHRIoaPHUFBfcrsFmJw
PVcEuoTeR2wznFN3PgkagynIwnsmoVP9aAw8QIkDFmKb1p1tXTibMW0gwXyx9AQGccaEl4ZtC3lC
cvodsKYSyli/vqieZ1TgglcHIXNRAaXwH9R/3gPiJUD6E0MhmlHn0hqb0fOwO/boTBKxQMIiFbDx
OL9q8t3jWBYhbtnYhI9gd49DLJr6/A5pjvd4sGqYZ0TVA94xiJwsPgQ97/uTBvWv/n3E+tQrHgNc
8pajaIgb8QKHhJYl56U6pFSrIM6bJruQsZSk45sseClcNml0Zn00OJrTK/nmwbM4pPF45k0TZIab
GixgvuTs3s0UfL6JkprjMVRqRLP/zuqX+9Hps9mNDRBRDTApZP54FCyz/i/frfK0Un23WwnJEC8T
r6qFDRY5N6iCFyb+hqtIq9sCXivpraoHKVlhY1XwVCz+K3t7ICGNbnhTFwjlGenO1Mm3FtqB6yre
F112w28nqroFwK+/3GAbOsef9HNFwNi16d5gxzEERukK/+2eI/zbtnbJoWynnob+Z2o0ScWTU2l+
f3gP3Q+budo315RSRTEdGIr1Q/pWVosoFP6b38JedPEDYwoFm4D9Ro/iCPfI/6DinFm230k1JmAQ
zE0lIrPc4jwkMZot9WjSaU2bnubu9MSMByClpeC6LOMkHWl74QG4p+G0M5Xt8LkOQXUmWXXSYaRS
FNuoVsN7HHa22O62gcsYiewSxN+1xVBEtVJvRgm3Jw7cj0puSQ/7jCM6WrdvNqRrw9w1iPa6XL29
dnh64sthmwKtLb1oluxzxYRjIxH71FqHv9OT1kiNeqgiOCeps260z/Edy/KQ/EQi4DSUZRS3547j
ud9Et+7Kx26gpYxr2wQimtaOuQADj6Y7M705ZLThY86bX4nxbpoWXw7Rvs6eOtps5dFGDbj66XjC
MrUiE0VhEh1/ltHH4t6f+kejZ/ecCz/TxP1cwyfYIhS/5CdoLrGk4dQH30mQlm6FEKGt7OrX8Jxu
V3C30iP2nw3hvRknLJ4UcuZoAN6/4XnDxucW2Qh5yVTReQHWIGjWIRA/lkBLkDJ7ig6f6ZNC/Q0o
C4B15XqdtAuNCrRio56QvlML5/gO0oriynEuvmgJmamZai3rm/H4iui96mWsi3kWninATLBN0DLL
/XTpejvFnA2A4whfIzEnQx+a5z15ngHuu4yhQmx5ZkwILcFNt1cbvWJoD8fD8L0MVk1Tgtvs3ru3
W+PvjBBK5fIbmyBAud15trjbAA5h7BevRFVWdc6oMenbnuH/OT9BfHCTbHzRUCBMWTI67M+lR9HN
PKKuSOnP5jmzQdem7cXcTLeKaqSFDQdOjUwvFcoOAxUhvoW/BYXhO39mzJ1niuu2fKKAWX88IEfI
ibUwfPWn0bOEEQ6aEzRZAzGaZIgCcTGeZLZ37bBL2d5NmzenbMDeTL7TrqLgpD9xOc+02/Qxv6St
UOwHuZ+WfQop+hIQ+dlgkRG4nLRDiXTuslR8FMNjsC0ATIcJ2Y3bd+NYx8g1LkSWMN5LiFnKZMkq
+0I2LnU6YlfeaJchM8vTbHLRYzz81+LbUSme5kV6cCNJGTEKxi/zG8tBt7PykCr87GCOIBnfiV2B
XXbFT7LLFzXLgrfxbB9DhjSL2mSRWsTiFFESJwXJv+F1MSRRdxnGcdMdsa1azUkkIgmfZXAfHBV2
5tXOuofY1OHFN8pzhjRWLOiSlVbJevHdwPc4kc7YKswLpnaTXvdhwuoHk7EuKBtN8hRGN9p26htq
WOJYEfVYg2HAyBu0DeQtpqaSl5mT6vKXeRynaJL3XqNC1VsqdEnBVCPBIjK3wQ1cZVK9Y0kZq6WK
0mpQJBNZ1mWsuOTu75peRI4QhwsYj8I7JgdNWEJq4f+o17y/p64+HqQ+6uGQ3S8Z32GhpqGB2gGc
2tCoge6tET1JiWpUfpg4ne56LYmZgLi86BkhjthcfrWhk15CGxT6HRdfNSBdEXf2BNl2utEZCxzY
1lXG4Di1J4PlFC7R7/IGFEFBKCtNs5qiGlVUKjEz0a7B+f1dcrrPSCIvorZzVTq7ywHc3lOsnATV
0C16r9E9pvZ437BQE5RjuLT4I9iPGs9+58CSaNYzUW4DTWroHgqQ4785n4/Qg1NuRkzczHALW32M
jwEDcnPiNjf7NBJ5PmoKW3/TuSDUJ5NeKzcmaPHC4AsX0Mm4ML0PJeI6g4wYKrwO3YbqMxhM4AC6
Z6KqaloOfK8C6weUhT4uDhhH0GRiHSTZLg2X0nLTwBPS+xL7vBrporaVacgjgDRXLGAh+5cZkYAx
WYiNXHUNldIWlb0qkdhKsV/r9HIQ1beaEaKykfA7iJ3R19XZ7GaNAao/WKGXA3BwD1INd9KGs2B/
+JWTGQ+NwBnLuRpPw4UCoAQ3FCTCUvidYAYNUmEOF+IHnu1pOBfSiETLCdJbM3hBj04VZ1E2HDxO
If87aUQ/FEqT6SF+Oo5pHwKs7nEgFX+Y4SVm8e4MTAk+Ke6KAe2O5buYNR9rCUayZpakp+3oooaO
zQQKwCzfVvcnzfmx0l2B4cfB2qSHO+2b3lhqHULF6SSvLmjkOW1zb9E7jJCDFd43O3x8S7hBRt7M
xQieG3jiFaFiRjTr7bNJc8GrobemTqmED7BWfn7BXPwgBCqM/S7US6xQDX9rxgxoJF3YWf3AiDu+
J4I3niNM3ZWndxq/DL9FYRHJeNeVpG3nEc9VT7Lqh44tZX/7htHF31QCNxVYt85p/yml96ajKOnj
DFNT43lgKZ/E03nzmuNeNUgDD+mN8Y2QLX2sxHAlc7etpH0NpL9T/vWZipBx6acSqGMx0HK6wgZr
s43bV74ciwwhexA1o+agndzM6PU+/GNd/QdKDGN47LWLgaCzUIFEqPgWZW6lYNY2wkfncMJuLIXR
+7PTRH/IRCo4i07fZunf7RIGZ/xopVeaMfvSpaUf+b3faW+6KnMbxa5GHaBwh5HLzgGbWI80/J9b
h0RsDZOz6EVPd3MMi2V6SSR7oByiZmB0qspXZeJ7ViL5+TrHFjsDAYkzMMMLImaC0o3xTCMZF3/4
1S4VoSr1ZvABvkzjHvfI47jp+5deRLFLR3Sr3Ibh5XsRDBPwhN6rlHIfY+zpu7hOE5xe5dJasQ6V
JDNe8/yznItDV2oRjjwSWeY8t/ZsHhlqE43ukd7uRLSHfS8CGSQ=
`protect end_protected
