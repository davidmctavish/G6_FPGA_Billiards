`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mABK9ttjnUgS3HNkzOkGSjmIPWvZf0pxvpH0FZJb9zBnKKzXmpWXAdRyQjFlPRaq+yrtOWXU0VQO
aHYKmwiyGQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
C95QoYUXGR7c67z11LkrkIpMM7hUQNjvUoSlr+44YimUsocU9Lj9Y3gE0s6YGHvsH2PlDt0t9u3a
j3TXshfPtgQFyw9wk4aY2C5DUSVTzFF5+TTNPLEm0lJWUEvXxHXIc+6IW5p/IohnmuhbwJl37EsL
fX8Aciql70uSIuE/M2Q=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GaiCtiCdun/oCWOc/AYbWVXKz5jVMZoR9/cpxenbwgtAmVX6tux2TILH0PkiB51TnjiFNGEtU8WK
hzHUgctsSXi3mDYQUrtsyNpjE5u0sjtt8dE1QmffopuN70FdnIabefQtbpDzTHPvR+rTOzXRTxjB
P6Xfq8xYYGDOU4+txqCdCReGhBoLp59tmuE2kWvy7k1hqKNx1ecdlVQW4Kh92g92YKEp17DjcR+H
i536gDNXiJL142Ml0k8Cz/3i4vmNqJMCFSYj+q28Qoz55Myw1KoU4Q9cNjqx3JQuc8HZkogw7ly7
tvrxLd94OSq3RWbnrVG+jVGGakHPqltrUPZPxw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aS9RmUXKMVgbNwuNJA1kzu563EUslTeU6qZHSNtwbQkpwhxW8vTETfCUTGUgKJVYveV/uqu1kP7n
05Y85IGpGc4/CSp25q/1kIFzjQQk0KSd6wdrzVtyjCdKaTHVA45PSoGF5+61zFX7fXkKkbTyILlo
zE+HBsaQCWbvpHLyGUM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PVgSjBlXBcPzuRRIGyyVFobuDVzhwU5TMBTET5YQ1gpF7iOr5HThIGplbRtApMTWRURAvQiE1zd/
UE84WBBI0g8tyZPWknk3Ni+mXVmXHZKUVqLPhE1u/MplnWc8KVffihNei77viOFFMtex58OfAU5p
EfEImyym3A9L3aIQ7eb5ckikWjrja7WRGEf+wjmCxltdlK2V+1MXB9deNkgxUCeazzvQ4ef/2m4Q
6npHm7yod7FIY0cVOEXM2IstIfelWKHZT+1UzLjNTCvdMNT+jct6Vwkq0JxparKGquwE1i34grAl
FefY5nWLE6p4uWuH8PbUmPRSrpcqY0OY9OkjSQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13136)
`protect data_block
2BlTJGUITJJGdjl9XuaIzlgXyvNs6GOWcABgrOuk9CLySjZ92SAWOUBTNf2RQgW8A70rUGdkiXyQ
apL9QAdKXz41v8zY2+BJTuxz3dMLLQepYGBPp4AqqnnkIpceV6r4cIY1FvDEB14SfNRfA7Fb/tzD
8z8KqHa/ZpPq2Vn+WGEpP04+gjAxl3e8KlJ0QKPZbjL75xEhr21+qdwJrNAUMtr5a1CUQRikcIjc
lEPd4HtZsA/FdxXsz74GkpDfX3ywXDVfoAGxs5PLP8xdoLUWpfA/UI6ZYhQIrADN0j5WlrFATnk3
3JKsYW85Yn5ep22t0Qj/QaF/Bw6oBXHJ37gOfw3bZbzE9EeZRQnHr9ogTQRksjwv+0dXFTyZh8yc
exhpXPXKpPgrp7DEHaPN2pzy5TFV4u/dKPKMG4ycoZ8XUnCrATVW3pfJmbqZwIww7u7eJ2rGZlg9
4uTyI8700TBhq6g/MP26sgUp0nExxBTuOQ58Mc9dV+4108gPjoNxntGcL5O+WlVm+BLuWEh/7Bns
npclUMrIpLQlYucharTI8e/gd/lPd0MDJRhqiI4X3p5jqXhu031ac9b6olLR0PSbMyuNCdTn3z/j
JWNArqgU6k63SLZU6TEQtaXRPJmdLILWu1VtAWl38JUkkxH28yXHBkFZ4+S7vfGbMRthn1MCp+Wz
iTsJeAgatcDM91Q+QDu5BpIvOeLvCekGnfh7DEtdqNbAwoW7sxY8y9pGlU3myq/qMaOdemp3hYkD
HgVji7ascPT4DCjimBFS96LDxtEgH+P2JmmSjCyg0VIsyl9/EuP1tF8lmrr/uSP/kzaCgsNAHnA/
fED53upXcvz1wIoKcCKWgXh4XhYZ/HnXn6za5JtR7YXA43fkPKoXsXVC0Y77N1hHJrkCYG+xUPZR
BlQ/WGFU8RoI2CROjYsvPG5IZ/GrPzyCKr8zNogQkQF0XFspR+G0hx+jCge4LiytfTIBN45Y0iQX
XHQkt6F53IO/s3SdUv3mbt3FsP0ucKLrilfF3SVOl+7TfJfEzQUTXqC4Md4sC+orvtif2ndsLTyL
lCT0W4cw27Dz/eDm2Ab3v9Z+KMnI6SaYn85VFI6OKPTDTLJkhGdzuotgcJHIoOJIiHfYpqD9nB8m
o8SOvmmo829dhZy59h1XpdoS+jatFtP+FxDCzzzVL3Ac2qIA1iovwpsRjiKPbQ16+wlAXv9WoDJO
UAnMAkW0xpvlZRGq/B0VotFvOa5Nbf861OWz1jKHZtE+pUcDs/RMjEVYDqmi8XmGiCbdSuQ+zfi+
R+XZrqlkBLY3QPgZFMavcsZRxBVdoRsPoqC4LnUJQmSJWatVIQGCAUxoULIVvk3aFPLdxJEI7AOx
UKhHwoV1nOxQ8Meu1OsJsIMqwy7J51zIJ9XOsKSHzXNLTU9LsFWbjt0IkWm7EbOLNpDVu+mKVmUf
+UvHwu9HB8Ikf6CcCyHOJs0n/W6J06P57Q+b9dOiCFdY6r27fbrve6X8+whD1/Bqd2Tl12Prm1oR
o1Ilj7gDbr9yIFF6rpGKYlTtEnN52Hgo7yZGo7VmizkmP4sIOdidLHzRkT39P/w9yRgRlBuH+OVN
dZjttBMPNzckwC+X++05f4qyVaT12WOfjFkL++xubvaS5+A8lbO7K/G39h4HUWb2H6z+7IieQqJy
IJYKsuamB0ItCcqeYDSPp8+y8dABXllZz738E6bnwhcCLFGH+t1mrbQp49VGa2Syib5uDIHAK64I
wx6G9s8iXE0psPiwXenNfAVKLUxkY7AblbMm3AwzBz/bCmNUsCl2KOAL38lpvOauX7/BxnOHg7wh
N9AGsM5DxuPw+xAqrE4Ug3J6D2jdWlfsRXBki03jjDHqRWBjGxE0Xp03Wg4H5lvPsihYPjiZ0j7o
E6L5wMaWVGzGSHApgK4elLkXqIz1hBs50tqNgGCgYnIH7Imcq0vF8/jFh5BN8ocY3Y4byHw/Lo/e
mQI9Ho8JzftAMDchn4ZetaS8653DuYD5+Ltnm0/Vu8etUkhELRzY1W0KPtGgQhvyNIsdyjgMuJu5
atMQBdupW+YS3HGAFkj2PKHUYhfQpy/d9IJEWg7f4b/mGOLRGeZ+TvqxLtXVZ9moJ/LBrQfTUsPe
SrlC3BPsLdljLemLVYdfiBTkP9W1kwC8puuJl5XseUp/aMZfzi/OUbMJXTEdcCjYVQ9rwT/C20GK
iEKrOFi2JXZDRP1x2/4+nYGvAFu8fzbqyR32SeRtTwjjGAWO+C6wKdrAXnorfOUyZFai+aXH/blD
Xq4cfwX+aPnZy8vBp5J6mR0JCKaZ46+0NmfhcI/hI+GGnx0sUTM1FobE2aQjcAljAYVai4t1wwo2
cKnQPX8eyz+pKIDcR4PjqExYGRBK3372fXa1UNMHO6rn9oynUFRg97KMezHGOf6EcaMh8GtLxN61
kBaWXR9nuPx2f1cocLkwLomehR3BmdH8ofIhEeS9lfx44tjn8uNHtJ1JJ4b99i02GA86BIs6Mgs6
7zP+ScB4n+WFSoNgR5bu+o9Yu8JK4FUuRY9R3yyv2d4EWlwUElLa2zY9UDE1oO6YL9QCbmNhhbLB
ud/CD9NQO5fYpz0XQlN/hBeFdOc9Um5GeRQ6mQIgRvvgOpwHAfLWzqdH7LeLmuSh2EtLES20wF3v
ySOz+Qxsw9+z9oC3yjQKckpgB4cnkEImEZdVw5+7wIoOKXgaki57c2N5FLYPlTjoJ+kHlUjS23W4
6f40WtPRwu5r9QPob3oMOhtScfW5pr+1PgCfFtQrQvn0dI/72BdTKdmt4L21Um4jea78lxSqSHTp
vIm6SgXFs5WbeuJg1ZYAQ2ZDGYRdzjnav5Sfoj39FfgfEq6caJwgSuQ3nXGRd9Y78zsaNqzBMNQ5
+uVJUSPqymUr+AHCBdCwJ2CWdf+rf7j4DsQTe78bXcfwU+gv8Q7QN98zQKC+f6dnVCqCqNP/01DX
OFZwmoj0oOSkuOiIYhfsOLaSie1nSWo6C5ti18a78pTEVs78DOGUhO1OtUb2qSFFHWRP1SA4WZ70
juYSWXvDthPVgcn8iVKdRwbxm/eUZrxrIc3ZkxVnmuJe5FJr6tdfANt07SXOPkaTjLTYlwa5KfMb
ERFDdOpSm9zDjDC1beAUqHVCjhkDUnxGOUOYLeO2zPQQSJLsr7cZ/QYYE5IVtNM83XneqS27Pb87
aTSX1i1sH53ZHx26se7B6TtjdECiREdxAfOuI8ez9+BPutsuJP1XU6rcV8QRm3PXtX4zkHyf6SO3
tPeXkCO68GMUSpe3VFQL02OR6rTheoBcEOTdQJwTuBzF5IJaJYh+TJ5Fj77HhkIkx9e8juQ5mPfe
eH+W3H2XL+qMm1y2M3IXlcv3MKSdVMUf85lqn/8Uc9KdDH5BOdv0wGPLIpGZLeyjxXPOf0c+ry3t
B7rQ1fj7bZiBVdwF9SsjZZaJISY2x1rnxilGLDRZuJTEhP75VhDoY/PGocCpdRVUtchBuTfOoXMo
a9OlsEJRty3Oz8TqBDMh88J2w/4upCotkixhiaA9XQXGt1appeWXwAlpknkEj1NigP5IcJ8z/juV
SCGbe9KgYGnsikz99kQ5jDbXefSu+ulvCCReUqlL+7z/2hBGcAvbeV1EhhP4ANdMl7QEhT4fSfVj
pihD7L/IGJL2YJ4rShv5JhhxZZKRSUjJ60hVfWfz/XNCehPCLwqCY+NBwWModAsUxu22WkwDkpvw
6/FDEmGfeUtnw0Ie+VbYPW68Qzvf834Tpq2A94pkiHVkTxodGG785kLyl49/SWfhNfXVsiZuCscA
BOX1R+fOMnx0Qii95kQxEFerkiiu2hVbBcCSYZ/14FG/71MD2ZvsreerMNxwL7Z3fzTW85eaIzgN
5Qc0gIL1yzVC2WtAzTaUlwZfsGmD+q/qHF81o9ytqpiHidEAMpmWVy5+n++JMojF8UonKVRw1kJx
j4UvCj113JgSIfSj33oR9n0+ddNdM37GqWA15u2ts85SS3MFAIepqp9SInCrzofYQeJ3umtWBoID
Z2ZNbkY+qRbAhkONmO8ctfvBUoGqzNnyEdTy3dQNq69QiRO8IZbjLDiDSfu454Y4d3O5o5+RoJGo
2Ql32HPp0LEC0MxaXNRE/qh22KVvRxk+LRRmhU43yPsVf26xGXnvZjGP88Q4cdMOW2a842WnKQNW
D89SwhlwunZGvVPEF5ieKQ1D9vthkkOOwJecnaGqm5vDW+m+w0Dww2GA7HtJUX54EuebqDugGtAd
/sPhOEAXPaQwCq6s7GvKg/d99+0JmJXHL4WurZnNbhF2O6FjLoiRxpb3bS8XhaDS0NdUuy3CuHOk
NVuVotcpbnNGt24kPl9ZkB531YdNbLqBKd3BQAo74ZEOMUFygxl05/kc3PBKEnV/4FoMtCYZ1rrK
8wKOTupa2lgVNG/W8cbicZIpKtA1yfEhhkLRkgW54p3KUSKddzH3zu6FjR9h/b8q4UOcasfwYwOu
mluvjO82h1jH0ZDDyPAffmzr7RAVQbHkXS42fdl3LmuhBygvqjD98JJQQ8GSLELFxk7f5glRvlpi
phHQHXTMZYO/CHxCnVJZXI6YJ324eqbMP+JK9sbUVx2GHvHG4UVtq95yBJevw7SuJhgMrwaMsal/
fFxw4+Zi6gsqyfD8WyUzCo7/mqlwfs22urvBVYR8I/tqHvmPtac+c2hEiH53K1AyxVaH/kMqDStF
vPB5vzCXB7ziBi6sXnVnh7QZI6FWglFP1PwMPYOep1kxeH//LorbeGMq1ZWTRj02qq1HAu2SPYDn
OUnhGJYPYyldKeplbPG71OEyTlkMF0DGxpeC6lWZ149b4lPdEJQloxq4RKbRtRueHygZHLDjjC4U
ZcC5mlXYEbyvYSLJ6mQi+r1VaD41gBMLy3SVeZ7BbG+iMnI7jtC+f+95xVrtS8vqwf8Ha0ZNq5ZR
rEIphWJzxpqIsvKOzpwgJOkjs7Thsm5UCyvv/2wJHxG95Cp3QWMTO0hyjhT6b8V0IUJeafWZxrN6
3Up5oMYD7ToyZ7Ec7XqFMNlQy50CULa/6W/sbk5u+A40eNOs/cxbQlEAH1XXS0F7RXa7k9Hrm1ts
h9fqKPCPR3aIxK3oRIyGKT3qpdJZXQ2QKMWHznABe1mc5aYt4z6v0CPArTq3p1ctgYwFr2Upo3Vl
xfFvhc0JXRvEgAwpH/I+xVpw90Ed3QjoGrkOuxNkR1oq55lvOBT1AB9lI6PgKrpojZbh/KlbTBlz
nLiLIn8ihgC7NDRV9JjIvFcVI2yDQZCUFNw1eYz4e1cn6kgpJwiXbERD/h4GdekKFLudnxroVK3E
/qmY/mdqIq8dS+T1VaE2eXGN0DzPZIc5X91jBn3LfKxLButVoR0aPEQFCQpMgz3soQZgRtrh+eRU
xoxNjeo2YbPbLLCODZAr5zUpePq5h7xR8uJDN68tBbcmpHDiF99H1PBVaFPbPeyl/MAK3l3+F2ib
+WG/ybx0Fug2Zgmp1+Ob7IHTTqm0SWmRdcKjyw7pEXpyhArgU6LdL1jL7S6JDOqdrKj6YLKeU1ip
TosUMVUS3yq99feVLlNfb24cDEuq44mgBy5dQNf8VY0Oid22HclivOkKeRz0UEGeEfHWfL3XFIDu
PQKkbJJmVqo6sMMPiR1O9illHw5x22DOaTsebbpq0lbisxt5BrDvZ8SqOpnVEWAAb47VmHdsfj9J
zzD8OayfeR9NVuhqHUaFAFuXmDxbzRW8DRpYsXghJ3kmyDFv67lDVqDBL/OkGHbmU9uxTjAE3154
TgHL/nfnle9pvsg3kFu8pKomQFZxdaeh/orQWPqk1WZha2HmFgz1tTslN2HUEMachd0+BBXZg18R
rpsgE8oay70my5omXZ9rKh8SnQLMrXffZxUQCfN+xSpW6vycqdK4kGZLmMmyFkhf6vnXmwNnJYie
hZq4Z+hnrgiSgAd6w7VSMcXaa08izoPNUoFCEuEzSBkKX2Awlt45jnSboK7oFakwaSYSsO++Lash
Y9wBfnA/Ss2VPtYPeum22jGc97hVN9lXf+PW5fyAzQmaa/VgGElkHosSWL3lzXLSA6kY8ftjz+7j
a8WCftKjsrrN1OGPyn/ftESDUy7P3ma3YZrmLSVVHiCTNzug1DsdShLv/jYR6OmKJZqY9Y8uNyi3
AJum8dWzBsoKixG/17YVLHh6Vurbd9YuDM/QI6BU8SrPgfc7dHHC8PjpkwU+ma8XvmfF13ITRQ51
vztm8a6R+CtgEy4/wCzf0bFb8Yog/YKL6p6N7cCQ0KyBaFp0SY3UWtvTh7e0f3VoZB7/JNqNTiE+
7WuoI/ydJlFHReY4w+6lQncaUkfo3v86QZhvoKVPkrxvcIp4KZCrufu95ohXK+Vbon7QKKTSiF/R
dMTOxvySKZohlRWNkFKRMSAdkTqtfMvEpMacBYSNACX+jyCYoj45Aj6u5tmEPVWrOVgdvenPBkem
Zy/i0qxzcGXAaMuVz6qNyfMVhXGRjr+iNNWXmnVg6Vp4otvCm3yIu8QU3p4S0SqyT+9CT8AVqhmb
8+WqRKWKuLyWfBgWsJAH+oh7NKOp2dopYWQFHnZv6Uq1HBqC2UoKzU/Rb4ZeFtnO9bIp+ZzmH1Sb
HgwxEU1r3f3wtLdVPsMkzGP3xw4lsEJHIMUTLEEGqxIT088jdhzbeRya+WxG1BhnFJaORTjDtFTS
R5JVBUbrrYakidT+o8eXOeEJypaN9HeAeAn0jOSZWt8abRpmfYZT0Qx9HcHm4DW1s92CfMkZh6o8
WrZpjBK9/WmDrBGlCqIl4fKJZkXAKgjDn27EA0ZMPSNeu5NEYhbE9tM3Z6dhgcxgOlBhIxAiT7Jj
yWP+2tgEkLzUQHNjAWOK7Yngwt3KkFWA2oE72lm4FA5OGpQPN8eRSEtKkzt1hhxgi8z3RshsyGLw
sK7lDGxuL9V2yaBbdQZeATWya+AgNk97XR3lWUM5OQjgZQJLl2khwR62bdFoaUsjM8hzMx7GucOB
S06Mt8o4T6nwm1ZrGWfWKvihJcv32aZIuhLaJ3wHfhUAxu/COwIJU3OW6teXjonDMJK0uNNUrJWm
P7er/UQEYqW0hU5ASOEG3nSq2PeB2KU4JttOUQ2KwL4hRmXuXaGXe0dLuCxKJqhhb+60EpyGvVya
Usp6Ih5ctD4wdyr4cg4UfGfPZf9fcGugV86rTycEFl5G56eaw7GVarBPOUI7uD8K7dSYo9XKQWtC
DaFTQKcAj2/MDVBiUZl4BhoGhhtVCe6APwUIQrNy2/J1z65GCaD34CVYcwXry2MtVubt/y2UDtsA
t0mnW+8pqWRxmKUQHIHuUhW8skEnlUIBe6rB55BNknkVx/1AaVWGHF8kZbAJqhnz+gjivoRvMcTt
4I3+99qd2uDbD8UVQR1TOxRdeuOC3NcAcgoX4PyTAqng3wASZljb8Ybgs3Zqzpx9kFlC3Tf2fFhR
/nhJ1EfppIQAU7Wg7QJQrwWl5/yK5IAJOtQKPSWtgRIb4o8pHEjGBh5RLpcVoEKcSMigwkhr/Vyv
5ukEMydIagjNfUgdfwE49FwhX7CWJPdacraj2wKotSpEIJl9fVjJcpVvtB8vx+w4X9vZAuITrFxb
KcSVCnEYmKG/W6xMwn+LbSTsLt/JeOYvAbWuuz27xvSBbtxMCGe0Z+Ye/T2oAJnnQzQMfwQxbyJ0
VQteEdGi661KZFO7kYozpvX0PRgoceIP1R818JlyXi/qeidJrZ8E9wYmP5LqsT9DDbS3Bzn6A4oj
yRIOGj6GlWZsEyLVddVfOav6i6jIARONne9fqcwl4wXlzE5ELrvU94byFBrGeQVq7UNIIendReqw
jXwUqHeLt6Ghpu3i9/UL7wTnxdrig7WHD621aWqrw+rF9prXQEKPJv3n4AXaUvCCY+OdjuCb84Ru
PiPygvTYomEWTMETwKKFBsUA/PmZhTMjWwPPxGNi4zWPlkOKyvnwVG9Qy1SkcGpXjsEpKpLBoVD+
+Bp2oozJLBxc203QPG2KjDyuEi7M25M/qgiRAsx6P/E2eWcbC+VjNekIQDwI1MFWh+g8DJPUIiIz
CeFZWlgn+rBHcZxOY0VxTrjIAZFu2O19Pemo+U2iAKaHRuuIWnXimWI2hZd72pzROOfzVBh/Jjw3
69KPSiOcvZxm07l710gaGtF/gT2B3C4feUuoO9saHa7l06oOehapeI2e258rLtbD/SYRhmsYXKRT
/2iahhM3oiK3V91oPE+EMA7b5/g3nl9eMv1RfwTutWjWGlCZDrLh+uMspRTGfb8BsLhBZ2f7MBsF
dnSPaAIQythNAdrvObhJWBufB1GlckTVaHACpohV8nkB9u2J1qpcnuUmn+Vs0kBpmXHG7DHei3Eg
WiJ57Epu/zRc17AMFnpoN7N/zFLPRk46m3KglcQXSIx/GrZF7r9gdOZq4SYgrddfesGwz99NKyAz
2AKy+pe9It33nEHkPjINfysIrVdCfOFTojcvQtBZBHxVtYnKX7jmHC1srls1KlQge9iGWxEoFu1h
+bAl4qgycAUGJr5sNguLciEGCiMpnd7PS68HueJ79WEkgO8VJg3ts0SLNyroF/WMUX1IX0LkWgQY
+U7ZV5SsQPWwHDDChWGR7zYE3u9NpkKnP+UOYVtAuk0aiTPOt+E89EOXGa2N+5/psCUtNoouvAUu
ycri736EzqUUrMtSjnckJKPMjLCR0Kgf10GpsllbwoCFOMox39vDVyLV5K/GDEHhbRN6B64V1NG1
iO7clwKp0+WLR7eEHiT+x6oSBNNiRBK/5aXMs0ts18vpN5Rr8AhzniALRQ8OtVkqJ7T/ln+gUPGM
+XSPXrZiYhZRHY6jY8tPfgKdxONM8p0pmVozX5+I+aLfqD3kGNKgldPKCAhpYsBp1QnYtPdDwqZw
T6Pm56d7PlnW3AoHegabxdRChvNK/UgQUvQXZdG0sfTsqucf0XC904TEDCI76DE1+3qqzj31XPhE
xz24p4EjD7kKKw0uHmfMlQ/apVYwi5EFKXS/5faQulo+qeVareTdp1QolBmLTM4pElosDSu5o97x
MMqCxJMoE8qKjfegGLnjBaHFjoZI2jJXupN6QxLb+JycmfIOZ9Aq7eeeMoXeHTuseUxVJDXiMA5I
WUk1Tz+TkSc8hWVQXuRFBjKv3Ui10Xww1H7LyGBOAnPwTI3eAVz0/aNE/OOwHtDUua0IkAhk1EVw
bOzBK/kO9/SHTbL5aG0KsU2ye6B7Rw0EMSFhRpv9jWmma+kQqCeRgQHzRSrJcqNnqRTa1PPX4L1X
7OoAS0SDyDNeyEoREvVJdAWteb2A8zmUi6j9BfpjVUt7jj3AFfAlQgTFtbvnN1ikYhLuWUtwR/O0
obKMVlEKtGKrHF+5ikQ5TGQ+8oKtOWpQdDucqagBvme5j649fhgjLhQNrFNaKavsIvZjUFf9VQIu
JPUuW0fb7IVeftxXltBSlHvuLmcd2h5qxxoHv1DuyWxsgRoh11nq8JZ/5Zc9PHxCFoNc4MqBBZ9S
qHPB+ub/eeSBWRPn28K5WbTIc3o9SDopIRtktqadJyUFF7Rt1Fpt+ricwx0MWVe3dO7UCsZ/JrcK
zA0hdj+upyaP4Rdc0Fdrxcvf9Koz0e/zV2gSFfiQthJelEXb07YIQfQvSBqkwsvh8l2w1mCLQZIU
ZpX3n34PF8sCVDrXW8hkEj2EDci1TBOR/krAwLyR/gEMJWzmVXtIhXg9hWxZHo84E07IM+ZZW7wb
V+OFtTxYppto4U8kbdl3K72YzAhSWaOBJFHpsAMqjKh3zPc0tBC+Aw3joIB+w2kg8gR+5XrGU2RU
j7Av8OTLYmlaLBwmzYQCmJARLjcTpqzwyzqO2pi2oAn2tQw0FttMNGsAQzGE6UORD/viYXYF7dBO
VH6WVodU7wNsuqENiVnqWbQgtIb8j4JXGcVpKXDUQe2zq3L8jrFyP5SjeQGKVOeup/QdSaBXlcWG
5T1Wea0ULKuNKMWVQsjY0N8aExHH33tL/Xn+omd0y39T/pG/n14YTRkVjAIOWm/l2d385zbknWoQ
CMP36jGLZGrtE7RUrUzdY9aS8VjYKaw+ehuibc9gAjetkd4c3U4BoTQApVIKaY44cPpC+ysIU3v1
7sFWSRLDmb0N5x8BN6mdY3rPbZv26J1PRqA7QDqqjZaQ3qxZ1hOWzRO0spL+TSR86HYp8ajVdnwY
ddRj2kyV9BXWoO1qW6dWOou42gODly0qhDi8s1rVeT31n5GWPO3YtYfuXEi0YTMsphLzZBLn74un
DbOp3VWa7e0Xv98h8eqgEktL79101sfk31BdPr2GNaPa7Ae5XtEELng3H+uVcJywi53Ibgyqft6o
ZSxkkfacGr7Gwvmnv+cYecdfJUNtXmVpkxzENgU43D/9lBoVvec989OPCIDfz/ahGkRuWhJqlP44
6wYrbQ1s2d2Oga+ppKilmxzrlwoSP5B/3l7QVTfi/xOp5SWWqSp8zisz2eIJp5MlsVH9PJc4Fll7
zuMZBJeP5tF/Px30BpxZa5tc2v7yEisjFjaybylGuNjMeOXETMt6HWrjFNOERXU5VTB/tvOib/ac
W6U6L6AxbXL/V52PY+AZjJUKlGkPbFQErqUDO1GOSsudiaIDwC3xqyzKhd2rZ5CU6ytCQTolSeS3
Xpyu5He+tMaD7TLM8Ov4JN+ySWmy5c3c/BidNe2dSBzlRmgN4vM2KeosU85Vvl+CV9bQupFJt2M1
SrggCovtfRA1vKghqChDTaOvwJFmc347Ae4SV+WFyC0J3Uircgzyfd+6QmDDMzZ3A74tYaCcZr3g
giDacAdRwoGMG3ua/YO02wnb25kwRo/21Ybzp2dDsqFhUNfhPLTetEZvnht3cDMR//tjlpvcSxND
7toDYOEOPMz/tN1FZQlE9QKHDePXwQMgeZ/Y5tkWcnhpvJ/6vI28oU1mmgL81R1dkhVPS8//rXZU
9qhHJZk/uo1SzpmULlIbOzE2YW1GgMeUbvqFU7KpkRBSoZyOC6c827JEy5XHiWInkVdObGF1wJm+
cbV1gBnrgSp8CO35l2zU6XSE5h77qBThmk8iEmWydCXpJzee9MNCN0DiOkAGfNbx39zgBi5+kwbn
4wshv45nNRufOQLRCedBN4gsZ53S5NaawB3u8e6x7T4qi7XDJN/mlj80QLgpUDsD9rvrneZMeaHm
4ObVaJUKTADYG1hhxnORMN+tobW8kX299Cm/2TxQmLaKSV5cMhKPJKKqNOrXzwjs1+/NB011DyaN
HaoOG8yH9IHITLMok9/3yreqUDh+9/STmtoCwMwSxCAoRngHPg6Fs7fkC4DXQbpmsNZrSEfKcPb8
KfD4fmuRNxJG54LhoDqJVK9JyqFyIKx9w/whnvCdLW9gma91f0LeRhrHAPZDmi3ethiytZK9XImw
Eur1yrx7XxIb5OttuoDMLVi5Z0ehV7+qBHnOTREMDG2cKSUg9SYXMQVeQHrLPbqzQkA668TZTUkJ
EsjAmHItTJH60Y0l7wExJm1ABo0KwUJOktZm7RgpQ+QnEbh1qe2P1j59t06VewdGqQtMkU/hgcOB
iEo9EToPg75P4d3GSmbquuzzbmRyCNQRXo9tYQHopPP5lGlfvM2n9AcN3BWwDQmu7xI/dQxWJSDO
RBjO2/9e8xPoeK6rB22iYKyZe/a8pePEP02uzxM2xn8nyC3l1WXTy76m/dsXMLUZ/kEBmeHGj5P3
WX1hrFT1PeUcarbMKlhN4cQetrkGGRaLlqVeVGV5BsPvokn0v/wKBr3SlYehcyaCfoPe/UZQstCS
Z3vMyFbOjejBRnOVozjEJCkNVtWaWadYX25ShsjbXNEPqsnLUUAIDIdSeW4snFshpyzpn0HRI3MG
61PXxdIS+pQdDxqXutmdI9DfwX8rMpBawrywKPv1yl0rIgtdtWj1V+5KdwKVhNktnMkkER3cn1pp
epxgv+e+ttKHULxSLbaU2hmqcNyyOseB4N0FfZkUVNoAbwyS/UxKGnRj0lSPasNaPR8eniPAZlTZ
ZTetYsCpJGCFdI8xN5X9U0pmhR6Ze24mfl9UUDaDZiLgwuggNyYd6q8POHXmzeNUr19Jv6294/G1
+Ec5KyNPKSyqUt1D0HExczT29ZJOuVJkMt+wvafjJ60kxnSI9La0pDAdgMxZfxIvWe0zOAOa63Wg
4Ycl2g/I38LSgt82+imkjCQjwWCTywBbllVCIl4z/UbTArrEQGJJgPqI/NzqdJRX0X9JMhmbxfua
TsnXzm2RALzDS63V446oEiauI1aj9xRFLh4Y6FiAzBOflxNQtiRHM2WcwwJfFfF8xeSh0ifjkKkE
0cn/iQimJnBz5y7VRlgev2+zQ4XECEb98reAFFNMfLXbgOlPKdMVB/EcgYzxunSqUxQZefXAV9hw
Fkr8kRc/EIb1H49HZRouJlrHukOLNqL/L7wfiiHhHkG4Aks9G5pyd8j88mAt3o9fy9C2aXFiRthj
5xj6kMoYtbzNyOyX/FmeKYSemF8LZIV4t/9NoGCG6qQL5wZ0NguHnsGgRcZgG/fi6HKNYoTvXJeN
otbIUdlMUwBHaMH//AaDyEERMbgoBEAGTgbCKhW8QiSit9NhEtt6SAuWnLtORnvfV/r8ZK2cRGke
D77W5JjBYojrxqsbQVNm+jrdmNTMQFlBgPYth/FmZO1QPPWO/MJtmXzyFftYsO2YbQZWk3GeA4Yx
QoXrhnfZWYGiat3CPSqv88rz6iL4Z8q6ADonn3n+5WjGuibtr021BCYsX/mrxq9MPb5jkEqSOGZN
2y9exn/BRQcTzp8wlFs7Z/04rl+R+XIn5D+k1vN+jU0PelyL7wn2wItWJA6Khg5nICBN1glA8CJV
ru/xOwxM72L/icck87YwopgBQOvwndC4KebRBcdfdXTJ9cdOxtMtjc8EJGMHBxgGi5WAJggjkA9S
VHUyTJHl9kKujI/vOKvMoEQaxcSQNS+HZoILQx8WH5OBY2I7XF2Zl2Ywayc1eWsmSVxRpmS4rjcR
tG6STIXJ03l3JrygSBQqX9vEkxbhyux2LP+2Ao53xqB6VBBbMqA9ziNeZOhC+AKdhASlxO7i9TQn
3tdRywPC83DAKzxOXsdKxDOhjKL/MzZUxlZtzdDtZLMzIjZKci+jSTk1R7DI/nf+sv6YV/RBwWaG
SqjSGyNkeuJsBFaVjiNsNL/wQUjxwxn/s8SzHh3cE7uAra6CTAV06SixPEwhg8gjBiUecapvMq0k
lV4G8ly7Kov2eTj8J+k+HmAJGtAnzdj0sHpFUHgcNpiSzpm0u/B4tFopK1XQEbkY37Rd9wrfGlFb
3SygG+qMCoFJ32mNOEpsShxVuOXrLeF/ZEn1x7uxv/4sxbZxv1vY79QJYWdW0PSuSuncbg/DA7sq
JkNXxARtJ5/bGmWJxuNSfapy0PsZlB3VC9XDnAoMqycolJ/KF/AL+HUR6J9Y5JqNmJwSbViGgBGR
FZG3MP0eIxRZIT6ScjxbDPCfEUd+vDR6UTZMYQCw9cbkjkKJEgtJB0HkeV+MjlKVqA7YaR71+/tW
013hnKAvrAUcB57iQapF4+0ULKMrBzSFMWzJeeYys31y2qX0ctVa2jTjCx4kvwirQ6CXhODJJLk9
ewXwHJptP3iH4XYq9u3EHZ1IZ10wA/FpX+4nUdlE99+Cuz2YzcL+jcnMtFfYq5NlQVfWogTVq6HV
IYx5QoyQGEuCGydO5t8YVOoPhrgK7z8HQ7CQDqIX6NhN+fau+B9fE5Tye3lcmaCDEA/YE42KCy7e
/nt1WcyNCwNKtC6ii2NJgKb/UaeoP975nxz2MCjvnTwtaDOZFegw2yz/55pG20wDSCMqgoWuYA/W
LcHBR8lzURyC5XWkL3K3Eq827Z5m2b16WvddlrUDWWYvv5BLKc2cFY2PlmZPbL7u3Uo7bODSaS0v
a5T5YjV+thTdogfKSrZmWZjhJ+m91YVRf+8jUddsyNQvZGbQ1rFm5H3x7ke1ten+/fMxTrMGgAOL
HnCbHcpzu2eC2ExOoPsqQ+OPZ127WH31vFS0amGRDsM9zbEYTlX1QdsNrazPrjWYHBuyiXvM0t8A
Xw2F847aLgq/WfXSZlEEaBVJgH001KM0Z5Ep9o64S99ppnH5yHY0aWiCLodRZ6CHvCFGhxb0W1IQ
DWTsR9QRBR+mmSEE14Ppn1pfotFWsL7VOPiJ6R7LAF9JBHk3kj+Ri1g5CJ+ULPGCzfSnv42IsKZn
DaAIptU2e744uEwj5z2bQEkGmHgSpvJHFnmxqxd7tQBOoi5boadJ3zoe5qfuuhYipKWScn+wkJXn
1MEMTDXu4yMkVU9ya+TLsYrcS6Ne3I/eNV0K6kW2Obw8eDNdfF5nW8SePmfnjH7A4PMfr/if4r0t
jRZJoKhqvgvGB9jt09r1gNmTsZ2GfwPZO9ix2i0YCcBFVT/nx7JfW+Ch+syKDBOF/t06Au+hi1Cl
fkG0mS7P9ct0t9Y+xIGa8tCKJfKpyeosGu+5CiyNQsEXsltmTB9dRNa+5ys+RZEWp44QruUJd9ow
yiTeby1VH5eql6ROdA3yuwrHSb7GD9esGkau8DizzFSC9Uc2nQafzGYd0YO7HeobBV2W0DGJwt/c
CKoLrAyFZreXDVUNXDmF66rk8B5zOTs3/mD41mqGxzz3FN/vKqn6hzRoO8cFKHgR4MIu5H1jF02H
dRBwvXsdliHx2USNMteDMriKmqnY/OtBCu5aFeBwwevVGmdr+FnzgUAqq7tiIJc3AerTzKZr14Ai
rCi64Z08+0VFLT42P01yWKbhzFTlS2uuJnGyxhXMSwsLGP/NptPKgZ5Q2tqhi61xgmlkcQ/9AQ3t
nLoXlKuqqsSzPVaLCmZL79+dDffnQ7FscwnOOhwx/LveaerMhChG4STTpGu/rh5Qn4lMkU+kF5Zk
K/ExR5Mqy9XKtPQHLAOOYhsAb2Oe2229R/cxvNyrpAP385rcPdF+STMvWy779qodzHFTeL35OQ/R
Tsu6SOp3qGEYzbRTKQcV7TSyWbk9TDLI761bmkIOrFYStgPzDJnJ9zJmUIYoAO6EnYpb3v9mKKj+
JO2tkMHWDDsfgWtQvT3fsvzHOYoOlEv4/yYbrw4//LgnQbSqa8O8zvSr7fpklCMo0TZ5Z/XAGXwx
m8HpNlFQ97sqWYapDxM+8u/VAXHGyok1L2OaJL/VuFn40GicZlwPgndlSMciHh6cHMHl5tczzvrU
rTyukf6ab6lp6T9eZcct1O2KYy920ba0PTT/vzNo+ipWuREfmZsE+oKjH4Kv/VeA/hokUxJYGKtl
PX4YHGdxKbJsi8h1EIaRRwbkgRtw8NWLkHMbocAMWHvVkczf7g7Vu/ZN3R/OSfZfaV2RO6+7vFWl
aY8Jp9rJO89n7FV+oPLvC0NbNA9DRqhmKlCrY8pXo07XlnHU2+LkFOlxHNdIpaqlZ7aIhUpSoh0N
V2hF+SHauxWl97t0QS4fSuJ5C/p8BpdUz4YLK8eFJsNT4svbQsWCgxItEjRBVdoMo5RE+AbrlAfV
TRLdoi7PU/Ovw6HL3kYPb52odZ4HcJ0pKsA+WH8f/hJyVLHRkCS/kQQs5d133rj6ul1kJPDmkCbI
EKKNHF5t6NYHx6dAzV4e649MKJ54Mg6G21QQXMGCg1dWVoINrKBavrl1p7Vw/AkIVkTta8aYsUdf
EWjHDxmx4Zd6WqpttWNfei9jkqirTvGqLL6/q+aUc9agwTa9pCsuxFZDm8lX2hgT4OmKDt2dKm3j
CaYzohOGAFch2Rd7av5gZetg9Xp1k8HTXpLd9Zajfuy3LCh7q/SQvTZq0IbD5uNCgzCJ5bQ+SpM4
ko7q7Y2KalU104Gmkz2wdrVaSUxAOPwaTEWoWylZ6Y0FmNHibdwCvWkOP9e/kBQyJ5MRMzoABapg
91Vnx4a2j1eYnIUMkihI0y8qxgl9/6/++yohlXu7k0kvTRCShfWIX3PxkQHKzwFjuH45+/pXG41/
st/VLMGjtQUzxdfesXm2NFxjgWHLLvpawbDB2CturIzlh0GzgQsvh6HS/2CCkOH5vaiNdIlk5BQb
XpHLeJsgVa9TLkcgUH9GRNszG1j5NVwsnxl45FEdostx7+T+IO0nFocTJxXwrCfSbpviIEB2O52h
hU6irKOnnDOcwgRwDyqQ4DLZVp+byqgUlsppLccK1e/M9dZLEEXus0P1G08FHB3tAM8x5ye5oqnt
QUiHUGioDX56Nl/I1LIUMUt+iAdVf2pufef9ZLKEv4jdPn0jxDfPL50vEAB7qr4JFooVzpAYq9np
EdIAa4zA84gzdXpXWsUDV7bxjw+lhWtcS5C90UjRbw4bVczfXSpKextMvKnDBopy/eNcKQIgkbjd
1V7Z1kzHYrwsJ4WgOjdJ3Oq41+0c6gRrrbCq/g1+NV7l3xD+H/0Y+spT86NEIUYeRxHDL4qwGXTd
VQZ5sLtJTM7AK4xR/y/WfNn0n/R8fEqf3g4ZiaG94rkcg8yl0QmMSa9MfTouoDHNcf7iNlx2bAK+
ALICBggrTgzy1xPKHx+2i3gYBgv64Drd2r+X3V6FjHkkVNo/NJtNVeSYqcAnc/zeMZF4x0gGJo6T
XA7qzdPr1eFB7gWraBPrIG52URKHYABozW6LWB9bNQkzyPbLlggLkTugGpikkL68oZ1eIag/ztXj
/t6GEdcXDeF/nInvZiA43gzX86vVsBZDAUyA8FN7gOBgTohGZ2yFk5MooKiDkVI0tzg8vtLSriGp
lng1j/jCKmYD4ULYISX4BAAAW3PWzwaXbAQnpPGcYfr1eZmzphgsd29otJDIaOOOngrUBN1HZYoj
VOCT79IaFzYtUDolo04Wjnph1mHjNceRvXr9EO2lcyUmD/bycqcDv3Yc2ykykjW7qSlgc28aFdH1
BXjwFX3y2Ty1V3s6MgGPntKowAXUYPNqymIY6a0pmnSfJGs0mq3aczWBButJcUn1y/hfLrVhvl5I
UhyrAlMvZUsBV4Lzzdxkl8rsYm1zjC8thOPH3tG1pMAlv4zrwRnibfN6/KhpwlgpRgR+Qex3Z2Ut
y3la8z6YNei6eVTHq1y+FQGZ+9680nlZMHHbMvlWmlASMx/IyZl2OTB+uifyzjw7zvONO3VcU84r
H8TGlTYq+zgGz5en5KU7QVu4WyQhd7Cj+TlQBD+TnLh/w0PVWTCwRTa9o+ghHRLgQXK5syLEHsC2
19vn9bsaisU4z0ep3KWdDpNPrENYy9YxBpfO3vBGugMB5wZkzNa1aBWMjTKbHYof1/yLAymy0OxW
2/l+3Fjqjb0x63Sco673CU7vIscfyDpN9nFVVVBK9CqUTus4AIgvI5xx5YTw+LJaG9D33rkcrtAd
4Spvh5jXCNV5jJEzzxlPWfZvHCpoX6LpEB6dATNR+dE8VwcLHfWbM+cfJOrAyj4sR7XA5UstdBTA
hyT/mtSlXy+QH/ULNdZ0KOleiCxLYD+1uNGtXet97viS/E/POLhHdbM+lGEsE5xQzSvJDm3WQkDG
feAVuR7/GyJGKd8rdKFwwQYmV7x4J+udyDA=
`protect end_protected
