`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qelseV9d9bvHFTy6uG8Zr39y9uQxWlI4JPFDoIaZTsOSmuoHUMlfxtFbaz+in8/5Scrsi0DrHBRn
LkmnIzgBqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kX+rrFLwhozg1satUIQSPSrPDSOrawuFzyf8cDK2aRnz+nfy9rSTbCGWDjg0hoH4RBAgh7nAGZJv
3fOzdp3fB0BOjI5yR5dmsnKboOLvYMYN9HnrEcHHojQtDHqmp3xtFTOKGx0+XQHqa4OwBSOa39Gk
ttHGg9GGFyvcexgWpD8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GgbpjC9JZfbNDjqQddfymGpuPmqUYexIsynBwQYI8BxA11wZnEZhfbfOYKhxMYuZhDI+4kU8HAfw
OS8f3OE5XzpHBgwi04LhRji3bfjjc0UGQgD6nbXRU8IJwgyLG2+L3YgtZyRj3iUWQudTU025yIl/
w/D2amtnp26a39pdv+JDxb5P62KZ2QmuPLFS49iLTzhyXc6A1UVcuQi6+/KeK4kwq7WI9gzHj+K2
0CU/pJTaZhbO8/HCz//o5jQKEKAtOt/5mJJNJWNb6C+2iKvWgg60+i66+/M2hBBNsEFKB0IFyFqX
4xZvZsvXY9Ibz5XlItdoi8orKLWLN62+kJg4ow==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jGf+oBAdHY3Ic7TX3YH5dPR3KFjRPDo4rNWLmrocaNy1FRZr06bL3K1MdqX0cY0hy4/CaYtm9L5r
O012ySqM6vsnbH6J+RVeFNLfRpEimyU85GamecyG0zpZwjxSffR7T7kk4p50HiTlldYwxnfJgRkD
vMOxhPf/j0exM9ajTz4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
efi2QMOx4uEHWRasjm/nyel3NIfbyVaS49xTM4bl2LzqJlH0OcLTSFNi+J4xKo5nrE6h+o1SVExX
04DmeyRrCGZKiZANccjEp9codC0by1sZB9jiWk3Z7YUcgGxR0lBPuDY8CG/NaotP8d79lKagCgSO
oQYwh8oxHeUgKbTXWj1j/rSYHUXWYBwad/V3ChtzdMN2cBlTcz2/OLvbnbtQCv2YFyLsLkiyRWJP
JsXSQ+2EOZfb5iEPEKiyyZdW4GZWDjuQYnRFczZLZo0KG20TCdwUIeHoxz+kesev6it6DghQiNkw
moY1YwXLDpfM4JYnNas4xJvsboNzHwsSvtzChQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 61648)
`protect data_block
FPO/tscapARTGOtQbudxY6wktqbeTbcIaL51gj6gPG+dzPD/+c0PyeOBySGa8zFEa9AZNT17vS7L
tod52sDKDjExgREwiXaoFn+iXrs/ZGM++6H/XYeIwef9jvCnmHmqvRE7y9p8GGPNWM7ttmPFbkKf
GVeE+9Ll5wE3jxRxsQEnK4bOTFZxd2v0l42c95qSQDYHUJrqja9glr5MdjCas+9nU9ruXhw/4bEr
SaHRqZxEGpNDHJnxaRu2BgTjPa27wzEnyJyyo/XYC6B7BIWCC09ycnEdduSTbMEDFsdC+gmlaR/b
taP/AQ3n1/0S3Wt41CSTDWupX5OoDuE4f8KC+TPCwK1lLQQciI0pdudaDZtXhIQ5iC1prymdtYDE
UqpUfyswcoZ3mzKEnIX6nctD4LfzhVP3kHKBgAlE4oy0F56AV+CCW0Gjsr1qcWReRJMzVH0ZPgJp
nkL5BeLkyy+qny/C7CldOm3Aojho+yYj1nbQYrP7esYGlqGiegFU0ETUbOnlC7ud3ft4S5ugTccW
2H1qJCgxlSM7TNhu3NL+DpW7Hk8+siiNgUZDRnLld0wk1kRMGi2+5wepZr+WLisixfGJziwnjovZ
sTRld2hSvcuDZY8B/y427ayzlaRUar0PNydBCuCh9zgMl31o7qpRvdil59vu3b8Pawm0igJoPsC6
7OLSSDMTwox+uT62Z/BI1hdcON3VY39fZCp+uaIZ71BOJ1VsAhuulu2ZlOE/zHbEjs1nSDVQeo6J
3d0WgS+7e5tlvfYcFE7Cwx3m6ZrjrsH/etBtgWf4dhoIB5seR1URoNPP6i7FV7ll+5GherAHXncD
GJq/sRR0DirbHULwrpVFaH7UH/7I5LGTbtml8raQShbAPVOasmahjm6diouMiPyl1HVae1wfmaZv
TZ2CQRlnp1Bh752jWy3QhzaFfNp4kXR6B4tnKKFY95lEWO7nJ0oflMsBVkj7UG7XtOAut/W6S/oE
dTOCGl9HknZRLLKJmMQTec5Z50R8qe0BAaGP+Z4jtyWp1mF9utJ0F/n28BA3PNfGPik1q2GIKPS0
jOop9zPHjXVwQa28wTxc6Eg90A2Y3Yq8hfEsHZsg6aQgbzzNkxqC2TLi6OV6RfbGdPOUXm34AzLv
mUKuwALX6Qs7VFdUPdrqsPM9C1kaJPywVbYbXLLhyUIdWGGUWIj1Y8PRaHWWDipoJm7+G+LlPus5
HopLKwf22lrk6B8F92iuWBxxAg8rgEJH3tG7DEwbeKY0o08rF2iswanhM9J1SnIAxfGOiDqTSL3t
Qq2iJGqRkOmCS8Ht91639RfrCv7cW1RSKqTIlOEKfE3Ahln9GCNA/R3etxP2rugxYsnkLCaHFSl3
zJLI3/5Kgor/BnE9qwh9HsKWrBNf7ZkAqgC0GT3ZcZo+Lq2NiT5DgZqvRzhvKbh7R9Hi4IAQ/4bN
jHfsLNTeqSl9oQwv7FVqdVV7nOS7vX+5P+EEBZUu0GUT3WqMp6Af5lBsD6YENYAwjU/C5wvJJeIp
EDXFFNHeTYwClLovgZ5a7OqFCSKCFV/yXPwCyBbE8pysqtV137hwd30yShNaI1I0PAPZbxL6jhOh
jKL7RdeR47SsHf7/rQeItEVpezcwbdhZq84Ij/T+b+X9GtdBzI08TWqIJuXrhxl0Qwd1t03gLWFa
Q/xBzcnZRjwd45lrv+6q5C3BlWUErexstt65dtCkTJ0S6M9jwcf3CXMOBrGnix/QW4k/8YY/GRtt
qxifq/rB2eNFeBhtXtrESBHjKNt77xCfJn2NuyplL1fzTXB6Lv/4Q9VE6Sc/7ezkJqJdZR55M9cl
7bNV8m9LQinHLKZ+HNoICFJTBSzZqQ0VUjqwiCbzBUc+UNPKUxtOFu/xxkk8hSOakqnQogFgmgxu
sTooeqcSvFeF0TIGG3HCpxAUjn10KPnAlqbfnp4RGh5nU9cBgyQKBV9v6VQF3lY+Xfp9toqsa5NX
5ycM9DYrDWSTCHTR6qbr+dnnlsERvSYW3xSQ9vEgOabPDge5DV82SJF55d394FOX1zXVUxSVAPLr
EMwWUw4wEGyo+0XmLxY/E/k1iDqqXg6Lgm3XA8TLw9JVqx0N+yVIneXC1C0lXZSU6wPmLcMjomDZ
+JN3ZfYsbIoC2HL7jQ0EiV0wmb9HvtH0ZFWJ9rl6c6sV8IXQhgOA27ll8e3OiOWwxILQdEVYvCdh
cc5IKcRzmT9ieJeVO9zDEfFMdBdZOMFGAWrj5yxfnZSwt7H8JoilWwz2db8sIVGB/2YCSFDZntSm
M3FQzSHmLjoVBjMsSOZwRCagWnrTsoilgy5r1DmTLMhlzzSkdZHdNh0KKwsA31UHBTYW5gYNa8a8
CuzWWWcyhH3sNYcS9FiEwSMOrTJsXBdJNPztk8jOzPQjb5LYtCq2YJLvshtlCUTVAZpzNVygj6Ix
J56cxqqYWTKHfUmDiKOsOwWR3weRu/za7cfhc+B8VNzLSh+2yA++7uCjs3YjNNN/VvJsoX3V+Pb9
mE3IxikkS/FZdTcgmVnWkjsK61oW21vq2JBhejwIKfxirw4TO1NwxkkxDabiqA4w4J8JoqMMpN3s
i0r0szdhHE4kDL0rWNu22cTAFIeaNjZGJoSYHBboiIotV4z522fBbhxhs/0Or13PQillsjONmkwf
HZhCk5WCIoh/A4qtpfnyoeQloNkQQ8Orbk/dUaqeoWVE8tHrJM9Fk/SBkweqZmITwuMZ4UOeIa8U
YZG2TfmtBuINl3DecP1WGE9Lgygh2iPmUxC+QFaPSGvgCYnZ7cBOusdfj1eMzKcQvBtE1HSXBK+8
1UUvJav0hwsFZHaRIVbaSuf2RV//LPsP+scv4+syerbNL13eEzv5K8BNVXbVxkRLqf2CUFRe9BMw
UuiZHL6rhgrLzuIarPn33NWd7n4uKMGz+SfjfAfiqEsxPo5j1Y9x4mkl7ONZk1vzhosswb2SP+r8
sMqq/fQt0fwpk1IJmht6X9RyRy92y610KJKNH9TRdf16vkaKhqC13jE0VvVCea9seL3eevwsz/67
VtzHJrGpm7P4v/bDDWFa5Jza7WlCWH2dFFrkwRrMB4dvN+9xIN37I8O6B441RlDJ7iUxs50UvvLh
Hts5crmaaTyD9jpJZBQgZ6kp2XEcpOWIWx7tbFTDJLhWSB2EbaM41CE/15jpV5IR+Khc0PqphOaF
DZ0j85pfmsqoEF8I0S4dYIsmBK4t6rGHyZ8PE6QfCEmj9KBKsLGXMYUc362vJ1SngWNWj5Do5qmd
+05+6RClUruLnv5HsNHVlXuvvv+iD0YIfG2it1tzwJQAxT6dtRI+FJzRSzozbyM0jUiwTFXx3ne9
Xk/yZUKfEAkBXdqG7s2NWwDja1fyTWZXwJoJRwfCeNsh+6lCy56mR67YXCDYHG5y0FlkkBpa350W
IYOv1giNh8irTTYH/ZdHk5rIqBdtuKuNG48Cjd1hxx/vZ4+w2Ab2Dksgdz7vYVtIh2aCFjgv+LV2
4jYLjBogrn1vEvvHfQ2S+k01YIbFF8vDvCcT7ROutqETAHwhYZikFrybtRaVbGr/xpn/w3gUWP2Z
UhTtUSq3OO0mS1So2LQzsbIj+YkKlFzzIHHf53iUL4fEioKLjiLQJEBcdi+VpdYBRykhD9u5c3PP
a3q/5MnG4qf2p/8KZCZzrlYgMiK9HDqV31BdQaL38QXuXJ/+lYRSDyb3C4Pfub6PchOq7gVK9kKR
Jo5crgeLngDZ/tUwmcPVOsW88+Y9bDXAvhgo+EnFhA92GkNnZsnDARR89bOeusMqMDBRQcBcAv4M
qHenNybdyf6yBzFEkztnyHf/GUPp+Vwl/d3O7nO4CNTUya/oq+yqmVUv0Z2zE6CBScSAhQTyx43W
E6AOfVIyGqQ0i+H0yzD/2WF4tQ7Nk2bcsfIzhWrJuqBIzSYCh7johtETd6mRAMjL0+LMgQsmebPc
iqOAbAxuj/YFsJhBBZVGF5ibRrM2li1tsBXDhROJnSufzKldgr3YZ066vi4zp41E4WfnRNnSlbsg
GSt0BfVlVcCUqbQhkI/VC6sI9uMVZbWaNqObhXwa+r91XTikWgd2HaoaeTv8FT4iur1ZWdWJwcLY
sPZCCQsyrfMxVszkOrOajlPh85EpgIi7KdmUgoimW4OWTcN+wHlkdLPL2YqG3nM0OxrARhDc5lJA
3x4BCpzeaxsbn/At7M2S/d3UnssjHVFDGmI4Kvoo+wijnMZPJT76cRdOBkST918fyLPlGLeNXpYN
A/JK2w1ef2Kyna+/VXnvnQlYR0748yrVdW9t7fYAPJe2uGs6o8c7brxMAnoBQFrbRvSkTxLDGNAK
b96Lf+C0sYE4s/rxr23ZoHU4pk5iB2tO3ct3Mq4+lyADc0m6px6wPYCSr75zA/4jYQH9KlAFP/rn
bXAwla+C/T90Cl9TRCI5L1ZOq7zgZcS8Wh0j0OHESEwSmMn8NXrP6oe3BvmTT+mlAwPsGB6TecPK
7LdAwIf8/eWcR0ak8Zq3dziMpGVPMqu2iuPCZQ1JOcTt1O5WpFQul9tpA/PdlRH8KpRrnYtDXQH/
twDeyvgPaFOAdydz1QcKx6SQu8LxhNr7Ld2ccCWSqo1z0u/Mqq/kvkS63fZgQYMMLjSbOtDunXsJ
gNB7qn5gZLDpN4bxjIrglzuYvVulQzgrxB/Z+6aG9dylYAdx5acnAfEk29UjYJBVT4pGGNzbLoAY
8OqEf9GbBoxYGkHwT/EczbAtf9C8TfEWI0rOrBRRhNm2ETlZtuPgF8vSSiN2Q3GPCZi+ahRC9ujg
Jt4ZxGRFB+kjUeQdR3bQE9lXJMGkRzVxbRuWeYkcpvOYnc19dsjbslqUmVHssUII3/qRR13XsRus
vpCY8LMPCooXkU88vURjhDs0skNLClqTfggU94TOniZVnKbo0cVI21TXDF7Rs6sN+8yFnryXHGb5
YxrRzUBdsBfUdj0KRZylAYXzoiQGLZMntvg26yvUmRaA3G2U9MmHcmQKHZ9UR1p/TpUC+HzUhQIm
fSutlu0Rk8OUJBJ5BPwnbm/8LnPD1nyhlBGyXNNgJkk2SnIkjnbqXjHnEVdRLFyc56FXUmMr3clB
mvUcep1JTnu21++gDVPrvU/Ph5z3BN/e8sKtBmW4oxI+NZU/j2midJ/N/mEh+6RDjZfE09miR0bp
SsOlrYGwW1rdWosmqx3EjiXqM7TyCmv9gxLbFO9+oOWhSDM3KzXlp/kST5haKUDWhx2zPHcneUAW
NtT8oPNbbLn8wMnctc+5bghkyV7kGI+1ekj9ekmnE0/AYkNQFQkWBDSFrKeupxfHJU9nvu2JMvNg
Lydcp7nUe0Gbnie8Fy9bRvad81IjDN4E37V5tgI1f6cazwd+xIDREfSSwWnvIkrOS/DDIZElMwRg
KWQHky9CoVypnAkN22+3RfWOGR8Fz6nXcH3GTRw1sR81QdDaTjpvuVx6lfWYPRRB1Bw4oJUKQ1l5
gzoqqxQHNrPEdAfSWIPLMofdHRUc/DS/NvSoULTFU6ucSDptRM+RMoqRwcWxjtJMYzX3fn458Ajk
P1BF2j2WNlLshWdMVJwy9G0Gn0LTvlpWXREYlBqxvo0HyJJK1mESPRHIKg/7v3OR766nW5Gt8fno
bfvk3mp3bqj//Vj/xsL/2MBZv1hEoT1N+Y+IupUohtaDb25Y7h2cwAPfX92bcYmtnlCitGBhCuOE
KVCxj9ilczznI8yEwbTKxOIyPVwybpzu8MDqoIz0AhLXOUaw3j/refQ9VdpLNyEPJ0Tr8vTf9gEi
htB/QQJUQIDab0MFnVDuDXFtCgCQ97YgAGb1LSZYw1EAkNY/r1jpDT+t0zWmFkwyhhC+OtF2yMDh
Rc9DkKZ0WopcUaRZG+NFTBWG2NF6cyJA/j1VgN2ok2kP+JjzuoUGUjbax+tV841jLhQnOHneKuog
wOs9ZaIQZ1q6SRHg8nHLbc2EuzBbqvmBonMkTw0Frl/Snra76gE1O8C7R+6um1aVx6Wh6uaZ1Nsh
cQTgYx4oixRyNoHmedbzmSAOQ+Wy2bkEyoOY4452Uyc6LLGB9iLFcRLKKaSY34Hv3btWOFlBjMa3
Z+8+qrZvD2jTEfv+M0KKcKkZuESNMPkSyQUGsl/ZwG3NlWhtNUWtNF0vmFpMQIfEQfUbd5p1IYnu
JlEz8kFpq3MDSaUB4RsYtZ42dHS7796U8GkpT0gNgtP74VBwCPyfBXe8cS7vdTEGtc58xQdCf7qm
9AA8ii9X69duSiszKQ+7yonAcmdaqKGrlis+XN+WSpwUI6Sid3jBS3/6pqkArwFANPa7yxSLU9w1
tUPdZ6/lxpiMzHPz+Hz2jH+sOGIN5NNEf086px2vBFbhsLwZZemLQHYAeycosK33T8ZhL3FFuvBt
/hHy9IwlW/0XqSFEnQFIK/jaXO5jQ0cOmXW2ftT3TEmIi8guBx66uthKb2vTOJonNU5XM6G/ZA7X
wghbJZa7p9D9NuzGZOkdFaJQY9TkcH9uyAixiAAgXtbKH0CQca6YZ8Rq62+DJuLbYBii4+kGxgsc
RXlAjRFZWvzoxbenDs8neqEJNfBAF71wNoU4ZzN5jf7zJFnkOOlg36N3hD0UmLToQbVLTg20fkbj
IPB2g1I8JXS9C3FukXWAG9B7PLJl6ephPAmUOP0JQOJDCgn2mxy6cuGkCuTIQrRhedUWV8+yB271
NMOGBLvFnZAZekevGdNx71ePZU/PtiPZWOJospxkDUPEn0aqoEcCbudVXf09HyoZjqXWxUB8dzls
jxE45QmY6VlsV7Uu6mv4krUbnCK9p6Yv0v1XPrs3yrxifuo4Aoiik+MsKiKJ0NNn9slKZAZXQSV2
DjNxW1dcyCzp6RPBXHrt9cHztfvTaIBIYovFxoavZkWByqt62kq5U85EzyIlU506A49FfVTSPaaD
mqR/R+Rrjf5wkxf/9a9WHfLiCvkOIHFL6hncggfbvUxeKaLH1mxerYzz4fc/2i7Y6VaMIYzxXcCS
63yDZqhfTW4iZGmn9+iqq1GrBbT+xRk6e0fMf37dsLlIqPXpaHBlGECqr2cyqYZex88HDyEuZgIX
lG5iSvYUVoO59g0dsC1eU/gmJuS90uRGTKPpUmClDJbnnEMZfybtSevTigI2rrps23s4Zjt+JHvW
OL9A8+cB8WKdhFWaDe9o78bEU4ytdUHMnCIF0W/3ItDIz4KRF4njabxNLI3ZY/OXCCvWFEm1X1GX
jO0GENgqhgFIawBUiSlL/Hulb7AJyVo0aA39qdyfZ4mM5qqqY51JSYDAjaCiBRYb/i8lr0CiZRoM
qt9Lrcvg4Bods1KPtmTaNJYvlNZ2E7vxTKuKHI9fI6g1corwlw+8fnWrm1Tz/n7ik1gWoEK1ffWn
Fg3JYGp2XWMJmvDxrQYYprNjmZ2kZacT2+Z5y74HdRLPJx6e6xbkSLHoMmPOf8MjLfZuIRMX9J97
oVjAVbX1/dXut7LN8JmZqULPN9Nxxm0LGRVZsul+lWlqlOHqG9COXd0I62IvLo67B8WPNn0JonyV
n6Ypd9k49x+xmy38QNPlPmhF8kmid4fbPpf7NjrJWWIwnYHka4CozlVnfKxwIOJC+bhWm5OPWFzf
e719+W/5RX6RjtbfAtgG6004AampEmHhpDl9XhnNLsEAR+eTk/Mv207dqKMtOzLXqiFdOrmz9kv2
C3p350eSUaFoufibsGS6TuhrdqPYPxgkrebRi+1YXP1DwoC1B+OJbzY2Cl76K7FGQWF9rpWXnI2A
wspov5A/xg040dUrQ6oRBavSXXgIi15yYqnAs75jf3Z+gTmlvQ5NqoYYyRIl9UyAWo7FzE8W8V6G
E9CiAfJSf56nCAgz2anjlWQWy31kMZ6P/pwsKS06yl6NRWzunLTObbk4DNkdhLYMWF6Vu/b/P5gx
aWvTUbhCvSoZIXPLqbxVBLBXWlBrDPZ/80H89WbPaQkQEdrJar2LgjH74XyrFMk7jT+mRKrzdrfv
HuPnMgScUe8TQka3Edl+WmfLs//MtzMwJp/hOzyGVsqYI5zOhCMqBrtJo3OYrJS/qwIrT4Xt/Vk3
N1estttx/ApjsnQDBhK1ZRa27SiuaA0Mo1ybangO739QKgPIJRJNGrZUyecmte/VjFmi1r1gxRWA
N3T1b/ebgdyOh4RbnaGfVn5/NX+cbn2rtfpzE1oTIL124WjySbX21zUBitPHLN6JbUQCWoxuYwPz
tWo/3At8cs6xO7fPnPCRggr30GtQQIc2ah84gAkEUnpNoFbFSrszJAHMSSO3gjkXzw0wfEFwHbRx
vrXlf6RiKBzH8EOJnDJZz9lwAhnTX8GBrf/cD736c8vq2qcAI9Exm5klvWFClkYe9YVXv/ToG9oT
PECRzm7bNYQ2rqAgT0IrjqdgKOZFieUwRpEQr2MJpgUnO2QOEbkXDe94c6CP9OduDGhR08pJ+zW9
m91b/CsuzMoz4560clzwfPHHRoSMLRUH00PmgjJ2og36CkDaz1kb8ajF1ZcB4vZwWUGWZHlM+/Fh
yMN4RGAPp4QaXj3LL3bCEymaHC+SlFSY4V9LAeNQGAMbQhus1zYZjMP55Tlz533IG5TFiADDqWjv
1bR0ZcaRJKhVGj0BPpf4HCksDG43o9nBFKUpSF7kpCSdmDHeYFQtvMA/nKbqfWF/OmG5YSDoTV4p
qVx52ieCMKfiiSbuAb2esdOZcVwZzJPv8x0CuW2bgjzvM5xfLRZQfRDeSAD0O8WFYaV0YaMbneBb
F+k44rshKk4ypqNYDVrz2l8J7/qUcN03S+wvBe9jM8Rq3s5YGsjyycOV68u4k8C2Rl//2XQYKtCA
0rT6tzDE4GvUFEJrzdlVQ7aQ+8UxLOqWCzV7dq9nDp4I+0Xb+7C1xtxHhL5nf7jJoDN618eo4Zj4
ryVBr17qpaK2T4Tz0ZgcSGDk3TwrkoQXf3lqo3B1NHRfB19KuG9F29Zr/u3etn1G5DFOfc0PMEM9
+7azoyH6f9d/aex76HgwupIAfuOgLNmJSTLKQZ9FfL7rGTEKr2MgB1BsP9mZpi63dBAl1dDyph0w
h0BMXI3BXSgz+X08XfqaNpt8R4PZUIgtao1TBBEeoEGOL9ISv7934F43Exzp6iS56lYcyG0cqvmO
oboVS8lQRHplVig/WHFOfifOdNOGmZOEI8wx8mpJ80ki2Q4pMXOBWktdgU76tvuxZ9PwDNs1xF4q
/UHYWTlfEnVkOtqzjBs0L0qE4iowIBr3q9RhjzxBGCdxXU2QKwy0p7FgIiRWc+H2poyKLqgU+h8c
FkGKWgDKgDFMDNfsUpBV+zJ7VpMrJbQcPkpw/7mMj3YAxIdbk3GQO4nJRJaH42ED7rgxP1eowRYu
LbGTpLra7PVqInIGbHQV9ww7ItHvM9o7gGYmmOfbW5WLjWbDcJAjOl3S5FXND5QB8vXM+INau7vP
n2v5rFB0mRGzaIM88NG19kZpWuIBF1YKZaC/X3FGs18YRKPWjtjUsQgBCiCkHklmT9g/MAcHxMCn
cUrHqN9zrE3sMPO4IS1HmgTXS24P2Hmh96VMtpvRHdv0YHmkixzlGGyqv52iBX4vKu8VriKW+NLF
2EnQhdnIbw61Nm2s1VmSxaYQvG2tBMX3g4u30KjDZ1TxFOLNVX59h8OR4VlNcEVaifqEBR19P0PZ
LEIAGfgnCKhTQjSgaWpksE27aesGYkhueaLoSK+FFdAlQ5PbQB9Q1mCl9ps44MSqQLQkTH+/07pn
/MaNntIIhra7cvkU4Jm+HjdK8/dje16bHqJks/2zNkkp6oQb330nFdSvqCO2IB5tfadq9pCOf/cW
vl/Ui6F6kGWLYQGO2IJB7OLqcA/62raPL0OidxEUBPYPldh7PjzzCHzT4bNMobpcSQh5n406+Y0E
HHBQK3AJaVAUlskKbfGrbtD7G0DKHuwd3OBy2e8Tcp/mAC9gZwiBeWpEA4z5BpQGO20lYsMk4uNS
Ti835AccYTWF5Zxft9rlvVvWeJyV7W+PhYy5flffPbFFZ/8bzJizxrd5rIQUCduz9edj9Y729K7C
dl7nNDvEltYmxr1fiKHI+Yp47XLdWp/QiGDba1jBhukuKW1WAzukyEWD4DT/87HZTfsBlgePIy4d
YkYFaqagQ0j1OgW2VELVKU9wkwnPyCanVPTMo+1JqnA0XJVteyZedFUUbzVyvScR7nAhOyabToaL
ujUpfrxJTA9Ze27S402BD7MQgpYqucjjclI6v2BhH9jMGZBZqJZ0uWIj3btZvmyBF8MQakuHIz0N
Of+xKz3eJEf9fnF6X7oNmqegOFh1eYSCmCDGJh/AGDXSeiZKQvqnHpPZp9XqvOIXYmttFl4eoWeN
4njQKb41W+IE8Fxz5WYmWL8h25K6RVvVzGAeZEadYa+Z4Ofs9WGiizTRM9MzdqLaWWVW4SSf5kHc
2Sk9uQR2VGF92baHJEHuG/Go/dWZlEmPzGDuDTms+YQF+XScbF537giIC2J/qLQrmVlvmxSI2yY5
v4AkCbD5ykgQwWO4h/IyPI9ACgRWBS11dShl/X4TAZos9aKw5YSl08ti1+hkEWHWnetDBo3KDuTI
TOo/KdNQF2YJQR6e7i/PT37/7+odMuHGpKkad5jDALNzEAtLzOADSxfR4hxjuD/D1xHUYRTY5dJN
KRGvPyVjYdCNQs36SbK3rYpTXVoO3hVN4mpqYo0PqDrUHWA2JRVQyrK6mj6ETNwZFy7jMLXrVUYj
14o8mzIPf+YwMW8zq5eq6rWrbv78noezBE8EraJcemHLTGrRdlFFfWQ9I9LgEKD7OHW4IBbrstPd
lVGH00YjZ8215hpZGkAYyY3bLOtPzCZ53Dt/68tRcJ0bCZF+x0BJ/uZd/00IX44v/REEfG6vKRRP
QRsHLZ8KaOXBWo+uGYqi2HMFDkbJ3o2hGOnJvZuo022hV9oG7/NNyopIxwJa9Zy9xmDkKbXe/UpD
SX7GmlEQZDzFB6OpO/Aim8GG2H6tb8fEtIV8BPemUFRCgwYonXgEvuN1rrlWECY1zXu5uQDH8p8c
xlxrID2oUfiBiC09IEpXst6sDNwdxsLJL2Y01FDpyAr3ZZR7D/TdCOcvzoWb2uy+SevGY1N7Dp0g
gst6D/grVJMXuq57Cey9IpWCGfl+lIYqb5zmYSNjNQ6ixRyjMvATVFv2Ece0QgkDTLgDzb1TPvTh
0+/lXpHSvZM7GDN/P8sMZEv0W+kXOx3xfBGOg26fAXF2pNz1gqXhkTZdg10uI2HeLq7/DMPhQm7I
uVzD0AeQ3ITevu5iylhyFmGxGFQWs/4EHh4qAx+y6MgyG1Uo/zSjthL103IwsZ87Qho1zTixZO43
b68h8PAL1V6El0iFHJwAD9POFN+ohKyn1NqPfIBDypz5DhzffUDgRax/3dTAVvX8E8Rksl1yoC1d
qxhLu+R45902oKKluNxYDnkCcJQKFgvKigxUndfuv8sC3HSVmnomhxjdWzdFxJtjoreU9apLohqQ
y0x8nRlRfUmgyQtMS9ZGvebiiQV5Uf+l3ZeTBb/QkJK4pxTTMsyz3wdnzdJOdnf/YZESfglayy8C
WJ5PPSsAzgeCFftRA2lCLCilfotPmOaw5wK6VaTJ4egL18tOKhqapsfFrLHxIQN/1GrGuxwuqARj
RLB8IbuWqTjoLK2z9lG4Vy8esAUBNvqb2X1xBhkvmVj7ZzOyWO/+nweLZ7KTcOug4l2gqn3/CUnW
X6h4uNCMzaOxXFI0UBomK1klh4rDHgq3BhHm9lUGj+Xfnxmn/Cfo3pqsJt99f2jYxyGdPNTzuRnW
MAFmJnDkLzSE+Xywg1ct8ylJM+JRacADsLyWpsu/LnWex63KLaznlY/3G/oW4OxtF0f/TcdbLurC
Q65jGB/04iGdFf+Ool1BbSQjzD2VgHzJ+Ew+apvcL6NzwfJFBQjmjnJ6j+k18kfeTHwzBl2RN/XT
IWg4vq/kDDAjP/JHB+EoLf0SKZ5sts9pXF/D/y62NnFwEXpDdLezJ5BaQiCkc1yQCZwFB/io2eTW
mEKvs8P8uUa3ccv87JU0z/8+WhdJB6eqz8rXWVWXRWtA65ivsGGgjnOVCT1LjBMFtOpUbdKlcNkf
5P/yna3/m2h7a+ldtw4zNtzBap3w0G9uZA1dG79VDiWVPTV11n9kOuYS+MCnsDRdcTrjbBMcMqoI
gNG5qJLYKgAd6X82ggsWPh+MYPkTi8PDTsxFMgi6kyQ0/f11ND9niUN3Uui/PqiAuWTpEloohQ/t
jybxPle0Q0mhChBX9gKrd8iVACSfgx036sUKFm8YcLIuIKFdhZo7SqNLijNPlLVJGqZhwHCG26jm
o+ni/vZPdbbX9ArdVXG5bK4BmtMLbgWCMFLS4/iVh1bIFLu1X594hrgzxf6ZoCWl4PE66DDvDQxK
KzPoe3ccZZv0MQr06PhtyB0xTLzuaTx+bDhLXyoxbeJWoy0pKuUQiJ1SkSvWGG9VR8LpGXPLRLSy
Lyel520EOBtI9tP4bT9813CPtUYjrmYvVacMfKRMxUytnzvnicanZkHuZsjLQNbmRo3rAbQU7wTR
9BZ5tFAgql4u2IZrv7mx02iM/9DkS4TKZ/SQFE3EOwwoLr/QmA08sONp19Qx2Mxlv7mPfFDo3QJy
VbOLAiCxmtbLXIpRT2eir0DJbeyuNPdsTtPKTzUI/UUjtQ+yDgmzICo1VxfgVSXb9VDfp92wpDeN
jjlMrc5Cq8y90W1gepTGuvrtmT764Toes7a60PtsUFVaZMICXjyjgSpfd1ZQP3e22nI352pv4+51
5CXmWVDsv/WvED44c4X+TXwUVD1ThsB7eiM43Lnvh4IwaZLpYBXqfSGuUUL+HHdkgu+PdWgcRXuK
8oB+innhEoKn8VkPvIQd36fdPss6mUMmc3Ylkbwhcp2m1H6tycIupBbNBHLJFFaiQNMFict+RYbW
48od5Sr1b9gnFXYpIz2LtKrgSv1jQtGmnPeJCc+CwqVV09JKRRZocfCVk5neP3Of6D79Fw4KXl1G
u9U5Ck4l4kp8X/kFzdfLY+4HY15yavfin2vHYIpG2f0v3PDq+lAr3Hedbe+RQt0EG1/hTf71F7eU
FcrePe00L/Fq4+DrSiLEHlX9p1PYjNUi7W3pvXycx+nYt6oth2qD71JOLDNk6qs0qh5fFZeXwpMj
d0BlT+bSQEGbsqzapAIc6Wf6Nj2vQkgvUx0vox3/6mBJFv0zqDQZiSsNkg26yk70FzkjqWigQBiQ
JD1UgZ7F95CLzc1PcJd0Q58zoZG6Y51I+bn6R8xOmNlpOQnJ0PKj+Xet68fsp//H49NSsTP1XjVP
IbNW5Njl40k981BYbVlAEzed7dldCVoRpTFad7TdYfJCJqESSsEHxGUkaFLQJDAfIutNhmVdOMl0
giQz1GMzk4sSEGsDs6Ch0gz8uVqAfZPJ1jJMSrs4aTNCuQocQC6kN2NVp5wh4xyuTvRO0SQXEhRX
iTUmkQFdCeyvBp+Eq+uwvBbt1NVn4xC14IUNzW+n41xJbbdCEXZAwk62PGEN6FiqKoyPYreNGbNi
XSwTIQrbP1a1etfzf5IiVFFWoJOKyaqDd2fEs88VLMAOKNstD+wDj0sTFsbEMIyNoeP4XXcskl+B
36xv5BI3PHcnG1Vo+JPcJrWbCbd3Gbcu2rqgbBMuJ/u2BbqboN0RNCrcIB1HQ+NqVU3s9W0pJM+j
ZFyAOzLVsnfqRUb9j8cPFbgYeZkJJuXyZqvvIoxFel4E8p+xGzw9g1oZ6Zyhl1r8BtmeCKJpqD9Q
fd20lomXneB4lr22tTI5fiFRAVn3QPt3SCOgMtxQ5VOPwC6CxSyp85nFlNACS0Nj8xzCxD2Hb9Hk
axuGq0TkVsF3mw6W4p/LjcoNNU0pvD3KrIsNyReK3ccmIx/xcwY1zKCX5WbBM7KEo7vCeOANx1CP
HdEEY7oJvWxRNEtedn+6nntaZNAlzbgMZNJFhf3iWU7tzCkcuGa3Sz8CWOOxETJkPc+tGth0Koqk
JGdb432bmzT10h9iMXagD1ey1mvuBJLg5IVhIwPwYgTl1KCnXw/56J1U4wU2F4SYj6KliAY67W+q
81eHplBK5d+WW0GGaL4FYKMIM9Nin/D5j56TCyWRlWlgf+6teynBfVglnAthVOolY33j6js2+2jv
pu2KR3IrkjwWWFpbJtWx1ZomjtgjZxAhUvGxNWegTCv8UUPVny+2sXfgaWGbYzwYIYUY9g/ea6ZD
tGP2gCSH06n/4CIXz/itbGdPPEN5SDCNvqfeqM+37CZdyJuTaNxf8hR3cNGfKFEKTyz7Qulf3kMi
L+v+2+coO/1EY2GN8Ebn4Yltgpq20VEY/IS2aFwOD60GMTD/1dHV/TsjIC3PgLWqGId+dn3576AA
XDaUn1BOtipM/zacAoirngMO28lcVOTbQE62EvCW6ufhoK8990FFEEh7mbvnhmJ+2MU5GvshoLvQ
7pjPBedmaWlvTovPafwxQ8RZtkQaORpznjR3LT5uoBfo1DKbQwhWunbu4SVtQtWWYOrbiGJO3Qqv
CQhY+JNTpzcEps7OXvqdUTu5JfA9j8JnfnKETd6rWozWLvK6QbfkO7K8gO5yEW+D5b3e1m4Hr+9x
MKtzVbvSl9r+5izXtEn+7o1t8SxjXZCZOj/gW/wiPQXD/7eC6PAHa4bcF7C0xny8uRgwpGCX5jG/
l7Y+qwkIER0JZY4enI8ACe1M87YNf8+MvWq+bbk18LxRCoUAmYSRz+XwbMlB2zr1topQV0HbWtdH
Paywrb67jovmmTneyiRbojU9OR29v+diRU19T0h6DEq881aYDd5UVH+zf1kIWZwZfIKzlG6atpKC
NTdDDhOliAqJ0kMbMek2e6vO13fP8y70ClUuOh64SN/EeL4O5Wu7Mz0vdVOeaoPNNImnl3ZkDR1Q
03ye8nMLhBCiHARyKkTYQaR7maVCRycoO/T0q2YO03p6O1/7L8IuGF/0yU9gJyi8Zaiby2HJU/NU
KJe16s672YoaE2P1UFKMafRKKoRNhjNkSwY2kDvp6xClNq/APzlpogdenzxI54ns0siQCQ0zPamb
8e5IINE5NYGf5c3f26cTN31OHcBydFbPR0IOMCwK77cw1miuYzQoaxc+0wvWh5JPLGtX2QwPCcb8
1ODgGQmdPJDk0LlPkCezPjbDlRBPkYYT9OFMmVBzUoLdy8/saueu2Hp7wRI5pULr1Xh4HEMv7v+8
DS/Sro91X4mVT2+kNXLUgBxfU2/Wpa9qHyCHM8odA9bNo0Y4WnbuqveBVrWOBi3rTQ63nyyAi++F
8iTvZnsZ/nRwMr2oBNhaTfQk0x7AwpRjK7NSkazHGIuQhNSbKI9zCvHLuZ6OHoIW0Vyfcpt6/z4n
jd9uZTk2Uuo3Smtkhn3CZT40DWsptNBzfcLGl0cQIH/mZ/xwaW+g1H28gHTpIjaODTAviUxI/ckf
04qsSh806IluDMi7X9mQarYfo5cO0ZaxrOBVJrBWweycTrwpTtPItcDQmpaisgeTefw+6P35CWzl
WoOhXgLEiRxxtw5+RRMFZuYA53+75HlqWCswX4VsHjV9hrQ4iO+O/gHWD2vJFuimnlQgBUU0nY87
5svvtqpDgdaA6Gx/QYFyc2MzFCFRYISK2z7QOgvPLHqiCa/DoAnDM3lMcmrtCWD+v+H/gUl18vxb
TwLKnjzasyis7+xt503kJdYxIIg7C6MDRfzI5Q6vSWwDIA/H0/CdTwN95lLyZD00v96T+tU1ECzF
U+dWmRdggCQ3PDEWq3izz7rVWWmvxte207tDvQJkrvbAdSuYWj1SYwQtlAivSA0cBdjRorPT8Wsl
x6DxjlghRRGl3X+lu2k6RGiaa1nbx9MlL78P+crgHIL/Xn3U0Tz+R4I8sbZknW8HwYRpfz/XCmMe
hDvpiDUu7TETRv7qGPJIGUZF0TPeKyfXLbIjv9ThCn+TydgL8Q7zIWawEAxM7ONv9uczEoywSKN2
X6X6LyF4dOr/bDwvIA+rJZEf6pNDO34r0jA0BvJG0/xf7lZaxUzavoUr41ToK5EPzJ6ODOpaDzhv
JtzHA7NsVbJS4+85nK2pBS5QNkjlrVSGOgGxhnimpKcX9cHldgW5UHgjtE+q9+uHfhHvoUrDFPHM
og37+qRAkipsLXBBbIgBzMfILg3X+5Ws0cIemzkZYnjlDgptvbGQYmTbRaWD2tVvtJCLJv8nn5aA
5QNI9NR1CqTnNa+HPR3GCEMQW/y2kgJfIMYmc4ZB6pjzSa28SLf3jFnSFeEHSDViBda3zitvW/Bs
luhSJrtXPA5L7S9BdTf+/32Oda4/9TUAYFu6XjX4MbBf3H9bP742Bq0cASDIJPZoiFTswvSunEPP
3YOf8IgVpo2jR16ggcq/mlQU9N9ShH8pZ6BTmdU/rs+IHiP//Yab1MXVNoR1RGc8SVchUeawRspu
KqQlAfSmOCZJY91cZ0UfcvvGNMsAWyoTQoLvx73in631TTxT9SC9OdD/P+Q2Pt6LmwuU3I083Kll
TYT4PucyfbPTI0Lhwq6fkFbaqWqetVmYwphMIuLZ8bxO6+VvT27Zvuf6U0XeEDI/qHjswMMIAQxG
PHZP2I4iMHZQdWbU46RddV1xYpUoB3n0hPqSMdDpwwIv8XMbVKB2z2UPtwj9N01p6uvxPcJWVvzC
SHs+7gr32UmnfuFTdLypeI7r85mHOV8cRNyqFUbb0woNqbQ8zHhjmWC1chsKGN5s3jH08euZzu/j
HWNXZ7GoKRzMc+gHDz6MiiXlIvwAI+2q5SV2B4JhyPdZOY6WNoF0JxmUCNQGiceoVEhRjzEGZMyV
WQUnvOWnnD1jL9W0Ex+z67bk0yNSmpxRgNCYJHiTTfPQf5pNk8UJDK/2FgKwODFbdAEhVfMfpPVM
+P3oz2W2S9/gfzKstAgq0raewq00TS5Kr7mjRyZMOMXc1ekE27ucT6HqcXP4suZq8BkUcgbP8HbB
2N+jApPhrg6Xz8VzFs+yRrFy1A5RRaPstbbkDYWMGtnlI3SksonaSE67ZAFtum39ISmGqv6y2Apr
lTWsyP3IJ9CYcTAURS8WGGUmUtJn8cTkAVNCk6MB0mpY57TVAi/xuDQhkSAsnhk5uVgoLwjsMzqX
VWG2y26fnntk0O01JlxC4ZSQ5XhwW6tZRZPnex5IAPF/tz1bS8oWzP6Uw6VNmvlItMCWkCxFrfag
vqQCdH+n49ORzr1zUnvetHlXjD21Qu8lL82a4HEZ94pRN+YTslZUuOTYCwL93nqtFTSRw3mqF1T6
o0R46B6hQK4P4u/WDrgFAuslhZRZ32rZbOGFEI4hfJkZYb3tgdg4fNTdpFF2AF4fITCX3ZydKbwe
KUhl6ouexVhHwOsRCu9mhDsHyDMMtpVfO4iaJOxTcf0841H8wRG58QTSihFDaAKArmUWQtUzmwFk
1LiscG3jP+LtqKCnEWMxFCVX3KvvCMeQdh3zB3qnKWIiGi40hNjSa/hBDWswymiwey5y2niKp4pw
1Dg4OaVsoLC2geKzXWcvEq9zVwqYVm7N1IJEVRq0PVrgWqOvRT3gvJZnJHeCA0WBisEbJVBdY43J
2SW+XKAbQ/IMfrpJ+X5xHghfHbCwVmHSL1y2XFOrIMy2Pgwb6t2RMqS+wdtOpb9IS9vDxDgmfaM1
AT06p9EMdzpJ2s2MMl5tDa662Mxf8pYe1QdQEDc3WHy5N1mL2D/bqhhALNafA6aqlgTD3gOa5uIa
bNLt6houbNqtHPZMY/8FSQoCa5FBMkUYQQMn0tQxm5NyC7HIOkcS7s66z3asHEpG5NA+puYGTKHN
uqHCUBuG05esXV6724yBe4s6hooCL6MgSctn1cxsc+ZLfXxS4pVTb9JNra64oh37Qr050oznDH8Y
AbMd78MFykUs8D5ZA1yaQAJnQsVfXMaQWenr3mx1n5SKUoHTvxo/b0IKA/jMvQCyAKQPBEpfq5U1
Hxzt/+y398q2LJwF3ttmDgjX4f4qhUkrHYceY5j9j757x6hEiJotrLZA0Daq4zd2SJj4mzGUc5kc
pS/lrNsHtVbz006OBTWs2rj621zy8SStL/bu/gcELWIwZNiOpWrkYgkPuaQI2bKCXDccn4BfztAk
ksAhYFAV2qIP1mWR6/YUipFCoDCSyoQElsWaUmbDf8yaUfkB0ewxgTVH6F3mmQ/WfD9bSJw8vbuA
2PvFcwPwoSqwZh8wCP6PmLI/hNjL8m3OZlCBv91uXXrFt7xUsB9zPZmQmIol8BiaX9eeUKAH6Mc9
eatI5vJaKCA/dUZWw8QUAU+yy94BuLZbVD+01nOAQ28AaF8on262615lz6VOYXElP41OgfXrHcgi
0Q5/SdNKYklRdIvLp/Sr1BfpW/4Tjx0KqT7eyLOMu+Xih8gNB0W39sgl/fWsEl1e9wthJ2Tm7WLA
5JgXc2P1ns+1Jt1HM7rPsaggv4cb3P7gPDuH3Uk5wyCBvwsi6B+qvoAlH5lS/Amfu1vk85nPY/Bp
bSE34ngE6ux3RNXW5dIw6jM4DIXa+Idd9sS8qk3i/XO7V791jthwOxVhmQZYV1SCo2fgkAkvqitw
5+chhlAMmlPQsFv8eH+grEgbc79NdMBjImIfZy8wkZ6kdof2wCpapf1K/1wgqaDLzSlqtQIhLLe0
nj4q3tFvbcwJetts/zibcQsVZATvhTG38+2JZvh/K2GXRRdxXlnKGinSZdqqPslJgZtQL6yo4Yf1
Cg1d9maIr/GIL6hvnS7MzRmg9r3D8Q1xISUh7SZzzCRzFX4md2v3DnUNYoCfcHTQlQoDIN4kh171
IzaWQtL2OAbXa905KAgjhkpsLKblGKXNdYiLo7uVp8/hDPROSR0hOdCXf5DBpNYg5WWbcFQPMhPA
Yl6agpdjUua8vBwpJJA/MaStwp/fL2VBBULhX7DagwL1wjvX0NjAeQe0FP8/rDEv6PsBPY1WjEv2
Co8S+2qslqphHnDLV74EJcwEUqyhAv0JvjNBF4rHcVFMyOASU2zwgGYkagXtQtyH9euCrNcUOA+o
AB7MciXhgvvnWQ4kXYeA+c5IAEVRJYR3CmQknABR5clsrRHFcrFCP4S194oYOOwNnnXJDpkGlz//
o8cSRQdxGS0scF/pzJl4TjfcRLvxnH+XRD90BUt+LGdE2l/wAm1EZRjfVKtO9COw5TUIRo1UI25A
IdUbZ5svLxgkPolkg9skVlsluWI8BlbN6dzDFm4q/NmLTFEjXwmYjI3Z5fpUxRwuWFEOYodL91fE
uvUKnH9WuKq9ZeoRu2ESoSTtQa4lZ/UpbGODWu7tp2Hba4g6Cq4ZmXmLFt3vh65QQvaKgxhWtMR8
U+YvyLPFxBUkQg43Ny94jLpIuiByUyh8NKrNmr8nS3JQSj4FozZbfYtzCJ9nwwR1F3oW4y9Dqxv7
+odPFMpAV5TxSqF0+A+97McV7A8M5sDYF6BwiFTyT4RqOE1BVgrbaO8bGpcVNef6HtVEXskhiVyC
FTcgDU+oMfiNTuwRI6Jmsfhp3toPPXpR56fgjevd+kakzY1hxNTQxjtQqYdkRZ8y2TPCT3Pl+opF
vGC/RW/hYsRzLzdbiVBRsE6XX8RUUK1jfDF5/mtUdN9n49yMF9tuGcmLQAzpcBkJYItnUiDqUdlz
0239Hs0MMxkjvropH2LT/bwvSZE6K9rMaX8TybODc2auL49w6dHFSyZwpdk1JNbpHsssvnsSsS8x
GnZXDASlqh61xXLVINV7hDaWm/yig0zZLexvvH/MAwNgOCB5+g9U0EdjYQ62bvvWn2zLW/zakP1y
JwHU9tAi0oqr3GpIPTY4Hh88ilFJlzS08UcKhT5QU3XLX1ieclvj7aKRNqWlIcumzoFqiocPWHkv
03A2Kww6z+ZwBX26ElFNlKXIWDVj7sdpGDqr3ShKCm8DVDZcDkduIrSZ9IteZTmw3Cuo6Lihs9Fz
Yq4hqg0bjtLXfbaVPuN8TfKNRvIgqP3Ndy2gQKQD0HAlUgImwyYnIUN9X2UzMO7xpG4d6bgiruRd
PHiP32ny+v0h7qoYGjdYHOiXPYt05Cjk1YuvZL2BBAEuj8CrdoYfrZrsY9akDuXigb86DqTWy39j
j4OVsRxOXRIeqDy0D23NnHkK1PkZxkpWW0gB/qfzoTkGrCTCsQpU5PACQkRrEQd1XuzGpVMBqhBA
r9nOb1O2XOEwFWKAFbp4R6E00GU7PhHVJrp5sx06vQZipzpV9AML1dsfcIvoeLjQhyCRtJ0FnKvp
p0jq5haagfdwsjjtpqSEkndNPBPecjy6vhuxaqirSjWQNJAjJUf9gyiuFuEbheaxgyOSTzSnsm81
5A7jIZnMdOq/TZ7RKDttgqSiB/cOulcSby1ksiN85PJtY7MD2MO9HFCGZeQZfJQltOpNsI8gIenA
gHuLXD+foHquBh9QGO6jngB6GIB5XeStvcA3Ph8FMIZEqIIZxqvhLBgvPzHKESPCFidb2iAdh3Ki
tqBPZjMQleS5dcpxlmYD1ErOI2E3ZrZwOZlzbhVtZNjCcYd6r7DwXQuVms/t67mEil5vWjF9odwL
CEfnI4RBhMXVV459cRR7bMj+Agwn4ZRnZgRLesV9hOVMRTJGvvXKtn1AxJ6gFPOJ5DNEO9MM/nUv
mSreiX/IqXGPraGKqMsipUGo+L8NMlDgiNexitBQLmXiM+xgz7medfXk1P+5oJsS3K4ZeiSvAK6g
4lchc8jGJtWxQVzUpu+aR0xpna8DMIqoNVK30VP2KhyFbm0HZ/OxMfFOLjM9lLcV7cm4fCafzUd9
oyFaj65pg/G4KD+Z+DiYqdoDHJcNt5sxPd3JhWuUL2ewD89sqP6muhgxfvMUEsoBPhsqEqqs1Mn/
6sEYo3aOgfgiLK2Ym+0TwM5TqsslYHClrlk1LucESYfAqyafPvTt8PSMwqAUt8VA38as5D5UIfQC
lqe2DH/URkjWmD/7TDzDrnqQeau2GC3HmOTLmOIjIMZ2BKoz6d8SunbS3eqhRJUfcysD94he+eM2
JP0mxr11r4thvdVtc4ktYqvEXwz8snZXnWAGxV9NhKkFqHR8y7W89zF3fBHwX8xPkOu5uWcIVS/s
kc+/avNdn+D16asvBHCJtxtz7Pv2CYaAXhJKKOyYaaFhJys2/WVN5tx0iYhkpFeBbUCIaUZkSW8J
Pc19Y9bn6XN/avqO8gKBk5x46OthqWKrxFh2brrFf/w0KWQmGWbPAVPFYlZpi9PrVpGZYBoBK79A
TD5QHeYSesKyDRzv66JMPCMx6+PSPzJUsljJji06PVyISHNxS9B0SQjKkNrIazBfkSyApmblhje6
iZqhVpbhq1N8UnDSNCnSP8AsGkt5PdL6jFRITTthiiYBUl5Y4nRe7DoRHFXfOUklPbGeGtf4d8Q3
ewC357Aj7G8a/+gEmDYpPPi7rJJ3HgaVGQUNWipuHenGnz7/yVu8whx/zJ935VIORV0RppIKg9Nh
guhvSrWfkb6Atl88HMDSJHqkDvN13qdkXNJ3SURCMlI40zqnzkOyk2kQ49M+v3FGXq1oQEOt9Sv7
PqpUuldLdpCheu8RbRmuXVj1gkicn8pTW4g5+BVoS9FJn4nO2S/K0GGtlH3YB4cc2eKNVzwashbz
1GwzlHlPYBl64RyMKkQB8FxVRPQ6ZtiX+riUn/CEfatU/UWUBJhzaF7ib4UVyqhmi/ApFcNlNdWW
CrcqCFz2SAOsmPEUaKVeAUSxgZ10uLhjjTWAemMKzHFUvVWBz1BHIn3sixx9ehZoPLCBUERarg89
j/qg/OEMu7q4hRH8Q2/HYDeau+XKj0V2r9mpEMcNK1Dp5j4p/alyI8LamEJl5EMeeEmi2m8BfEgf
4dQtmsmAevzgL+BL7smmWLZIymu9ZijAIh7joXiOrquWEcWI/RUD51dNZPA4CEkF2KOPlzX/UIvV
TPcYe92Kv510iZHZPl4lp1e9jhuwN1PW/nHzYbebdCFJsb+Hi2FuhaqTwlof4E/Xkr1bhRmqwobC
8hVqq5l3BLJGPaZirNYmuMsdrn1IoX9MzD9HqIbhQfI8LLWB9paR5sSG2wBnC3pG8KClHBsJx1ri
vy298H2de13xNWCKr3NW3gO5l7U/xLavyGX0gUNRG+9dIg26wPsZvqkGBBFACaK6cXNxiAclB1LR
ce64sqwJ1LjEgcAofLFUqXgwVzl76NuyYBGZJwiakiknFOdZa8JagsP5iGSUBLAsDQIQ4jaFA+gq
3NC1B9lnGrZffzYmW1C7WofDprS6P8lEDoI/zWtUm6KCWXcTDxqtPW2h8nnFp4Vjt372hN8651GQ
9kaqiOSmFfR1prcE9TkI7mP9wZiMuQWPrPnbNwxA5jUvW/jS5TvcEjABQpfVOtt2ZKx1mBjvNr8u
9FVI3WWgyLs8yv8aklasD/7oCcMU2rEq0fDrdvIC5xlDfZ0wD6d+cQ7dg4axwMxjBTqtaopEWJ2G
1TGEkqWeBv7tzQ+WxUEpZpsLY8UDRqi8d1zD0PAQDaA6z/sD5MS/4cF5z/Lxr6AyzA4taexYr9w9
qXeZ6TCMY6ivrrc3Ww9YeI9TKTEwpcixpDc90A3iIXZ8JXCBMR2vwIYivi+5A4DPz5DaB8uLAZ+O
m3/Qqpi9xyrHOsTiyHPhtE0IjvA2GH0EkHEeCFxuOLWfbnjuUa4J644C24Nt1GUTonpu2m4DJynZ
XU8Pn5nmGOfNu4kNd26ngukIo/58LpEdaKwt7/0LUqklJAB0jtcH9QJDmc/0vePtF45gzEc3jLPG
QWOMMNqIDNMYIe+QK45aVA1PWyCIhohzoynB8bEUOgy6OboR+wUW7eeydv+G7c8QcM5H12Oskv8G
opyP8ne0smsUkyjtHSyu+hQlvSuUzFm2Oo69PzqGPg0/57fJdkAq+HnDwz7FrUOhwaM2K7sxVmEL
zPZiqYYG4E7vddtebp/0Sryf1Ou7lwN4l7IK3P60zzaj4lFdt1IvSAA13prw2v40ryfgnmKvYZK1
lD4vLW2mg7paDtFa40xFICPMj+8bmDgsuPk85veRjyNlRTvcLRO7hnaW/6kSYW2gwZ06ZoKROX/Y
wE2GiCc+khbFUUlxGC7+ipA8pdRnVc3HFdd1fAUfge9R0Jemi9wLzAYqG8V7zuESyotZvWdIMCrC
c46RqE1u0sd9vTKzn0lx/9TY+dNVwHEyRkUHB7KZbYhgDSdcNeBvH5hIdNDcVjxWVUCKVP0Mge3r
gHT9FXZITGu5Kgj42+9SFUwNq84qc8rCLJueCGADGzFpbdlAk3+thG9o1mD1dPk1xGtqmpgLK/k1
ocX7gC/s+98kACd2vQ1C15BcadTo+5lu4FO0bdelJ4vlhe9LUW2EWoKaPjlVydeWCKp62TBK9MB7
5b/LdRTaxo5VTz1orDsHa9+ta1jrfOgUdsN7+MnQ43AFKqY0LdcAaMBPIzS5Rara6O3wo7HjGC2j
FrKJ76K95N+n4JeiqmufRGZ5EpreIyXPlQhb8+cYcXnQi3zPzu3A70WOCB8iXc3FFyJHbAl/i9Yh
+wB+8nnw+X8vAQ7FGIUBIXLU3BGks7JXmH2yNS6p7B14iVNTGT8LE5oV2WKyQyYwJT5BDWBz8c2K
G8hNQubsDjqFmb0mJpM5jTchlcpL+gDAUOy1qftPpt1P9PVw1UeNvuzKGD+a5WzQ5nGRwfasqNNh
EYbpXRIeIB529QhpPdJQZPk5hEDDJfqCZrhglgD9yf+4v/ajXYUwyRJe2dZo3BxjIHeN5+/cjozZ
tOkptjF0IABy481rqpq/eBcIxWzQ/TXwf73n167WQwfuP2YkGumg7jc0oPl/ERlCAa7zEhOGReT+
JkG8tpvyyVOWm5Yq5/pUYLkD2ZameqITCj1113QiDGR0y0FTCuQBiysIiYP+IkjZkuB18erSzmtr
axFNsmizyXloEYfdzM2wq0DD4V3Fa7BQBo4X9eoe5ZIVax+M9soWj3ufCPWyZjw4rM7a/Ii1pTw+
InQvMXmsLi0AxkkWYxYAji4aX2iH6Z4V19kBrEqpHyPsF3n6fs9KTPJeC1/ZvOfLqsGTojoCEFya
bftBVbLzPkGB7BfFhDnjdKvLN9s60K4ct47pIHBx+RvXLzgkKT05Dc+W87yAVNyigGCfTf51BIUi
uOsSHcqPNf8SunDnZgTIZ/v6AkmNOuYaOFD4XXAbO86ZQ5ELGlgU+ixuu9fls/jG5caJmVA8GUXb
awI2LdzjlDIR2izm/Y9NPlhyZeMGAYxMuIvsJg+DpXkuyArDgi+1uYBpwpQX5oQ2QKpcxSDWLA1z
SUUNY7vQuVVSWPcU4BC4D8OCPCVA/GEip7oOfxvNWb+HKtoQVAI8ElzxJyrOMebBuc5Z9GtrLbKb
hfFtSrZjiFhWd9hxfSWUtFKJ5g0Mb2aJhuAxSihttz8N82Oibc3dP8BF1BlFKtIYcYQcp7tY5SeO
Wn4G5G/t43a2tacuVukATIjIhAF/9bCX3Tih4zu6tuPCQ+Zc9HqI/CTn5RINZ7UynEeKZVkMoppi
4rRMuH3w2n/muIJJpyNHPHBAtkIfzsGumy/mAbZ0EyRFmT05jPlJkJjGfPwS6AddySKY464duaEX
uXLHmiwVXvr0lC+vdT/lNFKWKTcq5l4B1HQM4WfK1wTbCTloCz35yJYU6aXhtwSeW8RvC3TbjFLQ
MaSbh9l9kww8KhSwJeWXx4lPdWabBXS/uiRr1W3R82AxKRbfCeG1f8nVvmHxmPW6tBKovrpOnYx8
AsoobXU2mvtMu/Sy8MM9FZ5FwFyItHa7D9S975DjhiBJoBRnYrD7Dgd5I16uu/zVvzIq2DVTDm0K
uuWKxcu3cPl/IeLYNAYvlVhWxJboLIDouS1XL9Oqc56BI7NLYykfRMV+pNvsTKLGvDLIugBFzgY/
6VrHu63SLr7m/0iaMVG3xHcTV4ZCyQQkUN/k3HyIATjQ+6S7nXSQLAX/ePeBcewEcCU2ZZAKfPCp
qmVl/Eb/HhfWi3K7JWLauI0ZBTv4l03xBZmOIUSYf4h4cJLqhgkJsggZvMdaiLiT4pB0jkFKhRUS
R3/IVQ+3MDWacG4bUiBxug4WokzRZ0CWDPRqT8hOUgB6EcE2nACaJuVu09NLbILNvJxIFDACn7cU
rzZ8OgiohFYscMwYrDW9l0LJ27/0yJokQjTcvqr5mNEob1TiWAOFbm7xmhO+IgOxs2o8hkg1YiHe
iALP1fMrw78BqV4cb+YG59EtPT+syrW+GGz91yQhxR9RYkiqTXzCafkxRaO2FE4oAQCAk3nMzMfz
X+6/l79nfJXpynCQXNXM0Z6+uJ3wLuySfnIsKqXw76jpDnpAJBPUz1jmOHFFWQ5gkFvJUGM35G6p
QbwF7Qulul/qZYyCR6ETB/LzSyFnyAbCrw3GG0SJyBHMeAmuRkY3f+4yj6AO20hoV2RXqlfRYjM4
lJh2zW+YX1IedJ0W80E8P2pDI8jt0IhiRrlso4qt2rrslAoAaL7Rt8mwdMu96xEcpRbE7050iXjS
PVuYVT/jz6WMKsIj94SVJJ5V5mSCp8DdmiflQKR8yzqp1iDuVNisRRjBRsHyjMMgCEvjcHOS+0Nd
y4DukXRN7XW7NtXHmrjsH96XzzEoX4JKmwjrA9i1+4E6RuVJimNsZIUjhwZ67x7G1C4exVL94EK5
AdFAE/zldiEeYOlNYmYaiTi0wiAZ5geBPATF70JUKGQ64clxQM3QhrRO7NW8UdWjf+K2puw8jpiJ
wVaoP9uIx7oPlkJ1cFjmydHmaL9woqhDbgTcpIZW8oDJzrP6SD3D4/TlQWyYjXuASV0rKjUnM2zE
SKU7cMIITWGbE5eOgqiHqjKsOp4KfnA1CikYqkf/wqoAjAq4EelgBAH2ds8Whfz4IEeYED2G+4nC
qfIJ/gGUwCCCutD7YnitoaJKVYXTKsXpCh6slwoSfLgKrE8qXtXpHY8uFlEyjd2BcMzNbFKCJFHw
nM4LdGoC5YTi+lbci3vJGxUbJq2A93AXyJ7jWMHy4Hl6lb5fIQ6BYGCKRT5iOownpiBx3WogrmvQ
ZgvAhlq9TKTxUhAOM9XjVnC68mgcbubMatBLC21dPq1rnwHRYgdNf9Oo/vkCbqrYHS+0e0xKYbz/
NXlEl3tuTB/OpNccgI0KCTAdgzSUXrAGvKM+S3JnSkDtHfBNFXx1T1rq5PShAHTww5FHLjpoPkW2
/UhgP90jKHy4wGQv5eNw3oJrUow6tb27qjSaIcCdCYbzeb1xndET+uavH89CPkPtm+zHsHrQUYwv
GCpYEU4zt1C4IDIiPd7ZMh+Nsd5Kch8pdHZPnzAVBVf/AcocIrGBLY90BDKnYv/ww2OFGSpoBTDT
O/eDN04G+VAwUf6ybx/UGuUmHeODZ4SqYUmk+sQ4tzTcsAnEllmoIFHxF6fkgHkhrxjJr9DToU3G
LoJn23MxqqZgDpDWsTLZMQt27LeeYYNwCE/rTAPdvmuIKUbXZ9aZEK2DmNZKlzcXEMN8kR9i3zA8
dsX7ynI2yfS5ivq3bNkN/K27az6ZwHYTa/BtE2WiIQpgOL6TRM8CGSxEj4QjqDD/s7fO4TqsJHEs
Em5Uoafk9Z4huZdAbBqINryugeFF+jXo69E9F8actpJFZR2xjy5pAF/dUT/voz5l4N5OCNDPXgk9
F9zJ9SFFyjjkD2aLUWoi61nwQ70t8tUL2Iq5UVXiW2LjLSgsiZDUup1i8ZYwFvGZtbP+uOhh5db4
i+7fh1BsCES/9sM8CvOWYF5bKVbnobzxP8POxzxB15RtY7J+3MvDhXGms/6viJ2ZqH5jX9l74KGb
v2gl3U6f1vrsRJxpR8b9Va943/yd3FYMfMi1OHhq5ZGHzbe1N/9ebTyhJa2+b28vVW+YYAdVppzg
V730KpnIA4y8I1EWL8nzb2F7Shyi8kLVrclEtnjOB2FVrXp7kl8Ty6uXB9mQwvjz1bWrbGH78FgA
GgwzHo3mkqVSRMd2L3euTOx7cln8rVYaDkglERLxlMl+SXWfAL9V2qzJBDIkEFsnogbUpa6GyBAq
tFvjbjLLeGCK4G4NIjs/iqwHp9RcWu2E4P/WhC/iy+R8GkvftIkHEI0GmjPDeOH9F9zTxerTDsFt
8ZueUXRpF/jnGKU5E9143W7PvhGMmgtGGOja00ZkHSst5nSN3a6ACwQu2a0gH34kGf6XgeXjU+ko
3AuSjhvUxn0ua1Tm9vbxgIOG5e8h86ylQdqPr8M1A8KIaVXxCJ0K6stcroJ/JyyAkCvcKk1MiNxG
1hkt/dnhTT+xNnte+c+i3gJCujD+Yszv5zIfEI05jg3u+pu16dIPW9qEUKMJ9mAF1fKDbMbdwm5y
NHXpYCMi7G8GqyMoj99f+jMwtgRA5p4WfU3RXXsznYitD+eH7SJz48vhKyRzCQUBEia/ZjWKO4Ay
h30xY0nTeoM/dAYCzak6sDKtf23WAJpt/VUxRDrQWDSr7fJWJe6RJvTVzXNB0QwtuMbRSoQhuY/D
PiyCTAN6R+pCTB2IboMZUaxA70gXRqh2V+PI3HmHk/1m5FCK1nmDJFmpUO3fFYLJ56SmzKOVwdOa
9xbd3/+0QmbNFoeMyDzHhev0A8GM5AeqdhV23tSy2IwCZtqDiveb9MTSX0vbiBAEt6I4Y+1zf+ed
y5hguh1Izfgavdp7gyp2+GTj6/pRbfTLllKc5k8ukHKmHoDt6t2Ii+i00kSOl+vYCbUc6rsZliEA
GwfbCnPoEloT2ULXSE3VLo48BrMZFScUzt/dXUJMV9naDmPbScxX07GQtt3NDwUO/Aj3+Gmcfjrj
bdYhLsYimhlPZGK2D2szMzJ6qHpQYbFk8eojjX81b7RXnV9iA89UAUt+G48o+xRuszvQ+WPChdTz
+UUBwOqH2kKZ75syjKSRreF2mzTbromIB2nrXKwmwQXdOdVo31eI633+he3Rs2DCAIQWwtbghzjl
LlGYXLYbkT2yFR8pHQb/P5COaOfQ2VYmGvALWZSckxcn8bzgg62UyEpNeUiTmgqEVFGsgE1oDVxs
5pvK8tUfpnVGTnJlqQwDbS/lACc7mrF3YY/CBy53+i4a0OzpwMX99RlWDb7xIISXrxG+77sCrxCX
R3+XQkKvqipG9+hN0RrGoZDF43O+fwiJKTXSoOlahNhtNN/+Yv0FhfCQSuBJNFDOiQdcU98TJtqe
6tV5kovcmDXgMatNpxvcxzsGhWEzWJUApHxtTgoUlPhrsNUfI0bTz6DH2Jj/LwswMliCs4ySJkao
fXZ8KK4VwLW3EAqDRVduY8Eexfi2Jn9brjfl3sTZLO3LmVKPNIgzFIhPXA42zCSOXHBm8QlRrzy7
SbdI+XpLagLTOcITICGxfXetBwU6zakh7jzKPzC99qmkUymwGfxxZlWBa3BgdCOcDwyH/WEIUs3o
MK/5UXbTG11Rd+GLpJ+X1a0FEbyEDYEzhDrxq3aniEaI7ydQR0QVuPjpa8r6w5xjii2M0FeqEJ1I
TDvcmCeEGAhNjdLXb2kIL/WDidRcBrthSWugfBPZZiNFLyzdSr4tnIbEywSu7BRuYJShySawgKwe
zhEIPbcdajSAQXeO4769STGalBQ+kgKO4No8GQ4Iql57Skqtdb/ZMFX8vog0/Kwg5vyV1AokKHGO
Vx8Gh5kLM3l6mft4gdxz1Gd5kscnsX/fMhgkJbJSzrUioc491NdYS3+uJFgUzUyV9IHqTsmfJkUG
Qq185+1nHDCdxBpVG+VW9z2BTV3EvhQsYbkjwBXqwZVUgseorwDMoH8eBaHSWehcLKZFf9QHB9HW
8B6X6Z91Q58Tk6NOsiR5meyAvjhOhf4S1nS7ePGNiN7lWLBgBV8O1kgAxBE4FxBgWmT6s8/qmpy4
APP+ldqB+E5Aq3ayrYpopzkytfKPqYn0RWknzodlJEAaiaZV5ET6x8uyGrRb6cdA1lYXZIki56ey
oNi+YMuGJNfhf6OxuetskbM9u1SOOmQn/PAP3j1vs10ZWogz+5/9DHAmK2zT82TsQYsU6Jq7EScG
jglW5CUBorrbbt4pGmHYkZetmTskgWFqyCwto/M4Ny08AEJ8vBAhm28S8/85wOTf87+ZqwW1/7ZQ
efz2TceVMHhyHqZqHz+S37IdBA8g3JtduaRftTOckts5pgQoHRwWuW0CBX+wdPa4x7kfR1AzdMfD
vuXAdmDZmD2zMkusg9tF0pkt7yFEMe6ZhqqR44s2pSRdoAvRZ8gri2bFSpZ05bkoIbIcYF45JGx6
0rmu+VYSKXOO06jCv+yp42Ql9zaOcjMcqOtT3sEkLZVN+n1+nlovEusMSmGW1Nojv60rRSkoLnUz
4OaVtJgpBr91OVk7vTpUXOoQNGHMFffORCZWZ3r0Jp0vhm6+7q/PhgdYJUb3wYs5Jy6FJJVrzD5G
vggoaVN3mye1iSqtSk+pBU2eNITcwrq+Kfepvc+K3K3NM12pzryQkrQX4opYghARkAVa8FRJVgEI
xTY1U9e7SGdQ+YtK9Tn+NqnKBYGWH//XEzWaZJ65juAtDGTS2clP1K9kW4sKRZfNK0ToKYVdm2rF
tlrQRsmaRD4DtRf/4O8VlE/AzfQQUQDpV2/z+AnVO8GyL/IGDFGb/uxUDren9qrS4uR/ZcpXZkf1
WzMoX5Gn+OsRWQSObQps8Bej6WqFfluJvxxra3yMMDzqOsNo9N1MYnAA90msyRThXdXkWbSUzJyz
KCw8JbmwTjVTu0JDZ79E6ND/S14HH72KM+LsfHCKWsun7zQH2ohxS4xbxi0IOKQfNgbUiKG6vqN/
H84uxoqgJxqt/bBjNtbECeBnfr+lk1jEkKbE/0dfXXkh0CgpvnJV//E/TRskiVvSetGHTEihZQHG
3NstxJSYcWG7XIs7gb2xKHP9g+RLZuZfGC8WgaYpf1Yfa36ZeG+4Kdo/BzzPUc/hPFRGFISM0YbI
n2XgksVWuZa5FeW81XJQkUa6RvmnzevOUR0K8WF4h5tn40S5bSeqOwawZFPLzfE1qgZnc/3qvxO9
waXurNpC7VwZqrNabTpCClseFKJgJ9wsHSPgwmsznVneC4gqox34S7/5RuwOWsAuaur4EJKTx7oC
ZEjV5hOWDILF6EvBDMJoQBBuDioBgaN3Ij4AqWkkjSfhb781ceRbsb+F5kZxbGL4cDTh4/C8OBj2
eUL6zFwPPAV7gKOtUWufCfrE/76ImupNBJ4oPzHD7ePNtCgZo3b98sq4SpMHzWy5j0c21ld9zg8s
H98IaCWOux9+nklWnHEb1Ke3u883n7gy7x991mRZuC1/LSM0+QpdyAxEtoHCPpe0gbaoVrP9uAjH
AUoZQxn1WvwcTJfZsZ2jd6VGGsFfVC76727zHH0O3hsKcUfPF4QP1KTxhr1mI09NJwJfIFbtoFYs
ul0zeihXXlz9AjqAxzrvSM4apDmmOxS/Q7nzltK1PI3qyWNgsTSil9FqvdRpsuqlBmpPDNbCoadE
VDYu4m2hOk1r7d0lb2x9srmhrWl/KQR3Cyhl6tp/1LouG0Q3eZQNTAmzNoDw/xJstpP93F68PPs5
i8nwmsWsUe6qhINhH/8HLKvUTfcwMEVUpOA22GqndJ/RVXnlIIBj4TYcwAre94c87BzAPOIsqcHI
xgA5+DP3AGPaDYlqyZCB79UIg/hjeXfbbTHPfWzhTjUE28Mz80PccXUOaHKOs2KzXLNJGNIgkE/i
ljDI7Oq30sxavAFUYWLgXxce2IDX9npdfu73F4uC7Opt2zJwlx+yCWfwvs2ZddIaOb2/RGpC3+EX
jHGxG3umiiaJLrM88XakL5SxhGRRLn6zix20P1scIRpRPu7vNYy9ITehL1QWyTQHuGpNIhZ3ne3T
FdWe6BUIpkamXtc+TLZn6ItmSdH51ogTrwg6MSlPQaL7UYN5Z9z3HY0xWjgGi+fcM9fK3XBUv4OM
39Y8qA6BwpSzpHygLe5hp1lkDUt2IKUD/Z/t87OFbj2uia47dwM4hd36fnqjUe6fNAUEYq31GyQ0
fmXwOOjtIpAtUYRN+E9SMmI62Js98DPrqBQ0Z5deffjBchBRVZgYAWfLYI5qmwajT4XlrHD+jYAj
jbEb30sDOLxmLfo+q3RpEY6SggurPuocB6ioNZEyXal4VC7J/Nx+wrfVHoYC93bPrsX4TrlmxvOA
NpeffeZ4AVmp75xWV4+KtV1us/v7vcofeMaiTY7X+GHOnjIYnDX3k2vJLrrflFA1iorg6+493h3G
gdkMiEi9zadkEf7zl2vna2YE/NAXdARpNXZQALaLwrnS6fe3kvroQEHQzFFqV4VYJbEWY5dsYN7U
7wOw4mpNc/Yj25eQnOcFYV1Yz0ncJJoEyXKP4whLb90KsGCY6pIVx2sI5gFaE/yPIe8a9y+XkIwo
9XxEiGPKv/Oxj49JsXHzXxri8YQnY27BempshWRLJZBE54b8FqSY9ESrvBSWIZNDu7roaZNHaP0J
2LWj7Nsd4Rg7n1Iyu4c+CH+WDF2XvJ32b7o/fcyXESirmRjMlTlPJfFFwfFXpUS8KDVmoakLnwwv
4aSu3e4WmQNIShvqxLhOxTD+E9OS4FrU1gaowsnMeuxqQL2hYR49JlViP3lMPNmlCypVT5IwSEVk
JGsMmnh5ZrUdqVBaNIU1ZNRIoRwJcarIyC0MV78zMa2crFFYnfYKO9PH+MFLKT/4hxihWiaJVWjj
H9zBfMibPT7z6rPwKGMDhBXsBx1h6USBA4Kv9aBYT/qqjV2wiltZ4BlW01mwhm+ZS9Mfb5JB6Gd1
BCZn2JGFqAdRnW72J2e5k3muVW7ShCn7LIabFO7mGj/bWmAt5+4SPEXnSwJDFb9SPRKO/1WnP3J/
oK0VIwnKYKovvArM/Lo8ZOcLr2scMLlcYmrtLeSAjw6rUFIjnRUqjfX/YcRDuyTaPtPvEC/HD+BO
URGJ9o1whNsyn8nyL83hg2MJChXPCa2Z4AGcXj7RaaVwnLYuIT+1PrDkVGh6vU6HF83WCJVlspLn
ghh7Zy6TMwQHQ34VH2r3E3J/hbJDj06lSAHNO1RpKOQG49bFtt2+qge12PYAZg99mLL+wuq7eEBS
8Q+23c42w4IUjvUV7H1s6eNu1ruedLhQ/eHmr2ukPCf8/k/A8TGcpTNcK/B7vb224twZk8UQ8vHh
A5GsXH4ks9Y1QOmuXS6OR2VWQW536TDY6100JfVAOudIYjCNRqvTMwbEDABsbcnYpxqvSr1S+YPW
Q37NBimPdzo83XTDy2haaLw/NGEoML2BeSqyWCy5+DfL+Js3B1iY+J3vZWq4SIM6SmTtKApNLffv
9h21eYG96STVuH9VW2+1BA5Cy45Kew5sZIOqtKjoEBNthXQDXYgcVho/7qDicT2vGRj92CaM+wvd
ww48yC7nx9G7srBJn/n3PJ9JkBqrWebbHcXNUdpOy45Q2oKnrOP+X9+piEpq+0GJTdPhkdmbrpG0
h4AxjICPp05kCZstj3q783G3gH7YQqcDIv8GTFwIcHd6M8g3yi/nLcn0Nt8702GCWNPKZEB2Zx+W
PjmZuYoS0FY/V73SBsW4mq7wqESozf8eg7OFjeMjLG//vdf3nYu8zfXYH9fb4O+4CrAAD0i+FJrZ
bC4eQgWEi9aBVzZhNRP0bClrw0ZLV0VArTKibOAMpWALPKV9f1Qwr1Bng2NY0o3ySqkzVrszilGO
dU6B/9tL8Sgn6hQcFGQBbUJod9tsHYYYXoGFGU0lIfccFOQDHgbFwrri6UUznDbFnKEVWjPD2Pwn
HRxY7WnpxYXlx7KzVSTAQepO/qGwflver6gavsicFUEjiD1oKYgOT2z1vFCeQHlz+8FmUOPMhB8g
VGflMd8aNykypBCGy2y0qLfT5J2Jl8LeMK3Txt4WX+F9k7DXQFHwgwF8q2QpJYkjI6zLA9PHgnKD
8aNHRJGojJZlxLOwEMjWsi78Vv9LogjiOiiNnMzHZdmB/fJfjSVjD6gd4V0gC/BeKxzPq2FGrLD5
i66einlgXdDPMidH2MPABRuQYyvLK7XtQTz0GNIoyoFnLiKQjm8w8YLIVHPh/Tsen4RL5N3LTuhQ
DtwUsUXyPpEkUAjMRl+ZIwZ/6zz0W/1F1yUN99a00LwwKUvMg+LR4sZtVcY0kExMhgwJasV1Ok1k
4w1duUeDB871hoCquyAhQz76ycleqkEgR5ssHyM9J1x5AtEwgSYP5YxXXquVXDVBCzlzZEv4PVCm
NSqKygb4xBCtMaF2FTQEzG7+6iQpLpjscQ2Dj95AslzmmXi9CxMvQUJSStFWbQ1hoHZl3GIZ/upY
v+iuB2Xwfkbna9ELH/m0cCx+XEd7CXawNbp06Oo3twjeC79JAabRCshjO6IYsJdLuWyv3kjeOaMs
J8e+ONiYRGjJiEyP8MrUlPJFLA/hgGGiOTlYcvjHOn7pSRx8/2dzmz+qjCtEQUIrFB7zBsXOCr9s
I+8KyqceIEAjbBEtaWN/KgN5Yzn3/P2W+q4qG9g+tH60rLks/UkIivlv8h7/wmo2lN18yo0sonPk
SzGUfx95HctLk6olFLOUvuh12jrosVT04vn0Fke47VY9eN6O2s7crLKYuXSAfE9drrG4ejYMeNJm
3VuvNl8rhGjHD9Kuv/zZgUO8BinVDYj3wi4Vy08Hi6MMUYsIdrFe8HG438ICaCEnAk/U6L7icYnJ
9fgmYDDqgOsqq3hSrpvVEK0Mch9deMuUsImzPWRJsVsUAHRsurnPY2s5rpSdPRsZLWZe0VPCRqsP
zvV/RxZIKvngdExsePrrp4DH4FcQYaHO3WHu3XhVJx6eMByJ+6WOJ9LPrjSYqSivNvIxlf5S69FA
AtWvySgT5dk8vvgTYx9j+En9rKbj9kcUi94Jo617mN/w8K/35/WU5DKB0cVs+nX4lbNvkHKMcpKy
gN27e6cuY7zLCt4VaPAQPyKr75LoJDlsYIrskgUvGCArwB5vcqmbDQxIB61ndBWK5PZv+jd0t6ti
CCjQ7GgZsLHp3deOXIgogVSM2OEoEpm6RqkQ2cvRw+2pFEfhWALg57PETYFYEJURLQLeg60LIijU
vL/XWUPNmriqK5I5ljYMZ6Xn2MbX3QohIXuGJ64NG/ogehooX3azICRDx81pd2FHmIVtD7jwk49s
hpezxC0OF3JT82aZ1llPWk3EMjErnakFrXatZQjHhs3piLv1tWI7EwYA3mkmVgRVybNxu2SW/3p8
8MYxADkCUt7ArOFtcVck1t69qVZkaGByn5YgeuD5ECYbRorEGNXaD9f2uukVw91IacVRl+ufNf7p
lAsNBgenPyolMgChq/FgrIw8TUSgSQL57phi67eSkfgNOka2sT3s4PUMi5Tvn7eGRCNFcCbiM/uG
/KEyTT+CUdc4ylwURQpd0cC3MP24LdoCVLYY1q7vULVtiTvmYFfQxBJTRoE/OHED5Dt5kat4+L31
U4BYFEz+93Bf8dTEshPGQdCBo9v52wS6z0tlTT4kzohksak7ZWur+cyP7L9127b7HznqoVNFA9fs
CZx+JbcU/tZMjvl5t/GZ9rO/rO0i/a+Aq8K4Agf+4nfCW9C5/2MK1+r61QLWmJ0FGWrRnlFxxPrA
imph0TPlZbisDNzde/BfxAfO7fAeHEe18hYAa7w+QAVNbbUGbIQV4D0Fhcncr1a3gzAzAP7SiujK
Jj8kIrPSYdFTdb7l1rsZ0sy661vA3iS88upWK9vHDpzr8v0938QCC+QOKa460PNbIUAXdYqiuspJ
HLIsLA66X98geLeTOR4PgNyVaLvQAfbzzb2LeTIfH3JZWRQcKYYNeQ6jM8U27QS9MyxVY6tJXISB
7p6PSr5/jNGMvwiBBL0/7y1zITfA6bywI2wOogL16uT2gOPm7X4gyQGuBq3mBZkecHSO7mCfTQ4v
cjQ2lkR8Q95636Rf4rjuHtqwVYGGfbIJ5DOnR6BJxIlwSLmzhGto3RZSunZiHHgIyvgh0K7a0M7y
ehVnMKNPi0XfjA7HNVrnVx8Me3RIx/8o6YgUfmxlx8Bz9X25/B2l6C/XBXUQgHKBpbJqvgWF1nMx
fUvXdpr5H2ubNfVqaVQHzTfRQZQt7lH9AQ+n2YrF4a65+IaGAbQLfGEGE0EOFFc9bm4LkU9l9+8r
SCfOyZAdrISbeGf94K5q7aURYTVkQpF9CPQwaWuz4zRwxFgOeshV2T1MXpoHqNduQZqYXFAyLsEo
w3IeTmuIdnj870vMzRX+BuS8yTdW5S4BI+sOdSKoNmGnTQuoU9MG1ZZRWvh+GXMWN4gbm/beavS0
awM2L1A6DMI+diY7LiwBsoY2rFnVIZrRTEJ04jyAQLE5jFHf4KL3bEzUodrEHihszGPduQ29pGVc
GryPz+nDqcq5nfezopZq2qzSfFZ21J8FDKenjNesxbb/wQszMNUvU11HI7NOPwljYmlD7nfLOZaN
VnrUN2IjECU/7uWmsNXBY3sh/k7moc76vDSaPDuRTbjc4+7eCjKmNhW701o6Aq0A3SSjwCU3NSAB
+dqIkAeUTLw7CGbgsYSExMkBTRl5UxIDh1odlWb/Y4sznFDsA3OZS8e/VV1DFFPss+7j7Z5PnWnm
KJfe6uay+awciOPiZA49SCF2Awl58MJ8jUXsj75+wK0mysh5MeXu+mF1QJ93/antjmKvO4Bjd2Ar
YAlvuIy4mmjOoNrRxDd4bUKGMTTIH8JQaIEwSoHzZDSrHDZFRuOmHYnW/uHVCDmrRcCVrXMyTgUL
FfsiQCbJm0Z7m2AYRTev84kRWKw+N4zXDApJ5VNlVA3oowt+Dq2FrQPP7ipXtr+7n9Bj9m+Pch7g
Okl5/oc+0r35olN2c/beUgQd0Vmy4PrQ0mvQzygoJtpvmGLauSn6qy5+py8qM6wXUQszlEYCGq9p
dIjzFaWL/mYZcjPSZUNjqvHguPe2+hamKbCYmRa1mK+AloKa9IGXkopTXQk2L9WQ69ZuEVp9fHed
8UeFHY8puMk2ACGwE6IqY9wCKfUgQRb2HtZVlR90o/J3UUEQI9wWLixPqdwQQhKSNruTbvdQj9Ei
sAMMKSX6V1hwoMgwHhiiwQyM2b2mdoYriZQUL5SvTF22GGyWh+LPoq+qmBS+QljtURRmBcUBxZbb
xQiDjViW6K2dcU51fQH+ntiZ8R6+HXJEW56U9Gs5vT61KHUZ+AFeVMS9q0kQD70CVorqJFxp+vCF
StAqQxXYLt8+RvSqJJwuyIGb09pJdc6WfRuHyjfknQwd5/isCtHpf5Ll7zLjg2tMdgEBx6Kk55yL
1a9k03hef3NKHs51qGgVw/4M3hPd3hlBGDhLqTAcOB0HoLtK9gAnrWGY2LUnDoydTnVZgRmp2t+2
kK1u9Vq5IQ5gLtE48xN9eQbo1LAomMhdqzf/GWhtQxwyLROKLPCuuuMaDWYWLjuISp24MCsVUyRd
himY1wZ+zezFxj021qXoEyVBty86nGha0+np5uybjiCApaceTKGJpmyH8N+CjnB+82KqH0Y+441c
S2zH8d7+jdVMxnOsBab45FeVwpkqIAclvKiWXFYDeznbVIwfx9w5Mn2j55xNNSBoFcBb1F6nX1Tc
Bg0cyQCEps2aupv4f/bRePzdPKzHiCDoyAWOA6a8f19GOWd4EC+NPngT5zfMKF9IcqRMr98fj9N1
g/1SPXhxlJcP7rfiCckDnqB55bMEDNHGUaFpVzebK8Ym6l0xK3m4/BoNim1k2fGh4aOLcX2BycX8
xdtZQMOUv+5Kz2ejh6Y6jMJZefCFmXMihqUWI3MoBuIoIriJPSlHOldwgsQeKrp7+ebehDP/spaS
dHGyhfIizJHuut73Cfwea7I34axOfunfMBkYC6OUBxK+jJIsENf3D4m9Y1hZsQhWzG8yKaZ+V7jl
UFnb42W70fMT3Efxpk1TMI1t8GL8SEfu6zU6R4jiYN3XBDnxcapWBDWVLGdGhKvEs4lOpLa39vaQ
XE7kL0Gm0HsldMEJVBOHpJL9QlfegGm94gazv332uP0vsQVabxQcWx9S1fG496osGHjGn0E7f8e/
K50AKQH5ONJ27qfywpHwgBl1g8mDoHZ+nnvtpS//SfxEREL8OmM4/83psIJsBREOsrds/r7M2bX6
R7lnEWw0s3HSl3zBc3yZrb9gL40zoL2utuBEbOvefDV0IfaX1lYbzQhcjztFUWCVLJjKinbm5Sv0
KxNgdKLLFK+e1PPzVlwsk9UgFPNMwiO4SJmFzJAfZpoyC3DtJQeA+UcWfggJDnBppZgV3NaNdhAF
KYpNTTlqYl+MyRjWC5Q738lqDhTmpekezECLpAFNorpFRX0X2da3/nLvI989jNB9MX2GCAh85U6K
NdjQKA/OzjIcDY/Yd2qO/NYKVYQq2qypZpBS/xPAUvrqpoUXINYaDH8YGHtf2EDLhBGAHeYXzFFJ
8Xotqmuh8exYJRfEPJOQyGaA/MOI85hZE/+O+974X3C8oR+f2zOgVlkOi/5ZgesGTilJecODWbPi
jBK3VSQbVnNjI53qqy/Wfz0ZeHU+Gt8wtIc1jvlgoiVwYgnfpmASquu7nSNkfRt1iILvoMwEJxgs
gjofAfR0adzlRstdV9dJWlLGZ93Qyt79cLJ4EaTpq8gkTKCQb+/VO/rOESimB2aZZJWQrpotbt5w
sEydFuwTsw8QI0V1HNTD4AdnLhJSt89h+jO0D0U0LO8bxHo/vHnFrTi0RZFQibW87fHdhUev81+h
/q2sQoYHI/r1mUbfba6+W3NyV91tEk8UwL7gOk+qk6CNBKC431EaWNlW7S5gZI5ELQhzamV5hcCB
4M/QslYE/NyNOobgicnZtvUehmLUoBmjYoTm50h/5m3rTw+alTYZxsOrDBQONxvI8pWb8LnoY6Qb
jSaIvWEIS5EpSclspMSOnsoe+SwsML/igSIM0bbrOicXlk/2yBBkkmh5w3njmU+0v3UJ7zDiy9HD
alsuO/R83Xkj9QCmMz7Vxb69dBGHL3WoSYu8BSWLlxJzVikRPUYDU5HihiTi0JAYYmtS6QhViMCx
erWzZDSFFj+GtVTIOC6QXu/VrDy5TK1xY9YggPZWUH0DWBWcfP1Lj7Y5wz/POVbLIlvX0Dpdy27C
z990Q7BZwaOvd3pk7BAJsCoZp9X7D1XouSYcWoJACzH6p8pVl1zdbeJupxq+iE9AmpEeqJ1097TK
k5/r6TkWrNr8ls5LH+dyl4gdRNDYoWtjjSoDNL9+nk6LWi8zj7Ht2UGB+J/QrLIFzUw6CIQCWmCZ
PA6Lx/ck/I/CMrjC89piSQ/sQefCYlW/vJhAnAphjbqm/eeRSK4t/smvSp+8suRcQ4L4B1tOwb13
0rI2zTSEEBzPC4IZVbsNBRp16uH5hhRzraLxoDy/0Q4qJlDJ/VM48qGWT9cJaB5pMrW2WfKz/HFJ
JjgnK11MHLt7tPLPtU6ArBQRRF6dPcToyWvx/c/j/CdhZMhqt0+/iU8hLDY5Wno9Bk+4rgA2LjR8
qHluKaoEOR0NQvAQGDcEWNVFMSQ33dCvuqnIxjVANnjsWnzbyp+BWL5PtpYm0hmGz8LaFO4Ftrs+
hWJ0CFsNQBe5OesV5AtRu8u40KyCkgbhX2X+c6DiibggB1Fn2ewaw+5NvSuPK64PSk/cU9kFElB9
HKup344pB/xHJqgEPjjl9IZp+9+zB5l8fa3NurjeJe/87gXQsm02fGb5qeK8NzU7rKBVXZCrAzrH
KYBtYbZITCMoc2Y5k52MgSWOgLKW4j1VCjs8jBUjWqFm8qnn3k4zgEVNtt4IafCDjMBSzL3mHOLv
SgP1q8dKXbv6dy4ZC7i00+xRRE4yk1ZKivdNojHKgtqfpvvvkqxT/nrwOvBt5JLK1JSBENuDumQ0
YrSzP5xbWtsHVJSVDD96wuHtkjmNZBRH0vbXx1RwCe+ktSfpGrvKv4eTDVR78OMKdpnzLSNUERT9
cWxBj/2/5FVJ+a7WKKJIadP38ycPE9tEomOxMZgh7DwvUw9wOU06Q4vSj8fg10WNywzlGc03iuSd
oHy0pgTa5g01eUu9UR+sBBCnp1L+FXI8KRynbpVm15D6Yxpxk5UEEGmO/HOWZN4Qn4HA55Ru4cKu
rYEGbY4zTYU7gkckbi+civS/Hd3oQM5382f5crkwClH30D70q55v7iu0lQK/t/uLDsQHMg83vEeP
W1z8c7JT0+5YSFS8xj7eIjXf7pZW0fky2KHj59teerJq7cOh35+W9QKslAg8YAzHEQ2KxqRGlUCr
SqspJP3KSR7TTCVr2LIYr/1KlalLqEW6aEuLwdvarwddXlkKyXpZrQMnd/b/MxXCqI3lCMTXdUO5
VPswQEwiCDwn9r3GseqjAsdsJwhOnIKWCBVRnkkujaaszgSfLlsdoMUWeMeFfBqkq0MoTaOPK8jF
C9UNrGauR+IPOaK0n5KjOjcFOOgQuVOTLwB+t4hHUcTAVlReqP/UnuYWz+cWQyRgiNIlsGoI1GJT
cVC7fCcXQUz4g1D6LqQrsqAJJ98SgGJGd97LuMmF6jaK29u4Xn5IpHRcAde5mT3U8YOWWQJp1goU
cjKN1+oiLNXPSvB26N1fDsQJdTRB88r+WOeMz/ZI3AbyHPeHXU+dvnSIHI69VC6LMVrYLZzMFhf1
bCKqPmtq3P2cZI4M5eqdP0+6fpCkP1vafi24m4mEm+y7MXJTVM19/JVG7Fj87T6FM1+j4vwjJ7Jw
6PhMVl1oYquIWgbB/cMLi/sVbtAuXRBy5pns+6A7ytMQlRzyRnbmoorGlKgEFZo1jmaRH1t75Ynx
Qe+gMeR7D32nBSgC7hbovW1s6OL+Vr5/NMy9ZM6LQ9Pdsd/y6Rd+jNpNrGYW0BPIWJZipOU+HxW8
Bz+HMRz7jpFwIOCKXyj1sF1Dd2Wt0s1qiv/jVfl/i46wXeVWkow6bzyB4ZWBv/LDpkFEaYXP6LHl
qd8held7CrLYQcv4R4Vy+kJvoIhdtQz/2KZr/Z5/3Ag+u1kpmic4nHCqbO35ToXcnX9SxOxofe9B
1IF0JpFTWGXk5yG9oBmfuhr6LWp4KhVD+gdcb8el1R8fatITE+Ei9AO/26c0jz/Mns4GY7LK52AH
myINXj5YA0UmpuveyIbQ7i6I88OrAbxfPsCYrymA9SmzP4GTm1UXd1Y1nx9Iqbi4CwayXTB0h68W
aIUGS6CIUwqjff2N0iA0G6tcawDvf3ECLYDzg1q0TT+c93RYK53TcrNYoCf0foKISZiqHKcXSaOY
mvkv9YWXpCJkDZHK1msq0Ek3n5qPU7i+Jp/sdlTV0tXWm1nncivR5+90u9KLtD0Cuk1mbBG+k0RC
aAhyPjWp7duuGdWP3avgr7CHOwND7XZxnbKnsTXMuy9WIkUZVeHO0Fm3+sYPNAo3Xpanihp0sjA/
BH6xZ+dnBRN40TmY7WCFLVy2HMUl+BFkXPVgEbZPf0TQnOtzJjBMUgS5X9TRYOgCew99k8P6hHUB
yH99Gy2MZ+6O7sAW46POIb+Haa4i4YrGus75YgUSImSj65rlxoqWOR6Hw6UHRj+1sKeZMdcDON/O
Q2g32Y7afKZ9MY7JGHUJ/mhYOowQ3hWtbH1zbgykNBT/h9mL3Q2661QRLYEWs9AEDxcVmEfuPy+B
27GAZ5bz7XgWwIf2A457Y0/cJiNKSS22MTfVIDchwH57oBxexqliaw0BpizrS72ve8mCwy4Qg7ee
svflv8cMPf1KOLYq08lph+lc3676+5UU0uNT3mUQWT2eGo2jkofaRdtTEAMEXdSEQDRg19d/Avpq
qW/1e9piCrPgy06zT6HpiPp4dvzMbkL++Zy1nNdSy3RXD54Zz5BzXNZ7lbFMy5JNbTGqg/vHLJeU
Y72SEe0kqBFyAyLgWYcQ/hH/yB6O587r4VIxBE6bZ2hxqWiibneTBfQpTnbZBlpsk1tEQmLgHjqT
6ahnWKoVHQ0LT2A+rnFB788lj8WTByCAWUWt/R0WSfwpNW9jWPwEVKGMyxyQQMPM6+S1ynHhTa8n
3YzbPqJ8EplKhxLbgOe3vmMJ9qyRXAehttFxDverELcRE0C07Qcz2PSziucIMaKEcpkEv9fAok/w
FErOM70yrDWJNrCBr5JYN+pwVGTFsXBHkhx1L9gFZAi+IA4+0i8imYDEyF2GOiO3TzONPr2GqUKu
DvNsLKXqgSMq+XAc2YXNsfVYG8LCrm1n9hiFftr94GGaHRIhKZ0L185dkKgWEMgD74KNBaKlPkwM
PyXV9Xp/sJk3ZzxND/3xCTbLDtPNJwLe+JbnPx/xh+Oaksu7JRkldAd+ie3W2+pfiZObkIO1Hf3x
379MChqheh3KrT94OIdUY4yTUGUHLS1bATq5u8j7UYjM+vJ806nsn9d99SdDjqU3c/2rX2zq+ziY
QuyRfNC/9B+iEfdkanoFDf7l4lPn/znkl65zYiY9x8v0NcGx+FX7GY3Oy6t/KhIF6CzbWXLy4r5V
4pQWp5hrRre9U6MC2XgxmYkb11K9yaOkd6XXpBdzCwupPWAGCp2mfqD8B+oaH8c1Sp1r1m+FTCaf
tHy/OtOWDIzsA9FsECB+trEtv6w7YnsVbOM5JQccZOs4tMqqd8gmBcApDd2tFoVYp9XUPqdhB9aK
OuDm8O0lrWFnjBOPhbzFbqb9nGR0fVVf7iijNhF9v76E9Pj52ok67BRPnfzDk3cs2yBSNRcs7FDW
o61vcI2FUOoFOoxd5Pu75PBokH50+UulW0/xG2IdgkQEzx/gE9Podi1BDd7M7GQV55nZu0ZZcT12
rm2Bcyq76A1tlVsHdMhF3hQQP2N0E8bGpAZWELyGZhLvNG5E4Gdowtejm/q4cZXzGuNVBPn67W2C
HngEcizkDThtmK8f/HXOBo79m5mV+PQz8/o2/X16IFSAclkZPdTMdU2i+YvxwnbKPfzyh3FtNp+5
QXlmcHqkXmYU1HTjQkHS7nVSksxNAXiMkzDIoScoLxUeOcR19gXkGlohm1J/hyeV5CzewKlh7tZg
+GBKwN9T6oUuuP/HmsiCPFWnR2PuJIblqB+swqZwZLQTZD2jbOnfIanYcRzuSYgzxl+ODDKP8X71
8G6BXwUjJheq7mk4izgs67Pra/+9wDScoWGYLwcKrUY8X+/BqjWfqKMz5cUs52lWzGxYVdvaKh9g
nSEXGG2q0d4x5y+Y0TEh5IHK/tFZYNuVd81hDT80BHuXAjiE3SDvkVUJX53Iwv1uqAf+UY2OsztI
gNGJoPIaNnEZnGFx17/Jsh7STVpEYXjFyoJitsKLRrD4Z0HvU20gXn9gNCCIXsqKriQ87pGXPmv5
nvdfZNvtMdHtSjhRbwpLWyNGkKpzJuGHiU/0NXJkEmdvEq+r6BKDLvnpoQuOz2+tDH8ld+7NNOr6
j+qnYlIirTCWUJ86N9QLCr2E9TC/rBRxISNMdpOVjQjhrBqTxjGDJFOcNiL5OPrL+p9rPU+NduSx
6oMW60FgyBtRDJKF0R5K/3VWXv9ZO4AQFdQRWQqP1pjiHLxt29b90nLrLvwQZpS5HFeizGrwcxo+
6HygVz1nMTvNLRY17dxeqZMkknlwMEfBNVkL0gspWitfZ/B7D7R1Nu+aEliBiOhyHUg3VfNIotAm
HdJhTd1hgF/tBvfEi6tESQOpo2GrPtH8IuAyXRxmqWaVnWlJFi8DORWUJJgjT4GCRZmU+guc8UUu
N9oaH/h/PAruIg7Nx8bbkJJh3jQC6x6BroS5AU5GruprQRIVti4VwhqgyEFV+ciQCtGlcB9n+9Gm
wxEnfla3LWcHZrzniRuYKkOEMRdOiKNok5ofHBlf+Hy89OaEhov4hb97pS2Tq5l9LshLRuxOUnwC
j7mTF4iXmZVphRfX7wmZEL2+hY7AwsyaguUpyXbn+KZW8jxuwyENbqjXepZFeD7snTJMGBZsY06v
Hn9lEQPmaRKEhicCMKadkc21TjWzgNNOP4F6QvPrp0+i8Y8hV37GJK3qcGi8VKVUtc73qiGlekGa
H4KcE7p9tcIHx5jvvEpWKyfynwQYsuLTRfHQazqYia6K60Z56PuyYIQ+vCEfLBcie877OrdadMwU
FswcZSGikDHACKCfu+lNZpqPTFtz3c3zh1a5y3HfWbbeV2H7n3VPGW+JBgwTdPH9aSI5c+4R+jYB
zV5+DXB5qXPJOncPrpciBL0PD6XFZDUgImEG9teA13pZddD0UbQGLHniAR0nDgXfgqOFsTIX5vEl
+kORE5bv6qWjr8zj5RmHga+AMsaRh072N7MOB5of7Umq2SisEDP+qWN+MHY0Wm7j3zSsgxiK5mes
/JrAg4lkINH6tuaDR1HJqbD7potLzUGD/+HW8UZRSY4RVPvwblNYu9iqb7zM15puNfmtSjfvHYAL
yIOwKBuHj5oDsCSbxjjyQ5bLmkD74JCl/3IfyD/nlU0yJGySgqfyyBbwaP+RKRvjpYw0Ua4QzA9X
xz9KL00bs/lhzvQ3RtBFNmMS/0OP6GtM0scFlcYpYTncD81RjJxQzIZDPVsePJaD9cAtkPcAuMGb
FTuN4/fzPcQPNCmDpdQkeSx6zOwu5eLuE1SN6LyFg+ZP77hEBUPofhtSXp01zkdjJWWtZ6VuxynE
oD6yLj5jM3RpKcngviuYR8HYNZs/MGIaahNEVNcqciu1epuXwObJn+2Sc75QSQln0xEgPR9aje1J
lSI2F81bN25XP2Rk9iaPnxypGNgZzGd23ISB5WC/3uvMk4qArXnt7scXgdt0+Ki5q6NK3QIQKOdB
zjtw0nWaroATcGdRfI/ugqxYhLig7HOwMdxBV5bSFQ0Gwth/39l+lzKQ6NWLymF+OaNkqNcKTsu2
ZeVFdcecnQJBuV8L1i82KHYZPtDkbbNdaCUfNlITMmxcj7GDf9udE98+Xgcuqnl7v1IBvPY4pmJI
0Fu0vB9rEzGNJwPz9eMkSAoO2JjafL1Np6Wtrjvf54SNwSyuRo4eVfMfpdmYiDpvdQFv6ypUDcZR
26ZqLCDyYQrSk0NLIzVpq0tEnk4M+jbm9k0FweeQA9hX0ewKwEw9ZPW25LbX4hLsnWb9xMUrArGl
82noTOJezknWjTU7tYEueWHZN3Z9HY7ZINx9lUq/2gsazlzA2gjs1+52ZkSVPuH9wS2RZEgVl1rP
0kzU7wYW+ZaaRbOJPu74xRWRyLu1d7wHng3Pd4OqDdmRNn9/s8vblR/O9FsHjIa1KEpF7BnoMHUj
zBych/5Bb7U6Go6ktGuBl5Yiak8MEFM/n7qZprGCz/AtVGKgElTSuKZ4tpYpKSYivlxNDjPaw+4Z
bDrmTTp6L3BZxio5PwFdfGeoY239sH58HuVrhQNLp2NWwIvve9sTWwiT9SOMb57uG9rlDffnTfdx
U/psbmiZB+zhRDyi00ouVXpNBzmJGjB4H4u/qayXuW0JkiBeV7FnPUJSRpNi80qFeKmSxkcka/OS
+5+DN8kXU9l8K6Umtab7hTDdP7PEjIRuDj27gLXKseX4hqxIX8kMYm+3rSNhzN30HT84Tm3savwe
wdQIOdXXshJ0DSMe7SO2z/9B8x5McJ+EzbizLdonuW36rmDfnSxC+/sHcN+vrGFInuCS+d+iZFKX
j7RzuVMODORx8Ebsda8A7Zr+pppdPK81EQicl3/LK9zKbQJKDVLQHYjuB6bmP1szZooFmZbg1hTr
vDXo3faWW30c5tAc6mPjkrc+xT5bZK5I04wGIodv8X4W8JFw/hdKLYMASvquJFosrk/12JvWTP+g
y0PFwBAq1ZANTk8508v0pnasVw9EC1U8exrJpo8RzdlQan6yisU9amyWGDz0sqsGLd2PQqUIFvDm
zRQ4PXQth2GFwzadK2Ex9oefRPbmHOsk+8Cy+lqB3sRr/r2uQH0lqx2W0qkQGY9uhWzwE+3wh8SP
xjNrgOhswTze8bMZ1QTBQqN1pxI1QWMxmCIHXV8mCkPg70Ya6h5905JG8/ZWxD9h5+Z3nxaQKoji
/GRXZd6+3pij6ooAHBcDVnOxOuLZLb8dkwy1uLm09eg9/RvmySgMyk1acse1HHpjZFWvCDih9CTw
ogcyDJwe6fVFDxBRZ1Znld/DbCETJzi6YdyaeZjy7W9u5hPQNaOG3eb/p+hF8C39ceut1pZSywyf
uFbstuiF/2CK8JQMF7LcBUDDrnMuWbkIF4Lg79vbS10h+HbhXxiJTD+mrj5ZdnemA+K5hUYlm68R
shVXkFK/dHAo1ZSp1AECqQEM3N115Y9Ogcq6r9wOsk/18BRSJiElZtFBriN0P4K/rjEqpCujoU3U
sUpoa1eRBY23bNZDNawXauqWLdP8ykFL+AREnD5zBAtyQdCNUpNpA/34O9afngo24U9K0M98Ae14
txLAcCbwOHcU0kviNM0dHMpSljEGKiABe31iP14jgr7zkg36Qrx6TQmVpYMNx2E5L6LMuQiUUQQb
J4kUCoX6OoPenXLGqUKLTrMpz4mW+FyTHHOI94Wp9yC2zHdHSCh4XFWtLNpvoz+3ugt2KWp9WUm3
7dP3z5unjhux57DUDBu8Q/7oGGfB7UXVtr1uow6AiV6p1fyaY1nNiH4g9LyTR5cxisMo7/Guh0bO
TxuTwzyM74G30IZRkCh8nG7AUKUOd5CCKHYal/SLUFpCB6AyVvVxYH+pPZotyCcnFxiI0jIaiZSU
rZX1Ve4E3yemshuR9etFBcbKa9eFPpZmgTYnDqYrH1uTBYypncUca8J2V6d8+PZGVihU2n4q3FFC
jPTa/5O/oE3C7UHHvTJfvnfTAS61JbEzMQ15VOOw07PFH9zKQWmO1PS7U4lKNOun90xSuwfHpwVh
hBl/D/eTTyO97AWK9ermeAWCh/cXYOxq1vQdv3YkkeqG4VM8pQxVFv4zsMF2yUDwzOPttaNfOxjD
cDXXIZFrHQIeaxDDPdW0qYtBSBajj6aqUSrGo3hnlxVWStWimPKZyNeeNSphrF3SdXyjB1AZRQiY
JNtdbdTRmyBu/t2NdLqGasA+ifUafk3RSBr324V+baAaYdcQcnS74JtfR/gYNj29zkefWMTjsYQx
QHy+7rUyrKV0sJjE9EwynB98cQ2Xmpqmm2OJ4dK2rQy60rR9LHHq63MXpauV3a2i5EbRlOMNZVrC
ab8OIOl+4Rh26nEYoQAW7cXt3nV3hFkR4nq/cO5CyBKalB57d8SZt/a8/CM2UfwE61Il18Qmk6mR
1NsBfoYEqiw1UI80fKUCP7AH1WI/IkUcC3DleiA9uxi3ghQUhKIGygBxptHOrVGbbtHdlyh05IdA
OrEAJOxmfLMFmiCXqXQz6BzfeP/KUF02bpE/keVnTjJo6yRuyWtBmKp8VMuG14JVNkART5xdEQ75
gvBJd5zoaVjYwHIYI7V9SyiEZp4ILB9R0lFFGw5HUgl9H+Jh/GjXdAbDz3pQVBXm+hvE0KEabf6Q
0OctQ47tFxgKnkPtY/ffraJMsS9P6Vsrl05fyfCQk5Z4q9C+5TWf1WmJo1qYeQmDMzvkcIroxFjD
T7SfIRWj1sFZ7tuFWHY5PKuZw6kYXK2EtFRM3/vj9/Cmq2fgE19VkmoYqx8tC4G6j6AxAKqz2tyn
e4/U/ImXe3r9dwAgPMew7tasurhTrZ3ZZJPckQzdybKNufhDXtUjFRF/Xvuh7/Cchx4vHf42GU9E
3u9du1vMvPUvM35O0J6LNxMsvS4EReWFLw8LMMR01r41wbpYu7CxzlR8DXMxwCh1aFDV3ELLjolJ
RJw0esdHqg9+XDJ7bj4cMjdurPWBCHqpTCQeL3hVn6pS0PtSj/N1x+HZdVJjmI0wOHYmtH1i3IxT
PrxUr/WTKiD/nIHqyTBylD9Pv1CYSJ0tr9rS2G58tKfyHYHjVxCTCnvt+OX2hU2U3a0wtQwgDYPs
CWUctixld4x5H/DKBpG0X1NjvsTtBY6px6V6Hxmnf0pB7SP0YgIRc3/0zmFabYQ3XwMsmyZzgy3Z
IBofdvmeQmt4VAn5yck+d5RtBGtFAUoYas1nnrOBskXTLcUJbBXOs0ugTpKSAJvdFVoa3Toq4Ay2
o9nx6qvNevUa7CfdKLf5OB/UdYhm6uso5OTXkdqGD+/7rcqf1kgizTeeRYR2VEIA0lZwTsPkmnNk
8gbGODcfbNm22oK38Vt8wtC/uzO2finlTOVetAjVmuq4/mZCiBYOia1leH7JtnAbtcaycclIsv5U
XiOyid8PDZETroKl/O4OMYL/OTSz8YrpTJumONaEc6FFp1VxQzLDNamcSCeA7ZQ2Tb5pSKIhZDRl
oJtBoYBWm32uf1WfCYdp8TknSirK2RutogE9bhpxu08Br1ADYMdFnCLh4Xx5Xul9enF7oMvMtfuB
CmmAHexJvHV9kONGQ/BkBN5Mv6xjWlptR6idBTjCIOyx0VcDuTrsNAXjsl6Z8UQoGqmpU8YKXEy3
DiCWmfYTY90yhVbK1Rmx7QGwStAyCXNdE6Cl9po7H0sbN498wf+my40En2z2iHGHeu3Go7a4AHav
lfR63gI/cF+SSihf+ZcT52S258mz7JL5jRQFe1PAkPOtRB1o15uK8Rx/Vj/CFuUK3vQmdawJZlG9
UJgcrBOSVo2tlXnRqKeivFkO0zy+6OsxMO1pKWkZAlGhv2zM97y00YlZKUUaENbuYC2KRRMk0XYq
t0I7bEhlvqNvRohxL85nrvLbMAYfo/36nEKaTCkokRdhASflf90lDtyqK2XV+8YtQ6/ggc5T+PQM
XMNNu/tEPDioj3WOdsgHIzZpEDNj2Wn9yVE2H4fA+QHmzryQPW3CSORpfSqgCQpif8re2ED4H8e1
SfDSazQ4yFdvvm5FQpxZFefH3FHg5rWoPyZRfro/Q4i4tvG5aUvj5QR48poBOsP28Mo/+wT7IUG6
MUxSi8UUSbs47kyLERd07duSFTloOdbCSBghkdZB2XLt7IO2Evo0A/2FLhldgSXW4F0VItEHzXua
Ia+fHnvKRm8owYhkbfNdgyrnuvp2J+t99bDFFrGGVTOGb027e2TO6Sgds2F7d2Qt9gKwi+imS+43
MzZaBiuL4u3KmyUyhbWXPPCL2R2EnIECFOBL5Gv24sgmBqj5qbgu21ktxZ013W752OzeXyKGaxO6
Rbnu7kJj1ptB1Yb/TrEAvJ8qk3dYSHsz9/t2kEL7WabIxv17Ocg2yhztK66HyfXK6SvW/O7nw8Ol
fw0ufS1D3BzBlfx29Ne3/woG1gxCcZ8cIjfIrsNS/cL+HMU+o4/P5Mwa5JOs0LeiE5fdq4nmyI7q
OsxnwxcQNUAHnYozHY9SkBiRIvvOTkTSJoa+6yurgdnbKkHyTKfO5ca+2yJEybCwmohHFaGCkDR2
4Wcrn3xh/SLARcIGzHDHbq2UjLXlh2bPLzzV9jOWSdVGfziYGNHOGS+MlkYlBRNSuBzkBByy5jbW
hgpcbpkz4/M0XGIRKs6RVCESny4CMbEmJegl9Kk2X4L/BThOv7H/PlQU+d6k3rbpfGYA2VC41tbk
p2kOnlCr1p6iAMcZrUZeJ9dmtUy9RNaxG2njp+qZc7OLud+KjeHjYSoJuVbaJ0wXB0AV9wghb9EV
yZJ5R+iTUYSPOhir7d542cRkhZxlk5aLxjVhrsh+LyzyHVVeuaPc9D3hz4A46OXzOlgA/cMF0hW7
58zItZNaFp/BlwDAK0aJxUd0AwLJuzGavd1r0/t1+ACz0vYxgVcyHvO39tWjweQttVSzAVFGV/fV
CeJzTxm6WvnqpLdU9FCWn7yKnhs6I45SA3WuIaYfipJ6cSzxEZi60LMxrtYk36X/AQoyK+Hoqi+F
wFXdvRMBqLNUoUU8NIsWH37ryE5W2hgVrJe0/8SebQ38yRi3/AVQBJQnJta1pVGqeuTzs2dX/zN4
v+5G41N82NoWFsQiOFeNCcu9O+cGvq2PDu3rfFeH7biPIPoQKmumnK2rBNuS/nCUH/WlfAtVEHYi
Kt1EoRuUTucf2FFkn216ApYCziTVfCjatrHGm2tcTiHFXyA+QN0t8tU7ATr+Y3f6RfugMl5IMyVq
okXpyykO1Z3z1aXl36gf5kyOKBIKDrQxDudC8q53xFjEchFrwxL2MByES3a412Conha7g7qWUUfT
a/9To0kwxya7LLhBoiAzkheeTqPB6BtirHuyjHZDcoPm+bbXSYNTpHboXaA3/H+UKRKC3qv+UNjn
xlDW7SqrNMtBwY0WMxKnk4RhJ6BVokX+83afa2lQ0GXr09kWQ9KKCF/2pYMJfssHXFkDC3IkI8+i
1tW7S/oqCSP8VSnUZbfhPBa6wc9jsiomlhqim9ULSNKNaiWfOAgMfTfU6ywHoz71n1U/y9Uy8Vi1
TevBSbr2ALC+rhkpHjKqHegZhsFXOxDAALPUQkYzM3Qa/280Q9Dotfoiu7I/yti9m2fplc+2Pepn
PIk2ON4egXc1jkNCceOktfrTlnYSJq33LJqktJ2dTpnyTLYCeeIU3vXP4yhPZ/92aGqZj2/OSRDJ
Ner1LPnwAEsar5ti3Bn6SvkpZDHHojLIUkoZxmp78nRz/oq19vvKHoeV35N0evKEsxA8vEQgH+IM
BhKm6mH/Qig+/DabxHfDNYP51jKUhGIDhroglhO3aoEsid45RfrDGec5C0ZCEk/NPPR6EbsSL3yN
tOMNmb9kx1vsGXWUfKBQYFJgcwBztMGkeC6n9YyFy5QUOXT+uxhHVL1SzD6iUaqPQ7/P9NUCHKfV
hy3DVVBWZwzuzy4Jm+6XKgRpf3DFgEwxLQKZolr6wXnd/AGxA696EPspe8TOP3N0Zt8W8DLN9LBS
TInj52GsIF9tz3fYvz7W/WKfCsK0SqEQq1F+zeSqEbmjqgdYLRs7l2oiO71/SPcGQkBwcDYDcd+z
GNYTuLCzsamTmcML6MXWSXnwP4zq2qXj8grgMzQZhsCYEKaNMFqP0k7c5gsf3LBn2IwFAUdZGzhu
zh46O/SFZg3JWGBULLLQAyAY1EsXomP0U+iHIB6gbjjn6CLT7ObgmhKE1ptWegAtSVmmA3giGOCU
nElKoz26bVd89183gqKGq5zt8HPSJxCHkcMFo83Z0E9Pb80BMHFAM8zt44CMrui5S25UFQ190KvT
v9KYJ/OXXcLNDbPnYMZhs/UWKE1TtERNvI/ZzDmsmT7w6vBcVwo3Nxlu2u1JYbP7ztkf0b1sYnwx
deMXLoYNZrMDOORpMQa6TCKuwon3gf91Gh5GB0bdaG/xllzF7bhbL5pr9mEpqANEHUf+X3rZEt+Q
cqoigyTrQiQXDCuFcyihVKVuPcYgf/a4MfgOOi3ZIPk9ze6i9FiiDp6EhYmsVC8CDmrgyVt7eJdI
k1evLMEzbcb513RaoOgcAvXJG7VDEHIcjr3K+1jOnzfHmMoJdDJiBm3znrLbVi5KQ0VFaIijiQgj
egwBD7Zr3uzhvCx6vrUiOYL7YvLb4TIbEfvrlwCAqT/ZZ7ErDZzKjbzTJoNoaOubHihgauLIKOG1
9cMtOrMuwsRZAvoYja2q3e+RoafyDSCiX4orIHE992yeI7nGvS/xwloGF2bXtc+n40qfBsJ2hUYY
QnN910cBwmYmSDgQEg8qZmKfESm0ydinxTfd5aqSM91a0BqfypKISLlkGbaz/Lgjv0H2ZJFRdcBN
6xAyHRFgvF7HQlMWR/iux269zGuC2ngPhj8KoSvNIJITFWBbI1jXoXMAncDskFEiWOTOxJygCOuX
5fSssAbvdru5VkEfSzAC5HE6VBarvmR45T/JBdnYozqArBJiTEyc7dpMr14EdrtGkdbx18K9zHAg
PtvDMbs2CfRldfTjv1uH6BP62pyTxfazymFAqdL2zb78u/IbyKZm0YmTlCaHnhO3hpQxtfWyyiSE
iGEwjknZCG4k+yiUw6X+/+0EnmwDyrq/f5+aNouIn2uITl+pOI7O6gpVZdT/ZpAbyRs8UkI/8vKp
PVtOyXvJ5l2zKXV9zM3Pz2+E0ApU6cxoyIKjn5FyNAKZDbNyw2gaoaUVvmZzBcQPm8dPYcusuNc2
AVtJTupD167Cn+VWgiDa/x8KzmD+UEQgQ+nQ6pxfkEZOsgC0WaT5IazYOIQF0WuULhJfS/Te7yZK
hqoliFhyMmTteGHj/7GaMqnGkaw1pIBVa5ktBYECnpmfA0pdJ0bTCsFH6Ngw0khB15R4iB1Zi+PR
kr1qmh6QfB8vQH9p+aD5Cq7Q0sixLgLE2tcnVRHf9uDj7puRXONYkT8NSxH8dEpi3Hk0iNNG0QU8
+8yPLGj7x8tMwcDNqggXX/FtzdzuJUVeg3voFWlhrEhe7eHmDVSNG6ahfdkfFc7udtTCRPA86vGr
vxetYyVsnLpPB7qQPE8DP2TNyBwJ8TkQOUeyf+k4+AWN7giTNR5eS64zEUs/oknWNOnt1cFJ77Je
Bl0qYrZr54nXCfjvXV1akFEKx961AQ6xqxObaDlFhgk96sbDZfQ2kCtYc5nJR9deaaj+JQ5ppDiO
MmEFfGshuy4ZFjQrdvsc/XHA5tN2DO7jbhYprPyrAXu7Ti9l5seLpm7n98R775S3/1mAxC9E3M0G
eb9J6sdiyM0ZV1B6NfCAwaVzbKBsqx8rPRsrD5Mj+uJ+9FCv5rp8z9g4flg/0xaTw7lPiUXEUS5m
/vT5o3LH3VnnMDy6CC9y+2ef5uRLDMiAHi/F1Tc75OmbUoHlD4975BOsSehXaQjJeH26t7fC+3o+
4tVP9QxQ6kXQKKRqtGLx3mn/BzotYrqjyr/rjNg43OQidCJNam+2OuKeTjdYT/UzSsUUCX+b8pyI
a5xXd787jFXKaL/tc7eILIN60NjqrBDiy/WLm1rG0CT4qnQNy619lfz6c1b3PCRII4hGmHrpWreu
28HgGhVKFMaX/VjDeQNvP5RAiBs3spbCeIcc8rrxTB/YHnQNYEI7WneeMDHk779zNkWMZJ2TJ3kH
8r1B+bJdHJ2J1Eb/Nec2yeAyLf3k7pGDr8vmZWEOGGT36i7Qj4PuN6I2nMlUYDNPBrW/Kto78Sfe
Jw3oGN7/NHEbF/W4QYCs0osVtZviIPDl9cXv+0roYL/+iAJFzZccwS7GKh7ncet3dfQj5h/YcfXB
0wKwz8x8iafu1Z1kSeRFRa8dJ66zMybyWH5q3x3vUhLcBzMGEpOmBCgV5YIgnouXIziracVAbxRs
nRI3nByBz+TrBqQL4m1qcjN/Ryif2bgY5krtDd0wMZ2e7C6GkmXC7Fn4gqZfCKnV8gp+wX+7QyBm
6gwBRgCMCJ8pzhVK6PT0pHuJTA7Kr/eX9T7FMWgmkiZctgnF0hcRsWkzG9Ji7XKMcTlnzYYqNMyI
UjEjQgzhQVPGsxomwsQ8ZbOJVZB2/gqeqamhtGKoSdQC9aXXjPibcLW8NWDiWHVsFZ8lej56ATiR
83aOhVlw0wWSF5xErmn3to9rVhTmQ4Ea6JG4zn7Q3/FqRC+T8+6GRSKH8YCgdSsosJCLsYsRsM2v
Irmdoi6coWDcVGpJfCFOY6ufYUSVpapHW3HEBLbVaLVJoYzoaSRBt4aUKd7Uyhsqvv/gTIA2/hiT
ZRjgkOf8CV3Xa9SgvCh8Ee1EGmCKexbOJ8fabjUX59VbJSqzJvTNXlThkdnk8seonsFq4f78z2dK
EDqEb2inyvQeZN0ly770IOoWsJGvtv3JZGo1Rhuy7r1BX7z0hFC5IB81tJkf26tmwBaeXtjs+hno
Cvb018zadKVAXSU8eDHjHRe9DeGUeXtVqeEU3acjzPcNny6OD3NIK6ECrd8MV17HwUoszcyXTHXE
A/k/cd58v5cpEc4LGl5LqAP3xRG0stHSUvSECWCko8Gnvx37rX7LAmOv9Wtzey0em7pOoIs10RRu
cbxOck5EWJow9Nff+uCa9A4lWEmlUkIRSQlZip+EnHg+WdKujKtRhYKOeOUCO4gCtWIXGTU+01ov
q1wtF6FZR4/ZUTU1+VhpxqrhoVVzPaXFFpLAempXmeaDET4xObmjf8fEpPncwqiZ0ajz0tkn/Ksf
JPxnGHorvj+tR0xdH2Z5Qs3jn4OM7jfRlfMTXFyasWfZ/2pGE/8fcb/E6JMvwevbKyR3MW8BwZ7i
ukglvs5/FFyNMF5N+seg3t8rd7vmrlNu2bEnF89cq2qDXisjCL09WFiTB+7mFrL+9zLSXJ4AczNW
wlATZyfY937ObDJuPcmgRF3h2NICp9h3rNcVOoW095CPZWEz2qpNPjw4Y4BaAihNWvfceQKz7NUy
mc63XpjCcyHr2vDog9j/8OL9HwzC+TY7htPfIyN/saQUMDSKJ7rc87QFdoqkfVUXfBJyl71+w+fv
pYubjA/YoR5vgprXijObwco28539Psy1B8XmBzzdwpVwqEuHb0uS9qL3SUSDkTvz7aadk0UobBHh
dlzvI2yH8yxGJY/wG79QuZaqyP8PfoTVNFpvxlFCxpXC0oVbrzU0IRimQlZg7Nh9N4PFjQSP8Uhl
F+gqZQSUCQApw24Q40MC05e4zzHOzFklhJppW+ItMh4CrKmCLhM8hiuKRRMeLqQRUCA5DVwxKKix
94LD1RFghLas+GlTQfLmbf2iu77RAqvLVA47O/QZvCHys9mGdUu5CdnIMehsLTamJcHIwndSB62C
11tzrxswo0qU7y7P2OrefIG4xxvCH2Et8SF1sPG5RhmaM0qEez1n6yP/aWFMdoSDU3j3o9GvdUdR
1rKg55sYT5jAj85qjA6R6S3K8V3/bLyG0gnaHv3iYJT0x5sACe5dW5JNIMWslVpbd+IUtVci6frS
QYMXW5D8e9Jvcimxk7e1KKZbdZ/Uq26FrJpsGS37U82ALmSRLO4Qa3noNj2JEwEFoA1x4QjLO2Ea
qih5BgANbGSfv1c9fNbnog+qnZleC+2oM6oYylSc1wXomGI3P8x04kOp/Swmr5bZwYX60wLrk0//
1boJA177N4m/0dcKeGrbaKd3tBRykydQQoLjvse0uBlDi+1JpcoWVtqYR/SnzyoVldIwyrIHuxAL
Qvg56gb/2ANs73tJ10qG6OPLyZYI86E78hMDUFHe4DwcX8nqV22P3lHu/xpu4dv7npcxoJjbyc16
JMb2hgSV+oBhCf7lIIbvzAYbepWUhtv7mz/znCGrw3f/EnMJpl2WBk63g6OTvIMaxfAVChip5rE2
6a9wdmneCJaCO23tiToNnHk0cS3mSbDmx5V9qBrvNdtz6hRfaRmSsuQinlt80/Bk4aQmPn643pQK
LYPDaE0bycdPPVBgEebc15505XXocQClT9BlqC2aY/bTM0IH6bJ9bmOAmYy10P7FqyZI8bqBnwuu
v78PYWLiKYzEGANAc9G9F7EwhcF17wKRDWKYRM5fLMgFze/zefRCGsO2dYI3rw5WToJY+fSIvmn8
Rmvg3QzUFqpqpnyjA611gLEthPCyFBaqjfApfNH6c88jVP/2JRTUdp67+T3OAw5zy0RT/cXJRJp6
kn7rEoa2UvcUVVpuw0yAL87YptiEcygWeRdOiklJSCndAysg+WAaDqqEpQgssWdNPc+iKEEJ7o5r
etSSUslKACxMSwEyT5h5zXyWcjgM0LG37JX98V0sfhEIES9JkS7rmSi2xkocyaQc2yEeqN3/Hl4O
nlXcZCRUD4yFDRV6n7hTk1pO87kVIGrY/wp+5/igsY5R3uy986C4all7hkOXa2TJ6Qu18tMaDKaP
zUr6RWO0W+UmdRK4gToZMf7vu1Tv6/cR89moVN589Vh2kZM19LxeOi6HnHhJyWxepwKSw++VMSDw
yGx0EM2n+lSQVuhjwJe1WZ9Rpw9l54iu3b7c4bn8XZL1bN6utF/SGgk6mXH2HiCC6p/O14G7KLWr
Ctrzrc3RomjHtiXIjpQ7JvottwE8/ug9YOkou0TXi5o8PMLt/O8hRmFpJ/jwMQbkYBsrQ1lDGaNq
OPevigz6wWgaRrl1oXTHxq4V7sdfiJj13TXNtUyraWZ3d/B6RyLBAakC/fNoauCD7k2nIfFf98IK
Wo+lsolpt/SrZmu2YC26qeKDV44OhfFK7zhWs7yjmMbXmTgkdtjZif9Y38enhUNwtAqIexcARPN8
k/vRCXamuCh9JTFFBg6M6hkROTrEi1dZccytu/CN4QY7Fagh2cjRQ7740mH6gvpaanxT3z+5Q6e7
OokfzbChs7v7521xFbZwj/3gRe03jE+9n+0rTo8nz+XE3tR2CilUieRqOiYk7bmLep5xh/L8kfFD
d4/LYPsCQPslOUOcepV3X5CPMVB+3k6kVJjnf7r17i2uf/n18RgGh7i6FR6iTyhEm/eKJ7TQiRXY
c5vTNYNZ+wdulDGGxWOW9s9mXfbJbHNOXjIhuvpAR9pJiqlzVvz4/SOgY+u4MCIKmvsskmSKdt1r
tziQJCuI/yLI4YyNZIERjjFs92X0jWbbFR0pRfLSo/zV5+Qtk6+d61Q8gz01uxUbC00Pf5USwQvG
vxJ0ImZxrQbSZ3EKqincubBSMNDX/F1z/wmJ7mcwTK1FCBO2vbg4qgaQHuPb4YFZM6JJoX+UKVV5
SxKqNq7vuolleg6Ij8NYbokujhCUO0zDsvWdbW02Gb53TSDwDCWF0mkHfkmwf/xIj8T2y0fVhGzc
v9aX8swXp6mhn2PXvSXlVQOy+uY6mUrbZxGStl2zPOIlMCnCwIIYM00GjIZ2kGvK3wy8eX4aXI/c
Cyvgs6aBpYvgv9SHkLfmxrJboSfZO1h/Yz2UdP5lQ59fsD2v2IWZ2wOCExbgd6swvg7qkIRbEpwe
9T4P0UeWHVjIgwHLlkmGCq/rFtZod7cPhWNbsCAwdIcFjgliZf9XkVIM9KDglk2mOPJb55d69tyv
mv9KQY+hIkL1Sksa9APz7/T5PYnGbdh3EsQmweTNk4PhoqPpkNGHaMTTAXGjBV7dtObzQhAIahTT
5kt9TTQKKcyX4cc/Gvww/v1xoV4bdlwFaNGmH+DcECQllSrRWFYz0N7F/31HUYEWoPWZg0s/sFp+
7h7FUQcDseYHfgMCj24Hij7yqrEsvlE79iVZR/xwJ+egbpPe7zdkJuiugxAgIMhvJ36qSRbLYyNJ
wRSXGh9tuoxSATGG8d7FRmzCdDpbl9G406qIiPkWY7B9ucnLF/XoIoemtsk1wce39r1An2nGnJIc
PaFz+RGW94VC/vDxdsFDV2BMf5f4nq3tCwEuIrDKB4Lhf/4p9WBa5p/3vyC//kj4HcEmsnVJLAwW
FdwTmWpGAqfLH5g7TA+ywqJlMpbJYLWwsk0hkJS1NyKWHZtRqaZhOhLHGhfJaJFu88d+qVRqsfm8
TEuLvgYgaga0yo2Jp746hPeQ1ju6qwljqsZ0uxHtF8P33urYZxNAo4mMbfNmSlLD9dg6lzNs7ZFo
j93bnoJY8LGhEJNyiNTknLbE+tbGojyHWNE8fCWuyFYJZj2+uTo5uhcZwf9rpkWgc1XAWelmM4RV
tVLTnVnaZ5kVmXIsOEUjpJk1rBhfKNndY/AtCdazAV6xk8Hj5Bpw+mEJ6hn1HzdDFOIJtohEn2Bd
HAmi0LHrhuIUNCbVYLSzTd4pFQ4XTE53uGZv0xBWBnlz+CtlabJwiU5R/lwYgGEUbmnz1UEg1XgM
zo7wN0RaLSGDKWpSR2kkpFO+BgpX4/v8Dkwyo5xwnj4A2uqbyxV2uQkzhS1Z+xE5EshWd49aOkRO
dMPYuudhIuXgG9UD39aBe+gqSX1K9ARbHyMoMHUbneZpM9bjhIZZjDXbqtxa/e+S/GKmvPzKdpYR
0YYVq4gsRflaxxkzTvi0ik6nSYaiWeR+lSQ3NWS+Z6KqsJ7x/2xuf30PeJIqImnod9HXzhyxEvrU
sBYAs3NVzqTkhIUoq3nkeeJyruqOdO0sb55l/2eeAKzFWBUOLgpP84lXqMFspY7wQghQ4kGk5L3u
dTLxsPjGAJNZjMMCLEvEE2+CoXciyGjiw20CxBrJoNmDAWyaZw0ZYyNF33G5XDrNPX/bIl4RJwUu
4lr5VOdqLZeYP7x8QHEqKHSqvxiuqLqtTCvfJozkHvkm+wN1Qeu/+ipn33zM+jgzFGmKCvNh7sOa
YqLOr34puNKbseTL372oNKay1y5nkukVTz6ydEQ6paku1v5jnXTAgRsHRINPQKbF2RTZOqcrK83H
M+JUPaFpJjPy2h67OSVslobRRBw4JbpghW6W04PCGMUuMqZH/JPmGRq3CrJ0BmzCO2rr+vYGcRDa
SlLSW7Q9i5cPIlWmV/90FoJaF6sYrwgVRADiB5EP1x56TjcoWpOGIAsupFPk3Ey5sHk4m1r3Hgjx
q+a8fV8EGF7EfzQrMc6k8Q7F8UpGNjHjIMSrd8wmDFBSZWUq6eXqGEkyRY5loyi0I3gNcp8Ut37d
UWWcD/XhDogV1rgXm9Jp1onYjIWwQqdOsZUy+MqeWrmbGdT2UP3sj+8YwexirIpgnmxRnudW5J4N
BOHtjMUdtuG4bPk04JPenKmf258PigjAIr2oy8YKUVm7QBQRoh2fxa7bGTWQaaTGPy2gD/QgTCpb
8tkgGCK87EOV4jdVbSwTHS0YWsH56ELlZ674c429rTS0Ss+A1y2/+Jw81qGRN4MTIoxCgeU5DwLo
H4FG1LTJmbVYmNEdKV6IPNdy0m41OqR43DRKrgVH0ufzTaLBzO24PTiJZuqiP4I0fHpP2VO51gIf
Jw8jpZYF6yAY3s/NG1Bgig5eJSF3Sl/WGh9ZIghDbU/szKCtK+AQtilV7gldvIUSpLMj62xngI1M
1W+GRWBQAZldGcEhe1+bzRZmsVQZg8aY7ap/WQzG0l0Z9N4d70N/uotrk2X5ku09LyM4B6jgbmPx
zjkUqJrLQccnne4PO62Qbm5SA2eByk3YgCWopXQQKYosqhhlSmFm+L7UbE3Z0+GAYEC9GJztA+F7
/nqbfoylJs8Hve++UhfetZLHOD8UWnqdaYvpeJjCSiD0h+Z7Wayl96UK5hN3pntUuTBHmZlyesVw
7XLwNWOBy5ShNtkYsJyKISIgT3Hi5z/ylYdctHbWLqaGKNaRDhkTcZzs5/bCLq9rUNv5XFEOBuIG
J6SPn545YET7ahADL5EmaAZDBxihsv1KU2+e8sYRAYZ5MLbDM73xsgMHHidy1SaBu+nXkEXxM69T
CHNW0FrqV+BonNhcBA9YGoPWRME13jzPfrDMMMfEGOv5FyTtdg3K4eJm3UWEE5Kx7jmje67Mqnym
/kT9lJy71yl9mVBZRU1wEeNW90phwVwckBz05x/Bi+nVW1XBaaXm4NYS+EQSZG2fA1/tQwwWo5xu
jqLYaAjnWEG490TuftjSrCXW6u2QHC8ItUMCqEoBlgRgA8LMgfOgeUWVi+Bo6yyGKMWSa4tyBVxI
G2R4yVEilmM7M+vmZnsajxJO6jMGQeVKCKJ/UIVasmnfvTQr39qzS0bno+n3+rU+odkefGiL0MYN
e3kmHCLZSbzvi3V1F1YAjZ1Xlqy0+x59vMUUsbyNEwc8velreAUVFChRZ0Xpt4PYlSmudw/ilWQT
GVKsApAnURgIXmh1xPwW4mLT9KNEVZe+6ndATyHjrysZR9D0gYd0DiKabKWpAnLlcueSPUr9t4q5
z4m0qQmGQ2EUVb+o9EnsS85a3FLraVsHRmgn+KNEFaA/pL4QHYqIsvhSpF71etC40Z1wVSt6d5L8
F3h3IPHRZKYfRqQSlZhyPSDTSt8nDiY+YMuUBXEXPRvitTSF6vbyJ6i+Bto/HePWUa+3Ug+R6aI0
AXzUzCgCF7yYRl+OyG7uKjUe17Hrsrj4OLzxYTLtKC/HUmpTBewiQiFIQ1UAuDsWuWTdtxXmtR/4
Mruckzj0m/6MmMK+VqAopO3vwF8qrEpiz8cheGTw5CqISRWWaI3ffXbf5oBHfqk7SJ+cNoYADCn2
trenVWoBX0CLmonl0pT+vJSwxlem+SxhsptTdnjq7kbCO7WhOOyKaST15kiRnMqJ/cfjeQI+6a+P
M9qZhsGNUZMGgjKm88St9mr+tC6ZxLUFu+az/nuanpSgcMGva07mZUQLe5c9iHA/8GrvF0CVM5ji
1iIleceQPzZj8s/92vx55n8pcUWn++68uIALIyk8+5ChNsJ006PRAT4raKMd+mBq+yOBpkFkVHGU
gjjNbUcqNCVyN5g7uiRTIDPXbXhg+21vAKdbmUS06ytHINrtEboP+GQT8VpzbuZKN65KbmG7HuIx
UXCbkarn/HTiPTF+OGaBCRlQ9LejVRrocRp/QzE27NzZEtALyyP4re3qatjN6rOXD8P6k04LALW7
Hsf6eVaCTDBoNt2I7BG2P7YUDHwfpcJdKwwTWMdh5zeGNpXdjOoD1Xt9pvpphZY5xtGfM2C4cBd3
bec6O0h0LpznFZdnWwHhUao+0bVK0ExUSlWGTehHZCMa/U/HXJFIPhnIemsaWMJq0Yx28AL5ulqW
R0nzo+KSO9zZkXgCtaQPC2ECymSskqtCyg9vu7q8th5yde9aWlDKOvYjtXeI3EgKSggpuTKRgBpj
4joo610n/yTYK0omGlN/J1vR103G0xqmtPOslSt9klDIlN5oVmYsZzMXy5ywlyG+miCoT0HufYgh
q2ryizBwc8a2sphEVVAElHTcWF7kB21l19IhOa2ReBUJkAt3lu7wCh/wH/cbbCbsxNm7pXjPAocw
tk6oGEFqwcOCdQX8Cs8h9IKfsLsKn+fyu+egVpYeJybopFn0dxxJ+5I0LVLeVVDa7n/xrMwHbVkW
m5LBOnGrF8XoaHg+cYClTPh7h8LhTam31NUWaAR5tQ3mrQfAtjfwBzfIF0sPH0A1Bn6JdQticrz7
/3M1aPwkxM5I/765DUTJPgbvkdNmlPSHEhS43l6Jg1vKb2uZ+ewhmi9pjhrOTboLGU5NVKXuMzNZ
vRW0KMTyExIo2sZ8ZOks/9E4uSwGfWGJvGROUS8QsN87NgrIrikXNrMCjKHZ/Vpp3T3iVhUg72aO
muSacIbXSObSNJq1fRAEQI5BJV1X/VNa0uHjnSsCz4iFvt9d8/RAgzBRkP5pj8XbRqCYIhpVbIAS
3w32bcV6B/EEWYgVQPwJE1SCeQEUJoT6DdPDX0lxdIGqO8n63Cvjn6jxnw3yAMPwKvdJINOk7fqf
Q5LX5ejFV/ZKJJtot0AZ+BB72AdIbWIuVU/DQujHn4Apq8FA4OY5Qk7wlI9EnQx9bKIQyvx8MNjB
AQTb+9tM2GDMzkWtBgr33L9m+US7kFuu5tXnNtCYCCYDN5Fhfq73k+q+q7MFAMF44Cli2aGdTIkA
l11wPavo3VZmSe+S3y44aVzarZdZlmQk6G0vqdFD+ME/ql0bHM3cw1C/EjDDWl7KfAmKALC9ZOjr
K1kvjPm/CSclIQwk549t+mo/Nl0GErUauqZw3kDQVsje9cgEiLUaIYTLyxIWnwsIK/gVFX66isYs
k3Lo73lAcTnQ8Gdcg1mx20sEWQuoy7t1Jy396xPYx/He5e26n9wQKWsYnrDZJNdKym7SXvfwuP4c
a/i5CZKlPyRYaOHC5kBeF50CyKrUkLjpBhmGBb6eeEB96SymYulJz68Rpras36ZllcM75SoC9aIn
kM69b3WD/BJY6sYzEaI0LEFafQFH27ZMfaEUm6NAwPcDfEveGthAeeU57vgYh+e0JWJEX5BLiy5j
k8SlB8GYLvWAxqDY7wBdFvxILQqnNK7XdWqbD1GO5IquaQUiak4lMZ/KOu05XBsq4Lia4hiYWlKL
UFIF+FrqKtd4PfN1Kn0tKfTy5He8VfX6MCHEOm2zvHBF7uVaKXGeLtP9ohh4f811YcPdoLlQbGyt
5L3pOXYavzt2XnfsPIxhAvcSZuD4CorLJscC6a50WMSpRnzYyAQ+jtuaAqzi3KCeslbPJwdN2qyu
N35Q0RYNsTqnWuBbSr4+jo3ZWRsrh6jkXuWoVUA7v9VE+xLd5+eAcQFaK1Bbc/BTXCpr0Fn40QZ4
cfKc2P5BxiffvCwolrqgFcawj4z5WMCpOdtQtNRBkvwmxjAu1fUpm3PEBxi7wmPoxJ4tmnfDV4By
uF4LkTR9POWuMbfBOm1SqdHAJ1R1+dDfejhfD1Q/1bzlVFjY42oUZZihmau2lgApd9xvgzhVIf6J
jdmqoaMPVPdrt9yASVmfCafIcqOqVG6oYqTlTPvUG+eOB7iUak1CM+JeMkI+b2yWRFnRh6iq93VD
90Kuz01B91K7sOtDxMciJB/gLc3oOyYaCi0WkKViBsFhpB4dkX8anzUQ4bsAYDadWHBIctUTajJf
Ew+0a9qbgp6v+gy3C48yGCoYFjK/kK3uy9jVXNAy6UeM0r62IgN7KSc1RJdsEKsgSuHaGBxeIHjR
I2RkZjapewYNkzZxuKkdtFcIcDQhmlbv87q2k1dHBeCuqvlpGxC4hCDPL3Lw9qN6TwVbe+fHX7dE
uN6DpdULpC+d1VO8kNO0itut4L1uGBSZascwZJLIydWWW6CwHIj1NkuM/IyOZdaBEdr+WQ7M2TzF
awMsdv8/X1TOHlx0SCJC7FTJlWjxGBNPKXAJQh+BpVZjzk0FFQ6ZO0fSqRDg1idXKja8HmEl6Fc0
SqvTVygUiHALk/PtcJOpwZfLj6+zzUsnvca6mQcvZGtihgEmcVAupwF4+wDu5Gm+6j8lzQr8kXpx
q4AGGnT+JFMgkpYeuG5NG5UFj2fgG8v/Liu/WWVL4EHPaa0ys3r0y8lRM4KSEHHWj7Mxktt2ChKK
z18CuYL1Eb7ydfqZOUNVuQrvkeLrNBPwlB//W3MrQ04muOiq9H4mLXhfhHBoBoZ1c5iWj5tyZbSX
5m7LBR+boYD3I/NrD5Wi8+OotpIBbSCJPt+Us46I5nI7Vl8iN973F62BqAnw+5gry501OtfeY/SB
XEqPEoPiWirFm2cmtI1I7s83wj1kmukQOCh3yx0ZVBGzQzHkJppUfd4dBFlpm6P/QpmRJ6ChJgU/
T9uUi3iO51f2CDIw057+uuswSDu//JsDhZlhKl8Fniga0qdp5W7+RRqaO/L4YUxqkCkTyL646R9p
rMdVZMTirGyCsDTZ6i3ThqeHgTy8W4s+sOoXqk6gsNgr8IO0h8ID33Pp2ZAgHZ5814rs0Eif0qUh
zhjaEtGpnkefyLr6kLPXZ6Ptxyad8Zxy76RcAqQ/uXxiyhkk9VanjIWmRGU1KHbPg53KSFAXxV+D
XZoYU1UNKRfk4rt4QIMYLLobyvgWqU7iPdPhIqsOsP+dSDCNPtBYullwvJeRaH4lLdU42Azv/MKc
pEv+Ad+IPAo2kl2njm+78Vt7Y3087tm1wRqhuffyfmzIs1eh2qZiSxRPi0LbJkAcZCbj0Zp5nA9t
JIdpIKqSlJLB8qvJYujPS5b7i71w2ufgTRo/hrCAzNS48daRtOVDLpQvSg01W6K82pZkTo2HX+QE
PpFn8b5GcF1ve0pIi+BFI2TPu+WkpJvOGNv1Svi+BdGJqb//38eOkZJtnNkZqx9iTLOB/qbARhLK
AcYFbri1JwZYOrxF53BbZR2k5b8/SZrX480J6VALEoamKJEJXyiPhNlPbLIbFlnLw1vU4CT1OyMc
IrHYr7dQ0cu04RbxnL0s/B8rUcSB07YUG3ervtDpdy1bQuyG57vTSSSFGyoHQ/dsRCCGIbfw2JUy
u6r7M+ABH3alfbJ/cNTvnGBqbFlx4WNw68v1NBIfIk6tU1ejvv/LfOSa0Zsx1mOIEB93ZlCg21pM
YzGxUtvI68w8CapfxyJgBf7pP91JRZVVTbaPiOhwlKrcIefuggyQrzb9GXxufbj+PZJxhWdbIUEI
aB7+UXOK/R7eCSje7Bv7ekuk3IK8IhIBQ7owbA1DmChuaveBz3C1s8LwxaN5xqZaOp60vKbwNzcN
rwT95kjb1lCADjnaviTftAFypilMrAu9cyjCsxomjTk0PTKK2GMXP4CAZxBxMNHLrIpVVj4npFMi
MbJq72tb4m89UWZejk/gXo6ygsaDghFw7BbzxQkFsoEsp5UZB8Z9LO9mJvq1S6ODuXRI5Yo3UU1l
3v8Pb7wlxoZ/X97BmnOoKctEhMdh8riAOfoq7Nk2YKJ7oa7Svela0zX2EySOvrX+BzLXK9MLEkui
/juePCaCeVbnP82jGDF89xqmeiTGhBIxqpV1Q4S8nDja3B0BJARQOF1Hgqwo4w3KQw3ezc7TB/ui
hD+84TOhKk/Ey8PSr53ao51rV1MeLHzQJyS0bz477hCe9WUdSNG8RN1yLnKjmVqWvODVYdSMdFSX
3ne1JSrgxHdYzgsDMK+mifuTcKu95CdTT6XeVX1x7hpyZKmdmckFpM4KkPb9BiaKN2hyxuHXk8HT
aMALrPV96gJ0IX8C2INB0Hz/eiqn3aw+tb0od4JrksHpCyP7uvVO1uAcLk6a01Dk6SrnHRx6/JDD
X5nKzWAI8/pqSkCaY5HxpId0Z5IMa7YoE0jH1p2amm9n+nJSlz6/xMeS+9wDCewjo+wSCPEQ/sTA
wJ8KgkFW27Zk3aE/Nq0zTF3wlu9ZY7eDwmccNnV7PXXqbSXfUl6AAkEKGtOviiwPzR77VohS/X9/
gXtNgXbClBU7rftwp3yuzt9vraPltQSzlxMLcO5PipT92GJkj7YEeT4N8JEIZ48jOjTjG3Z1QwXW
dLKQ7zYB6i20zKrFrxpu7F8t4hfUZbJgFG06Ph5B8Yn6XVoYs4nosfBkv07RqUn6KAGbfvWmxum/
ybqEz0Guqx2LUWy9C43G4bQBkrqM1HcCys5iUqj3QOHsF9IWCWRzRZylUYigZVfE3yJRmQF4E4Zz
Gk5+dEouwhYXXcNJDxUZamwAi9nLlQTVHuBEDTuNsaewe8H5NUywuIj95ktAfYhbBXihklXzDJeC
pGi+PJFOjyn4PrFp+7tc139ThN0DxHI5BDFTJuUpSt9kUKCw+j+fUhR9kolIWNxWKbZbyO/9GwiA
fg6FeUSEOcbBCphc2qaYJ+EUB9uFPadQSiZ0JicLnBZZn1rRuiwuhwXIpK8Nb3UrSahayV9g9Pex
USDMjrOKeDlEgqWZxOMEOw+nz77ukarUKb6gjJkMc/FTgx+B9mbNB9Vc5wlOfmWCuXQlWTwHYdZi
HTPzr+JS3qQ+yYLtzO82JlPsakZCGvF7YWMz/dk3MRS602uuaNKML4sTmI0nSI5LnSiEhJZzytGV
xMZtHJhdMkAU5NwlPBzDf4iWYhPLmJovFUX3OJfcck1cv96zd7p4nsjQp/1F0KLNeThPn6YEotLS
IAmqPvk8N775uFymp4OlXAYcphayZyoBdudO2nmv14IRIMLcADqJyPdOY1yua5HOJP5P9Ji8SisL
dwPTskHgbQXO9REzAo2Ump6x3tyuJAwLcNjY0SKKNNq+feFsZ/oIwIp7k3Ltko7PXwNbyZwR/iwr
HO/+Myt9+Wb8zqejKL4VAV8DtWhRwW5WbfyIAUKHJktRWlWLqiqL5IoVTuHQiDnqFU8WdPlN8BlY
WiMHT6hbnyaiHZnbA/J0+CEmhBLPJkn/SEbNw5RPnd92yXAPfCirh1WHPPw6OqO+hkg+crTbXLeg
FX3oF1gF+B1TaIrEFLkVsaCVKHdQS56s60qtyi2FO64A4/Yvh3FCbDJlHI+hgW2s1lh5vy4QSeQ5
gaN+aI/TUYo7RTZG1dMbYkOrEEq50rBJzUNoFN/HtdSST/YUjdUOIaph7Q70vfLnt7UV6kA77cd5
WdtaHyBUHE4DUX6zWWdgUGLbV7Sh7zJYv6MS/rFwaWckCaBecchEH1GbAL2YHaNXDfinHV/OzwZa
TuPpYITd6JB6jYlWRzdDHn6yw5TvpHObQwB5YwRlhhfkIiq1l5cA7LujXJlqO2NBdtkF8kBdTIlx
Y9Wb3Fvc1LRLBp7ScB1+GcO+t6Lun8UglfAU+UuqBSy+hHJ/cvZQyJGn83tuiTHjLvzW1SrEpAqS
mD7mcdKSUfkduVJGYU1MmK/LE2RUT1Hj7ghFPlw+W9TIkXX7h59waOGn0RKap+3sNex5IrzXLGo0
+u6GbB3uX7by/K4znbIb5cFm3cu+skCPykcY0wkqx3ZdnwyDbVH3+1DoWazX+HUTrjlrDkLozTu+
EDUa+iVT13Kq+LDWILjSqnqTcACQOnikkwFjIFBzVghJpmD4oXnT/kSNfSFLsJZOjDOHLc2TfwSC
nZWQatQ1IriSASU9DnTfZAgIAcpIyI6/3NAyyeqeNeGFr1UC1M9d6vpMchfzBc7n9FizIvypEOdo
iMrmtqPOOway6tdaOdf/QW3lKe5HcbjLu+zAqrKZ7dv8ohsIJAx5YT+If6Fgmne/nV3UtV7qWPxw
qYOWxM0NfNplo7jX0JMQN4XlRhhlmVsrWEwwHthMtlbUioC6pmYWmrpKaFHn5P0Tandc6dHfpzrN
gJ8m/UcSZWPil3/f7anjBEwfq4fZDl7ptJW09JKNyrYXqjoQUH9M/nWKpkoVvbhceCZNwkI46Cnb
fAqXNbdX+0wAX+oaFKBPr9QjCYXnnaOUQb7v6KsZYh7WGeAV0daaOsuuOECVm0IJyG7zK990+zND
cQCelMivtury0BbyJCPRfj7jegnhENcVZXfq0/rSZztyluumzi5RLCNHJ9qq8P4r/sAobNSmuKn6
CO2U/ptbKNFDHRhM0Dk1g8R3tEMearw9jKcdwpqs7IFXrDmrejNmqAMZqnMNNLjr2PKBzuMQXw01
EjBQ6sYBj2WZdf/pVEEySqV3g+dUnco+wJTaOhPWtaw/KmccMgDslQEI2+lvjbRUHsVZqgR50HEX
zwyLYEd4DnbBXSxS/zv0ibXAAb0uLeDB6pUq157YyA8wpyUwlKmUeHoKGcDnJaFRRa8OqeOkQ5df
Wo/TBHxUvMyZGiQ+WHiy0ky+ErwGUrW8iKc/yMQI0ZAFXM9jYP+2L241puVlEw2TgyOtFLJiaEJb
cDv0FJJunUIStiSTtbA/dhBPZvuT5+cvAHANcXZdNvF3YOl8Vo/SK8mv3uFfDSa1KVZ3eIXafWHP
z1gyKXmurxJxgzgpIdt/9D7FkIqa697dGfQy0zgInvOq4zAg4OCAkVUO2uFuc2AwHgSdVfnNNLUO
LjnwpIudSH+bAzrgZfT77vmA1ofR3UzFab1S/bENrvAl+T+lpRFYC0N7RKA+1gxcpaiEcJAKfKfO
E/Ki4O03QVK5xVr408gBxjhKJNs8CRPocncis0RobK/3ZozvOVmhNsLeMoeLXw3w5A7CkrHJ9SsM
exndG1bjoskSImhlf/nBXoldfmqQDm0ZPrZemTOFhQG88AIBXFJ68ddsUPmcECazASWAtVhJQCJe
2JMUiYnZzkwPpimgXcN6Qlkx9o7WyhoV7eOmTZQJQ5Wgj1Elsp1FBtwaUEsjvBfkWfryY9c9+Huc
OMuDggPCWfKrYKvYiHU8yUr2EvL2rnxgOz4IRGKiM9TCDqnQdelcvpepGGxx/MgHgyPFA7tAzd8I
u26l+NcUGM1jdh6sNCBrfacFvBpPNGIxuOhi3e0Nz8IFBV6LKE8SUewCYZJgUYPscrOGDj8KdLTj
qZlOxInwSRQSccwX1Zk6I7u7kTws8FajSVeOFHl42W+LjhHtuw5smSUW2L3nb1lQHRSK+K1spN8Z
rKzDWLkqtIBeJzqkYWcQKMoNrRfDqP9oWsX86hxt241jup97c1apJ8KHHFRzowAAADWTjVGaPBut
bHYF6FJDj5Loi9mLj988Pj0rgunJn0iFLxaDoo7OgsxyT8SmvYKBxQJc1T/6h4e9jCEj9gtaUdWO
pyzSPMmmEEB9wd7HRG/gT3IteQnmSizvBUnc1f4vAW8zpPyc1lwR43ao6vwufXApK9M/jE2CuC2X
wY/JeuG52rgjfZeQcIq7UnBQRfKuZ717eJnEX86s9LSWB2ntyyo1bO5tjUqfWxjCnOHVnHI9daZW
M1d+RcfYRFuOSCMKExEK7Ub6z7Im/8bsnm0x3fv+S+oF0TwIelJKBowObvj6QJAjx6GAERh9pTt3
N2YhPLIt8UUCYOQq568OpV50JlVjk6Xz0vSD3Pf2TUVShasMj8jnsjG2IuW8TZp8ZB5+K5r3YJJG
IdTAH0e1o86EiyTQ/IyqU3NnGHVF6jbTw7bARVIDhLJPHmp1gfDio6wB7WK5dL1mw7G696aiTMTh
K78mKNtfu+VsqUlDFoHr4G+R6aw9VNgX+IIdFFj8H7+GMUx08kOtpJVDUeGf3da25hgW7rUEs5pz
oAcdLnYDnMLvaZHa38SFH3w3GMiUk2hAQ2ZMoVR+PrD13WraVHA8bn3SQtEzzGDXFevIm5cOn9tS
qvXejslUz/bWN6e5M1ftkUHDg9fOHM16+37rv1Vxy0HTsi60DV2vr2J+0pS3nyBy3v17t8KIMXVG
MljuvxBb0oB3kB8Md6yF54HI9v3t3ETo9HVin2otnnCyf6UWI/tjNm7I+JcByoW5JAlJh0WguABk
nyq8YSJTFAdWlAZfuLMfOoy7xTHZZkRjFqZ64ewwH34R6uAS6NfmkT0XEa/NfeRuYEQbe6YKBsaU
r46DhO3tGbpjrUwF/RMsDE8/tzLkhuASidq8Y0NXPoMvKDnA5lXVYtgEeeQiFL68sAkcEFpE4a06
682Z4m/8fFVYLGKFRO4W6RnyAx49iaxVtgi8lxdKiOfs2Mp+prtuGoi0uvZ5hMxokWFWv7hhbTPW
+6KVd2WxIXLqyevb4Ji2jIuY0QJ2QqTXJ4HpKPdPqtkQRJLZfaSq6x4vXTWRvwWjOiT/Z+08mwyP
Rax4eEfPydVsqyNxsZk9TmoAyIAZF7ABc1lkQpPCUSh8YJGIeZayrd5M+eLfRfrMXVWNxtre+5q0
NJdTOse1FNQTLTzOwMTrQXC5ES+dUvctbFGqOxQR5dv/N0bgCgFEjIQHbJy9yGBS3RFsvJSyH1Qi
5o7JOVxOCEd7iadxHtaoGui48yDPj0IAAAriO+n92VLS2Kuf10vpCYGE/0HE8D3iaXdYXBPbxam6
WWdum3ENiI0364Vtu41Z4tPJRNYvLkVY60csb716hB/eBIYNj6kfjWlFkl9OVYudiv0Pn52EjdLr
KOY9k3gm22G1ci+j0QJUMiHKxv4GnFNT8FiCSe+34fiaWKaPoPuUlR09cpshuEP7VHhNvgMx+iVu
e/ef0gKw+12QLjA+pmLCXW89iK07zh8o2zSNZWuEbQXdq43oatDtfN3X4D8X2+xciaMV4CToRyQG
VnmrcmMqO7FR1EQ1uVpFqK0lxRe06yp6YiNEO/UPaxCdT5XTM6Hea2Ibvwvzf00olGa3+gHU4AJS
Q5CexpQeK6SLcrqbl2JJ4fjhBb2qVSK3JtYuHJx7gxpR7+aJPtTaHXqAYvu36Mzpx39FSK6H5y9R
8+9S1/zPGrQx7g9LaB6aRxFw6rsM185Dr/NIl8MYpH4GCWkGtH+mOa/9ztint3Ngi6ivAoOMaHzP
zPFaKbvKN2Wh4UZ9TLXMqv1NvBz2dusENZDDWQlcSREaRO1WFUeCPADavJsOHmvK9vnzoL74246k
2bo3qYZvCaCeZus3URETcmY1JHFZ36hRPcCSXp691DLIxSN7eV4QtzdKfB4uhI/Lajv4oAGE8HD3
of0AGa1/j4cPCj8GHZx/MczJDJI+DMuVYuKLme+4to9ajxHaTOpDPCc+Ot5ajhWT6IEnilI6O8Ou
FoBmbjoe40CFOVILuGYgLV4K14EtadDUrCnouDSaFybL5tCcJPeqTrTxi2t+7T1mBTOc1ymeQWZd
jh/+3Uvf2NkeWndHNfpKxBXjgwtYpC0rFzGQ5kNnSFly8O6DraqKko2yrZ55i5v809Dq6PzFAaWW
uQJu6AUjVA76Qu0NDG8k0Ly6UqaddtKbkkgExBD5FhSlVwcmYNO02OyKSwRP8/6edTEepTk5ApGF
b4hYZ/mR1voGJt8h9M0tzFoVI1x1GjT9INYi9LjObyoFe/k76aQkb53wulCrk1Dij1chTgEt/XIP
V+913srXqWLP584sMv8C/YCEO0zRjZLJcu/AkPdXEg04S8lFe3sF3RQeEJI6RAH03gFxbgYFCYY7
DVLk1Ns39K7slK2X2KabToUZwI3+0k3D1VRxR5NflGKcM8+YnZRJAG8BPSmKZ2VANCkXIbpLm33s
OcArTe2HPVJmWxBHXtJvNDh9Y60V48ZZ1dBPHPYRcVftxSYpGTWcqmYcK8TdfhzF80hSGgwHZZ3v
iLP0VtQ3EgmZZyhdYFWkgCpB8TVV7K26fiZ8qy0C+vY7N7nPJfXOv44YXvaaoltZPOO/lxtUx2it
0tcMCGAh2kFLNdxmRDSsQ/Jvn2yhbw7+eS6JnPx9/x4x/bs/ROXkcoYYs3aAfoHLm+hstYZgbzxy
aDeJkl147ML4fsSdZy8gyKFr9t/O3asX337Ki9wxfF38PiMIdaPlT4reMeG9UlEK/tyQ3CNlXhj0
Wm++7XUZMjgn8aeCdnTD8g/3NREeZ9mtW9XQiFFgrS2kNJiBZuDtCuqtt4zEqJRfkExq+XNxKHJH
gh7HMl/08x6M1qSFoX1mVq7IsKLsTjRO1p1R3/B9qiy75jDUejr9yRHqmebjqZ2H71JD/VWFecUG
MigZrIR2YUTbaRTv9dQwXKng5aUNw30xav/3sJAcwho5Ayqo+PSN7JlXI38IMEC7ms2kqP+vmeJ9
SCEguAvLUrVUljqqb+8ySLSTBHX5RMLYU5f+T1wRw6SCgsYciKvYHQs+tdMwjJlif6Muo4iJrmFt
CMwATQAAXYSoOULX43UqzpDsOAPHPd/oVTgslejxZCZkQPWqzpvzun+vKeFTdKaLEOj6vnl2qIqb
y1S0n3Jx1OydxkMzwUmXLMYcaKeIej+Yf05V/wbJ4x7WAMai/LIpA1hSFV0Ci8bVkn3n/vgkZPwz
u04/P79/lFbHEx71CIQzRxE11WIyXXKQXarzvK4+jEXo8szzvinyemkT7QHUCiuglzGhxALRCfqT
XvwQGmyc0w6UMG5w2RsQYv7zxHIlhQyvyGYDREAZ+8XZqwOGdhkJ7HHHYoRecku6iIciLblykEsQ
NDerBlCo3Qtre+yxSEgK8+r0P65+W4sFTIThwj67vf6O4XA3ogjQMJUIN9x958OyRxwVgF/Xarwq
Y58rErgds2+lVbP4P+hvkK735ag9lmQ+IcZO8y84YtbImpNFh16yE27t56TnMLQERYzOulprOSq8
Fft+3it0cZYN5whaX7MmQeKKPvIXN+4ojrhMLjwgDrOMrpQjg6/yZXdyc9DbiQbgLLjpAbtfRRGO
Ova7hEb0NSJBZBVyKzaf9iHWoJFGVNEEwdrhIdCz5BuxkuGe0948wS/IYzLmq6ny1Y6qyUIBzBSe
CEarL7YTVJUmMfnQn9EvOw+D2px2eZ8gRW4SviMebLKVwcwF2xcoQkkTCcIz+OiDt3BUy/H7NIav
Z0CvqfQH/Q7xNINKei8HyfQlFk+tPJ5gQDMZ3KAifVpGAQwqQgJw0Br1ni9hDIfnvdgn0ydT0kf8
Ol1dh8IpW9hs+KIjpR67N6q3Sr/0SaDaWmZqRPVXKUo7LdGLV0VqyfhR/J8WHEXzbbrINs8LQKt2
CqiljFo7/dIGRZllFoJ1843SaZKkt+ffZv2vZo6nghmUGXvUvAdfMzb87Bv/k2LKcA/6PuqmXSJI
zxOVnmuEtrY1xIxyPqxsfwMvnkdOyQ32KXfeQuK5YxlecYIh0l58zxqDGyJJMVQLjYSXU76Ap/UJ
I2hcyUbaU6Y6j1b3wYse1lwV4DJ7IGYyBTXGnQm3DAkDShIQ9l8SKk9of6lqfEZW+5BaPWQrANM3
hx+PCmb/kTGBFJhGDXa7XDM58yos/fbltUKQBIwSWy53Kt1lf1XrnXM+2HORUTIf2e/dxp4sIlw1
pRitggIbaq1XnGCW5wLTleBUT0QcNx3Cvt/5h+BpiP7ttPwLVvObU8P9LmA3tlxi8N2VivDlCH1S
tAXbd2sqT37I24WmPnHD4vUzo7qO/bPUO+Mi+0UAKFIMsyy1udPpQMTHid3IkgHgMQXFalkpZDIk
mmfgIoH1Q3wxuvvyjnmrI/AQSVAU3ADpy6mrhXCxFlCh3Ox2pCvimimTN8qkTydnILdBECGX4fnV
Ng4uI8unSka+abV65xAonB2wZh6DihPC7TXr290mzYz8DsPBW24fSQO0O9Qf9tdWocP+NwOxK5Gv
XEdgs4TtBmdar4kuIU6FgFZa+D+/iYNXyE6PRQTif8Vf0mMvV1WSgqmwhL1RYSczzsmGM/cRL+LB
DAvC0kURlC1/xlDHuNgr9Iu7XZzv7Msp6rbDA8UpRdWgsDhVGCmV/yqh8Z+KYXLhylzHoT/4BkJW
lvHSO1U+iHl4hXSlNCYrBCZRY7wR9ZbFinIrDDDqWf+6XNElMF8I2mlcVjJSCkqJsDQin1ghWq+4
P8yPdTGxlgnmhjKckqh06kLFHkUiMDgBTI5zRE5PZL0ChvQDU9/frYtmHBkTEO+XLa0WtTTlO8RO
vtifFsPzdDb/414LRI8N4DpJ8NHgyr+DGxVG55YCCh9ppDwywQhVBkDa7QYs7VOdz5/hvMxJ1r3i
bV3djTdFSIpHXNhVN+gyrPajP1/iZxWOfFRDhj1+N4lJEU1ICZUF5T1Qn+5xQdeINc10M3P0I1/s
6aR6gTtlF2diBrHc7pWrSzDF5/TddnimFrvbApDs+07Z4n/xmXC6XFiou0PXsyQXOCB5ViPW7IPK
t1Sufb+aboGic1FWgTYwwFaioZARmR+rTv1k0q70R8A+xqSY2uBpsByGs9IwPG1TpU2GTvWrh36t
XSaJMXLcdtiFhisfTdzeiWlYvNS5jiGKmb9sQ75AHC7e03fXhNdOOmxex3/Van2FPIxJI9sj4l7v
KBFBdlyRUhRLmyI8Csuby3jMbizONrtKFlU40924RzJiHUoc+e7DpsG7tncN75GPw6U3jIS1sKRm
ibQI6SCiciDPtFsWbm7s/RjEidbFhHC6EW11et0VOWSeQQvwQJmbWgas7cd8G+SVC1Ui5AvVWSrc
SJ6QEcsBsOzq/In6WCznG82hlZuSKCDBZx0ZLM6fHqBd/Xh7pRTWnThLbV36OyMStvuthx10Wvsc
TIphBdrGUCDCsYFuF30FmvbGOMMD2K/7XaWT/cbeaqv6sAVnyd+Lft/1idfXiYCDUssB1GP+kESJ
/KqelHlTb8qMxVPVmsPy2y6mBeIp08vWiWEfAlmLiaY2ynkx3SFv7tDdloCmChcBBd/UfMzSziiv
RxlNXSKGPk2XInRZfL22/h0ik25HllFFhjds3x8L3P15u56ubV8zLlgkiWRYvI7pwXxwcSSQu7mj
HQSzeEFYuEifbEg/2ycaxuBHZPwkpGJVHYbMXa5E1D6q5+6U/NNP52vEQCaJ1jwDN2j5i38wjeBz
5w6ladc0lJSHRheh6sGtapQooWKjc5oOJ78UzNydDgdK+WomLilqLDouzGypluEGq6w7eSaPWJIY
9P2puPUBL5AYPVQjNUUNrOFoIgoH/C93LaPlLX8Z3PZlwhZ6nCuzPzMB4WPi5S6wlRzrI5Y/blZu
jqKhvY9IG6wxhp8KVVR7KmSTJvgLPzsYFHayoDPXRNzwsuJrytI+9FxgXYuVzaiuZsEfQfReIlbI
5r1uE3mdf8tArMBUNKGIc+DZP4sMxRmGbRTRjFjF/QepCtfCusH2U/QZv0N9vGuCf4QCgyEzJE2a
ojL5uMf2bKrMxbDpLTSA2NEK6Zw5q2jeKoD6SsPkigJ3Z/l8XRR7PRuB2xu+6wYEsFePeaZQRfdT
7fFvCHJkho6ygaRSkVRVNaQL9GgJ732PpEL4pmt9NL+j5QI1DV2Nq4vOOv++FlKRJw47OzW+2Ay2
qUoZkX2mMr+VHF01Ws/aQZqjEgQAljlSmJoUxYh/T6AWFpTB+P5tNzqi7rEnwKV5EuHuZ0A7Jkj5
0IuR3Ez78Z4oZDtasDmsG5I5rhbNnFW/H7ivauwJftsT5a4itZFS7Iv9zlavK0RzGWT6sgMDrnBv
+Vk2M45uGOY2sK8F7b/y5Omab44ICbPZBlURWW9hkfGGhjJa9QjzkLIGUoMF6Sn5K40RM27ROhyP
c58r7YTbHGJ52DDOnADqRkzsC5sVrN4/8emupy5YghGVVm6pJGZVbrbnM4MK3yel+Jahz6C+KR/G
0wcdnKf1CUpMgHPnp5G+R4BCfsAMWdQiOlT+2CKRFEZfUANnnDsK+SMr3TSqn0Rb7voyBEyVUtKj
NnqN0UCP+ZA4F9krHNvkZGb9ZrEsPNzV/rcb6M/0FFNCJoZlbmPO36JfklF5tp9gWD/ndPGlqp2X
K+CbIuaszAldUNVfRiuc6fwx4ajAbvkgE6YvK8KEPjlZZbyAl2Z6t9x1qDHmf49ENeU8q2xwMi1k
0d9aOX967BJJAbT22te2OvGuVT3x2S9Uhz1ykcz8KTs078hWu0G6u/351WE8QmuxgIBanpvdr1zg
bmq/U4v5E3OQs88gkCJkT7OvlOIqWbUtSTOTI9gptgaC52LYo1NXCjZ22e/fs7sf7+uv0i3MiO8Z
oXMbUQ735bCbrM6YG1kYlN5UDTXxvqitvYRYCsu3fQ6ofDV+XUZvYZHyK14TcKDsQMzSkmtnW6kq
1oIvrbi899Ub4YqM0RXvskEVhKZ+GAfK1/iYB7faV+7vinW5hHO11HIVCT+i1HwzEWa6T9NJft6G
vWkCcGYP6b1CLx7ke0XIXXVlvstd1c63rwBa0OsQ06DJCjQKeyKGFX+fdCz3MWdOTzcDj5S2I1MT
95e1apH/AH4rdTvnBcv3RI2mTkUe6j6pVZQK8kLWUUZ/MEY+tw00eaNivGbr/2Xq/ENAI2peewWB
nBujq7foqjyQ6JT1y0V3keIPHtMiCJLrzw/FXOq7eMX5a16r1L2UofDbTss0Db/f8zwPirSkYHPH
wulTpNNgpbj8CYgMGkmIQyynTrVKjyYyFiH4I0ldVr9NrPm0MGWpoDfVMTfnx4+bdzdkYD7/kDkP
v/dC/24TB8EX6mZGV4DilO2HblbnF1N4KfGUsGcugiTI3XJBeXy6mnk4P2r7e5lsSmxnlGoORb+Z
sZSbeLzZaN2qD4EqyDMbCP5NEJUhox1nDYdYPOZlsIo0D7+hiZtJDbCORbd8g8oo1egELgIpNIu4
DBRYg0fKMuGTdK6YELbZM3mD2ABvI+6CTKKmuaHJ66Svn9qQDO7BgezjdxUt6bkR0X67PO29TK4g
Q23I5v3ReYtMff2c6DyMYvgMk8T2tvCH8Bg6OCsQ5IvCas5RkGgapoPNet5Y4dCu6yJiXOPIdlN5
+8k+K8yNG19LbztMVYfRobQYqYAw/AhUWYOGGgkQTPIxsvgXyyJqLrbt4endV91rULOQRBORLWEC
rrW/byJs3NgTtLtK3u0Oeym19HaOFDwDLnkI+kVBB+ITKCq0kuJBR/F0IW5Ft8h06yQMNCOxi6Ko
lUtll/RSBzVtRTd96MHvf4m2XoHPTLf6/5D2QHGLGpHMw4uIW+2yPt1T0xDFI3R7zxRG4O4vhJNr
JA5IVmB0lOhr3Cr9jGiEb9A2UTa3AW8pHtrRxeaPPNKc1QoBbkh/IKJlvFYnZ1G9VHdp99edrRV2
9WFGQrX6HfM8yGbCWYw+mtRUwFBGmPHPdDrmyHVbAv2Sttyq5UZBcfj05T3ghQDkjsmy7eislfMu
nxDst+ukzL5t1OqvTlVHmdjLt7IOtdJcn+yTJ6EoAxl7a/OwVBdwXKS1W6x2YYc39eg/PNkLYrl/
22662sgR8XjrGZRGDKEi+QUjiNXQaQcgExyS0Vl6XZeiKEzzehgYGgoJt6vPWKPKe5Nv/lrUXL80
q6c5o48DnJwVud3fhLSeWId6ep2ja2P3KImsZF4dclO8QqJtOjseGIz9Fmr8uIgIUkijOJghX/Vc
wvJTS8814SxGIXR9AsG9dZl6j5ET+pzGwW0q2JhXW9SnpC82LS3OrZIHtZoRhBbeaMCObFn05/U+
al6HJglBL+9m4V9zh5iLbWOw0pvNpAInW6Mls+LEYocw1dTGErW6TqdadcEixpBRryA/VaPyRZIL
4jIQ+qhCEd7OZyPjR7oG1HJ8328VpUadNLFA0QXlGFRE8px+F15rrmwDLUyRG3vO/2QYDN4LffA1
kSvjH2AkYUx3dU6ULFEnQrPDjEjnNvffwGhrNS93UPQq+IloXmEkXgoaxXE4yF5jpIU9fPxqNiSR
GgTLN+6FISA4V8qZOnIWDAe4gG1Spf7Pne/HrzdqVZLU9fyJu1Ka4sHcDRafpTG2PuiDhDOtw3dI
01m1qxIPABNZfFvYe38or9yJc/yGC7W3WgzP8e+g8UOi6tBR4AldyMjUUTABauKGr/cNscfpkIr4
O9TJDA47uQaVlhiV05Sv2g7Y2I1RvKah07UmczJugyaIhtRpimNJXfA/bxTZKh9iqwrx/nKzAfRD
gpfBR97QJUqfRnv8bVOphfn2kQNm7in1/0FStNbKne0atQRJN0+r1noWhze9jGF1nuEluAGRtgnj
NItXdNUdVxlnw5TIhPGIvu9cb2DSzkutcOTW+GHbldSfzmk25FwZO4ud7yeflaQ06BbXkm6Vvcfd
5F9Pu2FCMypApukIbiYypTztabMMOCNOD3LYCZvJD3FHdqvmakpnhrGdciRhlaXTVVn2yGCAkVH4
aPVp1BUsEdQHHPBuLHDmjs84caZMo8z0gdKtZvMW1WTSHfRuB7QNI1pC6wsP2Nw0Dw098v06YpXs
tVM/HuyGxFiTJVa+rLlrgqjfoyn293FqzI+CmQ1g6vepCoNDRk1SYp5BrWs5hz7Z5u29h8Y0eHsV
OPxWFbkJcCpnbqIe3XEwVN+cg4KfsIElcnSC4+gOc/gwjjfaM9MrJ5B07QRE/QbkiANZ8QOXSuCk
GsB5Ilfk/VKz8jy3iRifxZyTnOTheuUVw0mC4vt83tC8rkS1cLa+7e5b5VyHeq/y8PRuLaF6voIW
FNF4H36xVnsKCrFmaNLfnBUCeCiPtvIldYzWTf61afF9I+WAXHg8Hf8BgyKvtZhYl02anxRPgab6
+c4egFvJJLQmpYTF0txzPL1ar40AxITT8tQ6KcCynC4oFz+FwMiXnc1TF5BiU1xBiwJFUiUBP1ub
KwFxAEDCQOG9sw5GeLUW1ykx9GjthZYUtuREyjggkcHivj+65B+VZtC+l7BO3/cxHhzcUXk/oynk
69QvgzY69FRhhsI/ZtZkT8mz1Y/bRP5rE5pCyfrl8iJjqBh1/lnzdJmiVEFRf91iUM/4RFUDqWDR
QOH2ldlrE7KwmTWRpgW+Zuh5r2o3uXBZQR2CuNIOxPDPbuE4XmxI3qGN26lWMZ/ox6FY+LG7UudT
fneKw1Yyqzl2Ng7qK/FeFKnncm29zCy0ohDA+zqq2T7SiYEjBOXeZ77ivIhH3bFNRSlrV980Pv5L
tlqAdpr+h6JVLXBNSbLXgbAl0HStNmBGP2EcI7TzMx6tdQ6j6p2oM31H4ZH9UKHSIbw4wVYRrKZB
m22dgyk2GYRciuUD1uQFNO9irzCixXbG5cdl3u82mLUJ8uqJtf0m+4O3Td4myvGJNxWxQrNvh+89
hy02/5PG2K4+pwVQpU0fnn7vwrrN4Dl0GbpTsodPl2ptDcCHJhXRUKuUNISvZHtRXp8kSkCG+8Os
AfQzmKfg7VFZneB5hbp7TIZQjlEHy/bHuNvfzaL8hc+Bu64jo8/Qpv8WQIAT3Kor9bSbnWiWYRSZ
FpUG0DeEnS3/+ksFu9HGM9Ow38nb4cI4PtbV1/mbSq6qC8gTqabn9UjVu5XlIzT3ggpIN6D+zBKz
IJCdNcwyFuAxGgxPeI1k9bswq+NVcUaFJPQPByAAKw4aHRWPGIpBeonCIENCNsKG5WcWxjF08Td1
w2UKPMcBP4pPeYE+RASCmbAC/88nDD7CGmzZNyR2C1Bu9iFe3/q4ypVzi1FojlybkGlGti7+5lQ3
1KTIkNWvzPTKvYWj/VQxkNBGD7TmormXmSdQiVXSqAdSbkp1jMJAJG771sUJtXg8QOfRJzspubtf
0KPcyqS/7hMpN7Sgkgn0H94WqAktguUGum73d9W58Pq1JyXxxKuRnUvYKx+D+rra+FCqaDJF1Ure
Dswxy1xla3/juWmAVr/XTBA2JxWey7fQIrcwhX0edKU8iyYXzdQYTXDekjbowRj02fU9c/f4q4P+
DRye4B7lftchp+ZYyP90mDJeQ1Fx1jI2dDN0l2ZCui6Wb+rtzWLhLguPplXTwL7w5QBNmdyXdk4n
4mzK/5SFJnKVxhK41cm2Y6yEIkEL7vbwYRJu/Q5aKGTeuDaOvobEtOkfbDZD3gf8N+rIby3Bw8en
mhy4TKaSH2AR3RKAS7k+yuyLtsiruAASDFyEGbXMwjbatG8qTbNVpvdQIgeB0Zb2PExwZQ8p+tvQ
z56y5qf3iCD8uZCsAOElJGtOJ9aZsSKQO03drIB2Qk8ndHeFr8XaQlWFJKk6YjVQaWwcLbrEQJN/
ULJAwL23iQg767wPSU2dB/eJRjIgfpwHwuGRAoC3YbIUTw/NiftfYBc83R0YPlpmtDjPrk8OeXt3
rn072CgBPCwIUjkjXPyPtm89WTL6YWi7FkkT8DoYV6VxLcWgyL8P8h4ob08DqtEIhrinylXCOOmS
mBBrj4rJ0tXGSdPT+PCNO8v6nTme2F+XUZuMjkqNU+izifeU98mRbDSUKz49cvAUSP7DCJGmh/rf
RJInNZm43PewihH/FlzDx4XQy39ZaAdjvcTKYMhgP6p7Q4Qz4tTiHwT15/75zvSjEsZEdtzP4cJY
1Klpie832uZiPxf4bv9y49EUEiK3N3MCS/7k7pzEbxc6B+6GJ7D2sHhhfZDk+4OyAE7maIwB67XL
GftoQ5wlolvi4addS/4WZ0kRYEe9HDBG2K/bqJXmJJ2TxFR/1k63/boPzBqygOJqNX7Xr7rFDWgn
0uF0WGyHsjYOsm1Vr95EISpaTSX2Zo89qCplG69OSd13jt0Am2vzI/JJjoLNpDdd+FmYQ1SvsHAp
rpVSA5cw9PPzzC25ew3h7jMk0tbydIOYQLsHjm6xLwF2n/9v2tDQ59oPfCocQQgL0/hpX5V65qyf
PkLDCFxtriGhch0QtDA7HrUZajJgnVyyu9TFt/7lGioZ+K+jc3f2NuB1VSOf7Fyk/KJ1G5Ov0MBL
WIFfpygUgsbevCLyl4ucS3wDpxjMqOEgKj0zSDXsv0m4GrtkN7x4Czzrl9L36PDOWiUu3hW39ggT
9i7fOh4iEfUsmkfhwBBiEWc6hAadvVMdbn36fwdL+Y/WENjzWmIJKT5c4cOFAPvhXAFvDl5hky1M
eJtlXwVCJczqHBP7bBpklQa136mxReUQd4kqiyBu6I/1BXvE0jh2q1OKy11xtY3ScDeAPj6GnQS1
BJeH1FjL+4oo14Uol664z99PytZCszIyEVUQ+0yh/51RLoOcdvT0uvGozQ8zZrzXb1MsFgSN4sU/
/sCdPIfEbxDkD1n7ksmxeVHcPHl2tCTTneq4oTQJam6d6flFUiO2t9kqo8AKxl+uI01eNybLIc6h
fzzsfQqY/upD0AhP1Yvd/Df+KXdnMoe+rFwAoQol+1YRceR9Jl/dnxrr3croYYeXvIDliS8HasPM
YJu8q2bAcN+Te6T7O0i28rdXHMD20SK07ODZpwb6RDB4TVhi2Yo4+cKvwQaSTkaIGR9GtHhVTR6N
tDRew3S656ms8eMvCLV4Q8LyAyJZXna9on1C2FL/Geq+hsyUqhwYq0koTcHKX07Mw7jFJ1VWd366
9HVas1kZ8GRwg3dO7IAgqvd7csRVMwW8tbDj3uMfDSTWJAKWLeYqpI0tUBBdnwur3vUDKbCJlkNY
hqqNMJdvcEuSGCMqVYLYbu2TFx0FA2eeFkl51J31QfbzSDfrfkLCbzGnmmbMUG4gCQFHyILld5ix
d6qQxX0yGCX6GBfJPFR3IUWrPQgOSgDRqpPj/LLyZbzBRI/2WePuTeolAfgbkVCiSCCCljqst0UT
xDCxcHOykf+zT3bVEaY/8EtlSX/gfbdG4PNUEA7PHZafTP89xxROxKOGZtOMV07TGfKjpYNhQKIu
iQcf0n/72emDPJDgI13TUKIK1iG4uPCq189dLb8BpyOVFzmO4WbDIeV3N5CtGMxqTSk9UIx0paBi
Z/BXa84olkEzQRYFGce/c8X51lLbOscF5MmgxFY4fuIOuGftEaP9AZtcaD63hZX2prm4tGVSFNjz
ZcgHqG3P2xYFAKWHAp9ncsVGda6PxaF8zhLC2d63dS+wfwn93kiYxrXIt7JrMDdzvQDWOqiosMDS
f5klDkQP9ZsdV4e1bJho7ZE5oV65HDm5o+4w8qCCCAzhZSorWRyrGvbqqMN36f7bGMqmsfalDIKN
VrIP1znwbupWcltbBvTttL4vFdvTUtIkOwbvD9JPSIDZKgen3ziM71WhpqiWrPotqHAZjKthlJNW
CXn6Y5v6JRVLDnMlYnZ54uArM8V5pKVNc5AmuJwaBDhIgE9tsT/tyTiROtLqzpzAwLPbCd7M5HGm
DZ6PIq4Fj6fZToR7hBMj++U+8iKIrM61lyX0nw+DecOn3GFeiheG/1SoXL7wrJwfHWBFAKUXMap9
Ljvfp8VFt8RAWO2eESxemVULl1qUlEAuqa0pxCipxRc2dk89/SqkiYQqXB26fDsIK+/v/kSIqD/L
uvKWMyFnhePEu9OxktPhz3tpPRN0sdyrPtvaE8rH6wnmv2vhurxRT60x6cqV1MB1KH4DXR+rCV0G
N3JfuveYQEKtzTKyrvew+/KuRUkruOjioHmPv54NGO8KqplApjVZ8VNryye2TeX6bpemCWtyfYec
iHFK5eRc/L9Y1Wt9nwN6l4PfChmhics1mRCoF9C3qPeZBnW27m9Hpcg9q0lAlwddkIzuyo90Xb+E
GFRU4Yb/AibbYJtjiUUwKun33KkeE7VGGozwwE+htlCNuwAw8DyMd9LgDUP2+SjZL/gINq3CHr+s
qk9pD73+myTAVD0rpErR41jZQdJJc7YSl5vjwzhIUlosyUpSHI/lO+YBKOS09/pWxz7QgjsqeGiL
VJEPfUxzyrMbKP6gBdoICkPkFiKL9GlUnAFLHFkV3G2WtwSsbxXfp8AON2tfzpS00LENJvtH3Wo2
uW4cq088Ly7P1Gk+CNJG7q9vxofclweyuWWkHse5mfB/zsHEL5V1c7MzrURylE9Wy11vjY+M6ntM
0ViRdwWYbxTBt/S3y1BXgLPTcVqBE/85pfrIL6I6VQxn9oZQ/fsZK1xdvVeIy82DGnbgc1oHjTnS
viDGRVbfIFL+Ohh+CMSgTS61LclpUZUYOPzq2k/q7zahGbpgACwws1iEqjJ5HQewwGPpI2M44aj8
hG54JtYXMJ6/xIcCo9tm7M5RaO533uZDsV/e7PP5CGwCMhdiOToZDPEkBhsjfHNSnbmUgkq8Uw7x
8vd82Q68xvMvITT9E9Pw4pTd3GEsz9lySyqgYwjMeKV4R3khgmVFnTXgLbTc+QxsvH4Am1qErWJH
WnFiwj0+8/v3msNoqsI9sOwFsA5mVZcSKY3t6vpnw1CKEazK77m/8Mmzbnvf+N5olMosW5vSUV/b
mq6DSiWTgyzbFbEQZTjrltX3IMOz8IP6ldMD77Ob1CjCXnpGJhXHp/s4LNJT2ZtA5y6OneSJczOr
Y8CABUHe6UaebrXd+T/9SBiACZjnYKlH153s4upI+7bBt7I+mRBozDbuGU1DAe8INtk0Qd+I9YgW
uL6e731E1OgI2Q2jORAbN8hUandxMuDcCuffRQ6pZ6ZgTAldxYLqYwD4cC2v0wuTqrobfMdIA0pn
ZUlAQ2Udwn6GldNe+2W8QoqrRIs2bvCZTBJbYmfMF1hpBqFmGCAloy47AFkpybWLDV1VY/eTIx3J
upGV5prIu6KmoHT0XcweoNYve3JMAQbAha4mjq1BnB6z083i0Lac4E5PyQgDX/f91OmiZkuydn4a
QWNxbV348bh6salq7AFHIISpps6aI8x9xN1T24oV5mesrfS/a5QK+yKQkk+ZGJHxhlKzsdUw7r2X
QkwKpK5JOM4XagMTV4SxXi1G424/QYJn4lwS4ydM4wNspWhmtZMWTZgq8XeF/MB7knI/ij2uJSZc
Y9cl99rgFSDfXH2rRR5GA8P1L+KxclGIPLAKtERoPnSyMnBRzf9eGY2UwoGWJ5PMB3OcqNBjP0sr
FXupCK4aHTfm/OowZMoC48rkcwsU5cWZkp7YVzsX2Jy2oLWpbvXGQLCuv5HWVpG0Hbl/yJPqVefw
OHpCsbRG/uzYKNkZRqn79WSc0l7B78/mHQvDMmRQq0czzaW6vvo1RyzqE/RAoUV2Pfzn2EPsgMTP
g+J4I8WeKYqL9OVyER9LnQ1XBQTsOtsDv1kQgshgpcDxPNTCU+ctPIVQuPd+/2zJnSAUKntjn5E/
ama3o/KvTg8+WxjoBUDYzWHzDmiUE38dp/3NmZWvapKq29fAIZ+IP/VtnBybTz7gk+xNT41dPvEP
LIci2uq3hIxNFf1JrNg7Wb9FKxpayuHJvBx3uUW15sPqY+wRhvJQVeRV8R1k+Q44sOzd9hx3nRkK
6UagPLKOfgdPW6AsQT/HbfdClTCdCZajZlIqVTt99A1K8qSr7FGTgOvBMtE7ob5ntlMSSHhhSKB+
/aXPHsytBtaWXVQMmVHRS9DOBaLrSo4gLkVe2Mlh2clNSx8E2DiLmWs3Xm8jBgDgrupU7zB00T/B
3OB4hlYI366ZoCkf3vMqxNmHZiOFkFFPen+GMLsDm9n/v/9DFc1CsRn10pqUf0iaHE55jcK/+lv7
3UDeY4kVArCPKEF386LXAKb0vyIxI/nsKItzWJIWAn9ql/kSyLtIOCYDim/gVpF7V80SwKntoB5G
hZkOFDirOwdtwtoclnt9bQqKtJFZ6yV8/4IkDbsZIoRcuSZDFKpzxy1sBDhhFaNW1BJCnJoXe3BA
o8nFb8q2oVndZJwlL6j50QGBwErDaep4xUKCXltnryMrgt/uby+kE9xA+69pmpoLML2mz0Kbo8Zr
MbIaP6pPSiWZfeXj0EOSZKrdJ76ZIRuLdMRJAEEsJDI6b4QY8LBByIMI6lCdZYVnAxewRE3rIu22
mZGhij+s4syONG9kuPf53rvf+o48+Ony3DbWorZt4HO5JsYyzXATpAm/PiSM5RVOC1N/uEwTlHMo
4o/zZD6nqcHfYjYCklZy9xl1ryX4AFUW8KDhDl5S/xG1OvkQkazKg/5GY7XaY1CLDqp7GXow/gVq
PFsrP4vVH5BErmpx0GR+5myZbrXKJx24PLnVgCX50SySkE4oTPkHVNzHG47KmoIeWXEm4YedRkod
iUI+/GLDe6Gs1IAPvUzcRWSim+EAAwiIVXMsv025QVCupGe+6ikZM+XQPSx+VhTdNecNBfBGr7C4
qTZv7nVh+DMJpMW9fjmp6LipJ18DE/wDbMohtxXtJQ==
`protect end_protected
