`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FpzFmER7vLmBWiIRffBXE4S71SPKG5mtFLtJBQhOjsesKPaU/T+y72m/x+mxcqSj7czwUhiV39To
H06PB9bjAA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W8L1NE6hMOv/k3EYkdq6wB+bYpqgyUbWLasF229OFhZ4WvMnaf4M2in0yThKD2r3BSuowl0f8iMy
K9h5vsJ6td6n0D5TRjPx8nL/yoRHwj9dy4Y+uzvGeUrFfYLQq4n2FBg071jzQGKg12ZW+B2Kxw47
z1JM+uUaBJbNoHxq/Eg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BLZAZ0IcyaAb71TwJiWMhXIb9hqcpKlVl67nX4oA184Z3LYGrtm6DuFZi9dmeyBDusgnpR2noIP4
1Pe6mgonql94Mz620j/jLoUS0X20LL+uxza97tGB0iiJoDvDfb0g/UvVHgFdS8xMvp05XBwHrdbm
0qHxk5bhpfZPjRKT5ap36IrKt7LbO7IA12HeuSl4h9Fb+G3OXli8NgIwm1rCMcugDuhId1G1I4CV
k/oSiSkSQtTli3t6G2YOlLirRxd22N+jhJS47NYtoT5Su1gJ+++wG3DiZH+4UDsCVu/4SmfRz+Kz
NOCnYGIdvP5PFURuHXfM6r50SrURHQhpk0ZV9w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ucn24gdPnN1kYbUbqIy4Em0uatkaUaGpAaMeU6upSU3bBzYvszdz89HsDLfasQGfQfIHp98nYW7s
SMXN8piHsKVGCDqmRtRSKk8AtaHhAqZ8zLHtl23NuZ9FGidO6VVHZ8jUeom32GtANmyn/keFwf2i
IqntbzMoaZijeqFJOUE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gKcHldk4iFiERv81GkDoDL8qunPDy4rrcK6lhG9tHQepsqxMWPROrjDJjAxGEZUD98XGq1CAqElQ
pbKR3spZ7YGnk1EWNzxw/tFcQSYrIrhjBzp4NhNMYU4hbn0pRoMzyL1EopnYCr3qdL+VB435jPMm
wUrEtPKCOpyEDmzyhHO+IzdDnSrSms+JawEtz1yRsfNRIGUTOre0D40J950YP1sM2HU5RAJnSeX7
/NgW4IFgVYv2pV9PjSNRmKa6e7KmrINnlELv8y+8Jo9i2JGf9S6P7KP6Ps/u/gd5PUn/Dn+LPSNV
/fCRnDTZvpEsK+NgMAZ8eCEBuEPGRo4yOsFr5A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11184)
`protect data_block
jKGDk4eEGFnr5jUGQLWS76WkUH9YCgA1aSLWZHUpYM6otVhx4dA/2R2bkiCAuSCZD1h93bM6Okza
wp/23soVeVlJXdIjQreKkHxgzoRDIt8KtU9Dv83InizDVOwTwniAnxRN6Ex9i2TO5l8rjLbtV2vo
iFi38gj+39ruPbqIfq0vNIB1jHcsTFxnS8Tn3FTaMYF6sOgQw9leHdTsd0vHDrKFrmtqWBVsB5TI
RDe/rMnwBKHPAwQh7go5b4yhbnJ3iSqrevoMO6pREPe1ezYc8ycN0vvpAjVW7TuxjK84PlTrGjEI
vaXXiFrOggsCPJJWMXw5FUjUbud/aquCrUpetqaF44ADLx5WEcSxD+KlVwHriUBBd+1KD7KkuknS
lwFi4fKoHBlKfkUc2RslRMTm7c8/St9szUvUDWYY9FP1S+VUSMHFmXRwPnIeX+iE02uJ3OfAX346
Rj4L7n8GiQww3NwXoqmYe4bywpS/+sEsE0R7CgzmM6gop9Oh/EtNh12lC2oSqz7+vng8NJfzhmM+
UoIcDks31sYL/JIYOSc+h8ox2BYVJpDXn6ZKUytd66+CqzdJW4OzREvVR3lRJOpMMDm4y9/KnLqQ
PbF+A6I/IjlUWT3muzJV8xeb0PPlT9uzskWMGtmRRIO8UF6uNgQkLdNTVKJGJqg4zN+mBlKFieHa
4aC0jJndg4jAWo8j6wdw/dEdZQGNrqD3QZb9cQGnhKUPfAuFHfpeNtHfKEKd8wEleGTFmRSPrHcg
oIqQ82f8EobJHcdezdqquoDWeZcZnkj2jgpCw3zeGNhOTKq0t9tHKk3GYdNIq7+rS8nbTlDe3zOf
dsFxuNLx4MCGKTvehBUKu2gZR81TMF9L2kInpPPDb3aOt5sowmU0vynoSdD2pDjmEJ9OgnpHGr91
dTgwbxjZ+77ANIA1m1TbGg5M3rcma2G8s9KXiSxbw30AEwI9FPH0vMNDF+48COaWz2UG7CLdShQb
1AsSvnqNmY2Jpi4wJdgiMbpqARTpgdQ6n4Tf/3Wd8cp9OWvVh1N5EI1EuRBrCMQr9w/6s7w0yjuh
hcLu7OhWnpeHQeojn2mBKb/3WK9YE2gNIPpKau4k3YSh5FvJDlS3WMP028kZzRD9gfPoKZnFaDxP
qgZV0DMWtrdfSPM+XuHg0zAjESgL6dlr/LNlkyD+ULX05h3h7tSQYTaR6AcUyC1wSNyoSWIE0k04
+8hpSTrAPK1/ftK1tMfm87NFH0RIStIptnUiv0ug76bX30HftOZoMb2XxBdonnhsrbf5U6TZK9cn
LtrwWXkzu8ZGPLtjHw2YVpFM+Rh+l+Jp1sljt/4twFek/wGo6+J2y5GvYLkvXKvCJ1Vqp5GWz7ej
pb8WhktDK13CkRoRj+MVaxnEOqqzj2ftljky8xaMOrfkWLqPEUjdgkAnqy5I89uP2xjKtzUrIJlq
7xnohGY3fyBdt2yyswIUZkAsaljLCIfObs9ANZ7S3/E+dUSGqTXQ+bFOjbz8rtEI3EMBCAd5o3/+
5LtL8Vlp85FilIujlxUfVsAyoqQDpjeq9SJjvGADVLtnkK49wB4O8nHC57VrSKm0DJ9X/2Ai6Jy+
qYaZK5psJ3T58G1AP/aft+D12F+dKIxjYb3vB0RWhtmOxYOP3CGffR2xpS3wzP7X1UPZPx6iHXAk
WTgS7LWffpopxu2PKvGg5nqKcjkucXuxPpUIb27zpWDbuHtrPoDFgbCF1+VFAmYTEvJ3heduwsDU
9bY8dbXDko+sF/SLCxg3WIOasLTJyedj1jO+Ld8wzgM+1ZeypZpsj0ENXOCMWtlMziDiPGKSAJ6j
KZwT1h4cQ9wDjf311m9KLzF7DQx4k6rC+4NUZRX3TXQwMB3qsVqmMX1FTsltmmstJ/r9Z+TwSozj
97r9GuHC8+gwL28r0nPCWi9fr3yzGcp4c5Bu7Gx/Ms5bvibrLhGfc8LBAIDZ1ospOuoIyCcykuhT
o4h6l4yZTMNJ6129xpVxaFtyPucyTsDTStzLDZDD26qy3bLL+STTYSZ0fgoD+KytoA9Fm/p9EdFl
9wsoxdLRpvzbRuYjy5SwndZWfiMiDG+Dfpl40Y/ZLAZkv1NQCEIqMxViLrfInlC38tP+GylNGoqf
BNTFUKb23AK68TYoOfzK5+FS73BncNedArMLuy253IU1wRWlU64nQQwPwQ0ldOWxeFgwEGf/vISE
lMAOeJbt6isA7hijXsFVUEwIUExcjgsWUu/xcNufRYTp3Ly7FEWyUBpKy5ZZBnw//RDQYNfONamM
Ei1rKk198BOWS1NX8DcP/rPOhFaHATOkoCteHwxiPCT8bk7baBxdmQvwT3X/WqKEXVeL6GG9hjqz
92WaTnYgBRXSTKnQWTWBvzcI06cfd4Nw5slYn9peb0jhruHjfXHrZ1fZFz/bX7jZ5eSbzciNlQMB
Ao4nQdY9CmKQwanLGIFUeDoeASoC40CbxUltkNTiFv0cPqp0EdvroQU1x/Y6/1XJ7PGZGziAiZOa
s0ND5Ji/5VuuLXPUUGZyqGutgjWyUc6k8BAg9UXY391L2ksk9QFXnRbG15hTUQSKLpZp+yJgbXY/
h5xGGVvdSme3yVIZn3TERZ2rBMaKeKLuLCR1IOK+wnIlVR7qFSTPqBiApft7d2H/wQT5+BrQeBBo
nkD5Rz0kLqhstX82YRDl+0594+xnHOrBjhj8+GacREYdmEnw1PrAi2G6thG3XFY2bZy0S7b1AZsb
2Z8FhqKNlDE/lX0RpyyEyd20VU7vI8JIPR+pUMX5uegveBzHqqKlitjkLy6GwyS1NK2YYryGLoI8
flg4XuV9Khjt6T2L74q8dfwoiqngswfDc96bvKWNhvBCeoqi0pLiFG6Nq80aWu0SrIyKD3DGZeO+
2KZkDUcqXX+1jF9SfpzVKBA/6ep6h4JRXPQOIPJwVSHuZ2ImClitgvWGRvDU85dZ6JMkJhRoAXy9
K5cXXxUaMTNLn/IxVTSX+Ttaf9iCyAyT3r4WB7FLZChiNumglErNFt21XTFBTFR7bvjezs8NVuCq
y6Iyar2qDgK3MfB0E47QvuGL0xzyBEmH9vMfCXVqrp7IJ+vK1EcM9nQcFiwO4h0KwHURg9IsD65p
kfNainf3btQBjtz7FVivWy9A/jI6krwEFYN9HoOhW6Q1HtJ869HQwIXkRnyp2MbIaCCE+K9Kjw+T
0SV7BvzazOp1x/vnvbvbkBqCy9c2u5KqThBvclV7goQsuDMKXJkLQJyjkck1a0cBRQOdSbc2anJb
lWXDC07ir422SoDCrrL6kZ97iAO1/A0mo//pNHisa5k5iXf03cteOaeeVAUWkex4urgp7pG1d5KT
Mq1233wXbHjODpolbnkWxrSkk9QT5qjKLPjDMp4sCqZL40IcjXF1vjAdldtyApD0pX1bXBuFUmE4
ws2paThVZVzYYrns4VpO8fcQAkfEn9ji6rKWAyD+HHldlhyj7P1mCA5sLy47hW1UHSNqecam6EjN
Ql34MvfY+gUBO4TM1kbunaJL6MF69iITiZ2lv9Sl60Yt+YHcVp+4m6N0oEsF0B6mxtkWewSIM58q
U0m/hmgMA2Iic59OwmXbO6bSjgQ5GCeLhwU5pwOzBM8OLtEW0FDScLBovyuKgRhh7CiONN4x0nTR
hGzF8p12Sj2EsfKz5/f7HYa3hqifsYwPu+XpEWqTXcZx1dJhSXRwUZiqUCjT+u4LDm6DMbHtHyf8
wRD5jPr8fBsPTAE5uMREPD34IzITV01RdQIykQMLtC3JKDReYrmKVklz3uXqH2SbwuwyVJ42nf6E
vQXcf3FUG+8gSy+2kMCHHZPhCPPoFYzxsJn0UQv89ii0+Ke//KIWNQrDeMu1WXSwkBAs0uZuTI0N
BrbZNJ6iP6Z4+MzYd/XYxYMiIT8N9DtgGNI2g1BcoteowT+qIqyY9lZ7Lo9j7IDru9kvsMT+5BlR
0+g7u5H+7HC+xngS4ILJTozsWOMOJMmU43MOAWtfN03DMPB9D6Xc83Dp27C9UF4fVF0ZEsPU0zBG
bF2g0oodSevKFLqJcxwQ7zsTsuE1a68ce1OSgMKzSz5Rsm8I79DDPvIBP1FRyivhDGhtF/cwQh7Y
TubbqoXILohyL78jhjfAW54ZwVisfAZReLRPRBHZ7SUmwe98sG9yrJVzbYq3Cwf6ZA+xRj8nQW4X
EL9OWxH3UIglZDNx/zWluuRbdjG+N7aCWdC5Oa59NjknViFG7TOZ6Nw8Wo7LeEgGWjm61QpBBo08
GTRV4Q1dldg19QhX6uwqSnjOWOXeg0sHWp59Cdpy0WU2IsZ9d/9bONut0NxVyst/HGaz2QMr2NNd
luSrNfrBISWrOLcAi1jlb4hkC13PKaMijXecWPUUb+1JpOrl6CEn4phDa05NLSmTZeVXoOtNh4X1
UG5w1ZjS5IkyVdS4uFabYtzlF/wd/6yRmdWATGM8Dzw33xSYmolZRVjp6YEXgzHvok2YMSxgERJF
F7FJUoe0K+9nPB5EltB47/mZY9cbtge7maE3jr7W4K/2Fp75JdozY+gC6/QL++ymzYWQ++eQ32eq
rb9gCW3vC3Nd5piSj7jsBfyn3Rc6Dqt/6PJ0W83aCoL6uWKg/+Qdgd7h/eODRlMNtn869uh4+0NI
/PU4Wa9WrMzpHm5xnj11206f7NZS5OlBUnT+Pj5zEABPQJLbhiHcQgaywBivQSSnNDwVrlduVKTv
yu+FwidY5o+uASTqveJPEraHRy3x0tMqlJdyLq92y/PIq/e1COn8vg1J0sCncmo2CTznzSMas6mj
BGd+JGV+TCDC71nGwRk6FlZHH3bmX0Z1enoba6rVZH0lhIwsN4/g4aQrNJqSf4ZpLwcVCsyMbIKQ
A9hZBvQA+Grde2B8rE8/9zDGquWAsAtcc4WXt/EWfNB3NjBJD7xlKMs+StH6T9E5Tkagah1zrHT/
Rcv0Qn0XquEebw+ryTmQFpOU5XplcECJ1agMlZ85sJV3HieptNzfHCBZC0BHPBgJzxFN+1T3P9w7
mefpoyP8xSA7sojtGZFes/4pb2L/F/zns1asuQ5tSRvAg5pIMR8wZ2YwSPQ/qhy+PpFOaEtUT1vk
U46cb1sVtKL3AUF6S59DGJTRaXIR2F9ug394e1582D0bTaDq/YbejFZnNLM13K1vIoWbo8sWO85o
ao/wFZSvoxOyKsHOOzakR5dOoUhapNAy+huS0QKRn7tM5ziDsVPSWabW2GfaqUBClQQbHvAsiHbU
aQx0Tb3k/EIDrO+ijbWQG983xmePkVU22NLXoI2NPcZ+7WU4qJIVyESY+x22ukfeit15KCYfD72d
H5bvuKH+S1V/fAI5RS/yWTMh32QdTAT8DNvreT0nyVPuxzOYc3m4gcJ9+k6LxAHZAjDYQ8TfR9EQ
z7rlG9IvcnNI5YG1nIgCk6LNwyfYaF7PFvJvGd+ArXhKrjNa6exi93w3U88rz4og2X1/v7XQC7sz
IGEl/5lzKMyRNltfZLYjuNlC7jn1AHjo2bRF8GAJmMkETnRfTV6XWPecrCjFbrYWyj/zdmAZodKE
ul7KuprcagB3AR+Ca8FuzWqhgoYKN9REL8KrYc2xfF7JenBV0gBXeq9NajsvBfRipGBRPtKH3ilV
YGctluG2NPY5/sQKRzc10Wn8CXqp5XhlrbBZpjTSzZhaDYAR4dtA1yamaxWQpa8CkUmBOdpnsfb/
D2G2DtIP6n0F2Dwy/OQ1/tmDU2UprE1LVgCo2dbdqdr13I6VqO0XIDsSJNHW3xYs1TBO4VSkohqZ
ereaG/xA8BsWKzbSKl4n8/We/QcNZ0wugzwLznqwAgcd9cHmWbXBfrww4WyPvP3dTbjHRVCrkLOD
v3eU+IGkxAoisS7DQIMqnoVDFH47xGtT9v7Kjj9kbBxSd5ZHyQk2LA1fezAnGS/hs1Zw3tMGmMjI
K/w27QeBdz5EwFT7DSxH34hcsg9R2zwz7/3tdngCE3RcVlUHikV8Rw71Jdb5WtWGgoicpE7+3NM6
jlOdQ8Xry+bP3moUtM/Hxj35l6JGR3UFLMqWwuGvud5Q1KKsb3oS2Ldhih20vvZ981c/rhdZ0tZA
+77KlQDCIizyeOr/n7C+jttpKxufbAU5t3o5kCDRQEmjelqYqYfnNdxSF+BxDQcxzIyGvPznNgQy
ObYY55THAZ3LkuQveTcbRYdLDQOm+8OAdNKPqFAcs7FI9DcbMX350Yz4BImvHiOMem+sjjZwiDFR
iN4bFzeQ1ZWF7lrA0EaQ0K1P3i3k1m4lg89uYzs3NOvvPjTh8C4X7EnaSmm+66WftCKseg4sGSWk
AaN+xGdF8FABrc0E3s7YKTMuGKFyBKaQ5mhdT1USfIhvhumxOF2HJ3IrUUdcWTUxP/heo2vjzc8u
+bwHWHZTXQmJkypV++y9J0AJNsaqPJHgNgReHLTbjgxji3nIMcdDKPlJXjPG3ZtJGrgog+PMPtxs
8FV9ilRd3kHBTGPJOHeyUa+mapNIG9IFjdkX3DSvJ1cy1KmnPCjS+yxE8HYugNEU+ISpGSd4ABPz
2jbpgg4AA+asB9lfWYwszlAjaTME29xnnMWONYNMT+1YsF0cE2ISLC02D+lpq6oAjdU2o1DiCK4n
jL+74wU60dIwEyVoiBVCY1NV/jQ0oVJiPq3kSPvKdqnWbSuoOFl2Z4e4+FDytaVYjO2RgzcY4Cn3
tcryNw97um1JY+8tWwq2go/e6aoB5CEV3ZQ8hr0beQg4uSTfsyKzfOdHqrmq+9yVBxML5wOcqMlO
9HfTYsiFWRY9kHU3VrGf1dOEvabHi4HG8Eu7ezT0nxzqP/ND98U6Z4d61eVQmGwf7zgKyRAHvhfH
uy6dO+IiWDA57840eo0LAp+pcMR2hEeD68cvGR1w9hk337TQuuhSR3tU+Z+WyPH2jtXu3diZySoZ
l0C7gKjPkBBCfTchs5fqEVWHNi+7YRqi8LZeoN+NQlpxUDtRT/Pv6VP2vt8EjShQJrdR3I8tc9xu
ZWyCT5o9zXtlfQ7KikJPkQLgA3lQuOZQR+77cjnvdpPNt2cnmSqNhJwUs2D3g7bOQ2ZN847JK6Qj
ghsAgAsC5LWWb8AxdzlihyDEyiBhMEprnzu0X3+/QnA/B4iDEI0MxqntgnT/8y9QI0/tLy0LlGLF
1B97oIlRc+xBCo7K++hjXNx0GSmh+bjyJsJOYZsrON2avJjkpgPGXxUTDXkipWc0ET/FyA2sqTLs
bOZ8d1yyyGfq3lshAJ7YjsUDJ9Lt/BOvqmoC7MG325GNQpaibXInda2RehQmzwTh+q99zV9bOQhu
HepsY2ohr+CfOSTQjhHVnVXEaADOSO4k8vCJtYScbkBt6miWt6epHkW9m4gUHuaOgwwwVq03BYW3
Q1Y3HsYW2KUTIjJkFifFIpNmEeZlzt4Gm/CAbq4eMiYppaXgHUGjl3luLUbUmzNo0fWWWmKOsV+1
k+85UPdCVq3T//YQ/V7SVHyTXXrYGWZi2UFCKnxBSGJfYaS/8BEBkyTaaUWJvbVNkip7VxpEPUud
IBxe2e5oKVOKCfbVClQvXdXH3StKA4BKQ6Dq9Fmy0UQ1pJCc6dLe7TEDA1LkJ8e69lUqAJBoGWCl
oQWp+0p/N+arjvkictYj4XUUrik5m1NB4H39X3sqMTVpQP37yCO9ptED/KDb8O1D+FvZY2haXWHH
AUqdcQHWqx5WHeO6ujqEiduhODwRyI/NKnrRJuPv+KRUsgFVDdnKPHeqbSQpXyT3db7NT84boPxe
oGR9KiJo5AOPEMloc0yK8WvagawL17lvMUoqnFM7iblwtn4moIoSqBBkbV+vzT122jDJc5dReoXS
TZD5wvhjtGX1+rReChWpC6fcRAHtwgTog+vkdig3DoPrNyphDJxqIoTYyS9q8GIawgIBI8/gFL3J
qmK4TwndkDVlvhLYsmwzTtrNg0Cg6arnSxUfX0FONMmdKTp8c+t5U7nWAXdzMzqa6SGF20/OnBFZ
fzF7WyCIoLd8/VIPo0umcGRB0AL/NKw3z6opC5madDvhEFjg5pub/u2Al2SLOgO6FzYe/nNBgKNt
daqOHQa2jCxtRL+2qIi9Ew5axzM3gbac6Kwf/2pCSTub0b6CZfuqtBp3rmI3dBxWALbE/7MqhTup
gtxVjmOLElCLHQVhX8bC0LgEgyuEsgLnzharrz2weakOp5pA6r4T+kgz3C19BxqXZFvqFYSU9DLd
H6SBbGYKNZNfXEfdOHW4DgX83Mf3sw0Ct8sLgcZ+h07w0+6gn6MIICpnbwTVlpyz0e41uDtVD6VE
UAawyXMYbvJuXSLjsqoFVlmc1t+aLP8D61tpm5sk/TsSXNlnQgQ68KJoKP2gOBPmHR1tTFQrRgV2
MPkg6yxWgv3dpkGIkP08Yrc+ntS2FyioD54EcNwDY81lc+3uL3dgmsYjC5v8X8oHISyW5airXV5C
XmO4/2vmYzNTjxo/zKUS9NK0+Dc+7elUXcK6QQA7WgY22Y63Pjz4y6ABIUDTB3W4V5AN+QDcnkob
IovCWRqNqFwjO8KR/6/lhjafWF5GwZQpdVSY7DbOVG9U68U8F8rAukjbPPJXD1sXLrenPZ4f7hWq
+7vKtiMqjPyMfk24p2MosfMMggeSvVQ1Gg08BkckmkBIV14EGLmhXzM7FAgwpKpAUR80N3ofOMS0
FDVB0OjCR9nNkXfcIVKdZEKpzynvXMNuokE3rwCat3Jg/UVDF9SpvndcctmYiaGKI2TC+ahBt82A
SFAXKl3V7mwL7gILqCJ+VXLoQ7hDvwUTdmR2OTJel+i4VDVO26asDRlTDfHzheVO9rNi8Ipdda1o
SXqB14+YCfO6O+CCy7EG+KN8Q+L3WYFbw7oVTlwveMs1lvLetvlqwV95uEeEPIFuC6QBJPQMj4Fa
IIOjBj0IZ1cImyd1SeMaDwJEZrkOvxHupkRGR9k2lGRMeBNl9yH5iVETAs5zDsWk8mO9Y7KoBbqm
l8PbT0f8YrVXwips2xt33QaI1QOWi/rDNlnzabfW8ZwsPs4zwFVQvIjWD8azHLJMO5srdpxWAzHg
d9xxSU1zv5XIlr5foOR1E5VetOhiTbWufV20Np8zauiLelnNdQVD+Hvv/RapSpEeDYh8dp5vqtPD
YlxrsfYhn7yVIoTvWRRRcyPSqoZsiJifAZP5FmHamDPvWqqAEaQG3OuELRXqN6FdfNmAmLCn5H00
+PyK/lql1+GQ2ZYzRFQX/LMrVkcy1tLJttieHXwqrHbHYIfUsLO2VkUM6UcT8oPzyOSFjoTgIXdE
n2uPQxuFcHx8CXpS6rr5BR2quyGZq5B9zBe3fFBrJt5m/N+P10vEDMSvHhGLuwr4XNE7ewnebMRW
3g7XyuY3Kl3hSvRZ8HQgoQljwU9Li390WA7rY1SbV1VauKnRFAjnawydU4RkP+nacY975/nWrJv6
fvGbUxkqnObKHKn8EoCtEDUYXadZoVLLP7a/d/oomg4xtVEdKAOHKaOMSsEWs5lTZZ85k+eieSj6
ooO2V/DdyZ0VtfQyO0swihwR6dE2QOWFAQv5+RarG+86AC+c+vx8vT5h5DoEMB9iz/k4LXXdfRwR
TqKYXDfeXSSwObdmFqiobLqXQSMFe1VHE2kQOXMTCxWFoBtu4vhH9n4lmT0ORsP9T/J8ccG3sBVu
2cggDpT+XzELHQ6OSr+iah7dJVGXjF2gBg3XozxOHMLHWGv54JjXoEiRv9ihOGyqBavyKpu8zv8k
f/pyi4GNw2hBWxjIEVdrB0kfkyFZWZA7CAoX0qvzM9+08TNdoKCpIFq63AWSHaCUneJ0BQ1NKRX1
tm5pqCtaKsVODBH6xN9vMUDhbCkE1SQbHf/dpIO9Xem8jeitqJwoMOmGfzm3sdU1SAWFLS7IbXyo
iituwecGsAJDoxf11MdIQWvcmr0a3QEvtYgBYiB3GvvC+gVX6EqcGN/7lfNIjG49Fppaws1kNooh
NkZIOt14aRZlkJpR4S5oVY/+ZI5maCS4xKvuMFNU4lRrFzS8P45HV1+aiCm8hTCB6lzVGIhK0IL2
yzebproYnF68Pj+HOH7tqjkwpbcCDPqqql0iXYU2G41LSaSnSLnNikF38Qwlrdhl2TAkXP0IXlX8
copoyvQDNy49lPP6yPgAXUAPLnTPcDQzkwm/wi/ZyM21E0CQmDsY9w5+brD5nnXp+8zm2tZY9vfT
BPeBY/AvCLxFQj6KX2nK9V60OVNkH2C6TqwZASbcRzpo/SiaEEaVFHI300etLoLz8ctWgffH0xCB
VFguvkfpzsfLtpqhBQuMgDG9DiTt1FP4jYub7KzGClil948qltOi8sx2Xpbfz+HE4J/uBTwAmx2i
s6Zb8VSy9r1p2rSC5e7DcZsDR61lV4EMACxzDQkoVurus/5cVOKm+ERATfBrMQJyuV4AML6LV6gV
ZsRLu3GWeAr88laxGgalQ2feo6wzn4V2K0PTfzho6yqT8s/OZh4wQ6fBpSM8JRIx64tA3Ip2aMsx
IZqYyK8rjHd0clF0qs915iJM/xfHKi938+t6Ut65azt/y7CbfnuF5v+6eq0AHoXkAvZhiuiZP4ZV
qXU0ncs6wb9EoMcsDYeGS3BJ/oxF0beJ/0Ps6ZnfonwzZjs2HINJebLQsrj2dH4LhlOTOleDPsTn
QColeNMzpbvwhdWKJofvnlnCfYsPmqNE/pnO3nyilfOBeTzEyPgHRvm5/UIA5eVsYvOk1SFZc/Fg
om7wpJWDU197DCaebA43LVK+LQxFC3guSXlvG06bhS22l7vK6d9U9icOOlTmRerUNPoZg6C2czbW
60AJg9Y/Ud1JRhmtxJ/ZI2Ng7x++KX9e2ZC1t+W/LNUiXRe9fXQrHHS9V8aRIjOI5ERoja3vkASr
ogh1cde7NG/rAU1Kd9k6s6JKUSWU+rjgEj6dHLnQ+qOy/GzSfHTmil39bD5kyy0cTn1MKgAbUIMQ
IrKOuKBFYLpzXCC7g+4zC9TfipzV+yO66r7DY5w8HtDyqlLK+hff/ihfcGLQEAn6Zu/FE37zc4sZ
8ycRQl6ye6DpkQhRnzACoprlTHRlA3MXc2i09eiPxZfKiAmRfe6R0y/aEl7gksxVlEIifSKvZs+9
oj7EwCvVhQ/sJC99ZvT4ej9EpX8klVKCBePYK0k6SS5B+9dKP1Ie5ONEYE0JOKynpeQHfsRPbpUo
XOlm/X68DtlQ2EFC0ieLIV7Jz8qrFO7kqURbaTtrFtSzTdxuu92MQwJ1iX++FNBSLNIHR9D1Vb2t
PtrZWJ+atWZofi95Sb3NFzK/emmJr9e8yuAJpQplZxMp7lsReuyGmPnn6+KLaNFvC68lxh3EmXOy
+tss0ALvDwpj5TVymLKbYlEzIQU2D/PerPwQZF5JhNTNcIr1IHuwJV99+gfp+N6Z4Wkid8EGrnOV
j0zGK7EdYANSGz9ck1gVsknq2fGPRJluUtuM5enpYdl6kdS1ZKhMBarhkF3+jokasBTk2Lyo6o6D
je7IjGMgVBfoSQywnvbdfn+QFXl35B7URhXZH8L6RndNE2qeFLm/3zKIY5Biko92JQ0Z5lxB/ziw
NA0DIlnDPzTRtFDwjN3RYznB4Gnxe0I1CuHGHdC4u3CFdITmYwoBiz/YFWiwy1W7eFaxfzioEcdF
I21bbITzPbcRM8CfUPe46vyOvq4FnaYSes0LE0MrzVfo54brlaLu6/It12lwatZSDx8IIdiVPPyZ
q74I5EXl6vziNz7htcXRPaAV+yLMaEBy9AUQRMJNNaoAa+0V3KRtw4RccnmsCDlXsrc2YG0af9ZV
b/9bmppu3v+JV23PMxZ95rNtv+j+Qr/Nm7ZlpUbb/KIzimJDJhsdU5ciqNcxL2X9ACvjovWY5rdc
H8efdWQD/wymzxU3KP63dVjMpEfSBIx99+5zgqVc5uud0Fo277b1eIVFifrlcqFbCPSUONqDLbgJ
nCV0ObbM9qu8IobrShHSYDwK9E140zrutaf6zfJeWYNVYOERAOl3pE/G419w36aGMXvIO9WnfDCx
jDGnPPMivtGagUO3RyPj+SK2ZPSV4VQLb3u3PNfIttR4g5dxAEdUz7IuSSUtqTw9/DXtABucKgmc
1ZCd87nHmR2HsaAAyqELCwi1Sl6rOeQU2aju42omv5T7eUf88bXI4mROd0yiZmOgeXjXq/F+HTu1
+YbF+jZHdgNHW8Wy8wApVh9lRiehhc7k6PCWKSeDJuiTeEfQhHAtfGq0/DQRG7vmT16sBApq+OaZ
jpru7jAlabk1LuTopYVHldUS7klJQ0LR6Xpyo2Qxp91sWnj91Hx12AReT0F6KqDuiJRLxkCzq9RQ
xRa2YMG+Kj6RP6RFsGpoDeCMaODAVoowuY9sTQTrTcIv95YE94FcXgdhe9qcfl9gghBlmGGR6vTH
7/Ff3ebmzhmxiKFocZdp0q7qC5LsHGUp9Qh4PwX9e+TvO8P8OpwnH3uaZUlvGs/qCEYB4bIa69RI
yjlFLzhQUnY9jevdQnPmpkxYeUgRdhoQQ5mgXsQp3Q+b0d2Vd4aM/iKix49RqqMlJnOOZSmguvSn
NPt8PqCwy0a46ykQZctllH0NBhgXTolxyx9fPWgeGtMV/HIejH/omxL5sG4lSTX2b1PPJYLk8w+A
NhBQQFCPf2379yV3aRZsyhjr+hTy43f59mvycK92RMAzfTzfQx5QNJ67kSVmuMEaepVgRlINr1Ad
T77Vb1RrlxERGzNZHLHfHUo11nhmLS8+U1sFEw6rp04BGFY+QOH5YLmaWwVxo7mZFIldMfTwWbGA
asUuEZg91mrsAHIhNFaYfJYVobtP3JiZNcSVnWOgSNezowZkNnx1R+hpcAm411ab2gHbVX4z+Ein
zSDWT+ld37So+ZpGAHcH9d8oLZoUZ8c/WGs3CE5flECdCwINkkPnA9OCvlswtVfR6hGtAsXovwHn
y2ZH5FmHvvVVtuC7Xl0F9ZXVoBmdF9ZtGU3RHxkU8zrfSK6nv+FS3d4unh26wSpHDv8Ggu0c7W9K
t1dqj3IDiew55vdt/vdq2igF3JmtM0oR1s1DGfpIA6OVkJbbTImqrSA9uoosnKFJmLAJ68oaIDx7
wNO/5d6nH4U0tib3NI/OB0iTKZLiHEwWL9xVCkPDUf6iySDylfUzd603R1sFS/12oEupcXiEElnf
UWOWhUWh0hV3emzYsT7Jp+lw/+bp7cpNQzEOcigDSFLXt7Kq7ackOypyqdCsJtBgiNQCMoanog3l
aW/6f2ru5QSq4AQBJVjHmuWjZ3FXVKUUBGEJNOAO+MWpl/28x1M+E6R99SBHQc161xf69smkPXqr
ZnefgAQRlcaVBW4ccOFNZOVkfUDXgApzN4jYRwMX6Eq2pTwutrnubIKTxR4CCcVK22Lmy16D6+Ra
tSMK+GL924/meemgxrtswq8vrFipu9vvcBp6Hd8PHmI/9v5H17ftfjN+Cparkge7wx8Gdh71DjnQ
OjcK9/t6fH4z9TBG1+zexOF6VM5QLHJnXOqK0+oK7ON9uwP/xUwGt0oWU9M3avPsXQlAJbp/Y4kI
Ou+pdB9ZpEzKKMaw4hb+IYwkCDhg9kRSRW82F7ts44of1dol76lF+b/nA9H7gSQU1VysqfVtNBUC
IkrYAMZElxcvLdyfXacDR9AZF+VwqRyjFIdUreIxJl7wkT5YrbFJ6HCfxb9/Ejny2UmHe+PmHuPw
vy8/f4lt6/aapNI+/G0kx54s5k4E/ohndi6+fuOmf2NA8/7+ElmPuzTl6RweFRERvKcrW4NzkFYV
xaI4GPAZORlqG9rs4JIJyYRp9+tgLsvK/AR6nUS02vt8vHex/ZAlOLNeGYVwTqtcT4uPytK3VOBv
nFKEh6wH/NmMdUdFZ4HzL/IL6E1iSU1epI7cXkrO/pTqJ7WgD+c87sGRZOl4IdyO9BP+OaKE9tqK
DWYDnExmZGYrvMfJjwKufBjHkTOywHRDlKWGcec8p1fIJJgLNRDfl4jkiPe0Cg6zu4TONXSSOl4x
D14fYrX7sD5EQnHlgDcKUMhYs1fUH5rot3yAfuQI9UBwWNENU3aj06b7dlY/x1jNPhmVdLIl6GVr
9In4gzfvDuts3JexkXGtVwNVeQ1pW2NeTlBgKdbPWfkaG1ONrgg9v7wqKWkT2wQfb7JUfenn96mv
jB1Y5kEG9Xf2ibMopuCqDHR7jljmSAYpMOqki5dVV7E2JfddY/XsJkQqCUP4aEuKaW6oeLaHKB9k
1zEx/hOqzN9raeTlEAXvjO2GAx74y/bhJSr6ITCld6+rFr74wiFuyNax+Zfz1+Owld29KroL2znO
SsV4I9vidP8mnVdl1WSCTcFZOwc0ln/QYo9DTGnLtRHCKITZO4vTmxWHGdL4dftqp9EvWseF9Rvq
svd1jO8v1XasMr+VynhPxOhdoepA//Ryy/xz7r8l9IX0kz30KbOdUhbNExJtdGQ8IKjj9UMArJ8t
nK7IgE+BTifySlxe3+4kazQlkfo0LOx7OvF/Pg3Y/3ID8IGwp4j0QwUc/BpnrRc6YwSUHW11ee3H
ptYPbF9f3ZIsnDIj71mn/nsoRD0d+BKinUTPidgNreq9sJZxzhW7ZRVBtfKqQqNRdg3pO60+2pto
UAOY6PAqSSsZbE6Xt7ih5vvcjFZAmbPuVB7ZJGbT1MUsGZyA3k6Z9no2VPuFDovGjLXP9ZLwrVKv
USftCzgjqgd4/zaFMu31K8vIfZJcaGWUALqKJ8sLnijbIKpU2DajYw/SevdmLWJTN+84wN/2OAeq
disTQL4pfkZUXYCiLOlTDYVsG2xG75TBju8YMa39Hh9KW3Vnora9xJ5fBDX/Z9yAMrpirv22Yc2F
hRmhtcdRnMhjvWWsxGvX2ihl54JCOQ/fo233AtynL97KXOEwoQGkAowNuv2P5WyWDegiVkz7/zDT
oL6lxJJPzxXZp5SR
`protect end_protected
