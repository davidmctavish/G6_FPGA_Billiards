`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EmlDkfjnericRINUP0NXhs3k6FoOztbxV7mmnH9pOaFcNKVDDbi+RSu2zjWyr6qRmwA1UuVsG7M8
A9xyFDfhfw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mvEq+zOqIsQTUeiGnwsB10ppFe6UA00gjFxgDQnltoyeYMbBKulvjgs8ng38te+wSVhCpLEHxs2R
8lUGd9G8ysH3/rxQAx+QakxNQuIxIK/B69UIU8A2+nVdt8XyHVguFY9lhnaCda3CQasdhxUVRU3g
PEYgzN3vY8QZhuel3Ic=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OUT1hmH4tbzVQ3AVYQJp/uNDOJiLMwg0uoYgECWEkTK2ZU2wqth80CWnZbcPrAQ1tEPNuJr2HbYP
cvWErbhsZl0/jnYZuUl4O9gh0DKhBV+6rAZD3cmQzMWQGPNCy0C4Jmz17a4Q7aDUg5VysiIQxCeK
ttm6I2+pDw36C6idBbK0VzivhQlzvGZm0OwVHZWPhmtnsZDsg16LMTDbTALz6ZKEHKE2MfBCb+vl
yDe2KH3upzWx2p7IbhEmGeSiZDtWWAKX0jc7XzYLKsjiwtIWT71Oh+QNxgkl6NlioqaBqrYOkLaw
ohwUvhnrN+wsWIiD4fDGdtgsO4rPtqkPvNuhvQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EnBHekLVCbYM+gBRUEzs2p6OtxfaVW/3MTv9P1y2W6z4VOlRqKXb2x1BFk7EDTk9VCfTRUzq9Vog
qgzz59XkoVOIbKAhk16v9KajOxERFNueWK6xhf5mqu4bvT+XNTDf4yyuE6Fh31WIersBpzCrzMku
Wiu5PreleyVvxbm2OME=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
toFYElCg7jIY0FzS0gX4waQz9/gKz0uM4/THXeAtz8f/S9TFEXZjRRXyWFRCnQsxVsNSVljtLtmO
vdTh5/mWn+6NRkzFPX7T2Mw7RPNp/ZVxZzPwNm9Hk4QSNuCpO+GzELYBaw4UyP1CQuCW697FkYEF
4R0ZpEOpGF6AXq/np31qgWUxDGMadVrFzGuyzuG8zKnB5RRbxhdhx0NAbImZ2h2R1o1Egm08UQbk
PQmXyGaEdBbKusufy266zby6MyBXmxkyG1IE8VPpoDnDKarfAYk7iwvG8vV6IJUcC2OpsT1k2vc/
W3D/os/Xa7pCcXCypGB8veS+7DuiN2PAE5fJuQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6224)
`protect data_block
zKsrmuyV85lRwAsnH0voObeiNjToKlpv4gkaz7gn6a93+XQMivSqn9UkjpcYUR3gepfvBGQlnFYJ
ej2d+jg5em+50d1w736BKUPkBvNYPvbLs85aBzrKKtt6lWrY3TdIsNkr7CyFC/ZiQPD/+kOGfdZJ
ysV0GPN0uZeR1lUFVw4tXsp3ud++oFw32BGgnSbic61EMEBgU+8NSe5yLS2XTr0EJR5dQUUcuj0z
6lp8ftlegjI1tVIL5mW/E66PMMRc/EIr1z5MdPxhAkP4PJ5lyZ1Bz7sx4wu7XGcWFaB/E40s+j9A
ixLHnJ0o08F3X/8OFJ8NiSNXdsniqyOuhg8JGK6Xeo7EtruUgI75h2UBJ47pWcZe2HURRkvbLxSd
Weubp2Xb6btgggvqmZn4GKBQdi+xR5CK/3PMEZkaXWkGa7is7lNlUaPCNd1sZGY4UmVVAUJrcOr1
x5kkv0owHB4+2o8pUSUPPK5LnCFNlIbL88Z/OOoN34QU9npPXmmds7zrb7QKdmPIDKDeApXb/c+u
pmFECmE2C18mF4+xrM8XPFNzyZKQnHE3Mpc+Z3qSHRT6n+cFldlaytc1am/uUGJ/887LGTaGhvbz
jQReanI/Ixp2o3R2opUUAWh0R6ujZE91wapelGbCUboh88W7D/xem6Wy381Txv8iOs4ZqCYyB7Rd
NEfhQR86+6Zjlk4D2IaOAQov3oKhbRckyT+HiseiRxaZ9w0/nPQ4Su/5Ygyw28iZkH9U0/ruNHV7
P8gUyLS8Al3olTDoWLDtk0tDb4xmX97eMb6B2y9LBF7KAMiFqfDR8k/Pz7SYYUtJMATAhvj2YLZg
lG0I6v6PgCYX8CSRzx8O2ty0WvQ9MKaV/qX/RNWtAC/lzkF/y0OH3W+lRolMp8qTxN/Q/2TJ2bnh
ySF7QjO9Aq5b6UduMblCXGjgMR+P5vhVk7FoM1RqLnHKO4sRuBhUods+fZItJr0o1sNjTEhMsXAc
6b+49ckAxwn0VZKTBRw8HlebVQgC0RYnT6Uw+mvyThrD4rziFoJXkmPDlmIBXzAkNCa2nUp62/L7
NvDQRyf2tf4mjSXNcIv4OjV7ETgFe0xJbviqZLkjcnEhoFFu0CN1NqqHwSsAks8jSYVHnX53hAir
chpHP5lqlFOVkKEK+T7KGMDW3o789/6i5ZUzELOG4hmoh6126aQ1kTHvZcKI+O5hryDR+v+8us3x
9zdfqM1HXb7OVPzF0CvATDZoTURsJm2ffTNmKT/G9ayEacG5hqPRSJI5sli8CnlBZZqsFcCK8dkR
j0o+q+skHpdKH8FLnw7mLnHGuQGwSTN0zCXMCTpjutKMm/SZdmNK9rHBybRQFSbxMkrtSeeHMaKa
vyn+hCnzfG938oyLm9hi/sMoCkqZ0MbLakC+lwFHB8H0g8XnZQ1IGYsOiyoGf07zeB8aLv+qilwl
Z+fco9ALl7r68dqMwPexSC7R3vatq5JOEI2gXt2L4KEg4aKI9bStZvf61wJyMisxnWkhEyburUeI
p8/gyzAfw6Pex0oG+R6mLLclpbrcvoHqyxU1iq9m2pUK+2+ftkDj28LdBtLGpX2oGMfxhm+GlBYN
CgbVLvq/yJJpUSA4ItZxiCfCZRPvGVlahBjXxrA0pYMqD7zPNdOljMFBjZkaUeYuNaVgcv821iPK
BZghteiHhGHfJpOqKuui4Vg9vRQ1AdwS/vBfRA2UUX931WjBXDONo74VLZvlkI9PnIoDkclCeDGd
z8VkxvPsYf9/qjcG25MtwmLdHuL/bkmYC5shP2XnHxC9ar8SlLTBBCrgCoKjw++x0lXdl7/rYRn4
0hZYDixNYHCUT8ZI1KqmlinYfc+JUpYu+XfDV1vGV+wIqijJ67wRM3LQUYBC9AVVLCPyTPbA+qjJ
ktlAfGX5AD/4f7fGn5CGIASWxqb7z+3VxAvLK6li8/Ac/OaqUrjKdQebIve7DZcR4/7jV47f2udx
2XBE7VJDnDXIGWc+m7o8BE1cmYiWG+37bOJH/pagCpYR9+Wmpz3T/cJx2AOgJW7xaIf93+bxIJb6
d49jE79G/33iFxKGVLAnW75Q7H8mBV5GM+JML/3WI1uAcfGBlejGkxcCCvQe+LtR9OcxSovPpTiN
F4lHb9NnCgAdWed8Rrkxv0OQF8zTuereIH03Z/Pj9myV94pyK19L1l5eC6S3cLzBjXbVn6YhT5TB
7djMet9cnmJrhyk8mUffQLVgmPl5zBwjUIE2wQSscRqRabyAvkf8zp4bsuJqeByjqzWhZx8reEBT
4yogARmoC9y8jZR0X6bqqx/GgYke0jc79A87N8Z86CVOsKP3hqN/O2FaGS8qxVTxiUReLqzgdXZh
+ZmkV7Ml96CD/2K9fums0TPxAZjQchYQB4Pk+K4oBCGs2HXyfFmV04HbZXmpwTUu34xfO3VFO0UJ
5Aflx24NgTMlbht0G6vDm6r6Ai0FitfkLyVoEEAb3dQsb5U0bwmzDYg29GGes1FIVlmuddXda81R
cWIMtszetzOUfnBIujBVzRu4d1R1Pm+pUFVDdNpW35+DfbRaUpjZs6mno8GqLi9eUWW1bcSzXfAa
KbSGRxFj4/ej0v7fGA7AumZ6aqg+E0u7BcVcLYCzzS6E3FJQPbDx3nLy9bi5xA4pZr5h62efhlG1
I2sPd8SGER8Gd8cGj51rYutDCMTU8cHWst+Hyi4dFDJ2CmoeEZLnskuiHRJ3sppyKo7vrcVZyNbt
rYUD/hTNvA6fzeu00EyW+MUBUHQp8KKcsqAfoy61YUghzlp9kz09GCLrp913MOoN0w7dJYq/l86E
sRTHg2xQp7sNtZ1971MBLcD/G9FfT78bcO9lKOU4jlykVCtcMSf7yUVE/Yn6aqcMX3q5B9v7YOxX
ezTMewjWkwicVClExGrNBVwzHGWIJ6E0UpyEWGfsZaQJpoOkXO50QZ6YWSGZAnuzZr6itndwJ7qf
GIV7JfErqA8iyKYKD9A4pjB8x0XcwYQajQadceZEuihcOIjBi4e1MukVZb6zbIjWcJdsKpnOmuod
fX6qOwfmLkSMO3dBcHooxc/m0v1ZoOcFzeP9acio4ZSYlhXEyV30AUJQLZtGCr/D0DFioDEKhvII
/REIYQlw0wqa/yHwmJI+E518UIX/IzGvhuFkkPbXffcRodwDe8eDrffqBDwR94us7l3xPxSswNs9
HWXW6Ckh0B9gGctSK900NudQTz0aBM/74jgieQxxQDcg1pxl0j/V1T2EGV5DGPubgHFkqHRKijZc
DDOl7vHxzHxtWMinqu/+kOLTt22OgQKUypSy8qDArG89wiTYS42pb3GnbzQ0yjpJGy1rmPvJmmUY
LIiDwA6puCiMlEzDm2NM1OaNSSmi21Q4PZMaeQgOx4APxwjgf+S6ifCV9mVsHqTug4lxQpmygzI+
25wZQSs2cuHR855UvRci2mMbZv0c/ORpJ8wTB6pBUqXZ3axrI/ewexL4I1nULKkZslRGC64wDTmQ
B8ZP4Qz/pRsONPZ7KuazHIo+5OeeM2Go3ij/r4y333xpW73RZcmxEX4vYwkuBHyfM/bGP5j5RZNa
5TQqgaVG3SsLWnBolNSImp7xObPXSyRYVsaf+v6mmbDs0H2tZDZM0hjAG4kQorLiAE4GEyFDsgKP
2I8cEr9/js8se/DexbTHjIzZK4MmDQpKzr1LwnJl+8GbSMctPiKo9cLtV23D6mYl5PdEe4NyW7i/
kVbKFeTtRyh7M8Le2kei9LzpKOnz4xltOAyPGT3YOIOnaLEdcRvtwLM6oJOTc9zV7ZjBokMZkcVZ
KA6MSGmexAfaJSWcss4a25J3OkkuBkf7VtP5dByF73UwlFSct6SJfnxT0wAM0FOjuAdgwbI/RLyi
K+vHR+ygqND1nig2KjLRtDwEGxYgAX+RRG5uXm3ocxUwFZvM2kphAc1kZjhxGTHbJgcw1sGn6X6J
41vC+F8Dfs0ozODcMeXCNKw4E5Yrqb6vwzU4CmGHsob/LW1GoAQRmm+6bxp9LYTTCes08Cqxo16j
4b++mIm0O6wbtmErkTnz+4VPV5sLSoScdxTTjBUYOs5+ifbKf2fmbOc0DHytHMdiqJJDwUD44tWY
o4nEHiGkhLkxL8GRoSv2YHiXMl7qp8WBKwUanYCaZI+3svBznrJm/sBw+rDpotEcN4Q8INqvRnx6
42MgGUusvJ57iZDbz2URBHrG4XnUUMp4mQU/Cte/C/naR6Z6AWQvu/d5SrM/2JkHxx5Woij9zred
K4KCfZJU9zs97mR/NePNOvw1VYOgk/kOhKu+JBRcpaOqJ3Bqf7Mfofvn+1azIntjHbXhAqtasgTU
4+RQE5X3bR1HvQUa1NTirYd4PTwysd/dk5fyoTLEIU6cfhQLuL93DKuFB2xd7XPWdu0cyZkwfDQ8
OeIaFz31nBfVGljc4uw4/noge06zJ10piw4l45rA6aw2W8KwMmhLSGWgvdfN8M+UEbd17EtPwvPP
K+0ZY4MrbMnML1nH3rOo+5GdZ+kpug4QjTP/dKLjIFhoAtfVBDniHJ1e4YFyNRLWk6iESWd8nObk
UAN2vI8T/8rUIL8/Y3m2+4o5pwTV+YmZPNeJ5ar74ofwBZuVt3RhSuwJigs7sQsE9n2NqviqhVFD
u48KSUqnPKRObHQRstYpYkFvZDPD3BQGBjxw0UodLT6hwYq293olwuhnIsQ+aZEqw1jhUbtZse0h
VjGBBP1z50kKb5wN5O1fRFIWtp1GxIRxv53tGJcAaa9eF6U1A6sFiX/aD5pgPwlpKF5tzhIJWLmf
ycB0DY/hQhGleaYCtlQkn1cr/1BkPRTMpDIwpDKQGjzWVfANW3v6w+jyQDKjab7eFQAyQDgv+sjo
JlZliWGqcJZ7STUbMZLKSVU+86sUo5RxviAdFCo7N5WOtjXQ/tsx+Rj9ZabQ7RQayHs3toh88dGE
z0TPpweaT5NfxRqRWy9/gZuZBJtPmLVOuo+VzIX4Z5p82DqQoCEIdKK9AW6dmFvRkmtWkL2XHPbC
M1iftZOBHBl+S7ZCmWEzg+HaAdXLOj0WyFY+IXPTxmgKLwr5HeigegNTCY6iYsNZU4kVt9eEBBNz
+IfR0cl7/qhS0T8xNSrN9Mr9qvwRCeALpnI6vbE7ksiWj0BBNm9vTR/eLZkOWqBE/R1VT0hqOu/C
XDJs10QXYBXavdszah4O+P4jRYUlL4IqMqum12v5b6BYfosCfHTsg28Qh67imNHFJMN5AYNTnE/k
H8CTpfNhJO5Z6WYJDdRSi/QUfhSSFAK+rIvR85W/su+AlG0y1coNaGZ1t/CXfvlvX8MVSIjscscL
Df6BG+oZEWuXUiyG3+csgiE2HPKSZL0sSyDacwoKrxG8Er+F7X2X+BzQ8jL3vj18D8kPp5V+LMpe
SC4AzS9FT9gF+E3+t7oS5dVn6YRukH0YdpsX6TRK7Y89lYnaN8lvMUJ9VSCIPiR6rdBapIU2htso
B7WIbW3BojTp/WEG8xN4L3AN5dS5jYp+AdBEwkEIJ7YN3v5SV41TZfkTkbnGlRLQrPVlm0J9YZDQ
c9uDQ8TMIjghqK9WomkmNhBJzlbKgpc4neQmaCYeM9b/dGDsgR4pMiyGZc1OOE0fzHIDJc9v1W1u
LGBvTgqEgHxDSuZhQRUqzel6gMdxLsbVXuF2+Az14rRVDmD48RnAPebJTnnyZFh2TpqvudHX36Gy
89tsVVndlScyJfvmCUkhmx3BzAeT4TiM1BqtLWUeOHzS6Qne6W9GvW1EXt9kP/noh55DHnYN6J5h
oN8ivjrupX92ZqSuDY14YWdc0Uw9xgsiT88Whl7Y62osVlh3rlhQO/QEP4v6QYa9jzqmmENEswkz
ja351h5nzD5LY9eBZl3IQC7ZOsCFjrBpOhD0V/wnWIyHqNrbx1bJCPQyRtZowDEcAl7imC/mx+Ap
3EfZQ9QsRwI+AjZZ5x2U9ArjYDY7DW6jgi8o1jTDRmmOE2z+Oj23h/AjY3WpR+PfvBNYzbgsdyM7
cvJVXQVvj1v27KwNVGzncHLbTCyNVW1CTXiUwWZkbhlcXjrngYtVuR7GkLgQlKYHblPiG7T9kOHr
gGFbJahizaY2QybsnUNnk5A22SVJ2i0TQxCbJNrXqqbYQMI3uBI4LDswluuQvZxYMWVvaQRPJCm7
kgyn42KsfYfJ7+jZDoJDai45/5NkWIWOegyBsIpltheB0v5Jfjn8Fm1sWV9nXOYNmZGwlrqf+e9h
8yFwsOaQVCIrUYNX3AtyBWCvSfB756JAgVtgei/99sXECcszOOXnWWFYEils3Rt08VD2Hvv++2Zx
jyP4scQ7y8A48ZvL8TCSeoBMgKMy0LFnku9MmCNN9zcUHGLjZY4x4M+NcIOQx0QkZ+PHE9fzWYxI
/61cqnSZ1ukjKN5iXqVRqEWhejhENxQ+3+wAnJ8ezp71rcnaLaFFl4XEVvNDi1ohrZfQg5mNYRej
k73/DxxqMqW/3aZdS10OFFGIC2clqtIA5Ibzh8m7RVzudc77THkYui0wC+lB6x3Pc7mfEKvigPWy
RNuo/W3J5nyI2Nf4+IbhxWFk8bfSEhH7NXdTLbWtXiLd8PDxiBolj0+PhqqbBiL8JEljW5PG2Pse
0OfKbp4qSqZfs5pB4pYcXYqkgbGm0ijfhL9CuKBXwT8mbzBATXJ5VRrngVUd8WEKyMXYmWmGfE8j
tk9oC3uOO0csehJWzmQn0MLEED2mc2dxWOsOjwxGv7HA4TQ6cg5HZ4QwtYvbCUV2YyZbvWgDozVL
TYcjNzy4GHk2er/fB2p3rAi00X5SbDKrjQqJbqhpWIVMxD4y22xtnpGjURxufIn2d5I1ROz4KRD9
jKMMg5HvrTJ0SeOqayB00YpJeqWu8Z5Ujh7PPjBP/mnT4rQs5N96HIP9hmLgMZ76rP3RmVXYNcCj
//faYSeiiK7wihJUMEVLWPY42x013kstaTn/4HpZPa3S1yrZId4b7tVJlW9Qn4Oggoy8KZIgUppb
HhTAyvC6HlJRzT3BFp+Wl4FNhO4567I5TEoDqCkCJRQfUEdw/TdPQXvPDDtXSUCCnstNEpC98f63
Dh3tBExnIzfKEikgwmrC9k/fTwXpx+bf757jQaQVwuYK5j24ipHZo5yACODvrYRbVBF/tqrXtfr8
x2BDekO7eERtMs0LzZNckruSF6hILEuCSnAOxwIs61wwDyceXCnh4aPgOT3qsXpO/a8YMWYa7+Hw
YVIui0Ku/9GDFV8OoqtKo8v7SKuLrPGNke7YUMQI26DVPpf6nAIZbUf43hz/sFIX5B9k9MpLLP90
IcUeHb8TZ4euG2xvPf49XY0kmNAhAM/PaMhKzu4mE71bC/BWeYGvW7S0kG5Wu/rXHw2f11cvFPHj
Vt13EfDlroe8ZGc9Z6LprlEt3KzDcq4/UpAJgiIhwoqVmwk/tA0lA9zw9ZAV3QPSGLj3swDvO+oR
zFWbaDTNNUBkRfE46LpkbhegHK9VBOpHkq89rD2rvlXnKymbJNGXaCZlTya/YUU9lQF7zN/ULHnz
OpwBan59l1eLZ98OO1bz3KcKmqX7DvfPJYKKB0ADfxAHdtLiayRCDyuUMDVmHlasLzq0jXKL3OcD
VgJezrXN6JqvAEdJRH21IdXaVyBrk74d1ftj+IcJDNLpCxUZtHHMUwy4Nhk7VX3ZyQCQ+7rvMs1B
FwVklU/ItSFZJI+fqVhTZmnQhiKUgau9A0JDbith08/i1sqEUKUM5vCDM3jdNykY2YjUyMR2pmS0
KK2SLZjS1nZ03CXOWMmF2ogDcQNFCBVCLPyZtor+SgMc4wHplABQYlaCPTC+TXLNmVVVlz47GjHy
8zCbCFrXaFie/g39lzNdI4NSEM9asGKXYkam8yztU6XSr4p64LLc7+GM9Gen2pFVzBScTughnR8n
0NjcMZS3CXKtCDo0oRP5a0i3svqEXkYm6MBciajIJyvBM8AAc1Wa+lW5LgnMECSk+ss4lDQKoKks
fifMcCBDMO4PjuOLHkEDlgQfQOqxRD60oLDrOojK5J/J2ZU/IIlljvhZAgQ9nwxpZs8Gxos2o0zQ
soVP8uc/fgmV4bAggYUpni+0XGPJr5I0wBAI76mAGLdX5Wov55tOfn5EQRSD5BxKMvHvlJbVOOrv
C3HGbzTDC6biXE5Avpm9b6h+XpGXd5CsYMdw7P4HJuckjG0h0f6eJ/ZshwemchREHVHFvYHSF2YJ
At4CuW74mDKB9aB7yu7MajSYb1FRvggeHhnyYfprSv0je8H2DPnv9P+2nPmXecuvFo4gJfpYL5Pw
ZCawFB6yp1C/V9o=
`protect end_protected
