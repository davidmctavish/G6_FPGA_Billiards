`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
q53PV91zSiMzafMQzq6bTTnhgk/4gmdrbACpSP2hbMFS915J9sQTvAtLWTq/IdVHKS1DO1hD6t7S
qTps4EcN6Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DdnSjM+idLjuNrTM4atgOM5uWSwWNCh3ZoGFxY2xlC1EDqs+1Zd4UGzVEWXWByXZCHO39JNtf+pW
MTABHBiDXPEuKdc9yMyOUzopvX6wyIT43Pn7plqVVxYsBqGocQu1i1hk4+7Ki2kgnkFRNOh4CERL
wQlRcfZPkPMlhkl0mPo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dBVYsRrjyV0l49VTcsmRv5zn+/z1dTsPQiLy+8tpe1XtszrEM6yAC5p7NkIPWZ4VELMAJUj5kk2j
UJF65hk9OZ49l8o1lB5660Ua0NbKnXKxoJZsKCPqK0Aaxvf/6lg3padR2+47QXagqAEdeT0vDFcM
b30YBfcERk2zPnyMojdkVd/qPEEjtYfuvWLcIy2Z8Is60WwSiy/ux59nhMCfSMOhxrNMAS8n7aTz
+E5H0O/KrqQ8N/P6aZcdYQqW0+MfsYFds90iCZNN2PDp9UeA0TeqI5DUim3gV/lJlfSKppCTO62f
ZdzaekVlq/xcpZ/pC5wQFU0vWDPnroTSB+Gz+A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P6YXpW+RnwsbxjhCG0YzxBZnsPLdlYtLyoZoWLecEtf3FmcY/EW/rWeUdBnl5L9Ty1x1x2Ghm7xj
+qMllqyDgyiqlVCpeOm32mvg0j9i5+zlGCRvpGWcCMogkQzW4SMPc3UkNtMwIEuimkHb1M9HR55w
5e8L0JJdfl5Afp+Qrsw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gPLP+F75vyN/2gShBF1JPgrtIjmacZXyAdYhhZP0GrFlCIFR86y711f7h+puZ/5sFNxAfPwZ6sG0
lqrLvmn1S0r7o889NqbeW8gk2ggw4aOAN0NHOVb6lrNSHHB2KsdMA/nAbftElMIapsLtJ4fBs/Vg
KU8yAgjmDB1MUI461FKzFuuidRDgJqEK5MOpGknHZV1AlMPB4lv1J+VG6KCty63ZEMf0N6bKuCA/
1tLRAnAyd6SZBkoF6mgGbN23ly2ZSz1eTSgOfSak0RvQNRyVogNBru0C8S+fNFCh7NHE/6giXNYT
rIVsBm+/AAKNaIvzJMJmWgplcjRMFgMxa5TQew==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12480)
`protect data_block
ldBAwWE18CgOw3YoBWNNCFirLlWVm1rvSEFpTcDeLLwUhzjdFj43MNZuVJGMe1HXTKNxbJ+MSt8P
syErsaSZKYFuxf9r62Oi+GD8WaZ921I3/9kpT99UqUBwSILSYP74VptePz2syCSnmB7DtSjmJAgp
a/mC8wxQ1vwJ2WF4Pl8kq6hkw3LefcoCMqAuJ9sXRRFspKjc2VZrDdlKzE4aGkm/8zMmusnE8iKs
KKKAgrZ1kJDgFNmqWJik4umkQLuUETBuMCeN3GJB3BOq1MxdQ9jfEtpWTcxAEGp7WISOS6YGjSMe
JLVfXluToqaOgT3/lPM1AocMN09nrZye+Dw0pWzxcnosZYpK/9s0GfUsbZDQZS/SuUaJrIg2+3gI
Xzh8iBmKF5oRi4JpCcWSvZ/IB7Dou6K3ik6veAdX/r0r9BQ2+2Hu2d33+RNHAu9qUVx+xJUt6v0Z
SFEwAwmWyNAhP/07IFdy0vvu2QPDf6WJE+ZGoi4K1a/b8vpoMCnRNW5slc0D4NIyJVvScABVu/35
HEbl5CGWBeUW7/hV+M8kHq4ry4467Sec1zgu/6hhLz+zmqNnJyfCOpncwgqXa1rgN2FWESsjurQK
kp6Gr9AvR1e2UyjzKw8WMDda8yZy5II2FU34Kt4I1iG5tVL+4SHtVOquxCIpzg8ofXfB400dxe3Q
B3thIjR7JseEGQRRTPEH58AOIVfn9s/52Nu5Ofct+pcE6BGvpZQcVXO7tx6TyIpSjD/oipPrHDA+
S0p7FaR3FbvkQr18bfptpARpN0EDdF1ob4799V7vd2tqgBfPqDHVMPlQ41CfTApar+pG4WKYWvyh
rfwys7LJop5fv20LeUw6o5vVOZHMLXMH3FUUsJWDiTRrK0qX8N03ZeL7gq3ya8ML1mI3dWVUxvSX
2WVII3te0V77XZcaXtP0wJzYawI0D0c+afFaAMn+JX99xJx3i6k3eouxOLAIBkCNBr2T9aMo6BVc
vkqER73/aBGo0mfM4IsDikYahVdLjTwMxyFlHDUuGYNxwg3YXHj4VOV7z9oGGa212lnG35dw+LbO
ROinUP38/tvqdQeUUR/Cvrt/oDUcrNMm7ssosI9CrQKe4hANCAM1z8DUkMwuGmQJmi6euMj7rE67
Np7vkJxRFuBr6+liNxoa0AdjQpvVDp8K50QuzOFICJwfNTqbfyT6spWmj+jxFQYqLbsPHE+bLJc4
Nsv0CrNbAjbJtRJ9/uEEGWaBx8aS78qIhBLDHkEv7SjehiBwiFLWfSfdlyFdovVMaphlMIykZ0xF
bA4XFGGvngJb3w9Z9I5YpeXXh3CgGDBQ9nOpTYmBh92ciTgGjAyazOMuLHKGHuziIzSSJ6YEIhUq
LPYUaZ6LGFyzHoQm90GET6AIVeXwZ3Y1crPO6ZNBStNu+4R4vrtGHY+DKnEe8XphorN5C5u5Na2l
Am8gkqnz7n6iaJC1iV+tm7Lp3zKAxJ+2Sy3t2jnDproc4ivbuprQ0UNqDjtwKFcpO1Dk76ZN0ehz
cUlPvyYcfOiqKn9Y+FqTakmavZsNUijW6fve9kxR3DXAx9FkIUKipWqN/dY4ISknYOlvedAmbTgi
Bs7/+554JrgpBYL2DyXCFmMQ+7RrH2SxK4NVqHrwDVkNPZSl07CCIjLmNUbdH2x08ljqJqTo1wBo
axq12PNfvKXZX/bz6egpeFCxuJYHakKjurxvnLdtBIuHPOJx+2jjk+QuXH6agy3THpMm06UpEdhd
J5sciJo4goVsZ1gThAoc+d/if10xqt/i7DulDIzARxcrjKvMZUC7bNMtl94Enyq6NrBEK/R33CVw
0LjH9qZGT2phqzZM9tFeXYuXWJYcy5HjpQaRmRa9ums46l5Bv/l90SLTYlFWrZGhFnRENpqULPHq
KYU77jR6v+Xj+xclp0zDTh12LkTAk5rKIJVW9gX5jKF/GnSPYEu89+C+I4LRk9sN8OMFLRvjn6Nr
zSTwgZDRGORnrqoGsGtgF+IXNF6/U7v4zBP3sVQEo4GH/2li6SbHo95Q4z0X8C/cQ4HcJLbv11zz
PLE9Run3in9C9mctXLCpeN0cD+vgiSXy29pvZ2i4pMK00/Sb8BvsjBvlcj0fIRnPc44Hczh6RU8u
tPDX2HmXXRwr/tFixOs1+gURKwYJpAbcB1UQkhJyp/BZSOeeahUow8AIhJldgO4zODTx81AZiQdP
A/C7SkltXrR9mY15NP3JtYi3tXcQLvduDIC5nkqpZE3+pWbFoYTF6qZRQZ8CZk6RR4crNWDD6DS4
TdNd/w2hw2NU7d5IWIMO9emAonVvqCxlHLzEjf7v9QeB7BJ89YUuavzYiVsxugdRz3qf+OjcDBaz
Qr2lkmsHmm90YokfzrOCKuTsiThvp7RsK0j4M2dQ5pF9Cu5vxQ7EhHrFQQRacJ/MWzi9DHwCVZdV
hFhy6W5zxz6c5kayfMuNqFuJ+BarU2elHKz6lez+rbxhqLWFtCspOHtcvYGr/TkExVCVsj4hvNhy
UugOshK06XbaMKZt8NdIwB4cDm9nJOwIR9zFMhOzmIDsu0W20K8TeG4ylACO36pd2TQhAQvUaZoI
2d5PE1cB24s4LtRlVoJtljKrU3RHz2HuZZlVF0G4inPU6IFNMxHapTDnKfTBFD0hC9lI/ZnSJEic
oJ0QKIp9n/UMYqpNIXc2TmSlLHsw7kzEI/+G6ONxIEWA6JnFznuewHc6h2CdhC0h7Yp9bUgg3g1J
crU0T2L4V/CpZ5VAz+p47nng5Zdq7CvGeg9P2bDsq/ZkYCu+KUSP8mHJIhLJzbANWw+IuZ1HCWXS
zglKo57Szbbm2glczsTTyLYwRLnPzhGR8pfqd4AVeRe2BNa0B2bR5RNPEDROM7I9DfjW8qxX166J
F8dKG8SZ0LKYs8S+o1fZAT5/a+acbDCuxXEpjQAY+DWmcOPGf+/MMSCmbF8oDvyvRnvRYapFJmk4
GPTepvuldR6gqNdGlNMiFZGvsMUP2Bab2W6bmgOjI9nK65WagYmJiLSP6iIq6AZUVv8cGPlg38Jb
qZhDXqQZ7BLRKIVLmQrbus9/YavrNXQNoflp2h/UipBA0/ACU9Wsh7Wv2waRho9VkL3j5tKYY454
70vudHw9BuoYLUoJ6P6ePJXaiTAVZJhjgaTUbhnEejwLkd6dNJqvj9Dj1dLRu4SD6x6gzxKhY3IT
9YHqbRmzS91ftBnxmLTjTiqdJz/BHxt1Fb/Kjnc4Cd8pUFx0vpAc1kD8N+QEQtvHhnbpNhs4Gc4d
5WlcR883iuQHbPmcYy0VHkiTjmpIOYzOZX8HteWFNtMcFw7CTWz8STmifjCIUSGSdovYcuwIFT3m
H0uRcK6Yq3yN22QgN5SAt4iOqoFl5pusT9RfQVjOu0GXG/S/zpvuy4yTTJcOp2daEhI1fW6xlaNV
scy/CG8pzIgKejhYkM/exk6PfE6ypbu1QWE46hKLSxbv/oDi65VxRo5z8o2pMmGqEIntQMKsvksf
gv9KaBb2Z5z/YzlujgSdIvzj4m1130kvtmzRuGz3fQesPTG+xpLm9wJA7JH5XoAGrSAxn3IIs62R
bmuvfsO7dUvO18fZBc6bVql9Pq1FTczqc0vMDcuaY6e9fwJJfOSsl16hcqB7c+eAZANu2+pWYxBm
YKcxgzyZ0YTlJH7Is9ruvCuQfkJlkq22oVjozypWviaj2Rgjj0FPOwktfXyaFj5WIeOMuM+FcmMe
wY3SHSW6VjeG2SIH8xzH8HcG48MZYOKs4kZbr85i9k+sQaskL56J6HDBrI/EhI5ScmO16OwcWF+b
Gr27zYqaf8zBioX/QClIdaZmaq3TntLrXMP80F3aMLBtI/0G3scdyjbfGvecKZvvuikCe21cWQog
7GmfEGaCToW8grze7rvYS9HVS7n2AehVVSYmnr6dLmxAWWMV91b+w2BMgw233gkysXdVvnxjiWT+
M6/6jdDaSzoUqcgsijKNiwA9fGjPEheCwoUxj2prKVpjLuPNmFmXg9rrQHOf/zOSKNVitACMoNfM
ICyQzAqrgeyod1khu4meW9XqFnU+FLzsNCBNEnlQ0CjlqhbXy10siNyB5FD8Ng1sbf/7ae674LUz
XQbCCx0kUwOgH3mFkSnFA8G9qLHRMUy0bETKNDLNRbsKgTvXFNpzirHXb1MjPs7PoWSgrj/4tz28
wT80DYX7x8UpbTFwJmyUiveQqBuVvjfRGW7D4VV2h7PRx1aLPdNr3Oz3w8a1GXrTH2V56kB+dvNw
btf2IR3sMygnvh9M/9MeGm38miOdAn0dxRCenfVQ/Gg128bLkmXXbwT9XkpTdfvosKtK3Ws/lh0Z
GG1GSQzoYrrZmG9r45fwdi7CFaZI+OoQL8pPaOEQHc3Hb2TMuwdJr6Xn5+TkOd32B3mz4fbRmEho
nijPnMdNbOSQM9qQFwa/Pso1E/AGnlJWsi65Cm+JU0AivhvdJdV4Ki+pyGSp0rgAzt9XZ8G99rjP
wdcyqB+b491tajXhhgUumJR8vKtUn6hYJWhJ+tYQWL9LdQPbhtetW+HJmPmfYw7ezRH+9c7Jjp6d
CHKrcbWH1JYv8iaWuswEr1PhSXVBffDbSGMH7kFskBzp+amxB+imEqxL73fal6f6HBHAJPpPLHpQ
ztSJ3HgTPtUZDWA/pT/epfq66jQfesETAtrsZiKiX+aZqO5XvtwlzEEz+56L3PydHRPhkE6fmtZR
SA05hSGHac2X0G27qzV/ywxgRK8N02YIq9kweLI0Jz1wy9YwyiUIYExGTtpAt0C2x9oEGnQrlzY8
O0qLhxDDzXJ/cDmhbqWq3TTJWl8TmeD6lAnUqB9UEUyFojcMjTm4G6yaVnebxtXnbcaFE5bIQDtl
oYz+PBAHMxFMFsLksY+Za22KOKP0Mh9wkfdrVFY9NdBu/jtAGcmOF6BznCh7A+KgBNBqZEIyVowa
7kvE7UpAYoBgOC0bhCtQhfKsLHA5w6G6tSckg//0QgZ6OLLIXTFJzDomURZNnb9Fu5hO+vrJIIv8
1Pm0mr8AUFMvmXpDd3WDLPtbRu8dAsIkZVlHE5t2xANvVM3+7+ACjfWcraZsq6CuXV1nv9DuuuIX
Z1Ex9vuutlJQ8C55WIxWwZFCuD+UBo1RtFyHlmUr2TlyFn0aHj5DsltSgjV8V5uqcFOcG6F9dA5T
ws0VQXISR41MjE/GiRsyw3xk+SJi/JMa1ePSazo2WSfzYgNfpLgSLz8v3yBLuVSrX0WR0xDnHn6q
YotP2sJoUk/tDXeku9s/rYYznZbTM3LASs5WmwtDUNgEbQa0QFnptc81foHZDiZfIPSMlYSCTKvF
CcTMZhHTP9NzuLa0eqbfiIfxD8MKCP8YBCN8M2ncf9Xna/z/jflbn4A/qReVav+0D6XtucU6a3IF
rJbPjEGVMXPLMyy+ngUd1YZk+5vaPOXlH+Zuv8wKAesqLWgvEYhbNuVtSIam/k4tcg53eQCnvAcJ
GCGIMM/MfGdmphRi3XyqNeVtd8p+PZN6ZunQlEyCHCpodWHAz2GolnUY9UPPyCxcKyHwqDMen2fg
ewizTfrHymtrxRxYeOzBEjvG6oN9xdmLBm9BSxn4zlrQ6La7+G+TgOrjpjwBJTukoCAW2S/4yISt
oqiIShKR/JzwyshejNPtLQ0083HQkeylfa5dIGJh6ZfehfLlpK5zuQIXT5EdKAJtYcOTl+R8/y/D
vb34j/mqQPRqa3cVQceJs5rNVlviKUMjlVx9gouX+cmEZ1GTyWsKcA9oNNohhgKUaWdGhTLsGHdV
J7llzw+3q7mmNW8Sh+s9CMGcrplnVKSAOXc8hBN220l5j7z2lxRroj4LS7i4VwYhZf4eKalgsmCM
OsRSvIgZLzQOYU2H/pOHicKGmBOA7KtuT/sfBMJs0asTM6JxYSSxCcTEgfJgZoI8cjc5TWGpt7ea
7lVk3ZUpm0J7ZWd7kAkYr4jz8TLdQIwly2gyd9Oa8ugpWR+arCIBLK9qXEP3u+43cKyeO7BkMKcQ
HRIVI+pIjkMjMMCAzcWiNyhBYDIZDkDMFZ+MU+eL6AG9JH6fu51PahPeFQo0dY4G78+NfgzvI0Hg
k9+/S2llKvtJPYyOm4svbBnCObkb6KQCypnfhUrhtoqeXRm52PEJXkjyB/yvFr/BWuDe02rIiVTW
V14NMaPedF1Im7Upwx3HlfuriPANnNgynHC6yo1mZ0MZZm6sC+vmSSBY6jmN3yhvl6l7cF90Q4tZ
qD0aYEVvRP9zRtRt2trCNIQ89yF/tGilwzpliKhhEIhpYDfRHhaLfeM3E58uPiGjtlByH6IK8hsr
5LXpZTXK9bZ/tnkP4mrP+KXK3hEcRtKq//nx1vpAbIZq6DwZp6zRXIk5RKxe1KldrTeX/f7n00K6
+9sr1zlU2hVfkxIVbCKIoAO4otasZnfC1UVb03fTo6h+/sA6CHI5wl8cQ8GbNK9AdP2rOl54rUYu
5PzR6RreOw6wvjBe/G6p9ak5QCkucMk61wM08XxFenEazhjNHw15Rx6ZUWRwTL0azhte7abXL7VI
thaP/ImeNurWSolGZg13pEjcErQUhHOCqGFoMjLIYwmzs54LPPYYDMMa7VeNXJKKk1ieNe7RxDDl
740VVfymSGqn4O/aZNLhhvC2p03FnHCBnfY57Qu67DJqrtUZ+30/twl7AglIxDNmdWM6Ov2PKrjT
8U9OfyT78ngPin/3oTmF0nZZ4UagoNChb6pscYt5ZUIm9SyAE3LaYEJ7Aw+ba15KELPUzgdLuQCL
dCJGbjOj/XA0w1WRJWIY3mN0+VDuPNzzFbhaWkJ8wb7glzfhI9HjkG4tNf3OLAAbf8y57mFQlPdO
7eQxBVPTp60Mp0pAppGSlIG+EuTLztjFCSiu7eW5mZtjjpasyW5gTsNfarNOcCBalvyzowt4T9oq
ONYhpcPFwf/rGC5w/WlTl5bCRNS5C9E9pJJav9l/obMS+XJP7dlP2j/eoHSC07CBiMUN9mPyc1uu
sCVB5x1n4giEfHU1MhnPZh58xMFPbYXMAVfBOJ5FdHqMBsz0MJr7+1HwByU8NFMkQ4fAEoYpwlHY
1ReicXYWMe17bdX4gcuMSeIriYucQSg8D4s2qsmLgoeodxnYGV5g5K0JgDJu4RGFACjcCCcWpwLq
edtCcmuycAbOtxYrnBfwU8ePsKxzN/QfhoCrqSX06B7YRvhgUESKmIc1j+klxDGORYnT87z1cpNn
yPiDcvQtvSHMbW2f/XghYwj0mYLBQGMco6Mpb/IBvVxCD00xvnOuyFNosMcGlr68mqBVRsKJcyow
SFPQUw4pcDsrPAj2Jki5vb/CGjgHRwVn/6Yo8f536yoMbQ/zHgQ9Sz8B1KN5LYHclKT/Bzg76eTL
3ADlZ9CquyzSmuBCiXPraU/5AY1pIINeVcDXXiO88y7LpKpKA9Kn9OvTM6oKJ6p3+Lt01UFVFvC8
ouv5CVINojp1nAJ3x96zHwMXjgbfhKfqxBK+G4C/nAS80qRPZx+8+wqk/BxM5h+R/3591Zj3zNI1
yqVz+35EO+FNqRwp6G6MTviPl13OVcXwFOWkxRzzYjDy+J9sUltd3HPjdBcMrTboCtv4fqBpJh+J
1GjSbPEEveMVu+Eec53ANp2P67tuDdCFx8b5w9mObSh4E7Xh5nByYLPQAuJkwPRpcGiWQpsY4VMH
QaxaDUq/RrxRmIpb5sUvmlTObK9uRoRvZkIyLyZTflnOQNkpOgECsG3V59PgfOpQK5yHaDNmgQVI
AzPUCB+iJqET1TxTOtFavHJ3xoLqpTVZr+381QPr3f0e44xSe9BwVl/JH/ejjjY7mgjiPs0R8v/D
yBtg95Y7SfcsoUtyOLoZkWklmsklyKQvRrozbnltCV06Qs4bgBQLsFXyEtR9tsvPVdpK4JE1wFc+
gzXjncxQNTn72+jE3tsKm83JNWpoABGFDBmz0rrjNV+31qRgBRjv5lWNXvp0saXARpVlRAiP/6a1
wICSMJY7bA4XTnUzSspzg0YGINJiqBXDmuWzygyC9bmlAL9FZj0qxMVh3x0jpBYvMco1fHg7QH5W
0dHLWn+dEPOIWj7O1dFal8ihxOovG1tHeOmcIuV9Mbwr7L/FuazraOZAGhvKCOJKxWsv5u8AgNkC
cqHxsgz5z80AMaIcyXEgH0I7wiEbOW4IBqARkbIXfbp1OweF8jwKVNBv0p6t7zAXLH2FzGOKUHxA
btD5cHIH5UXOeXq5ZWbrN9Q6DhR1PIk0CYUDQ/fvBkQ8xmcDIaXe5xAEzn8BWQ9TLYo/rBcgCdLs
JkFd1Gy6926b+UIZe3GXHypzgy+QE1vKsQQVG5KzD3HvdyPKFZl4gp/HWpgLtSV4901C5NoS2zsT
1qbe/ZQ/BSO+2z4RexSRnJ6e3Ss0ylRaNNI0IRthJse+43R+9TsdMRpNn1MXdJnzvkU0V3LKAg54
dZK8LtHS80Vq1USl6JqlRZNdng6SB5uwFtmJ9FimUWIkLb4ZXg84airKVE5RIIrUZutlLZt+wyJZ
R/sB0ZmnJlzl1AEHeBOFowNkL4j+Qxza9cQ3dKDvz6zpIxtU0NP5HpliIH7vBaOiVTOEp7ZmTaLe
p9Co8Jc2eJkUU3uLO2gG52Uve3W8dT3qxEw5NoelS7vLFN08gM8GG/zrhGULSkqul7ADe2M9OZW5
QFl1zvD7O5r9qX0Yr0OdNSMUBbYjXGZKXKLUdxxqV/UKaqirwaa79mDcNwbIgfyFOL5t+vAX8ujb
HTB3gkDdRmRGGYzFfKepCNhTXOfBoWx1QhTsvxh/Ch2dt/ij9cxqMB5HJBaoWVTaBAuV93KewQST
tMp7RuZMldVJOx7PSxU6YmKJZTQm+GX2eowbd4LQ5OuhbKKObGkpq6NhXGfpiKTbf9DzwiDpV14x
1SbNb0LURiTbuVsU7od8+P91q2tx29g25WXPGypfxS8/h4fJYzkLeX4XYJ2v3MjyBIZ7MmL92bcz
+5/5x+yk6cyrlnm9FAA66vJkOBG99CcuXykp5f3e9syZDWDBAWO59lXMeDDmgmzVrLxl8Bqoe+aS
UHKPSAqA9zEk9lFwRkWS2vcloNyeA/hIYnpovBlB9fm3TgFoEECGnmjApf9dmlS8fObThPG66XvV
AyCCuYCHg6StZKd1TFWXhvZ00/xO2jGfLqtVzXYUc/7ACBhHDQeSJtDemmU3qfslQz6/A55SfayF
NIMK6oYTACZfpvEaPuXVHvIQK1XK8Rt31H2jgKq6hWHnzctWgQQHbftczC9M4QUlNX6ebyMcI8eW
dwQ/6ga4R4Wm5ICl8lO1nwZheX6KEBfV1/DlrCaTHC7+MQwwryuO6RdxDB+74wKS5bQcUYZQh/0g
S7mAffxjnoqYCdlv6bLchul7pdT3AL0HfAJkJwYJzyertRIDrR5NfADcIzGMtJI47gG0GmDGo/EN
23qN5BWCN/nh0acU126vbZ1wGOJdb45qEY7Wq/DASjPCZywPaWJbGmTOOivg8I4eSugaaAWCiZQ1
yBDqWHEZMfGDyn8k3yhXyuaR3YlTVuAu3THZ1IL/wx3Sgsd5EgEe8KCQxH3EokFefI9w1YFMySFt
tYufR3TXe0MgridhHMFtYALVfJVjokui+qejSlJ0q4y63vJORLO9BA7GHbe8fJmhlL88cU8cAYjU
YGTlI5EH1JOJZFFvj+dofPZJpqu9ZSr1pyvNs3Sve/fZmB+PxLk+23t9QZh/7QqQe9vJWbz7rgNx
4B19ZQM5pKSoTjdP70Y8/6MW7klFDPyb0JQ/v4Ww7q7gzW8xQ1PHSyvs4pY4V7APR0MvyP1MwnhH
TZEev5PdtDManlePZonycBUt1R0nirlGyaqEBnleTrt/fC4TjbkdF80LjtnBnkIkw4i4QCDlRx/U
io9T6thh1wNvxZShhQink0vsqhSfZxxShorU/uSQfG3fXYU3ns3E3LfB4MHBDBTWNcEUHXGZvWRG
b1a5JfKcxQBa3/WLCfMNRx6rGubmw6uiSEWV70zXGaCfFqw44mSJbPwyWWVmRmrMJoic+WQovNsd
lozSump7M617GVmzMpDTYM32Cc9FiL6QMkiWX6pFvZ1j5bygVEDu0Hs0raumteudTza4qT7PCu7c
O78Bgtkchc+jSxRgS/MbwmNtRCFrU8X6kdUV2dAPbmgUOblbh/i9fm1vZzFFy0/xTuIySQbY2wsx
U5EnzO+CO/RmBdsFMBJNnrInacqpEupleFLYPK1xxXf7PX5Qdo7mOWOfarAYaJgv/hiarNrkBlWX
E6KPh8ehAebBjcRcvr76o/QMXPyw8iNkl+yxftBPpVcvjy70BtghpzRLYcdTP0FH1vi3HfykdTgt
y0FwuMOAwib7hLD7E4gAIY3K1q+VBI3s3SFjJgs1NcaLdLKkUNzBySHLclcG3U2a3L0ytHoYBFuR
2mz1Bv9teLrexVu443uSU+T4q/wf3phxjHl/0cji2d7UVTd7ftEpY3XWZJCyk96bWlq/Of9cnizA
J0ZOuwVJEemAWqMIXGPEsOSPpMTbkg2q84sEY2JQULu+RFo9U+KG1FEajfscdZ6ZTCViSJrKfOGh
p1mNK2Ng4Hcb4l0P+fabsqfrn+nzUCgBxNFZIpRJx/+lh1zW3tVnL8xJl2GjGi1jHK5DUO7VMdSd
KcQAoA3AcZmpcR+es0VFhJPbx2Jgz9bmhLNFe4Tk+E7Jwir1zkj9+pcdsyDKrPhKl50swCzSvY7I
DaYqBTGFMlaCSzUEBXJ0dC3ADhZug+eWCBdzdyhpZ/5ciA3H+9jDWb6irlsQHDSeoLqm4cwfTSTm
innD9GicgaUOGhrXGMZ9qnbV6Op8pDp4W83DCKDoUACbxVb23u+Xe4UpWBUP3w/sRByN9+wX+vAA
EgjDy51DOdHmIEqh/NR0vc0MM/ZxMDHVfVd+nnlyJ6y72AHcL0A7IcdivYu+LoWMgDJtFafk7VdO
1tpCcBHDMBYiwvmBQMGdhR1QGxf7QpyeJSsQ+IJy8otCJviYa0KQoW+FpJQZqDMntfi45+aC1+ln
yiaZThm1xMfDBv4V9xhvj0SasDuRBY6rsJ7bJ02D5QvARoz14sAZZX5zOytAoEssVg/tNAuhB16s
NNyUNP7wNaZq0QGGkJzJcR8tZdJR3VyXGu/nHRQecOSpUjZ45d4Cn+7cc/zVZkDSBT01AH8/448J
z5D1KlLAObLwG1QQcIEoPOLrYdMFu/lmMUGc/uI4W8vdJiUHTXEMiuOJxvD8mUgavrD/5EzxmaVB
Cxr6zFbkIUnDtmjbTnM3UQdtD5JwG4SfYAv86smIASNbrUOKtPFc+qWI6whfvCxqa/dqPNAXZDl4
KQYWshK3Fx9WCD2hY78QAIxIigoLJ+X9e96DN4FocAZq+1Uuy8fmmfASfPyszihz4kuyYO5m/N4P
KRn5w4Yijd2s5cOkdqr/NEwhsOJXDTdR0tJAhxxcI7QEAubLKABburgJ7XdBAFbIm7ohjV5Yb5G/
/8gw1jC/8Oyd/tMrgwmSojQJxl3VrzBny1gliSGWomErJe3956pVlmTsfRGMvf5t7sJvcPXI+CJP
5fE0G4Qeuh1Cq8DjK9E7vO8CMV8GPsiwD2VdwvNva+Yy+MjmkON9isx83CXzo1bezktzVDpaGvCm
5V4YVAjTwbdK6cOFC+kATq+Ii2Lh7Ddp/bZChonf0QP74/S3aAZI+nJQnvdlRuXJGaI4oI+dRZGL
oKjnHX+Nari1v3uaR6NUQrUB3sp18VA38Xa3ADPcMiqtl17sYPQxzH4G2zww4k4YXPvb0cINifRB
qWwSXGyX0Im5G/e8jPtVKWevV/q/oY6jAq6h9cKosolz6Kc3BwEZjUFbeSua7as67GbXx7JETcaL
jsGOCcDSazPQwJEciCqPnU7FSR2nmUy0eRuf5Gto5Itl1tSbmEBYam+3CDiv+DH/dRIQ2a3UTpgO
aEeJaFgSTNIIjSF1h7bHTzLw5UGVFNjyi/s2f+szlFD2ztrgsaitY+ut7THdD2RVNO9VL7caUqK7
CjVvbm1R9CRWOJiLHDw96Rk3DoPoJg7v+ntNzeIuzGJPkUMF3GcRJMgiDCH6zYmSxacX4VtT8SCC
cRq5ucUJXU3l3hhHRrTEXK36Sp+RVDm+GIuIxwV6mhm4ouNxBTzik/wgG8NLBJgKj61frCXXqTZU
DvR4L5AVU7ch+Be9PW6ejg14Y5GA3Gj8am/hQvT/1HJ9VtUf2vq6ul6qQUTO1hLjypPvev19/9um
DLAJCSg3EUZ6As9+1H8bxJ+/cSCoI0lXZuL8/0kCoJK62aObTvITok4Ad5KKnlXh/XX1H9SCNvS0
K9wHi/tYkKeYCypfXk7WuvGqwGiAJ8FBy4v917cAbwO+UO7Gk/Iw4BBk7ILfXLKHS7T+r9b4/mmc
wvHMSU/Fd/dvF0OWAus6Z235y0R+R9HdJSRuJkiArQ+GqTfVn7pGiYdH/7nsoCM/fi2zPHOyNuuJ
HoYFQ89janw5jiudXk0W7e/fYRI4vilBKU+sEMP7cKKOZ0YqjKza/dloUvVP1vT3RugVRkrjq1Bm
D205CzZsiKCdQIVqegFe7cuHZ5M+7kDSuMk5E0h2QVmiyGPb0KmY+V9/jknAKxzuz40YYtOKaOsm
HgQiqgA/2EEpH+dB/cCZKY4MIBPB5KKsp3SdlltSDSUo2aD9ozoeT6w5gKRFAfZZle/7Ir2rZqO5
0kNU2ETfYPivp43nE1VatE+BvCKEPXKjsTZVyII3okHzH4BIT2Y+0Va8pWczxMt/gsCULMaPXQ/f
/qMaFRA3jwdQJ84kwjmDmoDD/llK2co9Qo//lUj2DHCvvuH4AGUND/PfgcvN1MRYSov2QLnIwIMN
hWK5+tW4gY4mdptlaLDOnpj8NWlLcr0YQsg2AQyv5bO/8diW8GPCfVduzOlJRIadb92zzGsnCzhJ
WagmjW740v0k9VTzEmYS2My32CdYSUrqd4cKqVrvw3b8S65lwDTEfh2R9FUkikBePWuQ44XKG5Ld
XBc/dHFHMGwKjkC9vs4/jLGN3c/WPcRmieFzlc7WiTNW6ps/FOhuAzZgRd3X4qRbYUIvbNXzLV5v
1oT9Q6d3p9Pcm2e+cZ6yt0t5iq0dmm3sDeYADrvxQPmccZY3oweaU6BW+HgFiQdvR57sYt0Etlmx
nyZJTpGiDLincOC5ysEIyYqlnCEBk9gJSq/vsDsbVOWHnFpY5drPOlqkw08fO7vO4mLKe90KkD3R
RFjExIEwD0m1eRXSRSkavTnGhG5jNAKDqVn/cdf0R6j/PeJSCFiu74CYhJqmsr89jP2KZEo1mwy1
gKaphwDj+1iMyHvPf3J5fqnk/zK7jZ32Pud4t60560qVCbK40FNoBuHQN+h+GRgk8aNeE7mMeSUM
BLZIt2gq9KwBsNG2mivquR0VW5lxMCOVhSXWdW3ZwroSxzWtPDqIRePsylIwn08Rc6PPMonH5Ky/
FAgxzfr/memw+dAe/DDak+JgdBx/1gXSlZyPxQzZA0kHKtEXcacRIzuhT882Ef+Q1AShacBS8rSU
rogu1kKTdOfkVa8FA+wK1a3/qh9UBLeznhwvxmUUX6wvklkF/8AGCdfkvmg1FtKx7QVKQft7Wqw9
HYnT3kVq6N34TSJnwhfDYFnU2MY+/ZQRFeTVNlVVQmPg5bQ6Or4TYGt7tqH33R29ohO+UV+OoJaZ
NLn7YGizX85m42Q9lG4Dvq2CGXsNfX+LPXrOl8LqxMi9xn1QsH/QnzHA+lMTeZmU1gIdi0RBkVvc
SbjGY4Zhpa3PqfsL/Y7pQEdLwVJpf0NwpcQV6tDmJNWQGBNG5MvFKiImWFZ1+BIDZZ+jIeRPddto
aCT40c7w3wTXpHVyePEGXcP4Sf3gl4Gtn+eWaDJbQH2yF4IlfmExkWZl3TO3hzJbwz+mBbG98PNn
psEMhQJ9Hlv70D2ddwTkSXGaFRJOi1Y4q7hBmxEgAnQjWXH1Rb5hWKMB9WkzLs5GF4CTfkaKrddJ
GYhos7IuCizRb3WYLB6KkuO/ZVD5Ae+KwZnlqLLtfsgBNxbqoGqeJ1fSlVdtguAuJlrvBGEmjZHy
xYZTgC6Wluz+CE2jFER1NT/fxvQrsAhIz58zb4Gft143IULhnmm6NCW4Y4AjcMsrr3745ZAw5b4p
G5MhdiJe4QMa66X81eGwrHZklfqXeuu0labXjhWMw6OTJ20R7ZNlxqR6guymwAfqNoQLebteKXQ9
gqEgcoogpH7W4xKxgZu8RF8eAQ8ATptoVfrBIkPAR4vBGU2g5N48ZuOFbCdcteT8nKkiCsffy5nJ
8g/YWlLnZ7Y7OdhhOwDiGZYYV7fP7g6qWf1ZE2B1Kcc6Yu9NW3DL48E+YzUWmxdPB/Na6opIZPhE
KCVyp4On8NEA3EMRRoD4GrptUzO83CuoH475K09OKv5juNB3ij4ZmNmDIFCBT/+cKO3FWtNRz7lI
yR00dlA9yau5mTHZlf1xQfXAlPjTd7BlXAsV3FWZfX+OFrK0XMcHxfZOs8PwqyGY570NEVcYfw+m
IAx12QGz6dACLnMUt0sXKLGjifp+BGGOWHVUEHUMhdWMT1oJeZtpK/cBv0hwP7LUgMGot6Hq0x/R
/iieiuUfJXkLX5wy0HLtLZlmvUvNgyAqxO5WQ8p7X7mK7SQbFatbsOmpO30KDwGymveMaBsyKQxb
4BJKyJe5RD9rnYKkOGCWJrSzyeJSmOoPd4W20kaRf0GgKE2JWvh9R/oFxi2wWnBhZR6ZjIK7TB1H
dJb5gcY1YyWBtQGKQ7j20vW5GlZbWA/neHhwoGYiBWD9gc5CanzloQEhWb6RsDfeiSaqDaI9PYsj
N+RNp1wsxHg2x6B1kXLJhK+ByQO+1ymvEaJZipZK+NK7BXF5f+PFUTslld/wD7N8psLwZZck5z4k
BFPRYF4yN6hKfIRIjJtRssQ9ifu28+5Na6v++lv78WFQEeSsWhcJhs9jlX8CvJSErFsVQrW7Qi9X
pm/I9Go6mWLVxlnT80rY/6oD4DFUTAUr/ZOKdWsp+Emk99bkE7wPX6koInb08COrpLUgl+uQJnFt
qhEx9FOIFvDB9d3yG8KtFDQG9mLpeWYxlckTo1kLz7mNbISawv0h7NCWJUCF6/TyW/F6bpW8x+at
9xiv5vCWiyZO38crx0/8vqi4NRB5jLlJtzCVKNLMxM1a9Y/t2gyYO6r1gnLz2GQA5dDA9yrk+r0V
wBHEcKG3pMAJEumY6qBQ3NcnCKFgO9kuE6305F1bzog2MPQWnxAGjs2RxdHUd+k84+1wjf9wbMio
2M6xc16ruOfswm6htJmpd8HlaMis2i5Y+gTr34795tJuRxshou7nzJ5Z2tPwmS+7R+FdMw/tA4Ts
TK5NulhEqcCQUAvsbiJJGmpY4nyzxbJv1p0GL+gv5WlgLxwAWSt5Uiaaths2K6g4zE8uOqZ7i0n4
KK1WUD/rmgXZaQQFrCAfq+6DQqwzZ/CKywhz36O9kN13EHolNLRn7U2J8GAZJwg0izAZs+Jr4ego
4gzxEHnLbpwXl0E1HADII25K6aHzjRg74JoKevLOdUBml7nbnOy9GFA7wptIlJFxPFLu6fpgGCrZ
6IngeXbLuD5muql/UVzmZmA6vtwvoAwHlDLrWA0oGlOrRybs6cnW/43hjJ4fLjYlJ6r+0Fmwh/KQ
nnEMcKNR6CpTcEbVzJR0mH3MHDkfSzdd6I3EhEXeAKEAIMgZ5M8CWf783nqPvK8vzhGNXVyfXSKS
13H36zLqz3M5FdjqCxjPbLIn8oNhEm5I+g78xiaq01M39Y2jv+v4PDbF2DRTvNX5Kv5XdP46/yXQ
y3ebv/3eDiCKZark+x1VMZJH1hz+mgxJigI8vJqfA2R+WrJuEQi7Wf6NQATl2m612xHSjHRjT1I3
EMXmTbJ3tM2zEIUVOfs449bswXFcGtrez32Fu6n2XDSxXN3Zql4RQDWjLy2CKs5+ofjZxn7gtucv
AFr9CN7pwOQ6VCzqI04grCBnNYxco3kC9FKFha4xmDuisCMMg6ODfvU9uZBNt6NpS332ftU2x09o
FbXlI07jX9YCUJaUJhmhRFjOkXgR2HNQjnhzQSEB3B9cZWto4jpNLukAzPL/JUvf5RqN9te7vEN+
AfJjAL0ystBZZr+y/pFUarziSHeZcgH8xZvTPPTDVA2/gTEWKuBfPPHrO6CeX0LwJnbaJN4xHbpA
vGtrERZG6lz2H9LoztQMzyrxdFPwXE78UPDXjDne/zGfK56fLp0VsTsZYIlsAE/gi/eNAx8a8v54
IOm6teW8Xzd1FHP2FKN7dkDXwxHwfs7/v29mM2AzeN813XoKAIItRhiM83eamsfkG3Fn/kULSmsP
71IpDMtFiYxIkkZpJ9z0xUHRzqmFB+GVAF8jVWHJ8Yq5XiTewfMjOv1EUWtmOm8ZzemlTJWD07jl
mYOWL/8RygXGu7Y0uxCB9Cn6ZqqEob+nMl6DTy+caeWmlGxwqLDBUzkPqoOBzdrpNf+c6AphMsyn
r0ya9ce27a676ZGecH3OJZaaYSLW3dqTTtyYzBS6nB/EaFpf9Z1/5Pi4kAbVY9yWTVOoLqxaei9Y
Hak9+UlG/bCXJ89lYzeIQCzCsQq4i/YzasSJVtreyjOP6i9pCsDJBoaQjfVONlcsZ1BtByNo
`protect end_protected
