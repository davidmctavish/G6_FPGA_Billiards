`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eQVuMcIg+Ol9RIIPC7emGIk3RUdyJeetGx+ARXYNgzKBbRt5IOXtKxsUrZhQB6rop058cWVLeI1o
kgGBWavPPA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fXOPBVawDX3XXBdROzIiLsyxbgbCUwzxWs3dI/jSrw7Sxo7UoXNtHgEotYlhMBkMR0bNrlRsBb8l
Q8XXhwmvleZ76bJrWjxSt4kacqnustIjgwRPI+LccOeXPqZ2rhGcknYsXpIv43N+JPxeHYncYoq0
Vjt0GxwtXY1usDXigmY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lgFrvqFl4RgenLUuGM9769CdsWOdRL1UPndQRCo313qF6BXkee02ozm9I3tuuhciHvZXvmUQ797s
Np6XZDQPe80D+wSVX35SfdV0pR/VtlQk+Hb5gSjrZ40NjUie2ep17bJ+ACBOIkhpeM1r99rSyEPt
yS48Ez32EOP0ZfnY25d7kH6pM7mtZPoAtwmFjggr3k6ESEH7k2dAsjaGp54Gangwmp9nIAblJHnx
Puo4ehnw5tfLc2VgFccmSimzbA1T1GbIrkusyzzPM4JGx147Kl+wOIBv/GPhu/G7O3y6N9AQLiap
ePug2I2fjA7XJ1qujNi4Z1Y8j61UrzanGImrNw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W2uLXdAN4rpBtUSs0HG31YJbbuM9bwjKWcxQUbEzVxLLuqNg/mO9KLgEZ4xjlkV8WDRlmtU8WnM+
OxH+srBe2wE8m/qvPhwuQkazIv+sbgugedx42Zy0VDkNdxTKFoUz0E4qJ4b9OglH7qDC2+shEfPY
/wA1Zne676uHF2jY6Zg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ISxaWd5opFW0WQzhv+LeaDT5wFQOuFqy9aa8JblbWt8J3XbnsW7l+xEkQqkjzDXXx+rHtMaajogK
a1JD7Iw/T8ttJ8YyhUc2W5B2PFGgrurzG2XBPk0pxnAzQd76ItQ00J2wi73u5bTBDY5JhqBlrVGO
fErDPRH8KPz9hLGFtM7898XbP0MJCRsWcGyEmrM/Qs66De62ygyISW69RpM+1KJgNeiwo+CbqxIR
Y3WfXZQWdFZF4tEtTyEUEksKJq8w1uBqVuC9ta8Dl8+04508sTi3JAKN6saxRVt141msXJDYMtkX
aaN5JpGx/P78buHB2sbs5vv6FnKV4aEhGAPMjg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19184)
`protect data_block
+GuTWwTGO2e1Li+MCAgpsyeavDnmvIgiBeO+uRWJWAlklQovy2hoFV1DdvunzrvT5FW06ArndPY7
E3/5qMByw0yIpnANSrG9j//rlCsrdwwAN8kYoAPRipP23WcHNkzH8BMomMlz5IEIiln6EXHCOMb8
E4zw4cj4UO9etG5OzbdadZgzMn2rZIDJ1zU7KYNk9yDf9ZCFHszptfY3WJSj3gg3w+c9UVNkv1mP
NCDNnVIWPi+1v1T8dn2n+wgDLegIbJSxztJusGF6VQaJlewTn2BDEMOErRa2EeqpmhJnPyBVy4qn
mU9iE+yvm+f3cNrM58TEHgkzSap7EtugxzJ1mb+GmpK69SnJQlIl2k6sSqoFXBGKtJ4rSgkz+9ZH
h6txh8u6GJnAxHbEU2KZFdWZxMlESFutOyOC8K9s7ekMpybLBCHlrTQo8GXeVTvF4rxQHa8rCh7O
WOl0IQgmoiWVYtU52hk24jzxUZ8wfaoOMnp6uwRfFhk1Em57eyS1gRot2o3+ttwf0X/xs6EnyGRp
J3ZOv19UCebTMTeer0jL+uXHlVDBxVRdTMIWKN4RMj0PAy26vBQ43d5wo2suBqlsK5CNkTAUYB3f
iL9SclM3lpT24IELez/6ilP1YEkxd5bQJ7ca4nDwX5SfgWrG0nmliLyodZ6195MokO0FvB3o8296
2NC8x3148Upc9uRQhrI9QhTYU82NWMjAJ1LUlrzLnksv2cJDNDcSWiGqlbSikbbvlxBDCzSVpQyj
eMbc5fCGujvoi3nB84OuAxdDJ2BzKYG9kZqNCo+xiD68/fdBRr3yOjo5boueL1RoHPueIQezrbVg
PPK2s108c/eYPbr2YOOiQuRualv3KSNQwL0pJ3SLcw3zwNvjzxVJHYAAkad+lrcUuJro98RcLCS4
JVzkaM3V+lCjEviut8bkaZv/lClPc7fAmIQHETQvm672w4H5AtPQ9FhtJrqRbgnQARX7ZypaUhqZ
6xUBs8OX/TzNQdUqJOxq9A9EW24e8nQr2qdQkVUxat7Wsy8XsaAY1xNTctNcXLKqMvWoqrw+mkYr
BARAtbVjL+YBcm41KlbXtz6HGq8pEqr6Gkv9jc0FkPfbIA1sji905sU07RO0C8iJfULyfgCfbS6S
cr7xhXZyh9ndNV6sfRA/0BVD4JCCI+c7pHUq48z2w9cIJCZYwXe5zXMoSXxoUo1tkq4RVgC4yGwn
CbLwP/jvjQ4Qr7StAGf1noOk3oiFMvQJi0Y9YTfa8+7J2vUJjbWf3j1+PbHT8Ykj/PiFuCLrGc3u
MWujufYYk9UXlOX2cPNN0+KcDnCJVpnE1gYQRwb7ogywD0yxfpd7ksk3TDuH3fObK4Vmm64FqLqX
uqMjQpbQAtMQB+FDgkoZuTYtj8X/y4D25ElLqbK4YLsooU8rofj8eyVoI2X+03UC8zZIiDI79xym
hpQYS4pJ/XqKzhfGtoBPFY+HFNi80EdUXb9XffZUt2JUBhtKIdZMxqBDZkhVwXeC57RyL78kBKWc
KJy/p7yE3GaF5vBvDfszQdJizrmJdaE8CYTfEojdGihx70q0FMzGdyuL9SvMrF6ZGhibzKMsry6Z
vFQ6Ve4OfcZAhLvHpQQY2hHOBe3JsKNa3+e7XvgZ/dBWPzScAO+H/qp2iyylS4A81VknKLP4QEmb
3Ns7t+GMQTLKGAxu9AMtrMUrsyRhoGZxb1Z+ROdqmpPiqzKXNUlION/eVkD+AJ5IXWYbcNAyCJma
3uJbg6PzC4eHSTnuvJTdk813gnyty5chi5Vw5QMyzg/5iFSdl9VsKcRp+0fdEJLKjbfc8hHJNmxY
pmgs6oiOKHqgTns4/UYi0TNRTxThIYn3N94PIWBkutVGqUJOHmDbiitTfae5X8Cvu0E+zB+oahlQ
mi/v+kJY4N1AELyQ9nRbWIO6nYE5IuCriKDLXTnYwFF1yB7irjWWlTDPrqNICoQz16maykLM/zl8
RvwdAOG71Eauta1PQ1sRdpIb5UeKFRQXvro86HFc/aRpsVfoX177ex/HLzR8MVEd0suMkk0ttA/g
+DHvoJcQ0wuK8LBCUD7jrTPwsCX0dNvZJK0Co1yNWfN2gfjlIAOqQSziZw9H/tXIYzP16986cMoo
sCc4GgFbSRZFPoBBWWNDWY2N3DaxEbtUYe88MZH0HSqzHFbnupOrkycfOOFlr6SGfYRa+SKgamBW
Ky8k2KcVcUeYK1DyBa68c7NJtIfkk2MMt6ZJDKayuSYtknwpUE0BLBH80Gc5936kEJfOV4u3XE0j
W47q0MJrBsPgMU7w94C25FPshDnrCtZ7krd+awplAV/0tXMMa/3lDRmfqkJsPOO2jpw8d3U5cHBQ
w+T7200J20ILNEZil3fHF0sK1jsRZDeBXcCQnQUKp/JiH0Y3eGfUcVPrJfuhDAZNNJn+uuzQnPa7
tqRkeGyZG+X3m2yoBnZcbW+eaSU5sceA+sBmIG0g1JMxL2ydAXNuPsVmGOe+/CuJtJk9dffM0vl8
09qTUtUgcsY+Dvw0lNt4OrU+gfup3yYwcKWnmLPJRxJEPhTUDT7Xe581w695qf3oRQgJNu4DZ8ol
FkYw9Cx7m2Yv0R7PX53bS2epilZ/XoaeoVQYbDG9YzvJni96kpHQ1hPKgwTHKglAhRrcamumM6be
iMh6E3vk3BxsXoKjUqOcI9FIu4MFZTTyJYkwBZ+MURQ7Mee71RZXVZ3xHxzzZThD+Ns7PuCL6x1M
1VdfhCRGvEYe+4Z67Dte3avJ/CncJUCssNaruhXC2Auk4csZ7WRtTYtVmKsHmhk+bfJ+S4eLAlX1
NTQdduDzWPYSjN3hRt438Va4lz4Wcbe2BBhSr1lCveib8rtZjRIoMwK/KZbDgW9JnQIqKMhaYPIP
yNCt9gB+BZDBI/w9X0LlEfLV2jz/Mf7dEoEjjuzux1wcGsm5yjJD6zLYtMkewesJQfn3bwcwCj+C
hQINaiFZiP/d7ZC+NtnrXrpRsYGnitmCOVq6TkLnXtvGxwBgnZmeuqAe6Ho75kBAT2JpCqSw4jsy
tiOZtkj+2WaiD7U+B2/nKoLvdykIww4q4Fi83uHeqx1fRsaqCsVKdlcUhqTBFJw14c4HchEU3Jmf
JKSzjIaGi7c2pkqs1Cu3T+1bd1h1sYhWMBzKeeeuRLqHNM3f67ljXkCoO38c4G+FxbUxepUaG7CF
XUTFoKTRe9hIUjJNOGtNobjfoMjJZuklp+OuGqjUpvDh+V8zER9CRaJd7HY9OjK9ZWhU4RlKu8h3
HJb7bctD8iklZko2kQgw71YbTv0lDMt+6OtndKIXbmOv7sHyn/can9zr4m1Ie3gnIOCTGDrHPZUw
Dl6wKQl3ktxmakt/Q3ZdQGotr1rPlafJDS+r1RrIW26fcE4Kl/TRkslurTzbxwlC1nAshEIZ/xEQ
sIdSORMGzs2HY9ZtmQZId7yrKUhVsYUCoqXGFAWRYCKaXzqP4h7lesO4uNJa/kT/6UoSpcAA4IWE
fIA8HNtQ55GTeCbv0sNaefdchkPAbgWjBya7kCbncnQzLwPDymRq9sRMP39hJbsF/eHGhU2d5lQi
3CJ/TLKr8lcJ/meWosJ5vptVb1Zn4+Nr4ys+vp2kB/3H/N/gC0iAxkpIRH+K8+djkGqEQHDgqARj
a6MRfmj79YkQ644zZkNm+T3qVBUVXaRerMS0KiuicEhGePbSqCIXWNqvUSivadb6Skteb13q1ldF
7uGWcMH/tWIzvAoVeQVl0/raHHLSEILvWfJr7UjBOjKB0rnARDSFHmu2j8P3Ssq6FnncNFysQ1bt
raakqBT/3KjOyY5b7LPA2maJYHeUKlMmahNk1K7eOQZVmWfIfcCf44LHtLd5nRKXL/LjcQb/nIFV
z7NeLDmt5fRaCP7qKSprkRIXMaJtafYMLXwFPcVDDmQdBpQK7axymUSUQZfefN0+hdMvaVns7FYx
3UHyB/skjJHfrcEfQqw7hJUz8J8rmI5FjphNrpyOwO8azJCNRKuwIuYfVm5dg3sNzTb2AwZeR+Fk
E7NnbmRzmF65kfVRAzrF2WuATTEMtO9etL/2OvW6VK+rXzEf3ToRQ9pu/KHUUbMRwuaVTy/5/3ak
E68ry/Qv9PwGCRVHIYRmI3LKBk1H1wjsU2TkhPF0Y1s/FISHsEpBMTIzBX+U6+uzrCVRLJKFFOew
s1M/BLf93aiei2fhZ5xd36FcW89ZHnVYf08R5P6G8G986AKP/icE8XkurPOx2+SimlkZ9Bup3INi
6PUSfT513ZsnzyM94CYlEX4XYnzRcrOA1ptULJCx9cGcBbudODd1LmK+r1sd10HN/HXcgsviLYM5
9ApoxVyQ/VGo8/3tex+aseS/8rUXAlXY0Uyykv7uMr/hPY/tfZ8MdwlsoPhyqAPFBVPjP/F16rxu
E85HI1vDW2QT0TavCDofIhCkUxUbyWSb8lhTixV07HvvR+woyyRh/sROpAVNEXp/Qh7G9y2mBGSW
4e1rfDfS54FMvrqxovLW/r++IWaCkqGw6yaq+3c0ED3qi9cwCH9REQnvsIe3Gcss+jLQGLbCS14b
21fZZYC/15aNeMxRpzRJBuDgU9n/sVmXcwpcyHu0ait/v+T2zvU4omeCGgGviBe/BjLTKKa+1e7m
A7DPvl2DU5BYMA7RVMzkTcsaJfyjZ7j4dKxYKKPDn54qldjxFSKzsW3A2paxEiAdoawGrx8YTgv8
dpm/0PEmIeLkP7pFo+MDpcbG9I3txPFGQ5Q/pXHZQ3ikDCR9CJfGg5JI5LK//XEwlAmh0MhyvzRW
Evcah7Ksw8+T9/bb2DADjtupAXZyGYUqsSxosCNjLgYKHepZY4IVNrYublpV9mpcai+pgGVSEDTx
30ZSXyQcbnHHSTdWRgaSYChVca6yaEoV1+ogeh9ypORCAjohpSwaHnFImm38/yYbxeQ2wcWszrTJ
t4zvXr+Ol6GWKpEbxaNaLcoiM3K4o+P3AyJNE0kdjgjptlAYVEW+MnBkU/TMA/szuyF/LVhofzmU
NUEehdW8HFkzcoUTTsBuBWlxFdV4v7nORwdiIOO6AeQAl5DYJed7jaFM/f01uxVvqyfgc+fwPNpx
bwEHYfuXIg6rUJTWimbZl6cfVg0VlEtCvP2VVrvHUVi2Imume9PIFtTpHY2CIHWfDFGgCLog7FUT
xXQfySk0tifYIWshi/QteaiWJPhgWs7wzA+ztoEG3JYZtL4njt+WBhRq4x8E177mixhnauhSsUh0
0lgtmB0Q8pK8XO6Ew1LQucooav8G4HwuTBISAjiYxcJzojlOB/WmV3sF8FGeFHere7JC5GQGV0d5
nYdLjl1QsEM2dRCfy8/MJ3c2WORta8HgUDrjDhjyqUSyq4lkUAJiTrIQk7vMYU0iQO95pACA5RCE
+sY5Qm7xRDPJiIkejJBGCAHwxZ1P4PGDY210AKXTBDZ0coR9ZHOPJ+nuegLjCoP/xTotkLJCeoC2
dZXJr1Nb/HEKqRnDN8Q5xxebDxlbW/te/JJ7IQEYpLJvkOZzWdsv3G+bk9Psm/IfEIkox9xZX/Ni
f4MMnN/im9DNIuSvGKY6FaN8JZu2+sYS9snTBdb3Q/bitvO1+u1cb0BPIxRqXxujZFzDrKft1wdY
6H/GDd0Q6AEos4cA/6stb5EBwRBCLZEYoO41HsMb6CYZ0QuiD04vLO3lct8vP4Wu0/lYUyNv/S9C
gNo3sRc65t3BAIGDTE96kXk/qO3dgTtuRTm75haHEIhAoUqhNWLpwFJYOHf11XCkDFQo3ybW/d/c
n/hjbEwP0OhF5rpUEloJyuHCIq2e7hYkhRwS+RFu/GYCxxI8hK5Lb54602Qg3ykl6vy57CnZJg0T
i4snqd8N1asIa6N+5bP+Y1yvvGrHt76fT3v3VMkedmOV2FuSdT001PqZtFNNUWmiNm15XUCneR2D
D8ifTTmh+43GZoMTbgo2Jh64sbpVHJO3Hmbr4pXLj4/ntfM0ytB5kKpFCdtHPDFDWauI990jbSdJ
xpvzI63akU4OMpSLuYJlchLRL0LON+VQq7Kh4S3s/h8r9+XZcYcmatN5MwOp9Sf85DpxbTXllh8H
K80RNXQQirv0VwO/FbAHeu7/xNlCJJNzIQx+I140k0nzgputmJ2+zNC/Hg5Hwc9WwAr66L7nqNH7
6YCvLcUl/B2PXpzMkpXqHzcNOzb6+xdn5TRAhIh4MJAdRYjPbwoQh/0T9xHyKN6pqa/cVRxhStZF
m635e69x4F3KboCwjQsm/0tCRzsXTM4dh+bB0pCL+VF45XoiMpDo13IjnsB27rZG4WuOsG04LK2c
5nBDysvhBemkrIOtjXsTsxaH0iPDMFCiri3hJ4oQVzi/w2oU1obGgqasghBEp/zRQvwEmS8o7ZHh
EVcsqjPXIPJiwnngJ/gkb6JOPHYin/fTNkVlAzHZc44oDsgbSekCMIq6xgWGSRLCdR9aYtXONXIP
pZ56AWsaDerqrgicBRXNVzhRCiUx7bAc4Lr50efOLr59v3ExdLwbLyi5aW63EWQhxkhcF78r7hg8
BVJcW1Ni5vb04E/6qZ/M7iJV3k1njmhG1tnF1UNZr/XanFu+WW6D7pKYgallfGpVNMhSHaQtoao9
NkajMS/xbnhPbstjLvAm3AqozkB+zeIX/ZY3SSQxwH4n6CSrvJ6wetRbxrZ7bG6svj0GMuvWNwWC
fK8Z4R0MHOcweuKgQXE6cO4zCb2ZET48waLMVvtM5Lo2HlrhFraQVYGJVUrImzjZEbHgWpcoJ1/Z
EJkvax6WVPZJMxhSmIO6xeeLhbFRGv31y4fu9pcyvPgSmf5bN60vLJpr+vLU6nT3z6e3EURLC/H0
FYZvb/qI6NaY0TV4/7mNANpAyNm4wVSI2OKNXMHMqSEPA6IPwHwHKdNn07y/PdXtVPT6xrYx2/Q2
oGSMHPX/zh9MAYtBv5rmkyHwTSuro7IKOKk3mpPXvQoyGh1Jzynk0SBKmUDQ/PuL6g2XcAX7Is98
G3HxnNrUHmOvz5KsJX39eq5PU77MmVQG93JM2x5JAKJvg5C1OeV//gkZHfvqzphQLWPsHJBJcvVv
rCPoMFQbs1LYNSo++6rPE7oXcAMvGZltdkNdS9ouwV6eziT2+CQ0HE2h9Z4hpHbs7ZEIwqlEmIko
DNfJUlaT5raVcXupcgbuSbdK+xfdItaXpn+J9zMPh+KXZzAuWL/Wyf10BMAtVtW2gf8NWpw7xs7+
g7GT4mNQdAfsWY5gKTC+i474CJQJdlANWfM4sxNheqqHGPCemlJnyPn7nGZVfEgPUuUynufbFeAV
PNypyFucp8NG8yeLgDsz+mgSN0AHXqoP9OrxicbyqtaurM49B5BRyqI3SwrBa3ks0qgiwyulDoX0
NF9iXTxje9KLgC4VgRw+Q7uaElxpYj7o3iWHype2/Ths6XM4EwZW5C0cVLNUezL9dMSXs5i/Up/X
Hi5sLnhFdt4Xk3OWCbQ55EaUugItyK2rm4jSqa/IknRBTrsNZgZu0jRlOe5NhPbCfdfoDc2VmpWJ
f76cspuiki6VGwvg6uBouFD43vYwVOTPLGaItMOU5n7PasrYppgdBF+E0KKzJrpp49toiyVmmbOq
9XHy63YHJubqq14zPdeIZbGg+pAamHtHbPFdAXBAShSieKZ3csmVkQimdQT+CHiuZMzRzbEq4+aT
D4KoQzMV0zIh53oaBf8m4Jd6BOOFt2X9GsXrbHa7wnXv89FCn/REZv80ZK41f9Dsh4fCfeJoP4Fx
5MXKCGO5MuoMPPuZOBQT515MN7VHAXN+mM43Ojd1YbJuaUx8e9XobfbBJR1ec6o5L3EKYcBmfh3n
Jz38ijhSA1ySt1APmZytnrw1q4NTFGVkqJ4Xe7YwRjH+Wizj5IzZVJb5/eSFRc1lWIcw0epPdrdV
B2amQBAPv8NhIfz6g2ofXX/TmumCw6Ave9maETG6tUoSSwuucFo+Cu2s55xYE4fuTNgf1bO0KFTN
be+SYvOJ7Mfp+l7UFTl5ZBzZMI9OsfASQBPcxw5hvXFhoJMTgot/lXNMQWqhNVkr3zNdkNakGd3c
6c14Kvf8gJ8l9piG+oWUleg6GesocyYXTN+vbV21ZinClpOtygNcqLLdDId6AsHmnAhtda1nEhQM
g1Ow01SjYQPtJVpPnqLrGyc89XGmyiIWnT8JAwu6Bo4Myd6F2VLHfApR6/76Tb39Kqu6swAPHLRE
wI60L8/DGRqhBH/Q/hPNJU1M0StlFZ50HX9ankUIWIz6OQ/BwtRdphX5G3kUElnVQo9Zd7khplz0
0/aBSBSuR4GfG76CccpNM2KKqU+UsO1ede36a6UAA+ftrRunE2XVr5dXSEmDi1ahVS7VmZDqIeTx
u5cM4quaZ4A+7WVp/mFTcmQ3QjPwhcq2M9dJan4V0seEcfXHo7swF3Xfbs11yqhErdS6Rw+6CWj+
x7vpldihS5x67sAsWLV2wKYgYQCFrhb+ATDyC4YSwUn3vU/Orz+y6N5N9KMu9+WSE69avFa2A1ya
w9H5gC/wY/2Bs2niWu3RwAqIC7VJjh16siU6BL85sp4EaP1EwNWOODASCe7hM/QZjNv7URdtrcmW
DlscnvPTJSAXVmTItaHJaIgSUUt3rBiJq1cyKCMnn/LMra9U2o2+xrQeoP2zQDKxWg0Ft+9YAPqA
iD7K0DKHfWd6J4jtgGWbnnZU2ju0hfYk7nVDA9n1q1TMCg3L16D0sn2avEjRBzCrWmbkdDSO0vWS
4Nn3pnjyns2N/u3micBLIdDFUnfme5fUeRw667AcSyuGuzO3CmJ6xREcbNxXtCr3KlyXlt2oBLgp
XQT15gsv4aNKLpRUBVUJDz3CM5kcS6HLSM08Ost/A1OfjZvfC1IDj347dZ3ZnFNZVtbX1GZpHjEt
tU2+hRL6kYqwGlX47O5eVfWkIP0KY+qBXzNCjhZ6Rv3XQjlH+t7icqEjB+jkFiEr2agRmoXShzdq
9LA0EILWy20+wdhYvv+Okc9rNSQ4PAtJZslb0QIVkQ//aYSsZE4RjPVmDk1/BrponLDLxidyR4XJ
e2I6h3QPIMBGidsPsfDReO+r4qrNj6Z2v7WLt8nJkACjgQeUwGPp0xJviUmL0Ed8Mi4mOj6eKp3X
sVAAZ/TD77jtPPFCCEyqTs12PeznNhNwXwBFulZ95FCUqOlrABptyphxSt4eykVP1k25Yzjcd4QE
YguvY8UnJrj/uqRVKTmbN8mwGiSf5GasXAFYudsx4qPYcB1kIQ3a0TJd68/eGaaVn808IrN+n31C
vNCLT8ABu7USjdvKi3SSl6QkzKjn3RNCG3cMcMLGJz/4ISxGvNVIGVD4UAQ5Vv57A35uSnD0UZjp
+LcgtaDDLWbfjCrWl9KE+WMdjNTw7f+RY667Cx8W24MpH0m9LReHM69xQHEcFedpIkUUEdz5/dmZ
221+++qneHk1sZ2EI40P+qK12OvChifUKfGF4TJMeDs7v0LRjfjcZI52IK9ElkdwzxeDvq8fN+/f
5uhxMMNOP6bWUNUwg8u5C93engSIHlCGGPHDpOSlkpijEO5JuZryE8UJeZ6PXHjH8YRANk07vsTX
eZTH49pCPEpC2kUxj9dKQYajUU9+U+MSTN4Qwum3YhU/OEcYrBvVOv09+WtBzv4hVPF4stTfVZ5t
D5V67kEybx8/1vYC1bIZftHKCO1yR2X1kaoKJ8m57RLW/TIXaqPOIhBfu465YEZxNswTAy66Ujwp
ADN0fCcQQCMWX6/PcrZptrZ9LYrR2/xgsbi4IRICmPLt3E59yXHiBQUdLVvr2omsGJ6BE9di1cb6
aJQJXKz7w7BhR3mWA5bYWRS87l1HN59rvP08KC+Ix7d2uZrIH/9ugtzzvWS1B+sbnPThex9fif+l
jfGQx5lci+MKTEkmt/2t8T5V2zaKENYoDPLTLpnQkUMdaOiPFGl8dUe1iLaEQEFetgYT4ypJ4FoN
lWVs+vo0x/1d12btapu73ZNxlJxj46utVs3t+1Y0GX70R9m/mGsNyiWxxY0BkpT8eIQrmjAq1YDZ
Tt9u770JJnVR5cmPdwDnXK6HckCmBE+5VNbMUrQxjMrvvr7UAJmU+AquIT6BQCsggL/Q7lGsfx89
Q7pRQSM8JfvL8xhz1Tyu2jbOwMIoA18e4CFj2ltoMtIhRsT8DMlWyJcqKhvokeXp4Wl4S3q+ERx5
Px5myo8r2jsy+HByVgkUOqTunIDLjugjbzcVZb0lTUfnDMzN/gImeoUBdnHiiikFeXU6gCzKAS4d
CDt5nuhYXOEjQyAtBao4iZXH+/wCjBjcwWKuOIxPhc01QxauaYNbNOWV/9k9vOmyyXDbtuDzEX3W
0spsmbqL4wgVPbCok1TcXyriMaBNYbARlLe793lK4GgfZ4EGRqSrXzag9YbNCzIfXJ07QPRl/SUX
MvI5hfaS5bs1KvmehArBg93Qtbbfhr7v3dn+iLYLs6eOs2mftkR+apQcdJc058FS/KuLS1cHdufm
wIyF2RueyqZLinVmoEqOvf57XlZzatXgMiUhQSbAVYWSa6nyqb0zJLKvFs6OOHHVp69iMOtPlpGQ
Cfibd63CaxMQOBrhwBKQV+v2nJ9D+EdTtP6AndG46FVmGK5+/zYUWKDm1LX4qZ5/KOpfRFd/cOm+
4i7VSq8iwCO+hqVCt2myQS7xFKux/mcHW355cf3l4rY/7vVo9AdqBEOktY7ZNS2JWRYv3R+V49+2
OlMXs/8lE9rIAo428FDrSZJ3xhWiPnkCzBs5OnOAA4iTbYho0T7jV1cVc6+yavkhQDzk3/kjTfWO
5AO4slYMwyKLMfv2VOOn8EcJtTHunFa6fWXzSlR9l/VYJPOtcH6EHzqTTSFqtuvnbOyPql5RrpiN
XYLOe2VXc9pBYbfbFLJ+StUKgveBtx64DQzK3Ox4nkAj59KflffUd25RAWcbsfAVv5E1lttzAKA2
Tp0ZS1ykYOlEfAd2Uy+t/lPgI4ZHz0VRFhGi6ao4RaFjZaYVw1J9iSzmE4GU9rzrovhNreJYL/mK
IdLLSUmliFDvY/itR84kAlrb8EIzfvJCBXBCNNoPgUq791ZBITUDylbCGXE2cnnwk/hlsNWDWeU+
CeqEFV5wHuH2mGMhe/1L+10Wy2o4ienRibP5s6Ayu9ry2QpO1BykQ9X2paJtqoYzkJmIHkdijFfs
6Aj4FuqgRa28ZolHTzMjrq+vZNFhxGB+DXg913jMXkXINPC/7mNlfKadxxqsVPNfke8b8nl9rHnA
bYnNUDJU2Ov/r7DIQXm/IB+QKvJWAEZMM3KnryZ0/dV43NkOSiEcxFSGyWAufT0JiwyMS82xYqa5
zJUtL6u1lnD7BsTXp7H646qyhGiuJobhXMORQmFw9Nuyu7EaWKuDpEWDU5MWL8K7XdirNctXgchL
VsYZ20TNHC3XJHIJ4afbkjwN/AKUS+2VCaTzu3RfafGGZNW550ek9YfKUPnW1GDwqyTa3Ii8vdrQ
QdYbFRejGae8O8CnGlVsJk0wfCL2uK0vyLzem9rVngIaPHDjqcODCGLHOipEsELvtviovaOuI3N4
cim3B4Rjf14cIYB1ciDY0s8hqPP6N5IeABVX8M1P6ThiM+7msO1gOo3jQUxy1IbZTji1B/LxUH53
HnKqIA/VRsl7okmbtSUYPqC/1Rj1NCG/U4O44EK7EtYhE0Vvy7VDypAaC/nbU0PY7jcUecFp0Bjb
ek5TtY663RxOvCawLMv7mIu8Lp1ZGB64gY2IMcmCOJDMl2gB3WU5j69Kzh4rpkMQzPlK8dNjzXq+
f/NCPW7/tkiSHz/KQDyNCo73o7F449X9t9jcPC6dYvjPP5HL68iFJaJYwh2DaWO0Gjs74AZPWQIb
4I/9obGBlFAm2jWuJrU1OTcIO4ove/OhY+hineikXBj6qACrMQlI+igmTxuIw2lxriFHU/9CiNz6
prwgGaUiNm5xnXlRqO69SG6i0gbf/7GtsYuxY2xl1/GLGR9RZNXHM4lul+Vvfzzy9YQYjNXnF/fy
Fb+XWmRG/M1/S9l1JsucEAb1Srr9EMQ1kgy27/FAL9oHz16toD6CFzAajzB0k3ki3F4B8Y+HSDeW
qdvqlbjr5OOfQPdba/p2pIKf+2YsCuBfvi9pekwNxiihB46nWxWpaTF60y2qFHvRIReA3n90Sx5p
qdLs3mgd3tvHIEOWEQzNiUYD3eA6Az1G7oNNAHrEGUun1oVgWIt1Ayq6FRZP1enTG/haddmxJzKQ
cJJ1tbM5PFnYlD47AiAYHjAT3iFp90BcImvXq/oBMZhXkWKnbCnce+QhGJPCEqUJWK+tnZf7cvJW
pLaDj06McKvK6Qt+0juRePVJUSuPBZcyhK/wEXl+THK8o+8uBDnpLjIiPZ11UT/Nflna952rTwbF
c6NHfZr1fpXo+RC4CWL/burBIhGF48bU+5bpe13CkV/NwCaNt7lBurXk55/2crOnqKMMf1JZTxnZ
7GueeK7vJohQjoK0BzTjrPbwre0xPEp3TKigd+0RAuxVnI2t1XxI4tbI9zFyZZ0fXs+3+Ljt25O4
IYx0auWz2BePB593W29zxf4s0YSBAnADg7nJnQVW9ojYdnQ85jZVvGuzjAaMFk58uuuO45e4McUF
AmCY7RuQVwpCFEW/sHdGZRGQjCt0g7utr2CpMLZTj/VpK2CSGa1xuVq/3lqIRRevtcf28APNthtO
ZVBKu1GaBU85nJBsQ6XOwKM6Tucc8vLIbFFdMRWKsQiQrIY+RqJClhFUwldIX+gM8BSm75HhdZNz
kduvINTAVPOE7lIK+dQ91NeNSxz6boS+Q/cjNE30I/RyYWknl9Px8m4InGm9LeIlqfxUw50lh4Vb
J93y4/nCgaXhTJZbQ2ue8Yu9EG3YXj6TNpxeIEE8pu3DPbXErYMByg3FtAoWguMK+7vxj20j8Vje
yYhx9WOn1gACqx2ECKDDYFm49c3MQRto7WPnXnQ8oOJSQZDTrYuVEIkcj9PDwwPYvM/LNc0DLEDc
4qaav7P9TN0mUiBE5LKtOQycH1rvv118VY+SQ/9lirJXgjmVvjjcf23mr7WbAX+ipXEzo7Ovem+0
Kde6E8is374ecQd9+DSofK/32Hk/3q9krcXqEjnm7dIEFiORtt4dVa1IvMoAork58sHr8TDvwPTI
9BgKqgbF5AtNlo2jYPZ7Qrko7IU6zTr3RfBvRmkqDovO3+UtWFKo6TZJs/QYmujYZ2k5cSUKc4zY
t/i/eaM+SwS97k+xCR8+eHIgnqcEsyUoaHG76/BgpYo/BuTkxP72Ouir5aG0oVUM2P1hzNBe/emC
V1QBlyrhbRaYLTrydYXeqbwNASd9LTxkk+LTjxZobQ7Gu71EKrqWkKLeXfD1ALOLmsaQnLhlz9bE
PafcJJfSWxn7V24+gtMl5eqjOfXbEoKjhG9ZZZsQr5Rk1qFAl5bDpvpx/w0vlOr8F3v5YMYRNmUu
Osh7VMcSB+OlqA8K4vi8h1tg2+49MyFS77f4lMOboVbjjmsBV/dBebiO98pjkcXEY/tbBcO8RGXX
JizNu+s8fVCqXbPxbhhiVBEziJXKB39cmYRkbhmoPI12D+f/m+QFlWrCoGlMHK9lb1qgk6aFAKqK
MPoWmUMP/sGBB0hVzOkYbo2iV/W7aJrYBWozZjDc3PhCHU9iTP/C2VCTrgN6UicjKhvamjeCtWYp
5Gf1egX3oFM7qrlXd++7wgInHJdXtDaeOaxQxsj0owreS98bLaRKhZFI3qMq2aQ8ieqefyup0h8J
L/pp3v9ARByA721NfScI1e3/5Dcy5s1ayunkvl/UbYyuti6mYnVnKcwY9es0Sc7EbX6PtuZGhvOL
ZkXll2zUI9N4bR/driFSB+hE7ZedwNdPFIwt9qdY6PQP8Vp88ZjMYY5+XS61XC2Iu+uGOh1ezvPI
kD/Arfc4wDckKY2gtqCd/OsDglKPSiYkoWWGP1OlBHIgELVS+Fch/K7icFQ05s5ejBrz8Oqxfzyn
lo1JQZxEB7y4TeYc9FktfR2pHireHq3PH8gXyNGc4NJVRH58E98VKxRlH3eehPEgK8KhRQUUAWKp
uqbUwL0JPW3jkWmfGnm7WoMPlXrjdbV/waVci6UrGHseyv1GA/8CnxZliwa/5IJfBAXYEdaCTA1P
KHbyHMiv7qzZVLo/uFfR43XKJS6vsp5/BWnyzrne4lQuQl7AZW9hXNGd/wraeer4o/PJsJBAGmNk
EwImg+XAFBEqqWCJQoi2bn9uounPQMxqBrTycU3IlOUdGxaVM9XO1tQzv6rCE3nbzR2vPtbVjjI7
tBXGZBB/MuOjeu83UEpg8YGHb9ZbhjLul0She/N8Opi6UKyUXhZDVRHIUdPSFr9lKyoRHfYLsBlX
A1qHGhrYVEy1gdiS34sFiyFekQrz3dUQehRQdHhIPmZEsZPzLz9gXmats7CZQDJFSI8qcCWLDUEw
Qd1efmfEuncmhLgAsmafZ6rX4xggFOvudW5BbQsbv1QRumUAMsz4xTfKDTwaQjYKScrPh+WFUB1V
wbxM9k7uLSfzzATpHCqNrMMTHuGkzd49OaBT7R0UxgJuXgq88qsdrpD9Aj/xjUeUaS0ux9C29kfb
GP3waK+yX5sv/rZL6GyYinuYGymWZ51OqA1MNgWEBeydsxri34h+8RaxBNwMIkM3vxVBgTMQdVUH
dv+Hsd9FDzQbJfmBl4dUFMmMEuNI4QK49Uj4hiEMXWsmtJ9L33Wg8NkWeIJFSUbAGSQewonU3+1Z
Hn3bTL49OGewYXXn7lA9vIuXJqA++ek/GIzeBquUGV9FXtWKvEeMWkY7DEIVZtxjMs+3gQykRyRs
ORtCjDHN/IOxXm2pmesnTfnhkFamBOHLSEuZmjHQVaf3awU2GxyYJKnnb+nj2I+iq9/nNidScGBS
lcaMdGJbWslRpS3jPx/1Yb7y3sIJs9nQYo8Hr9cz/J8IUdBbLztj0Unk2T0QuzwQqQjJ+ruxQpwQ
YMwe/Ofe071VZ/NJU2CQ7Jtfyq7UjjpeW/t4szXMtYSQD0ohQSX1pTM+F9UUgEnZ6c4DDNSJk5bl
kLmM1TTte7D5EBx88DGxzpZmme2tJpNxxXnzIeDQLEgRSzgZMmVJQxZlJzE0yMYqwC0jUOIPKd8s
oalbDXjRbNgJObmJOi39LeJ46f6lyGrsrwQYus0dgtnhcNW2o3wczNxenupcW2as8DccCfNPHPhK
cWn4jknXZ4es30RZ+jYAoz3dIOt4lVB5GHw36jWr2szzz5ooYMi/16QKNAEksZhWCiP72ThsG1D8
Zi1sYigroaT8+e0pC6KvQPk1RpCNwEp8MTMNsmMNgy5IdHLs/QVP5dYjiy6Sz0fj3LGipAca2J8a
4banQc9fif0LAHirzePlWwJfRnsxUh/JxmtqTiuLL03V2+3D5wFidkhETxAXXFM5bohQz6NeUOtG
I6mb5BNArAgsbA0sermh1vxzy77BoFXZUCFflJAajJA/Fmwrmnf642fpKjdWTYGo19vXVWXTzJZj
bNWyO+3QgspCFYG2XzeQsBUCJAuan5n18gVYXBtRbwrB5DvnfTgeYo18SNOR1kHcdxDCH9Gv+g0f
S9T6O/M2BIqV1MscCDVTwt/PGobVapPcoWt37MKjFbqfwGhU9cPctagfq0oYjYPFKQNHTWQeyY+B
h/LyZ9Ix+48t+cydZ8ET9wusJi8voCOYLr91uyyrC8EvW55eFUrG/Y/32yei1y9w0tXfvDZ9zjqz
xgZrHOhlWKlY/VI/yYhAx3jL/qnoBxDoYc0aj7v5mohcXeaoYjp2jli3uetK6XmoRyLFBsSrbBbE
f9RUvqx1C8WJHIuwbNG4wCJvW6xKVdhHaTLJDmRD4BEB6ROHlUCjjoBHsX4DePUivMleaome9/sQ
u83UsHARgd6jeLs+ZSQ7gIzAlQ17vc7v8yUT/oh7VKwg6HgohqysDQL+Mz6k+6DrAOtvT/zTvh8F
8/hO0vnJHIEXIHumCoe60KehFwrVNvbD2/bROhD4r3ton/VxyplIzZ4OkfykmBISE++rx12AHo+G
x18sThC6xbTk0SlFjIoaXi0u5v7zF6vC9pIAqnu9qvsd1Xd41HpMJKWxcruDQo8/2uAV0GFybsBP
f4Yrdcs2RkZxGZzChhNJlSgLG6PSKAo0cLVYHQArCUkW0UqZBhEImLNiOjJTiKcWwK0VrrhErREj
/alY8bXNfqPIlxhT4ykcC7A3n1nfh4om0Jr8Xw0J5T121aeGgDkAJXalcrtYf4ZdMInt21oRvOjs
nLzhRPYjtxvuWCd/r6tR85H6hZyRiuL0U9J7+203kI6uxTWvBA7INOLoTsTAqiJDZO61lFnuj1ZO
dxA5ZNwfZsN99WCu62FZudYiXhvjOh3XlEwdpnc4BVne39EnDWqUGoa5lMNx+ZCH9Q+F8oIehCl1
h8+Hi+aVqP4zGcFZeOCTMIpRkBNVHhy2VyJpBXjwsmUwegQD8qAK4EkPCIefHknUeLaggximiW33
ltoxOPDUXKfRdPQ2XY8JLsSpOf48QPL+aUzGlK0TbC7gxg1ZG3MxAJvpjbrv/1QGyj7YN5QEj9DT
Ii+Rr8XTkOG2tbkwazK8KvcG8eSGib73cyZ8qlFX/Zo71Ojs60Ir6//TmqABT7mSXiuSHvj0jdz2
b1PaCbx/AP7apcWlnykodWQh1O1INt0iaAOhuGWqvNU3KbnmXoVJ43E4FbBSfRl733SyLd1QL7zk
pgey+Lbstk2G4oYLO4Vz+zz5c7iANo+R++156bvJl6mdbn6ih7F8CXSolrrPdaagTrf1rkG9ZEE0
fAaATFFTmRKszyGPHstNte+AAOXWO9wnocnO70B8nBmI2hQu3HY2jmJ92GglUuXUNTayj67uSD/F
5jmWL6QAEp/xdz8V5BXrligH6DhKwYAAGTgw8aba2xjOcGJxVQ8h1MTSO127iWX3e3EgpVtjM6fF
/l9z4iN73CBDQcjzQlpbYoaa2yku9zOIizaulmP0j9p3toRz5ZlrcBPyedb+7GWXDl9eQWacrNVF
tsK39hopzf0qiDUkgYLfNTtk2a84siNg1Twrmx1YuISwvr2nJfpVdaEDVqyfUzsaTS1puKV/UcIW
haZGRyt4OqSjpM9Hok+0ovi4KBlUO52Yv4e0bQUzLh7gElgslbajXyI0VYeZA2UY/Zvv4N387JwQ
eOh9xy/wdG3dIaFFgWflye/JnQKiIWGyRjTg/Xe8lUKg2vQR18Xe0Hzp3KdIaornOo2NbrzDO7xF
e8Oho9r0l1L5UrRx/qc8HAJqmeOhUjfkg6iNc4pftqqIl9gXoY8ZKsBTbvKqpox5ATAFv4jveoVe
TUmXT2+dMX0zxU0CBxRdYHByoSttl2K41Emvub3ZPxpwIc+wJtjAhX8zLecKloeyq64znQc4InMD
Akd5k4V/md/2Ltl5VUgysk6TuQL9cBVyGlwxSa8zik64Q8hHxCdPps+krsY8QlLUD4V0xhRh0nrq
aL1t+I9JJOPz2PBynAhEn0R9I8hw8SUlnAygZHgPJzTFukpBYMTyFIKCC7gPiwJTdCbNCtrH/MuX
D5gr7T27C1MLT/nfvUZE9OngeRXVUhBPQOrsBSVEfKiHrl4wuygGtGnAFNFA/TZSTQZdjSye5rfO
5lcbGNAq4HcdwbP6R/GBjfG8b8D53eOeBVsOhTzC+v8AFGUxveGSHlYPe83hXe2XXJWWaXlyyjLK
gz0n2pnHrO7W4fo3S+haVZgHgEnKbsMEIl3sver6itoke2M0RhJWEjglv+1SykqjJZb4AE7SzH92
TSQxCINZHTuuQsiMsPJZfBMvsEPhttO6S8iR1qAa7pz91d/uuGIu3rmc6f8MAvn/fNlktJz66fvT
GzEuyls6KeMu7l3wJJ2YyQKdwCx/6Uf796wrdJdQ+KAo942qOcuOTF7PLfZ9iNDvZUn2l+bfpMfI
cFfM1//oV2p7zpp61wC7T1V2iMD0v1rql+UBdGaiNimMdvxy7L9WXgP4cNJg/qu1lnSnRzKAcPYb
2AobOaNVNpgJmbsXqo3EJ4be+yHwI82jd3V+vsEBNJckVg/CMPJzCohgfioUygxi7kTRVbF/2/Qo
13aeOaRUWKVgCaueiIzrxe+qlFdbnqdMDbNaj7jZK0NX6uRFTXv0/rNgxUAEJHcMjbhOHXb0X9+q
Uo+m0FmsXN5p9AEwg0Rh6wBvUFEuxNzr9Ic0+egl55oq70IB4Tut14O3Ca1/gt2xsjusXlHHINRg
t8uO1wmtp+DwGLnC6sB04tT4vkTdKh9PsVB3AVyH01jETl4DTiF+gdJZqc5EEciFwL5tjEPc1y3X
kNc8NQlElxtZoiJKTDogqgQ7wfTlBWBU33rLNU43SGbJBbQ319Q3hb0DvlGV3YeQMuVGppt+9cqC
c86Z7zLOquE+EICwiutFuUjWXVrRUNv6wOCj4lRT+JdxD7kXU5MZndtbN2oTQ6EWnqktHbSww1my
pM4hJ+KI058PUtOnnmDdmq+Y33KqKYfbQiYOL6e5cXegnXkW1QdxuC1uFNUMe7KqLBcHoNnTERO6
0hbZvpsRsPai8ZIxOuLJUdwdWfKgRkE5MjUVjAwlcS2RPZwhQmDPNCusAuWftzqBh3LExlRkph5Q
vbQzIe8tBMVSN3wsNkdK+QP2D9sJCAY75uA/FXqNxwkRpAPkHOMdql9Gn9k8wVya5e2hk3mtar0G
GlvPOedf2HDQtfObaFEnRcGP4rH74gHa0JSp+lGn6sCaMYISILQLkCD0MZqdr2CfB1V7Ml+kkmf/
CM+ZHutUl2ca/g6mQ8tE94E7KOeZR4s9D+tTWEbeEajhMi3R4hmPt20p02hJ3OP94jRszNfLZ5xj
HUGXbH9GE6bzsgu4U8EzNCZTvV7KMU9PRX1wXsyRJjVInagvFsiZ8M4GYhJRZr5CBvJfeKTXyIdh
YC+5uXg7pgtNrzTaiF/seupfOfQh++8E5EYipUepXGMNzM3LLruncXpmxXjb8Y0LFiLGB8pBjIG+
2BtN5hPZQiz9iPB7h4IDywS1FkXwruX3FudO9bgMgKgQREaCBAcImfs1NIRyuDW5tfU8NMd0WzyR
HOFwZ7w8y5G+xFeCv5inJnyxGXAi0s9ndgnySGZ7Llpnk/9gDqTfypGTwTwAYi3r608zWKlmYSA3
obeBBq+BgOwEtWUpce5SW001X4IqK7qg3Nrg+OPCdil82Uu0braDyOjRf6DJ5f4PKBHIviTIJXmS
REbGSONpxU6ta7Vz3BsfrLc4PF4JzuONr6GenWpZzxX5l9G56Om3w0vuw4dmwVKZSQo/LJTYHdfp
HhJ/SfeDcKhnb+bz1+4C7wMqv8YoyFEOSpszAiahnQfDxL22vL+2gpR8lDsAWKXjnrg17ZKxSmES
xxo+SIVcRUIm/MabmiWpj0UYxfnSvVJl9MGIo7oudNbLstRz8AXgp5Ww+SynNcWxPe/z6N3UmHB7
qlGufQruevFVCZQNrJxcGpmLnuUjTDfcHYBHutydqq7o/rtbCIDuv10t1UCKr2jfAg8joWlA0Up2
fqEzNARnLEehrp1sQujTyhkXkJgBiBkb6fz12dj7nbjR2ws5vyz+V0NckF+ZTyp48d/sxXh/ZpiW
syg6l27S0kOVmx8q8Jircb25DrW1wK5j/lFCTZ4P3S5YN0SvoLsU1OPntrAtmOwk0sE5BPcDx+lL
XKq1UeZFMwy8O07vl5BCjtGzGUv+sRjgilIe/MDaNF6yfvTtIm62VMcw0rKk1UUiRCE9T9/Otco+
LUdEkSfi3RjW/GgpyOBCpKAgkKcPZf+DpiHMD7d5e5XYcJm5C9S48RTcpkC4UtrkXQ9l//g4sYJb
d6hZthSdcODfdfjfKWZx+4AN2+qogc6Va9hL33ywPJE2gB3m1+nsTA/UEmZQwKNryvwl/o/TOQiY
g2hlOvz+PimBoGbjc6ovfuRUv1hMiMP9UbL6GmAJMkmSHuAcVCl+V4pZjcKWVGC0npLJpapzHYXj
CG+7nnj2os85QpVHhJnZPcxfAtrZ2JAPEfaJORbwIbUleLSza3LhQY37hAitjknsdSw0d0ZDfyD+
lf+kT0OwBHcY/jy7AopH6K1DICV69jicS/QV9v5gsU4PmuG+pKDA8hhp0nLAEBHiNj4osjBOdkmU
LjQ/WUMZZMmJ+sAqhGA8mm/xA8Ule9FKDFLkcBzMjueTRAQ5MRBlfE0zb70Q9Uqj71cClvG8PTKk
pSF4e6PW6yvuOomXrDJ7og6CxQywTdhu+nm2TK5vdi5uMxYcu2Ymcnou5uXC2onUjL3IseLJBrf6
0K16ZqZBDJoeQo5xcfRzhk0O0YAssZoeDUplt3iSBDbboH0+qSnuaSBrzHQnAu/4KDrtdatZDUMr
vT+NpKrTbk3dYzLbYQjXEdVindu+4LcAz2qsYRrp0spKspnNuvH5j2DJOMr1IKFAKazjkC1y7Oxv
0/bbXeH3ynW874f/LyvOcOB1ChpNxqtpXfTySZr2ZxHJdfYFiyCzdBg0gjB2UDuntgGVq23Li3T4
nu7DXKLc+N9DfAFXdZpNRHwPdov7B7fDkPD9Hd1F9rvGfKEYbGY2RRaxqmzGLOWpIC+Z3jUumXJc
zklU5IoS2ushJ8pvxkWuVmQRqx5ZUulfBMgJL4HD5G30OKMuxJ8vQ5i0uKZ+9I4wDylEvur9sx4i
Y2mpZgXcHVVVWe76y/MLzZ2EIEp2BxN3s9aoOIAxnLJsmFSJuugS9gzS+3f0f3GBMb1m/zRl5hV3
qd7/rAO7J0kxhhc0b0OVSJL5tqgjzSs0VLJ6EXybpBXoDI2h9R71HSEfOX9V6ljAGyhrKEWTL+DH
TuU2kV4XxRu0Bkpt1wfeR8RD1S7+13G8C9BvnMvxYoaD7P05h7y49U56YaM83lftYuXDcQnrFJoB
/NtxiDOZjetJM1vAFQkRTF/NN/WNwGGiag19ivGxbV95H73Q5BzEcKZmC0mMnAgo0Fmp6NU7pzfo
5YLZ4mzi+33c+8xSgcGuOG7vGTt9hIJCDvffqn2t5Sa2EUqsRrrZCsxDWNGGKnzxv6T/ZOeToQK6
+MnT/1e4qeg5FHy3SNeZ/ZsqXCxiFrc1JnFbOGksrf6hUHdk7roaUwewQTna8XhVw/DbxpbnOQgB
9EMt0vlw+iiYClr1+2SZloqzxX9OQigJcKSvVo8KfbE9i5W4O2G5noWpSD9N55sGNLzC1vL6Vk79
GXogcFHtHKUDr6oP4niLFrm4vk6aRgqlllnjC4IYodO+KYvK+eFcQbclYfV466+18tUr7AtLjNJr
/ltciftw9OykIdX+9IIOMb32gvFtYeYkQg83qbHE/SSuRlfI6nNf/qyKtYAJC/RYePSiFgLPBgDQ
SDEnKYP/WegcTJQ7dB8Zvp8rPjv2L28xtUjbIkh9qfPSJrFqYo2wVkKmzFDGKF8UhC+zl2dazscQ
JIIDnhbJNeseuucBRLKENjq9ffheTfVX+SdWF6G6ta3BwqNJhSNCFFntOu2U0tXwfsx3iMAM//TR
BeJDXTFR/tjNVbYS5HRwRdMYhHP+iW+T4llP5f0vdtkzyT+kNUI6tO3ZId+6sYsN7Wc069az7ant
waSgFttuYTHaQeZfolecgJs8aem4S9tnKq4g6UW8bN2VUT+f0r47DETLtROn8A3SKRkTNNkerYe/
gJhoRF8liQER7Dj5P9nndnlgZ/zCjxyuHkbzwApB9HzZkV+CABnw/2kX3ktpDZmhJvEAl8an5DSQ
F4DCaCAS7Mr63ulDvvI1aoYuXtcQ43sYJdf6ft1/vOEghsXh5FMF9HE5l4ZdLzrP/I5//LQvWN7h
bKwxCjz4ct2K8/+V/rdsZK1YQg4OzTZjfD4Ie8JvOqV3IIw808PxBsEYeXevbSUBEpsVsozS+4O0
utVxaAAybKppMbzo+bPhfNfAcKtAAQK4LAzqqFyLMisUoquViiyPa7vZLrW2UyvVmFNdsNhw02JT
DHiKALMbueq6JPJ5cBk58Z8YpTGIk74piA/d/6vbImlUt537G9rj9RcMBOxXjILz+IJfOPkVQPHA
Tof4IJp3bNETceeV3nGS0mGIdyN+u6UqhZAbBiuTfG5Ct17yRqR6lOPEuxtEzujj5z/MWMUW0Qhv
zJvQpLvBpHmpR5huPOQXaCKkrgtXxrjVi4rZdkC+PtJHIDM6UWpPJykcBb1BfDZZxpKvtRDf9wH6
HQK76/ZOJfolvYM5+vBX4iIyx/yVFReyWzoj4GFIbDNhczYsHES2gZlumjfBMGYOd4Yq6UPlw8Z1
lzzEjH/lBXQVDD4YUAIMkgWSc6kIaMnD2mtpym+lSp/PjEzSxS4R5cK6T2IFrHeeXp+gcCh3Ja8F
lEclu8Ry+qCSFV1zm0OxhHmnsksQfKfr+//b5q3d/C2PJfy5Z4+DUNJUPRb2pfczn8abAj4Azkvz
uh5fC5UTaw0Fr4kaF0SwWU1lxxHVLujSDDzSTWy26YUAUCHR4zOMWjk0St14PxHHjamxrQvInjiQ
USpNPqv/QqhiipNv5pv0wLewe+WEZiauWa0xk2TBE+QwQGoX6RfgV+/3UCYfxTTTi/xKXbWvcO0G
T4kExoaZGzHVR1LPn3gIxNimWgQVsJgPkVBMUxFdStVdfzTA1WqsThjemz7yxAyVy9Eedesl1IjI
GjxlC4W1QK/UTPcsPOSEu3ZnfQZWTWrztVfiqNz2Pn04UULlysgkB2bA6h3kB9v5DFmH6MnuNSo8
hJB+8K2calEpkVIuqpzmguiPnP2zvZ6x/+rwCt5vOBum0dGTywducJJDoWQpGXQrI62MoZQeqnhz
BNW5gFzTgP9u8zA92hgHkJurfC8vKatW4wiCrdfq8OsP0BS+SZaXVFfstLt2hFyJNKBbRGAZ2uRP
qqB5wIpRnXXhBkLdOnPJpiNw0HeO+OpHLjaxbpL/a9Q5exyfQqMoFmVDwPmBO5tB6v2TzF7V1cpu
DwY9XsqmGEm4zSxk/dtqtdGzM0PDzoVLyYvv8i5fF+QclENNSKXGOK8g/Qk4D7djgou5HoNr06vL
NN9Dh7dmsmdqua1Sbl/DnKS71XPBAH6GI2ksNzbxnzjPNy8LNR9+X/DcBabr9KLT/WivQ0/3hFbZ
wcjnZUS2nmHKOeSVFvKaKZUU7mUSnS5MlsxYG+Hu1nqdf1yTZJKu5KmUN3xygyEVMEWelrSys6Oh
49lOz9J8jJDUG2NTfCo0j/o1YNV1KWfh8399OB0OARgKMkFPoFB1JO9bn5vgh61TxnvMnPRbHvVC
DcsqvBr+nJJB/c4bQ7upZtVlfnftatkcxEogwlWxkg5PPdHXwECr2kGyEUbTuvrIg7fUfj4sXRiM
1mG6F1IeVqscQCziVterhtbh6GYwGgnu3ryDOARxvkZImtcVuZ0BrdAnFWVp8Opinal8CwuHIYZO
0vnKdVPVP7x1Ujb62mAFH37DWBTfMvmXpYrbKvadToO0cMlhhKI369jMjujab61ztwgZUoiCllp+
F6MAU0cjIy2KMPh8FuTYASHzSLEzcgTvzVJK3STd6a4xolfG9TI35bNUMzwqRscxm7AkwYx2TH3K
hbWdiNbPmakhQB/axvuMc7FU7EVLmYCvAeVZCoEYZV1/fVNs6ErpBuk5SsWjMDmDndVc69Jhnj6Z
T/u4dU3rn2VIHoMsstHPGx4jZQYMxXh6SNQXO9PxYNVxAASfbNzMY+BYkRyhkqQg7gBZ11DS3MDW
7wQgJgYy4sRo8mc48omdek56/Bxg+FUcAnwVuXG5YuPidty2BtfIiUVYxy6nawa+TBsKiKdSJrKI
Nv7NGaVMEHWcrAAgyCGEHkU1R9pDzR2phtfvSxmGsSttvh/hR94pM+W+IwD1yXyvq2qBq2AMEVyT
3/MLZunQ3FKIomjmFTzX6W+ixc50YrFHskgf8yTK5qEJ6/Uh9SAMe1dV6N79ETjbqFef5jGEp2lb
UEjjlGcwnXuxdWIAdLBJOZWPG+pEQTNozBGw6qIwlwHMXAT7L1LRm9LYuIPaoj8hy0XP0ZGrunCx
gIePOV3CkTBHY1GBG/TKup1THFOHuWoG3JGMCRG8vXiJ2RCTM3V5UknQdcXies9QzFEgYUdtzLZ+
1ScUR0eTnrYr7+9mbhR31RXDGyjQ7/ufyaaUr2BXDYmhebIk6XOtgEO3VJc/Se44qhgQh8fdpJz7
V5h3ic2jyWWGSJ/tga4iKvB9+EEbRM5kJDn+kaIKyWHjZyOcjoGhYzNMk14ELh2ibyr7+J1FTca5
DyFoMvqH+ULZzP4QkfJ7z8WfzwURGxbscJuFm6FT7/ZAJcIFm6RtHCRFDajr6zlVGqdrvjCP2hkR
6GApYPSYEvMF3nhvAq74NlysGXFfbMGokuUjXLb4S1ZLicQ4v5EIZgbJiRBHlis9asPJSiN78WLj
lz/T4OOHaMePtbTo5LnxwpnZX04azp/8bEIN/AUrJnMhlF1ZID5Qi94oDjiGgpQqQSjU0kcX8dyA
rBmcMDRsOLupRNeumqAa7VFNnkjRdHabtao/mMr56bmRN+UIvlppY/3gNvQ/RqB2pLXj/DIwnEdx
MhMEmQmr/5iA+sSGdR4666WRYGFtLner+wS41UeGqDVWqWneRuCZUISQSI1l1TCg1TcTs4+mmH8Z
8ERALVPeicojgWF+BYuxcUjCw1Exhp6wMLLPYZb5FOsv+sokSN6yem0PgJJQVgxxGdtGpujMVUcw
buQKp+bSiSfi5OdHx/nh6dyIQW+DUDuUAkX71OdjYhk1RY3inVMuVkAAZiAhRzTav0cZGzcw+kCW
eATO9iKTeToEQM3RmRJOiyxOx67lAE4vK06jNVVpLNxbyi+gXfIBJilSsK3aGdjVfxAGw9K0H/Y9
NjZSQuI4f1H97L0w2BueexxAQPwBHCBd03wj6QFu8FnIRgpSwmBjFjMhx7fXA1A9bM93/rXna1kD
dSog03naa48KRXZ5k8zjH3ulvCTvF40w5nIjQKG8tJy//8W+bzIv1iRBCzrs1ooBxrSPSVWsEtsB
c8uZ2ox6mt4rPhOm6AwZWfXFttl2tUs7do95R7KWpQkXEfD0Uv3RtYz2XkZqLwGAHUIrm1AW59ti
IjerDBBrihkLwEMw6nzjqiUDvTzteZm3+2Pfp7JPjPA9+yr9eEyM3SQ/E8Jef9jTdCYzw2eOwnkE
APQgsXv6R2+is3aM6E1ENH0xkv0xSGwUKDqO3oo3HcTsIzMyqRnqSdaXkJt8PZRcbqf1OVZYj7aD
pQK3yjh6hnkKLBdmoOqvHYfFQMQDCnPTBC62rwDjNroyNxrroMHj6KLJDwn00EaGL3R4i6HlrVio
ltW8DSYYI/DkAwfQVyHDIZYuxeCqpmhfB62gf+pP7nmfyJRLuYs575ERkXTKS89kuwbZoRO1YqVm
JLhFy2fDzeNmej2AzdjpfgsaOHDP33J/p/wHkm6xBcgqSmhkUuJgSRQMff+H7cqeblzELjQfk9d7
xld0Q33qnCV7C57sTFX/o4wQO0aqA35wpFvEc7AD08US7YGxvz9Kjf0IxVqVJuiG7QTlul8D+2W8
uCPHXWTUHHT92EQ90fOD6hYfoIhmAwC91O0TivkJ4Ag=
`protect end_protected
