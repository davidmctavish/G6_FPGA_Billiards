`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HShNBWeCwbuaWSKBgN4WHNQ0Y1iLKMSWw3jbK0ayiEt9filvm8jCWigV/HWtAjQPRDoFU0sKb4dg
HMaIGYtg7A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j4hHL0EZG8xpQFMA56qfg2r5E+n21pRX+7IjA/Fvk7Iab9MDtJx8F6YFzUsejL6aPcy0cj3F2fax
Jafp0ZrvOolhhN8QYpYaLATSzE4S1DQLmIvKeSdhik3fJDEvpGfQ2Rm4K0fEGyprrneXKMhOEi4U
TZAx0qqqcWWf+9Gd0SI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XP7qXI1g9QqmmANQdMFoGL0qjwmzT6Acxuy2fz0LxUxc/lv3s8l/pOzispLTvfAXBRAQ4IDzFljX
kdxyenvLZ3KavsCgHIGPdUguiCU0u9kLSCHVVcmCctmhDLfnIiCA9wF+akHZlHP1umtD9wmNzn5l
t0TbE+SoF1dUIchS8yny8Fn+Ng4chxNxiZ627UwOvPWF4JwM9D9z3+RfIcYYOc68DGFUHd2AWnDw
YFVbY8qm4arjHLXC3gOxMoYIZsSwL/fR8C7135WcIoHM4SgyNPI0Z9V/DDmr/UdRcDFCwiW9jTUY
JRvCJ1v1VDqGgMriuUfprb6e//GxiojCWCTu4Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p5UQNkIZbS6/9hBE8fGfrlwztCVXNUk4DwEmc97S+4SYI+0iwU/KQKLevSF1/stg9CIIZcWBYer7
aDRMeJmFudGmp8XRIz+DfVlek8Vb3R8quJP4EgO4kYWbWJ6oFhZXN0BHg9JzsURZS/Nhm3JQURjJ
eHiVIKlnrjkei59LboQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UdoNvOswp7y21MBBJWmT/aRz0Wcp4s3vrTDNuC4hYz2ifJ4lOS9YI83O2uS7aJ1VWJv155eK2kvN
mHlhA80h2T2jnBTJ4MdfLk9Hbw+lkjp738+qRSvqX9XIXGfYrMBRthTSvszPrclal8FrQAaOSn+m
U2IZ7GOEs3jcSFiE07t8fesve4jMSe9Fy0Do1VZl0xpV2zZXMRxsKUf+XAEuJkPz3WY4RBlmHBHS
rJvKhDDB8iImp9P0LjMlQcuoTvKX9DJqHA4mLMfVW10WYSOGeMS8rw7q57k17k3wWNmzOegu9DtA
4queOFU5Lkrfwu9HkZdEIqJUqlB26q/CzpBnRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 414048)
`protect data_block
6P3WM3opyUPm2zcoDDC4b8ntBIZm/s2mIaa8S0HerHPVcKJ+ABByp9iY2Csks+pOdBsEIXR3ZiY5
Agj+j8ux6c+kSQCGCegdDQCIXbDj8jBtrYOCsH3D+x4gpxOesrATm4Qa/Nza84trvkalSoo1wAU2
o0IGkeAjTOL+zar5nU57LB0QBQL3B5FB3KHv+ZWfyCYV3zIE+FXj/ijGPWjpsK5U7aex/PtaoHuR
OapiX2kHa2faPq05fydLfsVeZI20u4DjsDbD1jSfsuzONniHQB0rY7k7sd6mTBfWR2uKzXYxv6du
y+NHInP69VnYL35CCCNoo577fEfwHOFZU8at5hTFQJGzVrdtuXDbl4T7deauqHbeplfUoMuNMLBP
JxDOSv9g2epcMnx6rbDZFpeFD2RXFX16k3/eqiaAe55hRD6IMlTM9KMrdGoZwexhpI3hs1nK50Mg
8Yo3MDUCkDVV1oHpm/CMvPlvYAgYnK9L0benb9w/hRTJrx4PGSwIrEq16fI7U85xLJzFQ4Oln2c/
0ltG70AalLCU5CxgcrJnrONO6FaloPPwGSyuCdcUVgen+CXxA8TLraeaZWxsH9UODKgj3QLiY+5q
xBZZ4Yi8Q1YTtvzbeXqR09ByyCJvtOgV4hlDpHDqC52wWJejmUZRvVo2ZaBd48zrZb3FBZ/mIFO7
bVmszd0cfEC+lOrDac97Zv4RtSfa1indnXT14yHH4i54MMfdHb7gcoU6TYSq8yBXDpf27ZdX5oqd
jNUlq0W3o0AkjevWc+DE9oD6vmStbZ9m3wGSiCuhUNo80xIU1DMak2gSmyHLsrEp2vregGFCd7ai
Xu0sStzhxdD9U5wWnXEeHyTwIGYNxXka4iZm8yVFisfNDxHIO5jXxE1TkGUk1G/qheobkHzrXPS+
NyBxhuwJwOwQ+ebb3MMqLFXLe5+kTLRXnJHbZ+uNML/dOls1Dh/7hoVTgklchy4IJtERaFP00lnj
/B7+WFEKDE4P1kuIBFnmCQ3Xs6+1ERHlZIid19cRmfzf/5IsDZ8OTtQUpT1XctFZDwk6XHXjfuCn
XRiO6Ph6qKTZHnyhFdzdQtkkvNmPdhQW9S2oDARMP4haG3b4XofkDv2dkzrf0+kr0511iuu+sJVl
jAtZORnWtrT5SS1nsi6Y9qrb4t10FWSnF4nDnNDgROFWWoz+XhZ5qw9GaNtPPLJ7ujobQon7v30w
LfmISWQkGBFJgbcZawYc1vfB0Nz5QiUnj+ziRkEouEeAc2IiqfvC95SJ57BzDo6/QOqAYH2Ou7jA
WKt2/TuCYi308fxZlsrM0yS0/dT5Trz066KtZgvCzbgxL0KEjlmtM82NOZ3kBujz3HSMPOz4fWa4
C14+SOU18IYhTWkOoF75XMxHdc4t448+AdtBGP2rOw5YdYEAF1VV/cpZwQzidtWvBoKCqfBosOMY
kov5AnxaYDLraQz00gBpM//CWP1BZET3C3udQXjhiUd31mYcgVgsWsfLGs339l/UOhESzIfXoGZT
zJvI2xMvXwk1niaROrxJAzohR0pkx56Vjm8tqH+XKcHxCGjlMtEVA6S4y0KlkBTlXsatsaSto8Sd
WREl0xkO+wC911eZU2sjOgrKkfLxv3u/WyUrinSDgZvJJXILBPP12PooPL4KxmYqkfqv8Qby3fil
hNOwvWg7j0MRUQLyT0TQ+xn4vyhTYNiWLCFB4ON2Ant5GOmU7awFhfzSG6Ccf5XB881PA/yd40GI
ezUpc7G4BwBVloiEc6YUA6DzZcPsh+oc3VLlLBNxV1OrntzWfoZl0ZFPoqFymPOylmIhThacB4oT
HDWabR4I3bNWdEMdeWHpU2vc2OuR/ArJTakrFiTcib0WQ63uI1Xgd3LAsP/E2xEMi3Azjmuxlp/t
HmcHd6QHIQbDBpmE4xgTmjY5d0DqTwYYYS8kaegk1UUcDZdPEY1Og1KX/gnoV9fc7kdJrlR6CuhI
wiftHE+HPAyS4sOzMlU+d6/TYgZm2YSU/9kwA61OpqExDfcgoId2u8LQXCfkjIu6wSRukWC9Ble2
+VQxDsMpEIGfSRWZp8kr7CM6P9ZWWHFTt0yhoEg+qfhdv0fkDyiI2mm7q+50vtQESCK1q1lYDdwE
mvPKtPyRRaDmPHP//bVkFCkjHaDIxasJpyw5HlXNGcipuB1SIkgoMxDbcY901Ga+sCmX/rgA1wr+
U8/gqeK+Iz1RQYkvs+XaZ7TJNeuY9T+J0jru6Ksl70WU7LzeXWt/bBfyC3dwzEnrh9EJb/nvc9O/
mqBpWvYtB5vYODp48FpDBGdjxyReaggNyCQzFkfmHiGFAd2P2WNtWwDXW2gmVqVs9Tw+l5u1d/R8
iNovi3aDfZRDLKxxEESU75KoKImcQp0mmS/giCnJWL6Zez7jCiflgfZmOlopAcWhkt6VbsXjzyFf
oHW9pQrFB5ieeUMfZO2ZpoYivfgPHREXw4DhTkli1pjGqGUMSo7O/C3RFyoV7GM2maVHj7fDVnUM
9JozTY7IyDYsi29KOp8OXUw9ymlqmvreNb3R0QHiU7sGpVeO1F3Z3KgNxXW8s8Cn916nBu/Yaxi0
Y13N73vfyo78e8FlCqupAlEDvxTiMfjWXja0k1X/bhir4oYinYE3MgeArBIo7fZBCDbBQo5TwV9n
1wiBMhbSaVMpnz/fo8s8Eo9aVgaVX9wAxfyHVn9mFaMPkz9qNLAmtdVDxXTkIazP2eWchf6n8E9I
NNbW/Fq6dMV0qXLtOpkZs13O4wm5e2oxGY1JL6FhaUbXw62pny3r97WDc3jnCqy009RloQdsDrO+
+yipLiC8cbGld3qwT/sdDwasAG9mRMIoM1jYHQS2f+DHIx2BNVg7DepVe3PTKENWZAPqfMGDxlVx
vt8sOFM5eStUuzR4xHnl0e6g61R1x6mF7eVG8kYuYfKJZLeMXz+nuOrnWNaDOfGbGqyeQi06EkME
y5AzG6YNe305JoOB0owheCMIPnsKcOLwXNH1t0Asos5G3YBuF6VpSCyjV5Vim/xcN3gsAS+fi06h
NqSLJhnVW5hWyeFm1qDVjreTMzNhKgeIkPlS9pCCqgl6CSxAjGraGUYnj0iawi13hk58J6/nZ0GH
9+eAXPOfSqEuxnfPbOMSNllP/78JN5bv7fgNcimWXW3mz2l84qbMqG+hmi0Bu8fiSzhcZEHa1IA0
22KpYjlaeaVq4VUK2pbmQ3hiSYHL5JbgpZRXv9lGDDytqZC8/DLNg9Kf8w3ll9PudRY1NFm75FKl
4sdBXGR0Ba0vODksmmj79AzNZGSqQ9NK8lMU45kKgi2cY0zDjjBqt0x3KLt02kr7aDUCYV2A3snk
bzn4QC6IOxU9JWa3Uaase0L5U8s42KypnKs4rNHkBB4jBWyXWOBCDitwY46r006K4xw9uYoXr5Gn
n8IF7vlqLkzZYfPmbRAH3+C3x6nWNy5cFuEruetuo0qk6FWoD5Ejz6ZL8CIn0vlEY69jh2fv0O8E
vastntSOxy/KDNgqa4ADd7koz4B1aUi1ejerXEpNcSCqeiirXuJiQkKxOE5nbg8Mwj02mIqZu02O
M5gwkizCylvZrJkhbt7e9m7U/L3zwq7uKdcW37sw8Hzyk3OUXPGRWijV7Vpjnu++bTCrECpjxbA9
lMGdj1OlmiPAR8bNuJzYaCasBoOyXTMai1P7Ko/QEaQ08PE9sIiIB1u1/6tWOdEqmkJspsoZDt7T
WiXdRm1P5osmLfXcAGDQTvW1GVjF29q+vYRopz3xkBHZR7UdiUGx+XQ0vK0zpr27cEcIWT8+KB+e
1pRyHANNTr+vJkFeaC2+xtj1v18WV0UhX/k2EPEz9f48DFzswE04o2zc5utnK2Hhg8/crLTHWwf6
KMrAps3YQUp0yDZJO+TNpLoqU+NkaVBZPTggSmklYe/E/Wlqm6R/O6Ozw29CSM1wuhkjUohv9D4T
g1RM16eOtf/2cYHX/Db2ab1OZ9oS+Hb2AydR4mgOLeJFqVYp5wtWGYqcIc4f1SRNqf+KjPuo5G8G
z6JJNAyd1z1q75j4JpAjf+WNdo/GL2vbxFa5z1tHK+wLfzl6aWegZnmvZzH/Xp0fGEFcVGBUyEQv
Wm9pC4LiX2Zc4XNYYCyhNVhwm/kkJshh9jhfLG4zEdnCBNeZ24rqjLOGWu9MgDr/IrMEZJ/TG7/y
lRrzVkCsIiBGVl06XEiH3WqHaSZsjzTkzQSqLEMkaRZtE9EjdR41VpthgEY6S3ge8Mc/cGBcqiXj
7IJM7wSLIuFT1kQiR21+Gx7dqpm+zy5SmT4sxLJSTdUjK83rxyomC3eoDRbz8imrA+fIqzwpPx86
gbDrf7ukwZCWP8AGHd23jX69iJbXl+gYwdBdcQ8Qn2psej9hur8tKoG6mfLrQjT0ml5vqPaT+QUO
2HzwPirTzGctBeGr/OgPnFuIcIh0b+q6ZuzN6MYm2kJUbucq3Bm/w/Q+fNtLnh14tXSxrlfFg7xc
cGaxc0e1sNmXGPkCAGre6u7EXglu6nM9H8dapACcZREbjhj7EUv2sS+fHf9w7kYU0y4HcH37cAwd
eCgRx+CbpO2WMqJqhW42M2qNDDg7DYmIOwlxp76KgMxUR5xj8VtyXtDYA+rffsNyBNS10poTaleR
eW2Xoi3AHDWoxmC+owJ5WhKQ67VtTnJnpjHiTJX4Tsa6KQKO6UoGQNAkkZDPeAHk2ikWGoo/SPBV
CLJcvHnsjWkLGgKxmSRf9An5rCpIyqIkM1UUhTnIEAenttE5ihHTdpzbAPwD1t5CY9taI7Z7a+W+
u/oN8cYp85iwlk9w2HpEqCMgwrCLbObZfVkOovdeIU9qoJybo3dGELZYES2/sXb0QmtXEwQz2lyn
xeS1XkUsPlayYKZ/b70A9QOOO8YE9O2loBkerAUHXtCYQ4hOrtdekDp90hKhMI0xgkZFiag6Jz4l
WLwugCEc/rO8BDB5H/kpgZhOufCkgJUzDfdKlSlaqtEJrmey3BuU6ZgL+X1A1AYqfeEbXTfp8w2X
GLxiZKitdV2AAee0Sg4dnUF4g827cGMF5C7D6Az38j0YwrK4iE5sxIyqP7q6N8ehTlECOXHABoTr
Yi0j5prWO8gtuys8h5es+uXFfdCwT6SbKWxbL+8H2CbLU2C+IwgVvxs0XqIHbCq6vRYvdCPfC2lw
N8a36gaWHcfStOFoPGzNSRDK85E1axSFcwtdcIq9tjokNN1SMgZwJ7BBfBfuT0NMATld0cXnaWMD
pF6WT7feNDLCBKZ7fRMNZ9Veord/DgNm/oGDwbq5kLKcpO7gXMe35rY0vqackNVaszepQseTffLf
i9Ehb2JDYjVcXheNtfqOwfBprPF8NwLsT2vqcDXNRp+7DU46impvIRxfD6+S0XsZBI/JXyAGIzx9
QEOv4vWvLqdp7vgK64902GkfS0z07zMOp37AKEFP7gj6kfH7ID5p8yLYSTnd1GuuMi4oi1Cpzt0T
Kix/huN0L3WZVXq+YfROkxZY0HM6tgW9HDvNcFpQkq64YwfrImE4P1vc0xgodeHoF4CsnnhSYWcc
GJyEl0S4lCNvV/O3/xaDwIbvt2EiwYyuXspDk85ISBqlwvj/qmj9wWH7FvHQfVFAWKGtRwNastiM
iK9jObjEffs19d4D78o2Nb1wwT9mYs5/kFZz4JVGurfBqCnxS5E+G/HPwkaLeuNWV3PvbplZEoE3
w9v9aJPpOd3m8S1brAIDLBtEd2E1ISMwH5y0gKXUB7rfA0r66fERPYnsSzSU+7Z7GLJykFUyCXWd
ZtWXof1Bn3nkTf+Jtm8DLgdnNroXMvKkOmiXFOSLim4BfGWi35722+4F1VgOVGk5/FCC2GDufmzd
2beMVQXdxy1GaoLeIF99GvPrnaMJaDwWkl/2oPDwbcoPRfHTgXk/JZfHYSAQcY4/vOqZx5yN/6SO
v8JTr+j6Hy27QxUEugsBCZW5gHcQ0f88wtESeyWXYOO/z+7m0SQn8r4+SCSMOwfnTb6MkZvOHKo/
0M6c+JqIA2tXgGyH+bFotQLuY+3sUI4WvTID2uW6eTCfQUE95bt5jPj0nhc7P46uhK8Zv5U5s5VK
ZpP6KD1T3UtmLXm/0iAqployit0PL9+e2WJF8vkmx11jueWATYkPzk+mMSMUF2XHYI/F2egvZmN4
TnAxdhE+N8jTa3Zz+98DXVf0p/tLALAByWe3GBp+iGpYuPYAcXrIlkGnXe6VcJm+ImRJgkmlq4Wv
jf0VdRRGO2/DYqCotYqRGb+PdD9jTVzNIbzH28Q/CXgfqrRQQBLZ6A6ykFKw2HO0izRuI7uSAVeO
GpyUWa+WDah+qIfUZJFxZrigRixhf/l2b+JKRkgMFg5CW/2OjXtQriS8XGdowK/NcTtOGjk950v+
UkAKeONnd87KgsOncIuTIQJtIElcI15hdMCFQwl8mCjH7HaLgTaRWgnG8axjXI1WtoxUFvUCHUCf
mf4/YrOcW3gYYlZ+9dtSKYZpIfd/IiX06K89Xz8SgzuyFc2yq3tXY0c+XuTuJVp1olFMb1IYoMWc
FyN0Qi8gamlcvl6hbsjUmMqezlojBeMQMBhplfStIuunli0py+7j3GAm1e96Si+FNIWO+oXif/0+
1YlQygRGt8zZGFf/URD4SYtTDdIg+8Uo7x6SpRpRjTHHO+Vxb1nwcbgcF++gnqqJKRI2KJut1AnB
66vrHxEJzO6wggUjdLHVN8RjRDGEzuFKdvIQGTUOgeoJUJlLoNf0WnP0JAdKQZ58mk+J8/iXDOQQ
BeL+oVyPD1rkoH6Ki9CpO7jaS4Q+5AR2MHh/MaJYwYGHPniPGu2KgofAEQloIakqT7zvYu/7+2Hs
PRKLGh4PMilO6q1qwRgnDGiYXIWZHDKrBnNe/Xbk1girGEHDxIUL66+m3+J7qAKBkGb0pZqRiUgA
gDzdLV+egOLYvIb8AePVBhSFItDyn/B7EqkypOq2ASk626fmX7JyYPqMVaLAbK42xaxtYgztDdHr
0LqqrBnswsd8GRNBcKHYJoL1ZaqUhnmE05Se2O5PJOYBn9E9hl0kRzGweCWje3S/7rzBHabJgFoo
axIwA66cEYMsXlzH5gJE2Ejm8LWPBpjr7T8Yc9Jpoo3XCkxDuTF4FcKHydihoRysqsArLQHX6zcZ
lnPX/62ol5XWBjSbaYvghZaTvlZ5MUnRVzCyRUlGqXm3P87nbeJg6e0E/N/07f0moMjCb9s8zQS1
hp/kXOx1Ba80IDVl4X9qybXNZBt7jFNNRlOLZtlQ0aLCssx1BHTust7abGn8mT2WO7sHL6pQXp3V
mTBcQPpneHpxm/j54/lwZPLtIAGQwCQOcwvoDV4YWYyBD3Va21w8JQBByQM/jW5dqDAyhzdLgq0V
l+mIVWU2Kre5bS+YZRCHrzri0t67m/efy6qC1nV2yjF0Q3LxrghCPAkiwneNxHwItifwEqc6LDF1
fMKMo0U7e1F+0a99P8ticcI96sEKhe9xWROHpiGrefUTm6anl/DmNXiaNavZx33XZhmeeTPQB9xu
+SA59Hp30Bp6ZrxzB8LMzTI4hcGuepo1wn7gM8N+VpZW68pfkXA15+3smWSfP+GUfVNt1zhkYUPo
9242YA1XRyJQnf0od0Jq5Nsm+RwlXKzCVSGYtDKcTdFRjiONQjZpnm2vPayikRV+xP8syZ0e8TZN
t1mxQf9OPl0ZIF+rrJ5C8Sn1NAnf3hQ0Sz2/oSGtbxjT0oL4goQgJJoZ84vh8mToQwF18TBtH6GN
gM9k1SQUY9b76y69txdIP1En4ILLoOG3lkgOCdzUjxa99Xw4L+OE8cGpt5RI78h1lN2FDwj1lLos
Ndrvi3DJMQSYgTuksE9lazxKT8gYdT8qzxl1zfYqJRvbaIpHgIMNKcODvt3aH5Qliepn5qekD8XT
+Nz/p3a7WZj3c4He6P76lPfDabEw/Slrn9H8mOsca+pAo6drD0j4D33l7HCxDEL7C/4MXtk1q0d+
L/N7GIy/MqAQ8H/aPhf1OLl1js8iVeHFGQSvWMkb0H1kAvL9UnyYzX0UxQyqp4vQX4wIIuRegqpD
36hLcP/JsUY09j6bOkGiVTWBRB+H7k8HMJEYYzCwTX2zSuPRpf3DMAMjyZq48YLGV19zaERvJF9O
27mm6vecmsHW2sl3XhxTUPkIj/uskWg2R3UL8qK5kHtej4tvlnx3XPrWK3sd9TreY0GI6b5j5DIM
4XOkRNcznMLksDHusftm5zEAofqL/QE3+OlNt47twv64yjQU4AQxH4nr7yDv9Fh489Jd6G1dVi1f
6EafxezYnoxVK/Q0NYo/2Yse0PyKHSTdD/uVQuTeTNgEz3WnUOxkkc3yi1PweDWl76VJ7/7GbFNS
LYFfNJrflMB6psm7k7Wmxb8ZXHdCbiVouf+jgFZOuZLKklyfAfMDiUKA18LRt39DaqorKep6dHQj
ie/Vta01cLhJuEGZZPLYVXEpDDS1UsPgnPnVcJFBcXIGTf59Nu3NIZKHjJau3pCF2aahO0ujLEUp
subbk9qni/XY9WcNb1SayeGInhu+iJsov6cWSCPMR5WjQ2WStfuYEZz/gWkmo7kaTsQmjdJFsnpB
DsDvlywhsrGcTQp+7weOdZAL4u0MhQPxaABH7nrkNtWiYebaZdEMrP+in1CxBriWwfZmSaa8hLf/
Msqjeaq4Ja1uxRxkT2kpUiuIwGOvtndUXk/qytxr8NY7PPGjb1822XQWqyhm6BJ8ZscrVFgIYmQn
LCY7zcAKRHL4JIvLiAjyQjHaMr6sqvxjuoIk46WTzkjX3mjFBxcddHvNcQNJgSInIIpjF4HM3r0f
f1uzwy2l1suSrjcAOU9JATijCBmhguo9IMATc05tK3a6FelMkXOo7MFIuLbiZu9meZdMTDxhan+m
jmPdL/qgpgb9vuLsalimKJC251J/vY8gLorv1QLTLnnzx78m1nw8ROmOM/0NoLoL42dDAVJa1X7C
yd1KPFMOK6rmSlUdQiWZhzivHCNMTNeNmkDyCshfyd0lhTiebVg/if0LZJeK/WuZgynq74nM4uqb
guuSWU47OwenrKiCAfKEyuKfci/peAKLUPYuy6J6vuoavFOLKlMnY+T7VM6DUyzwy7gTzZNeiVEL
PE3tLPMNLinUUPMcWYQ7Mk/23Dv+Jr+AOl4HCy6b87BXBIbLpwKI4QK19sBmUwYtrLR5gLF0YeHQ
VqYJJAjHHPO5Tcqey3lPhudDTViobLCGZww+5e6yepJCVpMztQwybITo3eiTlq20Q6XqTyg+b1JY
wXqUKtKmN+bUWrVL4HEiXG1guwjzKN0i24JJtAi9DaQ0/e7E2egSBUuLWxq+49FueYOckKouqsbn
H+y6lizQ6YtvLOvnOKlBYE5B+UltIuShpmY8SgzjUjvnQAKYceKTBaarN+eWDqIGz2mCQbwN/+Bn
jHMueMvXPppvG4l4RizD9nwuNHdy8uY9fljsplu7t+H2a9+btBPmZV9gNonBPzBHVNfJu8ImBryH
kjM7qooEq9curmGhGZXsH1qijcTGN+XknWfP337+lD0sSD5sVcxVakdI9elhfbVcu1TTFtJfRVe4
W7UucBcIOxQjHfsv49dzAT7wlwVL/uRak7YTZCVbNUa01uRv8ggY78c0Akp5cVy8S+O7+YxpPEnj
0HtRst1DAz0Ewn0K5BDO0DsJJ2p6i7Hr3jdWfbmBMOlAJBmO5Na2HvQKVLNlD0m+B223057muuOJ
jUAd5kboreF5sfd2KBGlcgKomZ0cAL5G4VuDUfn4ISzIVoEdZiLbPdKFxnpbb99gKCByvUvFMFPO
0DrSyYRF/vAO5FC+MFOfAH+Uj7IlPKVwlFaUevsvQ+zWxW6EyOOqPCYbZSf9+C50IxIbPHHIcyim
08s7q4iYvULPkWQvds/D2KotoFNPSdNF6GbwhaoOGO2k6/LoxIETQF1TUJRLmq+u9dAgmJxO7h3/
KWRaPQ1VoqySFXLgChJ1rNRSXcnhPTHlXMjmu2EIe3V7Rs3Rwp5w6opkD38jrE0JbtM+JBjpQic8
zYrlHdPQorkMkdDotjd+azAfvVVWLdbmo+dTCWYutlDiGEOxwaHyZeiCIf6P1E8Wqmhk1CNEUTd/
7UA342JU0FQVE0V4BA0AXj1IhGc9HGZStQ7Z25aJWPqVzWzJsjAPHhrWQuDfQnvOauUAmbbuOI/S
8JSvuTpsMBfq2mWWwbqZ3jGNTUyw5dw2o+0irPCAvIrK05pjgay8yxZAoJxYVQP1v57tloJnP/il
wb5wLuHh/VlDd1rlPmosbNhoAF/IGEgawYDJ7MwcY0Pco2zeAn5I1SZ5f2JvNBpUq4ruNJsWCA70
DDVAy6qTP9WjvcKmlX181iWxU7oPWmbun3mDI1JA3vrQi4XXkcF5o/1zpJFZuPiu61LHX0aMQQsS
1H1TUliiNcpLW+N35GBxMgjeb1e9Sx6O3iGUSaXp/MQL2nUvc/5Qtett+ebbP97vexG+EzRkHbJq
SZDF8ZR8x4vUgrz1BpZuG/vZLox7OBenyf8Oooowpymj8yipHezSiY5DbBwS22Rg6H4m/gZYNpRp
/MCv7tUynDUwsb58DkkdS2rQtFURi2Cw1RKj5jEMokLhu4hwuSJIgifInz0hRBwhycNB4VZvJBV5
5V6gRyu3EsRztz0iWkvoNC8TIc7hcQB1Ifupq71SMBjGV5LGbKjvCx4inKTuj/ZoexXoYfpRSClj
kFfEQjupjXKXKP+oLTwy1L9Ap3gJlwptcYPtH/HIK4CTmDV8FgbxxpcC/zuzx4nhklmYZ+LE1lAU
ElXoBJ5iBjki/cZ5ZNuXpiS9tJVuFm3A59uXJidDLt/iR7/KeBXWF0GpPUTJveeojNQznKgOnd5N
xGQRkEeActILH+h61phvYLLlJ6apir6hGnlsVE918g6Vy537LAwUwopVsPen8hYco2RHjbMAe9KO
9HURxGOccgDvqVdIsInM3ZwONDrBjsgSHlPr6W+Eo3Ih7anTpzLmhdrQaYMRb2kgovRORrnSaI/j
auT/Rrfa5LSsPExLwzOm162nfFIslYcId+LG271dB+ZU83ozwTwKhedAmz5VZugSc1WrpNxM3U30
Vn2WfqVyP94sX2jlkh1O00g0ao6jw5vsNoIpitBWAhfONzl0MSgeOWtHbS+IBo57cNLnVhhF5xSD
6NsDJz0YY5anvDq0Kx9I3trpejTmQjucQU/CGhjN+oPVoskYG3F0L0EgMFEeRfPbud36XSoyiEnJ
+ia6IGZMOgyr8JEO87axSgNZfLus0HSxFvnkwlAGQWgaYJFQnIX7CcUPTJmTZWknuGLP8+h/XnT5
bPoItKfDUD+ILzGBEHItWD0/KG1B/Hcje9H/vDk9iWnQSMYElppe2R4J/IVLM3ZFSlCp++uaiJV7
SmN1aTni0cAxWG211ZQ2KVq57XUfh12xwGbYTweA+yk+LkBHOgjFgUhR5tx+le8FdWJBS+TIpwAi
cCue3t9SwVehs77/0AOZi7SQ3b49m36BBXXVtalYA5FWfk4NyhcJVmZACm29rJsFnv/iA8jDtkGP
YW8HPzYQvVzw+SENA6rTqkyf+YLh9Wr1mrgZermWbJsyIPaFDjYbVkyeqdtH65UBlqBK/xwQ6rux
4sWpd8PULHzPDhtpehlDP7Nq/FE0xDyYIW3LAfc7sAk+P7wy146X/sN4wLkhyIFn4cBsj7ZsnFPt
lMcA2VHDSTAKshH/cKlEQFW6Yg3hLBPsle9n8yzvYLSE/wqErmoQLtX/CCkFWVkhmZ1XcFgyeWbF
8oGgbqUZ7Xd0fKlrrpXih7aeD2Ip7d6b1QpNvHYOmyd7VY6Dx9cNUZF8zFDg/KPKZeVnY/Kvc+if
3Rag8B+qAXUhiL+5CkbaL4KBe/z5c93LBy+fELr1oVi0zapbKNgbUUc63opRQMN4EFgey8isClw9
KbTQfq74VXaTmXZoDCzvHEEqN8qL2JFwfPH/1f7vpE894CNzeEF6bRF9lzAz+5838kw4VrPCDjKW
lJ1PJ/nBcZIB42Sq+XPyvnhqW0rTdJw4QoExPn90O644NfX1QTt75JXTcdfjUHvdxVdsHRTIV5Sf
/oXSv+60Yb6qv8CFC3QT0no70ekIOcGKOG1VNh4LPNSNdquXjmuyBFOSOuXcW6zh2xJh5ll0B73h
3J6DUCb59aPq1ciEVDvRxbqJUstDv/5vVGtCPzqap+FFnNC6ZVoCH+AXnfxCJukIoWg+/q5xx+Q8
+gLMvC4A+dnWWqnCBK6BcVHYO7k3cuVaRfrnmi2dtXnUGtibUExyC1gTEvP8AIdAQEdKNtM22g5i
xHEO2OR3CHXi4FGq8fFCrVkw19SHC3vfYb+8E067wQYn020fSpbXhdfo/Ft23ya/YaHaHeRZL3AD
JTrgS21O2dutd+MsJ0il41S6zyWRh29XROE1QhZSpZnOkqi2NzLXvrHfgw5jhmcMwn9AO+kB9l5s
cHiqEO+iIapbMT0dWuD3vzuRX6WF2ESNtb3j/przbjelJhKay/B/qXEIz7cHkz/EVfHz6g5wx+pN
mtAOJcf7Eky1PFfS9nol15LIsTjCjESElZt0hGYR3EK3av3tKNuhpkQcJ28KcH9tDofKndW/y8zz
wIvlqaiOcfR+R2xIjUn1ACiy/RaxYptl1SA1MB9MxOsYSPAZtkmcSBtACmImzMd4FspLFyewdjAo
ocowyCultsaASAv5nU70dKTgXpdWPXm97QM3gatFwWkK7kcsK6ORPYL7cpdwEL3VLgAujwYuwsrW
cz3SlJ3TREhCq2AyIRxEMShlpn9QDP6dtEfXM5fNJyQfZE2kTfo06RaGVyx13xFcTIYSvjQ9VVpL
1w9EhF+icLX+eWx5rfzbqGau8maRAEYz72IAzAhFFjhRGNqgweZxX/eGlXuA5sCr6tFcRIszBG9B
AAepNe8jxdV+C8b2w3+CpTRX5Usz3EBnd4TlbI+2Ei4/AsRqEVG2Lt7tR6Bl1xxarylPRLBED3+i
Q7TNlNNoDTl//cKnJkkT4iLLIV/lbvWdfJknn/RuaSASndKG0NM3aLCJ0FkcY4AuED/d4GaEDigS
yBkVBu4PmzLDDGuByIU1il32EyMCu4wDDoNUpwp7mauN1EAiToqpSFHGzXKgDW8VbjZomjthjj1D
Q0emrTt+BZBVUm/SFweLDe+Bxgz5WVpxnCpdiB39YMjzu8UOa1NjhzSS0a+XotclEnc8RHR/KtUS
mTgrSZJRKOK6iuXpOuuNixutwY2EVkT8lHB4rUmjvclikjY+0XmikVtJOy2nH/nOQCHZ6Z+J8cOo
gwBxRQ+hEz6F6TSvIweJBh+nxY84HNUBIHqudPHeKb+1fKUntleG4w1CkqLMtRrMSsjzHLVdxaYN
PfDiaZpdTYO9CZO4ZwfBnbRCukklQRY5eb1Z9ut1bHw2cvkQtXHANEw7hk6qn8H32+YSKcljRQ3C
BLP5XqfmRfDGorWO+dtPMwpund+pu1qmvDlFi73utKj4AfdT43mgOvzoumpGKhKVdyaGa5aN3xTP
gqqE1joYdm0KJfiTbYa66M4fBCOOEn9Vo2yMdTcm/5Ok1dBKCMu75TgKKBKoYMdPUCZDzo06XsvE
cP0dwMFa3gqdHyjRbnYoLYBhdATgQSgKLl1Jg/sugyZdoPerop1hTWnz7WAxmNk/ABw6fv4CDXQd
5cvWiNRBqtZPjnyfv4eiN2ybAzXBCbNFHESWzlQ1vAEv8udIzRX6VwtXkG6S8ienLfPSkgefOKA9
rksx1tXT0VMcq6WCS3P5mJDNZU8HDq5CdQDww94GG8WbL/BhHlwJyGtf7v4oPosOiv+thhW46m38
3GMO1oH2fH1hIY44LGmjT40NlozAkzeGywd1olyw2paWs3C/bSrKyPYY1WuwVQZJtLd/Z4qpCtsd
l7gaW1wazoB6a8ZRniPVHIn5dWw6Ov5ZLdOiyBzyay4hknEXjcfcWEFsjepONEF+IzgVywWevzU+
QBy4vepASzzm7MiQqCVkXOlqTjMmcdyMjPuRzeOnjMcoI1FBPxzhz5gC6EAv+KtmvUS+W7Hy+ZJ5
HYeXldL/n0TQZKrbEV1qFmuIRaof7jzCc3MJZaqTe4LNq0NmvKkQcT0BBkZAWF7pCWzm/1DyZWKC
xicXSeENtjU6hvAZsNIM+whRL/VHKpjwF8OIhtJW3pQYby6wcIzb/Hzn5Bf9A50YX9j5bJ0W+0rQ
Fu5isgtmypTikfojOuVvDSeSxpnZo71T6xiEEQ/DDL5xhEjq9AsfjXTfUtxQb1YLwEYaxOIholtD
3AGxigyCxaKowvdSkFCtGZbRpbJPjBGkKNGtaKYSP00P4XCbF6P2Z/QJf9Sli+3bKJ4OPrM67iQN
xNJvRTXq8Gv++wjTlmAb+85xVvv44PTQJPMzbSxFyHXAIs8HQ5ItpWEzi44AkEG1rxerLORKIjVB
4eAnvZ5xEn+tdZq6O50t+danEwxwvQq13AyYGf+LTjgehg3dAWwypdMJox9cicCsS6Pl4k234sZD
K6VrnwQhktwgkCIAax41SzT2OEbaJ5zcUNg2M/j1hGfRQEzleM3yESU/Gz8wFs2qkCGHq4RFUPth
QAGfGhi8kiUUJ6Hd969bpXFuCy7PGCl98sOgBy9AYklAkzu1Ute+o3Yk2w1iOnMj/dYQgFbK1+XW
MC8vUyA5heMjsJLQ5DkXw7Bdzc8FGlgymlZiQeMN/ePODfSqzZyPlKk496BWmKrDKOrzlR9gy8F3
EjmoXoaUzOl0myj1WyHJJHxk0epvb2xXnDycF3H+9DrIuR07fbM5M3wxuesddGGi0Y9DvpvCIGrP
k4r/6QgffNnoqCKGi1xSnv5dcfGO0GxIB7jRxuacSv0/xn6oq6QwYcCFRxwS+UoOMyRkRqE+MyYr
gmu8RUV7u3onHnDCF1Ch67RMb1L/nN+dzLhb77ebnxow01/Dp6aeCrbJFzYCpcuUaicr8XTGMjmE
jFTuhcuBzsFEtbBk5VLaYqSZxFODoWT+4CBvXcov0uvyAxTHoLvaBIVJ0Cq2uQSIYGIwV/7PANzs
b0nTyN7M30VL8oFwvDsU2IuAOswP11PApzb42sxHvtJ81zBPhJudAg3F1XOWQbN5nxeLT4gkG81z
tMaQhRdRPj+HvcfAA6y3dDaWELHAmhICoSye+Aofv1/EjprcT4hQUOffbFnZc1BkRlHB5gb0KPfH
0JWb4DfsWV3bFqFF+kL3Zs5Jb0E7tmYeQm8gAIFSzF3AYgzwrv7NKN1iH/TChFBoK5av5InAdToY
iZVtBlBBrr3rs2QI1QxpNAuOXw7m0GuESqkv23UDvTUKQLYztHA3oNBDwLhLMK+jFSB1Dhmrfae6
ZPrbWoN3p9iZqPnuyNgHRnNI9PaMMNq7TTLr1ySNJEu15ITelCavxOH0Rt3/4OeMgvP4I2JxrYzN
JEs/DbCa3dZuEmDcmXH4t7X3NQeGBmO+Ykk3jYPt4tvBnDUZ1yLl9aeCXm5PudjlULDr+J/UQwB5
fInsneuwOGQRqTOTKnkJwukyT7+y8AjAip0vjoT26JJbDH9uvgF2Oh7y1j8PeIymXvlSgjs0Q5sQ
6HCOv92j1/+rt1TeSwNZNNE47IycExL8CrPON1WehNrOOvmJtoZ5aZfr8n8HRGcxeO20K4g3RWOI
FRYODvAXXEwObz1hgrzldAUEspD8zReq0EHkup9hkxBOk2qGDnRQPGWZI2mKwCTCzrqYcE3gFsnv
VxJS0xsarhTFnSf4E58wdR1yoBIEDVY7zo/8ldeZagtnRYa3Re9noEmMcCWym+Rc+RWc4DFR1tBm
DUykEhkfCLezPuO62CTvFhbkinbjUP1sCt5PvMG/ARZ+wgWn6k8Bz56oo7GJjrGz/Bjfsr8m+dEX
pqf3FaSUrOgbJb2zzXf7cF+v9L+aAmtXn1AQBpArwiJEcDypSWRXg3MeZlaGKDfkzdOuZEyjuToV
jjbkC77FV2Kyp6G13rFGOuSFejUjPPHZgrObUQSFiOnyxQiXwkHfTQCLLtFIsKeDf01ZGsMtsW1C
QiXIW8xNr20p5DFh96MQYJ1NcI1wXJxHi485NczHzBXwWpxuvAfIia/ghlEn/t45508MA3tPjRVe
UqL8j6ZJwwsaVHWKC8/eFx8tVN1fCAXDoQgiFvnX/2mItkRDUq7S04UEF2WQ4SmSccv55QWMIgCR
wI6HxHp7vx33Z3koypjCJ6pSbKBL62/UptpjSDPIVLQUURarjoa/2djdFGVQx6enPBlv2wub9DRR
ofwgRwPd1KKDGu+aDZbtjfTTbDc8Sydhud8HRVL0guc1acF1lGmWvSYUzYPtv2cx3Lnf+fkZogBS
eYzFUhK+80414TJCSw6Vm0Ji0pzuyRiQ5veP/rUli64NJCBv4pMk3VqElKeTX6YBwYn02/5mLGXx
CVmn0sgZEPVKcCXW+3jHbdtnAYAHLBcKCOdK1ns7CCNjac9EbPKawdcvWAvnby4kMkk+bDlpc2u0
GNmQHYrJruPYgTxKV/jE67aVizcMggjlXV/LtGP+deb8fWmg6yN4huK7y1fTT6RmlN0fByzexA+7
S/EsCHgCPV4zGh6dr0tHGnrfZhalMfB1HCKMl42+QvBaODVwETfbdiqFhKnATT42Qh117/OdxyP5
wxp3ltJv/Cq6DAMl8UTPJbBpgc3p4e3/vswsA4FjqpjvrJdkBj2IWW4sMpLLfKtgQ//dQWt3XuIM
grbXRJpGUi2qyKeVsN7900jLNwz5ThbMVkbvmFOQXiTeX7UcbEJ3hdHljPjSTLDLyIAYb0tBiGgi
Xx2wzRAOs982pStNTZnxQp95Z5tPg8KmWeKSvrup8QcnXtU0xkCOZYnKxrlK6WKK7S61W57k2FL5
G1pAtDwRKBUYOzVi4WcUoNmaKsZzZcYe0/ISSYPo2lnciNIkI94oUYIULw2YFmoKZfHllLfRKXCe
Fuk5jaNY+bX03cSGgjgioxSznTt0lvxsyWf0VPqX4D942qk8HNWHbJHEueYrJidKDMNznwVpNILx
SidbPnb6A8NrOAKg3Y/FFmUECTtRzk+Ca08I/pVhbUl4m9wnH+NohfKu5n8+egGf27incPh0cGJU
5dG8zAhzfIMa1f+zbkl+/SYEYseQeAMWUFNjjMRd6JnHf9/4ar1cC+hUZ5s51ruX+H0xFvkU3L6c
1oR2gcRIG/Rv00xhihlO8lBaxUd99PlwTXBCbgB5uev0mH3YpTsc4IAMyJUgGfCCnjTMiH1WLtHz
eh3eekXYJiEqEjrlk2HJF3N3/1X0eGscC5zgj44n2OtvkGYg4ktoTM4TUST9Z9Je1ZxaIetrm28a
p4zH4N233hFErBZzmQgnT2PVesA7qFj/ki7KYsRseXmxv5739R82JEHme86X0WL1+mUZCh07PzXY
NHzleMb53ZNh6GlKlmSqJawUPssOC/hywl1+UwzsD57o8n+YIgH4yKLnZlmCuTr9jcspYRPkFtKW
U2VNtNLzJCci5yl3CYuyVbP1yomVh/pUxuiMmnl6STcX0q1eQbMIknTffq0VkXyBIvlXDPIfbRj9
YQMHB2I6vKIgzhF2PhfAIrn+IdNtTs1FFmJ3NvafxbaDgIowPSWjQVpZEoL2JHTq4T8/0GGn2/OP
rHQVcGasC+GUuAfW9eYRl3m1QJ5fdhnOP6Sx+RvvCFjhIclgb7cR4e+jY9Pal8r6nfnn+MbsbFhr
k55U8vhg63HFhdy6jS9VAF5A8GzQIxOZ08d3TLILQA04oGd1/SadYf59WaTdIwucjhZShC2yNjXJ
QpdI17J+ye9PL4gqhH2cBprI54Pk1WWlZg8GWj2CCkGtXAf6nEpOxTV1CbToQ7SZZafmFcUNwD8K
8Q5reLKVUyiM4EsXJwiVkqngNRdTkpcUi9cja7TojNJScGqN+v7jTI9YRjpHiO4BWNdmTpgk8ND9
Sv4fzMasRbptWYG6ew/ABwZQyPvqRj39hGO4guBXBMOHgD1fwvjT25aALCfl5bJaxC6SkKcoekAS
O7jkMxDpdh/ki4nHq/iTMRjPoIGa6LG2IjinVhowtjewn9mJPOgr5QZ7r+kRty9EkTnFkFM30JC4
vwBXzRTVa2sC7gCxNi+H3ssSTpyfChAms5XDjc33MvlvqdKm1O2C/kwCV9LZnOpG2f9zQ0H3kklO
CrdKgoCuZevjX5vZD2cyAKp1cks08jFFCZyZJQDWjPzMyLP1LQ/LNYgfQt6VfItxkhevhqmVEZRq
EVfdlU09xsn7r0Ki4vSRO6Fo2RbXLLoMSJjb3dnRIr9fgSLG+VMPltUsMU0tnkgSImzs3nFHOx50
xa/HSwycWnNoRIrdZp4xO0WdV4Xcdd5W9Vt7Df7gK9Bled/u9AzuoXvkEd7kxjt/S/HVfQ3rKfz/
H8JfDko5kENLp6n6/rUbdnge4w/Y1FRqbfVd2o9p+ltU9TQYI5RSI/ox9UA+7ke57O9l/fCxJRh7
/501TJ3YNldtRNUREcl7x9LMlI9L2nO6gh7F4iixPC2eWuWM3rPNGXGXzxeh3aieNPqSkeXADsQm
wurhrIPt4g7nOmeqKE/nErzebCRVhf/iHWYOybYGm2g7EXsAd0BFdnhFQFAYQqXEehmKd/9eYmey
jKtFb4sK8P6kR+DYq+jPaFcF2YCfA6a2HC64rMWJTp7fKF20jxNiyYU6vPjTDXgUnz9hRvbfho/d
dUil5Twody3bpotJ9xURMGVDiM5fgfU4ctWS+yjwWksBe5dd1hm1IYYoiU4wHFISvDlJKLeDM02Z
IO/KL3xGNll9iJZL1tjtR2IKgoJPcySWJxbHsdbBr0Y6N9ffGS0w87hhm7ZmW8eosqoXlveEgvvm
gFe/WCnBs/ZnlHwcaMbn0hTEkH8TONOSUbe0lNUMkzDzOMDVOck/IBzHtD06DrmSq1o7oNygIY3k
DmKj+S1RZ2Ybw+FQO/TYM4ifCwNnDKVSJcD714EYbdJ9gR/COYzj1r73hb0jwZ+x4eWtKcgzhBhn
22ensWa7YJTV26V4L95P6wOhsfZVefFNMZ4guSSuGEXqHkXVuNIhz7hTn4mumcQoUP736rxLB0Ai
+BJy4ZUg5hR0dGD4M9hBv3itOA07ahVbTRwV8hzv5ziY+TTH89g+gwP/Y1rzweTBfKUrnVBuxFLv
3+qrM1h5XUiDT3YWfcXE1b3ClPGxlhsoZw7hCABxiJgX5nn6PJoM9THazePU5igtPr5wJEsPrb1E
Cv4S/zDy9MWF3Dl6kuwZlMAdtq+GfgcM0AOKVJHLVW/2L9Tcno9TImE2MBAzyuWU8FJ1JEPtNL5x
C2R1R0lkc8qpYgVXKLvtxR1lWR9ZRbpYpD2w3A5/rmxZjDphjmypkejG8G2ESHeetr2HJs9L6hRf
iCPUeliM2TpwN+CflT5ssX/MKvU7DxbTm0jjPrZxlHKqVCB1sRRJePQkDho82Slq/dPIs9e3ajny
Twj3nTa3fxfhQCFMbA7pfq9hm/AAIAkU9eUjqk8GcIJVAVOb3PxasX+ZtTExS3ygYUWsWBt/dUI0
GSOg674qLRUxEgzFQqIFBl56DSGATAqX892fErOjbBK2nCal3ySX+TqGpMFM5Z5/TL21TPTwU3VF
q/NVOWs4jQCJqrnXAiTB3UXH9Wcrx77V7ZXJJA7toeEYWuv7xWV/QaQ48PUr2bfTnbs1GY1X0yhJ
pyBUN8CyJln8qQNQdMso4JTvb88nh5GogsYsf2OWroG2srWu4fqDNuJWk1ijSvtjbN2tNBIvS0bK
DQ9QpYy2dSTtmlm0fc0Ikbzvnbl6ICJJAslRHQTVDq1d92yGQx86YVu1UEgDfot6U1QmGL66RJW2
tccPuk4xSip3zpOMoQIEvrRozPiBvTe7SnrD6zy/MO+4sLnHZcAM5ql17G9fwA6hGx3LM8txI0Nx
LvCE0ylT8IJjAw/vK1OZ6V5AAfqbekRuWYBjlqLn7+wiQ62edc34ZwvnjmGjrsTjOC9eP8AUhqdj
A6UC64R9lEMzPAysatWUvHwI90jvmU2MW4H56TCn0Aun0BAZpbosk6AqXWfMCz9Yzzn5c6k5kCFN
FYnVg2w9nAoBLfnmD6WmYx/QdHcveFZflMUf9/44zl8SE9jZO1PZv0e6XC1IHP+FH9X90QIqpAf8
7U67+a50gERDiZHXbcArTkmMLc1tZhDpRzV5vsA/Ht8ICHqEN9k3UZ6doxDt9qfOXtOOeTYmkqEX
3acUCYDUCq9SSQOnP0XfL9emr/T7FHaOjKcFfYZuFMZY+/RLsdrCbdJKKggv16QJfjOuHrI+8bfS
HPypeeBisjnmZpceyoIq66E0hv+1V3j01D5zfdgkK0NdKI67HIuG8juqpj//bHkhH64QQDS8VzN0
lwTH6jHDVkIrbfGR7joH+18MM2ZxlKCw9L7oW+rv0Gwd+jxyr11zQnmQNuR1YeIOLZcT8ji60gjv
7PrfPRwtFklGQfipbKXI29vAOZ2S99nsrn7iX36BCE92Z7eydcA+UazN9cvJLjyrqy6tDCqyAsgy
23cO7t+EKvLotLtbSUkQlcN1Y8ZhH/PcRiYjCKSuvZ0jRpyXPcV8E01Wg+fQler7pdrgEfQceeqq
/249Wq+I6QhZR3BUsvB53zx3hiXSLI2pSu00h4g4b8zFHJt2OmeO+nBjdWY7f6p/gUwGkv9oPTlp
o8yHdXKWqDN2jDShNCNsJbkUdfAxTqcp5CJ6J8s2GtcvTxBDCv+idCol396JqmAvJVVrGlQLi74F
JM/TFKAVlLFRCnoNlzuQr0fZglBvLdzYTjV0yUXLGuncC7Tj4/XYOz+stZ8Ppiav2/SON02cD2A9
1H/8p+rKoID1h/dRAAGiensxsOqfg3lx+EHf4LLWdaJFJsHitNbur+HD65u3v69yjBF6ABosGx9o
GSKPPyH1YoSvyHoGJFegh8lA+bt6/aDM6XBLFWfriaoRfrThRo8pW000JFO3gdXJG+teTrMcE3xC
5/VliN472YWq3CvQoeTASjqzJDuFg7u8urZOw66Perm4iyhuurtYZs6kpJ3J2xHmzD+/487U63X8
cuF18jmYIOjgHYAv0AX1H4kXfZVjHtpSInQE5C45VNyItqEuTsrQodYJ5/4rdcSH6FTVqWWl9QZE
jjV+U42dMFTmrXRmXdyR8lipNLWZGzuCP9JUUIxVy4wac8wfZH2QsPmAZuSA8zvLfjIr0CefvlCO
a0Xw1mzCL7E33rOB/JSwhsK9XtJtKIJDuCAZQEvrX54twe4BSiYZZWvGTg6boM5joK+LQ/AT6PFZ
W4wSC9Lnxyd95C4Fe3wGYyRptxWTrEF+X3PiULdUWe+eFSJSEjsd972yUZ0mivxzm92paCb8Z1cj
45tIQheVZ+jM19wKTIgnwfc9d6L/yZQP3EMUoDGsYfHszwMWLDge02BBFCXXkAQULoaGnOHdnPhb
a7l3e2E65fATM6fT0JLfJ9jumLvqFIy930A/YEuuq+0boVOVsu2XZbRCAKSLmvf8lavTbkhzeHUU
bdy8lc0sGC/5sSi4hBw1mYInX49FZqYYF0rd0eex6a77PG5f1WlFpP4Nx6UV8h1dvDX8Hdm3o4Lq
gnFcrfa3SwThV9ECY1F8+kcV4iMi+5/NX9wqhHgChKcCApFp77BilpbcoWmaG4Kkf3iYbZ2o9kpA
EoO1WgecSeDtFgg4hm9AIkXQ/Um0qVg51rWjM8qdovu1oq4u5Adt05owVvMXJw7s25tfg+bXc2TF
88dnfgwQCXRWUfpd1kFyKYB4gl07dQJrj3oA9HQdC6Yj862rXpvLyYLFxbo06i1SsWeIAjiv2ljI
aVYUvZE1MNBE4Zpr6Va0MwhHF4Qtq1Hkq9gTIUFq8+nDElvEhf/lLn9YWICdUoaTmhggl4SCInNY
Cz09ydh6lQsVZtNBT059w7KRLcHIJg9OTcZ2Ih0mYF/QhCJ3TwakVf2Pnuc1+jNHqY/nyd9CBrnj
9P77HohyXISZ0utLBkJxnUoPBju18bVEwxoJRWvSowah9juJ9ixFyXxQZ90gck5B7mJwjzkVsSk8
sKQB7ENniE74ZuSw617WNSCDmggC3swJpmmbmucJMQCdRUf4G8MSeIFZx++J3a5JxNltWQeeY1pb
bqEcNgwuX9/BcY6tvsoi81TNxs/lJPhDosZ69XTOvCLQHmR3yHLYUtGafG+kYX/xqPpK4FgszEtm
xzlBvUpytzbtWnVE0vI8IlJ+G6R70IPSDO7ItywQ9NrTTGWkNtbsmewV00VcQ5/tkYimVVWJXVJ+
1GstoEr0tKBQ38gXjPAfuaXRCp8WaNJTDfW9dt9UiFr0mN6sInHUPJ+yXM3rUVcmbiAlr4MqyhKD
/QCWf2lGgNLeUB7er88smXjLTQAFxTw8x8eW4fU9ykKsoN8d+3FcyDo1xqIlSwP1nv4l5P62l+zL
HAfUNqwDyjomjt61SjlJmbf8w1XZysmN6eR7cZi9Mt+EJ34wkqgtkIuvj2JBBkbW3hio/3NwfaaA
VA10uHPbCyl0ZKYpQcLlu68rnZm9BFFkxm4Y1eW7Crq2hKMIDjRTsq+f0MyDu4BRPW+sYueE4+EN
xwKNTChupW6Stwp5ISN6z1zXzDGQVkm2ZiukApugBdWTqu7UTdZpRavAus1bKSfl1mD3Gph52jpO
BDIiWyKobHHk+KzedfvnbssxmEuOs9Th67oqHZXyklPImEbW0bEx/0O0NKW5Py78K/c8EgDIEo/N
Fgjv5eGTWByKnTxcdIcI1W01r24mOR0ZoVzMdiHkFwWKmiONXT4MjLFjTBA00LX0Yamp2+19ZvvI
J94yZcFX7LaxkeUHjhNCgk9tMEwvrKyYAgq+etsnW0VKbFBOwCihZcxBdFFtbCimT+Nl68IzZJ1E
iMBlb8oVTol54Ae4SnrstEpYosvGknitqc4W25NaTTFoGkdzWlNUTbT2Gf0LaFxj8pBoYsraTL1h
PWwhVyJ7zNCICA71fHdZ+xaiEnPKFCBvkMzdEhzpBa6IV5oU946jOBkrQCy5eZ3xcw7Yu0ufnHF9
F4CsA+sONThxlX4vhSad86t+gDyhUHwinyQDH7cgSrrEH/xW3VQK8JHuIJ4vrwYIxmsvtBELAd7v
RnkbYfRmQYDTs/FLLW0b6ZsZlEhXKbzPr6xhkDEAQiLtnP1QSInXBqv4edMgIu7G5S0itazom12L
njT1JhKKrJ+ON1QGh/ZH53+aiZRfmNvOGtvBgSiPOcuZQ66GZXPuyo0iIt8WAIbMl8vynjIa32rp
bRVddfXPKqRQM1LTPnZLzbrq6hUejFBJ/FE35TfA6RiOb/40B+yvv2OWU5wkviQI5Du9IFNAXOep
NbMSHL9j+CwgV1ojjuXjdSKIQguWub0SiiRNP2bbrLFj1YVBs6v2eB09CMKEjOMtB4wZz7hjUAR5
W+ZWKO6NT7MvE5me7ff0ijck2f4rNHmFGeB7jgCIYFOZJk7jecD3xgTmJmMKHBVCmXIGmuclRK/M
S/FE6OO+HAMwLNJH8tN0hvN1bd3WgzVZ6/2P/ofDRzYaoFT6RAtMMl2p9YSs7swqwTPSPqhYWXf0
H3LwClBMhiHn8N5h9fIvZpkWNubVFvN0mFUlIGJkzcsgnDim9UdbEI3t5YCDDPsxAOb1iLbltQ+l
/e3fsdeXO2pfUt6r3Pfp9nYm3ZtDOpCyqTeS9sop1ylQCR+mJYzgmrNzFh5oWKWPLD4pIJKo8fij
BtVrhh7O5BKNpeKovCap7VZgG+pP5KUceMbZVI+nEcZmPrKR3arPU74oFjfKeWxhfVq4vLUx6ifj
+WjxpGmQawkAo0ZcllcWx+fevCn1zi0MhPs1ugVRzHC9B3ZJplBZGT7qkTjc8sTQT89QP9G3qASh
jnEaYM50QikYUqrsvQO6npoGdHjAYpi6/bsMyhTLeGNxLe/44Km0RBuynB4mFEO4Kblujjf882lc
yCHoYQQx9cOGtX0FkB1IDKBo0OoEe5KNz4b++QgknHZteIJbzP8O8u5kDFPYdJfb5yxShbUuox47
0ff2f9ceAsuaFTgX3+War399tOcqg1BltVKTC1iLiOwSeL59ToDjOqOiEXVC2m+6mVuq+MsKNJ9Y
82z4ww9a4wi6fubpWKfVW+mxnjhg50WEUVh094sO5njnWhVYTI9rz5R1PyJ+LSubbGD12zmzKPTe
93KTvmQC/isdJzc5swBrn0PICdvxrBUoPBuE5t+Fv76RU+CiBEE/Eb9Kvf3v+xei7ne/s4TnmwII
ONuPG0buNOWgoxc3KsGfmglFr78cyu1NHMYw8ODo+p6RCy73Zn0SYeQYm8OF3Vl96hcylVhcDwOH
0XJ9kbXhHB/W8wwbdWauSNtqG30qMQP7nrJ6nf8inmGNpCB++X2RmSgvJnG0JHAig4vlstXIjTVQ
ilsAGAQeWC+AkHp2QrYzP+YVqjj2ULoKzS7KdzkbEGF4TPKiln+09cPij0HkNMV99kla4Un98Z+a
ZoN+7bi8YMjzLTCTki9Y+1JcyvrTWcvTpLj5TWgdznBjNGn/UaJ17oX5cZGtvJTZEj0TJYQFFVPt
HvOQcIWlC6kfYuoeETzT0eGg79MpX//KemD4KLl0a0Sp/DZCIBOXeZxBibh28Zib24ls9yrt2V0b
kcNUl2ua/xl+kKdl+gU9Z1KuNd6eeXwaNu0f/g3Qh/jXC+Q9pgwb883v9hjBLT6fTYGolY4/9dwZ
QkpSAT3YWbqja4rfzgSZJrg1gCLaVoq1uBZsn7jwrTVU1STyEeXUw7w/RwT7pDACk90OENi7iAMu
qJM/VFn0ZG4+4PIcTcHWrrRJ8g2gCwzVSySChLLIExQRtRpQUxlFVS+eV5+PC9s1u1IG4H5hlnuD
owF5KcMcAKxoQ/NFNblXw7k21E4aWQ57UXLRHbIJ26vF4Q3xXrTgON3ZoesvGaF+gj+y0k1q9/D3
sNvRJOmuCtxcmnNah2H12oGh6GJ2KgdqLyHBmI9ptaRIbKHKjw1X/6t7pg+zZEX0HfEqu2pxy9FA
s0mkl7e1LtqKWIfDFkib92Sun+XH1d/Uf+UV6QniK1mxRwC3L9IIegvwjDD9xOlqaqZ1OPi1x8bu
kutDqLoCfSbU3t5eV5wCFoQW/7I/9oro7yn4gS9NzL8o4LOPatw6yEl6u5UMfZkOCgP84DNJRT3Q
dTxEYP+j5hb5OSWlxO+LbwP3QKK0l3d4QWR32f37zlQqfgEfSVNmdqCZVF9QLN2gmqpSKi+8TRWB
yxwSUwwR1qMrZNRUBZahbphI8CxhDcsFXqCwyGEWtqRW7BQZDNO3s26HaZwHzi3IvS03BPT+nz/e
IU81kRah+GXPU6J6fXqSamws9VsZyOn1jyq8id/8bsUDonEYDmLdsIZ6kbkPnGBsFdbUngf0f1s5
XKzCnb2AIanRAP+riyKRuMeYt0KANekNhRcIZ8vkaSPdE3Lll5eHB9SHHvW4U0KaRFfIUlcqyhaz
QsUgiW4SOVKpSwlU2zp3kpvoeihEQTNqsOvzpsLOsFLRyQ1k8Rq1RwvpQeTnYW9BxKXUm8x1Zj2Y
7JRRzR2YOc2CSSp21e4Hz6/U0H0nS0ApXGPutxZFRqbZVGHXFoEOHKffCMvUDLgQtTjJZ7d/kmg9
twiJ4a92EbOY7w6ITU72Tdhc8uZ89Jag9UGYXDn/9AQ+Zrm+j33ZKJdHeJh6liagQlL45UQkkwrR
dl8HhoDOIyQ9ZfLNxkizkJv+6U2ZZZOxsLsKVAoh2JXAbjp2ceZGjK/7EnA/+fqzWbx7oWEdAi7a
9FPt7AM/++6hQx/gysJg2KU//w13+vpMIPgetScwe69Kwr/ADKoSpcY2H9gsUmz3TjqjA1kERcin
Ht2jMo3vQEF/Xz3dh4QlDgGyRLNaIy3RpGjDSAzVZife8jxJOv7qmydQ4Sla3DTzy00l+rW+Rujo
TBP5dC6EK/x2cWebL32GySYaGSOrIbXNOmE1KCsMZeLPdqlkteix5T+4KqA1FNeZoFF+cqG+6q9D
fWDwdczcYfwjYX7SOKoFDsrGuO4UevAbu1A52QDZfQ9yE9AsNxJby4EFhgt7j7qvx6Mlxlo+ShMW
GdVlXaorro72YzHbnP3Jtdln4q42eO2oB++A8hV2WcQpqLBajp85PigAMD7ATi/59uTbMmBoTsL9
Rp7Yr69nxTEnNFZ9ckEAgK7y6OUndraeTTOZlt8X3xWQ3Y5xew53g7PSS2sAS2B1LjyjU6pxblDG
F6af8bC+FsOr0R6adyCPciJ7B0/Z9XILhfAk2lEO159IBaxgvZJJkAGso/fSOC/RgFojZZ6lyXJ2
zHJQ9bj45mAp1KMkdbDoPYtGArKwpDp2NPAtAuxVGi/MBDTMgwGqUtXswWHXLMIg6fOd/X17vwSQ
j/BHwxBrhL7+XQlJzqOMjA7mTt0PfwJmJ1drIAQOA/bNhFxgqYosqzmYLqXFQaKIxA/l532WqtXe
ypu/oClQm0O+incLRiMhP5tVlscI7k8WzWX5qzY0t6pdrNVKGbuyhiESToBosbE4psS1nzG9FMZ3
/fIz7bmVwe/iauoII6cK9qhGGvKoBj1GIjPbJTDhsh2aA4bJnC0oRzEr5alptT0fBRsO+3DsoAvH
Fvp6WG1v2FE6OrcTA24+ft1u+WVSi5GDkXagiiV7YyKrxYRn04s19mvcx83qCiqNjDZyA3CEDI2p
8k+iWt2bAM2Kie4IV4IhqCQZ8EkWPWZFKc3Rtj/BdTjLpFYWwmnDEVlDnQLJEp7kWnMnX+dnLbcd
FCbAsayn5s7iHyepGPo37kvmLrOW6+ULmn5t8Tmst9kPS6cPZKXQXn1+iTGLEBBVT4PkIWUY80OU
hmDpd172cjlnqqn3NswqXhitT66Cn2SY/txoJTfh3l5gkxTGLiwxHYSOAvwhUlSPq69srMhPgmoV
t2WcZ8NO+k6QGrQKnspDw2JPA5IIorhykhoRM8m/3F7RrRcXO2Xbmt0tL09aiIqVU+ROgCB5Ng9n
FM7ybGXdxA4cqXJJ9X2xwEAxLTACavYXlUachYCyVXrQh0YaExso2RrVV4c5iG+aoJJvU2yiVy9f
+aPlEYNKPgchNnErLsG6VrV6RwEGmB7MPh7iOPxLOi8jX02hMDRx0DT9l7OWGPhb1MzHhc+RZELj
CbK/ONaHczDwl1KbpDjigemqWrdhVIqNRUUchqmAQa5Mc1kCJw7jbTg8uxhIh6tj2jfdp+hL7/WN
efNUxo8eLYKdH7FeDbViJHhRN9qX93S3aXYKI8AA6ETVpaltIJsLTISysymYT6jOyeVeha4/+3LW
aaZQhlUELXrZYQBUN8vP8qL0e52Fd1xIiyQFkLHP+ryG0A8BcIUFtFdqlVuafB3D26wt94Ptg3dx
QSe2CLDwJUkBRla5Bzxkoh26eM3A00fci9TkdGVAaE9Vchbf6CC9PqktYPXs5Sp2saRzjTdpmmkW
UtpLTTwYTCs8aZhFhiLO6mZv+qPIFvyra627P26uCXJje12K4e8iZs7Sccn1qNGpESxketqr0xTl
O4ZYDX+xUilRYEkFJV8deOzJYgcWAQFzMmU5Ojv4f+OFCJbF11/UzMldvMin/kYGfsFVj61upI5D
daUoO/JbEeKbuRqsS81wAzAcUD2IFVvNPOycDGMCtuz+pjoxiN1HU8GLVOG4FQNDGyRRV5W15/aX
YYNc0TNeMaFlZsYGJ2dg6HJt/XN2xNv+n7L+4qd+wKV0+cTWv4gRItXLBS4g7xibtlU+B8PWSHve
1X0q9/jfPCfJJZU7zc1z2Ib7T0wVorx4EVp0jUCOxY5na9pHFSWRwCJrxTtrPLgutDmj0saldvaP
xpJhHxqHwMAYfPjpldp4SQxJViZxClTZsdgd6uzHghRWqV+cNtVHmuJ2suXalkC5SDydGGMQwCDo
EesWZxCVrZMXambGaatnXTEsoOSudlWEqCF/NAFsIAMakF21RjfcAYuKl43BtS2rk1iv6wMW11wD
MoM1dkXe2GXG9jAmMHR8gcVY3HPIq8zuZY5mxl07LsELS7wiEHc762IC3tgpdQ6CM3XAx77PqnXa
xa36IaXROMCXzobs8vdU3DUp1sNARqXIRz0mo2J7iynEi5DTmUUZ42NRNks7G7cPrebQAXikI5kd
1WSak9nMA/PGij7PWIyKnt9wQaqg2pkhlN2eBVdhHi0i1ynR/hIEreh7myDzvhVUtEdXkuPNgcCh
OAW6YN4CTfVDJoWqm/BbekkaZvvbIOGleehM++BOztYNvgnUVoT5PzOU88DH/eSGBreAklBz0sCW
NoXfmPzu9mH3oCOsIX/kCT6oD9eRJm4aEMHc9wAUvzchrUaQMe6lk35JmyZ6QJxtHBTdk05/S32P
BiMw3QOJBc6O6bdJRDxbc9sCotlYCmrrN544ezbvrwLokdFMwhFJV+Iq/miqfQ4kV1oPyTTOZgW/
3gORCPovBNjkflJInqnpWlG5epZTDgmbLtVTsqHVnBA3fs/+pryJJnJIjeuYUF4gVbDfogAx4Tnb
SQ2Z7JveUf+KMvozauoG+iPEBGKmRbFu1SuJluG/RxRs5GJ6cAM2uisQiKpq+jmXxzvo85Moi1Lv
LYkjawWynZW4ECVDdoowmecLy/K6h5ZHcO3A4IcOxNqqeuNKDSnlvz6SOgyBsH2ucNcVy3aqAyOn
MP6lDZjtS6ZonSOJA1QzHUqgURgpX93mxT8xagcVlMPPDGYxVo2zyFs9jr+jeQJXPXZHfY21qjgC
WPItqmQVpiWboMmBCs0TQtLgah67c/sqpCZp0hU5yNVjuAKELG35YqmeBEw4fipVyAKpGmaTfDmq
yfGWUn1InjQnp1mTkB8+H3Vu7MRo/I3QmMvXAnWU1RDelkjKgi051Tyr7LMbpIuu87uF2sv1mqMO
G6Lmfbl82YJn+WhxRDp03ZUfegqffgR7A3ef4jC4K6XjCMwdFV9EC9FD4Wvfp93aFDMoDdd8onPr
hnLL+jN88gU6nz/Xbl47pY+KkN7a90tzarWbHjEuAVj9XyfMkdfZrDeCFOjrhn/q4zo3jJ9tFx0e
ytbDcUdO5HKbPGn0egHWIC69YgSqEDetYPQ8KI1XVFid9rn3YyEN5KpZKXfO56az7xLRfpo2hhDd
sOCKZqDx+693WVI7fPah/8BkHZORSg3fQ4LfNBj1li5lns9y5ZUwumX1b5akqNkz00G4xIbqH3gL
qERy3W8q3sV4wqQ77bQ+W4gvMEC3zbWnwGIteNgwzOap0HN6xmxXCsAgReqH6ydSKKXt82mYRWvT
qYRKsquWFgLwvMf4/PumTewbKFUd51CoUJhPeB5Ig55CQ+O+gJuB2PSC4z7teVw+TCABhT0j+oNW
QoISe4ek3k5I52YfrmOYqkM6pCYqT6MMI+Vao7Vz1kLD6mB7QFvTJkpY3UoWC7Q4oxA2psJHLVm3
wU/ROPzGsyzSu77AagdTV8YVc4Ir4n1gV3N3d8+F2rtYPe8CG3RO9X/IO42XQLU/zKSOzyDxBhxZ
tR3kXINQPMif9TVLMq9hbbAQ/pmcEdBFB7gLpky7HALauGDp7H54pemsA+mkE97pdg3TN5tqEHWF
a3Fq0d98JTyOoB9V/N1ggkilwEfGi5h/iNKUi2IXD6yAX+9rc2U079YpIcRTMHQC1fhqsN+AF/jh
+PR3QVoEU4nXQbmdmv+5pv1y7KHvFogeqlfdBkzjfWuCF+1lCqIKBd0W8KkQmJRbK//O3wX7YKDm
X5WFj9G+3D56cpXcWqrGINrBIhuQBWVCFESjYGX54gUuZUOdtaj5T6DyouEWTHzbSVIGBYQQzJ85
IHKKMuQwdgH/c63nC61w5cSugoJ6kVrFur8H/8h+ePJD9ixiUnz3P1owhC4lAibyoduo9q+CIfig
M3PbZiFJwP6sYakM9/tYYdlW0chdplcgCDLDDf1IV7zOn04YsIkXmdPhB7m/WP/50kLmrw7L+l2Y
GSWhW003q5/mxoxTunGWYmztKo79DTM0OFlDpzWV7/O0Ua4WKnq7KdrhLZp9DF8MwRShXvzRQV5c
8+SNESQRCaYIiosb4WsiOtQc8d9V8fkRs+Oq/zuwJs8qtDOwIj9q91smXZ70++HeggxMzbLdVK8v
8cj+7XDFwSJiooHxJQNJAEql77Pb92b0+ph8SaRjxhLhJpQFpVeWCFLExusmpIM6VMJAEx2ntJu3
5DzWab1DfTmIfQSf34VYJmE+cmr0ygzRQ5JW4kZ+iXcPrlqZa9pIFofEFjvcJQ/HtwdqLBK/CLyD
I1YXjw8xGowJvx1Q2h75fGgmQbACuwca1tVDkobVauswCG9ip0I5ZZaMPFlSJzzbMOFVf4GcohF7
91IzbC5Q424mQ/wjRgq6pgEtSSVufwgtB/fLsNOgDJpKBBQ3zXiFFXzQeyK3UpZYNF6R+rg0kfNe
jODrRgKXSrvJJbqxHDbljVvBsZ6WiEP/k2Jn6I8o/GXqbMfEvLZjAEupRaah9uzFT+UR6rjnSKBK
mxpUhrYyw+bwEEbyBrNOFgKvvwZc7M6HcXSuqq7xZ4f1tnxx/bIgHEFMEcNCsn1MqxNZZUiWMnqy
zRsY9PhypWC/Xu59u6VONRTSjKBSiH3kQ0U14Rij6zMq15VWGv7jt3dWxUnPGUxO8DgsmKTgazzC
AU9PJIFi1niwcnwFOD61Xwdcks0Z7gSAt9KLJEI2xRovhgD8zIg4Tbs5lpPHsmLgX1cc31G165iC
HaUn++lO4e+TaYPj+soOj3R5H6KaOb3Vay1QR2Hwqo5Q7xlrZVKrrmvAaNN1kpkNZi5oLQMIlsW1
XI0pMCkPVctXOmWI2hjgdI4lTnViPXjup+qZOfI7NoHC/lTAQaFkd431b1gWBlibarDxRmUHytgS
liSt4aU1aebsP9ncJfJ6UMqja+gC4D5/VJ5LClocOPqZ2mWHE6enxEeZ5ATGakIaKwX0d+bnX3+n
v5pwWb/d/VhiAMTs1EeLcN835w8cKX3swtferabVpZLtTSvz4SgaLLuiIeb49KdLh4YZ+yYV0pHx
JHUmTAf7Y+UGBDFgyu5IR3yB9PLCn9jCP0ryMrXGb7ZkcLJQ8iWT3MoI4tsOtg9kbqa5tCGrzsNK
/JLsaYjCXpAQkGCdiwQPWACDRUtTt+zpCxdzWizEhY0M/K7tSJyDpRtSor5s2ZbVxmtknECwVay3
tAURc7J4GSlHiaKWTlhp2+DBxPmttELeLJUN2Ulm4CM8r+0svM2ofosHaPv17ahpQiIUuobsuibO
F6jrYmvhxKjltDzlKMEHCYZ6pgOpQNSprhSqIuboF/hblObvAKT48B1WkuhvBLtAGkPlEbaZni+8
TtVHnDfjJ7vx4ewViHIxL4osHEzOHZuR/QMg9MXOKJ/mPn92L/4BxpNfKuc18aDTRU2SvHwjrFu7
WX/2ht8EP7ko6rmuxZFbMkwQ1/YmDhNJyCCBxVHWJ49h6Umu2LtDZAkyweGn0J8V6hZxpHvBnVWh
p6PBURTSBLJsEXpnx/+Ip41PZ28uf4HshmxY7I+fYd3a64cgzBpSIHmKJJtcVZRl/1uNAP6wJqAo
98i7MFJfTo8n+yfQemSmkQPSo+4djhFJvRuigCROVNM/1SWK7U7YUAuTGTtYAbETyldYGJxNQz2d
R3q5bxOQ8c40Bfctz6b7mk8+zDAyYFJ8Ow4pbFQMMhGACtif+jCEi+xUPiM2P19UVAI6NlD9zKr3
B9V4RunFauyxsGiMu4EWv2uDao63aoG6a/ZHbQG4ROd0BeTWM+h6MyE+Xc3cgesvcv6DapfF0WqR
xH6McRmQ4pcS3s7kpi3gbo/C/1hgcJ6PeCNnehjr7QLd7FoE8/bFY7jyKw8ZBgnihu8YxL1/NgdA
FfdvMO7O06oNaxLJkhoNirCvGSl0k4FxxeyyeS/0aTRQYQlQ+DE3CoFOMBKcteirezOgAjxLZqCW
VMAwqu6HK1QoTRKJf2+M8D3sMzaudUBxIj8sf+2FWOwgalD6NDB6pVRWgnMCB89N4V6rOhmf7kSq
EMJ+YNTOxtKSwOFvqpeTMJixGDaoOOh27POwvUDGOrIxMiqNmI1gkahhXJKkjZfXSZmbt7IkWcYP
2eQ4ojK2qd3+CnvI4C5K0JigtKsWa4SCEWnw3dBgnzf0cvZ4M2w6a9jIcggv1H+eWF8rmZu9llw+
WmAs02yr7J1rjlfnlEDDLFB5+6WY/Ef1Larww+csig9qURKQBFzvf87vFm/xh7gu5/kRqLl09w+N
yAPBOIYbhMwLcXvSDmTJAReGcdrenonqq2yRQQ9nU+ItXFPTY5I9UwdNH1RhBpSr+uaick9jO5IW
U+ICz/Sxx+5kNLgAQPFLVRcdBCtjILDmiT1M+U25sPiJlJY7tJPTlmVhs88lfTyq8xRL4ZiVOZPj
W0x1BO0x/zdQajaJVLNm8nWIPNhPnTgoq/zCZJuEo/UehOs8G3exKOi1qXkZnDGR7n/V/XxlMc4k
VYK0cSRVOX89MbX6+cwTw19xPsook+NJv1yEKqXoTJYniFxlD9tC1HzMj1+T5lPxYb8mM0RvLTPy
xCTYYspSY7lvFywk0zcDlJ8kRD8P6rgmnDBy8TLJRcEaK1D/woJodEq9J4Sc3e0Zf2L7pKih0Uib
XVbybHtskjmQi6vtcGXOXR8+hAPJAXZlaSu9nbAD9bqcVwL4iG6AmqAt/NKgkYsGpanc4tpeLVuq
9yPaCpHm8p+n1Ol1HB5R7qcyZ/IlN0LLdGGJgTd3gpapt+qx99CLMT8Ud5agt2rwcXiSSDtDnJli
uEXlXFPLuFvZuWvTqyXf17NS9HPtk9UibekT9hxMwDiICm35JTghFwlVSYJhdNsVuCHPcDvQ1GUy
CcUOEe4zh1JlnDeR0H1GyDGudtq4tDiwW474YrTmEkdkGvv1Ktpgzgcbrpp7ufClTMAGBD91+tW/
MCwZkkDpMSYl7FmUNLWwmfYc7qhYCXft9p0Ru9o0oquZVD4knCOqi3oxo/oaU7QSCAIAoRXMudxM
I7d6zbXfspu8xBfb50HylfMEEUwio47ymXFzkg38qN8MDqi/D7E4d0Aufu1sz6lqU6wSyI6V1u3w
3Ca1BEkXh/5mvVNa7W0kOnXLeiumA9KANd5FAPjLzUVWa+Iifi1SJxaP2S6m3JiSfYq0Tl8Ar8pd
TQyAuLKmKdIYRS+AI2CxUcpc5nBO52R0HGJSognTn2WelB6tvsErS9hSt6O9DkKVrTVM9Yp12zod
wDDqMUlhZiguYetUnuY+5ysdMVlWRBBYDN8h6d3sRWcZnhdwNM5viDyI9wtqSb9Y+xi3qowl5Gtq
+qkyZmwSTjM1XKcwEHqJsG1xyrcrsC/HpwAZ+plndnFWN5Q/Kr4FLAvqTGRbhjgKVepcY2lo+Niu
KvZVGCTytf+jZx+rdMGXP/8cpQc0MYzY4sV6liHcjgOZAYqcWS4KvEdLD36mWWuh3v9IuMCShl6E
9paorBOZhPqbFdOH3bZXKwg2S4g8Q2h7eK02yc2kWrEYaS/j6APBILaVDww5D9deq0NTjnFZbakb
/Wx215hHm12NfPQgdC8paTCg3fJfOgU6CKvtSapLP9JICOITXoXPqABATPK9dleC8ZuOosxE5D2v
6AZn9Rivl/k7CEWf5XE99VkL4+8p0sZHYqdbPnJaRf43n0vhyRu6W6d9HtXyt5RW03jWiA0oTxiZ
Aw96dgEW9FuVE0P/wjV6k4Ezm534ksN6gJ0v7+cqusX9Z73i6G8dQp/K0VwGSgA+WwebJrOW2dwW
w6ZzSuUsT1KFAgXh9Y5GmNi896myTlvKTVQryEcrGBn0vIjLm2/gaJIJUDvgLU9T4DLzSUOym/Pm
WnOI6+TjQZemUov37ee0zzNpYIHJJsZiOVaaxFSr0jG/HaOP3R6hcvQixLY5i+FRJsZCWMmYzRwx
A5sIA1D4+e/JbElcOXed+6TZS6GXdwdEWFMgYTuZVyV24TVgNrElSN08/GXfaygMMxkRVmfKmv5A
gK7YhG9q9Z8ATrNA3JMGiar77Ju7Rfc/pO5kTnoLXuFu/5JzbW8Ii7aZl7dQs80/pHT94Ymc8RW1
dXCHnGlKyg6YHFZedtLtlCVujyrhvfRzpoNtinvmav5ngZXrm8bQTQ4F3D2IGSSFSazTU1wtWFwr
mN0O9s9YUXSLZasKroQcd2IuawG2zxpaZiJx8j5Jt35cRTOEMrGNCcG5GnOulWpMkwQrlMVbv4/1
xeK+WV+y2Cr/kUz+kDM2Rkf3qJdiucPC/02DKrSgnjdkQBcZ/FweWzrwogxHhXG2yfRq4QOhhGok
dy0XBFwa08JhWunsSYAyyNLuEpbOc5pBiRj8jbSuxwN1JVCbJs7PQeQa4BGFBcNkbQAtI7p3CXxs
aM2hJFFPtNOSgd+Yv5twbSjjXzOyEFCphsYfUZbmY8eFaUU4Ru8ZxMceKZSNuKrobmgb4QSWIyUc
gbrrWnTtOFgYmb9Dso4PwKkwzGDicx5H2uEmsVTVLJyy8Bqo/ITnm7rR7avNby1vYR5aqRfsOreR
KGPqrwX+S4oITOmcmaibFE+4RcXdtj+/heHZMF2+S0+ZfxKE+RHy/gltPHv1oNdb3J2JOuWTU2cS
Q0nR6cOqGwWQpb6j8X0wmJ/fVkp52MFjSPq2v2XULv/2MxKGx8QqWSHUib8xmoGo9lafPd5aANrp
acZYqDCeB0oGMtbqcYh6JFdmea8W/ruL+33Cb3JRFobKm5DvcanLeWrr2egoOmOJoFmyFT9DNCw0
DOQsqsAtFozS8Q+i64+WbeLNAu77VWktB1YpMEuYv2sVexIbwS9vfKTfFw+h8iaML4KrJrQ1lPEn
lzJPLd51Csh5q3dRkAIa6aO8KRI45oK0y2I/i/Hd6guAP0ww/LcI/MBpxrxNOSIUFvZ7tbbX8wwM
lEdi56RxJMUZzyVfjAesVAy1NI+SYRZVdqmopq6Hj6ijGRjkU9K+CmpjIaa98XWq5pp9KlhIQqKo
0EZD5G6BVuSch/hUnSDJfqWyrzoIQtBd/kjUYZ3KbMSPm9XFetkC72t9KLD0TBHyD+sDuvU+4J6s
BBJvTXVYPIUzFBPkKRInUGWy/FZ2DoBBDFnL01e2K2HUrP6cpXwk21+eOR3iTI9qTKDkfVe1Fg5P
2HmsMeMaHzdHekK5lK9F78T94tVg9kFATs+Cv31sJrPAdYfwu5l6krnnW0qB4bgIwB0g/oitF6zT
dy4Alo3rImy7uu7J999JJeQh0BHGSsJ1cYePf9tnVA6nstOhoxFmLy9cZY/OAbLXMThBaJnUX+vW
0EAu3xcvlJlx75WUczQG6RndVSTYv/Orkl2gSQDqYri3QIrJ1fDA+97d4/teqpSLoDcj6Rf7RGRa
uM31j2YZbEJXtGYRct1VDnCjrUBZxjGbRJFni73+F8FGT2Wgt14/XeCu8xDdoaLnjB+bbP+x07Si
ACp0oYphnNxzfj09IUYviEsGtAr3Y09kXYp7bTIqqBDlST+yQ//LdT3Vh0DAcVrA+UZeqjFmVzRk
3CWplswntapU0wm1QIDH4L2MMH2g8FPqkshh6Vd//ITNAdElM3+bdkCAf1ib2w5CGxss4ALaaZlP
XdBaF0Y0KDR7CJQ5F9aXeItyax2ydBSgp/fWOB6YW+bz+LBZuDj57VO3/9x3JnBYq2dlvFs7RAIa
KbQiYYD7vxcqt69JH1hx9I/AZZujsDaS2xpvwLfWOS0GsSeioA0ZFyNrFJ7pazAsIaSU8l5HB7PF
nKA3ZKo2HoUo82JKz9i+VCgp4cttKRnM0DXsxHyNJt/hctehM/FqvHfBVil+gIX0Weq6nck9Jufq
aEaDiKyF501uNyQ8E3hBlqE5ghpiUdpe5nfKOAzlKlwB8EiGiCmJO2KQTy7oJ1PTxMN3kQ1IOoBJ
Eyy2/u+M3Wm5Eh8a0Wc5+uOnlIdzJf3tHSVDKPstrqQ2niVcR5aljd49x5kdpPZBqwlONnyeM8GS
oT4KUrmoZC3t9nzMwgJoekph+KGiCR5OOl0wRdLItvV1P07zv4/M7n5CFEJJkrp34GECVbz+sBXX
fYaBgoQCR9IOoj+BFWkfKi2J7I0MIC/oTRf4DGSufSWeoULTTgwUR/zgoTNOUGAjuRRpz22XCtks
IhPR0lGIAnTRpW+RjMBq6fy4uqgXl8tfivqh1RSk2QBLCWCqAs7SzRZxM8xtNfJzsBROLsShFGR8
uiFoFyAl/KU3bWswrWtyFWL9BTYAZ9D/H7zlKAaaTNXY7VcQthLrCj4/FpbFdslc33tH0VMl7psV
oIz6HQrSAlPE74wJWJBVpKuZ0+rnToZok8ZmB8jG7bksrJPKXTQy7EH33SHiiOLAvygtTnKfsQ76
eRvnKga0okSAZhufcG0O1uKIX0CLRGDAIuPr7tBBNbbl3ctD7mLNTr+F/WzzBs193Kuvr9WUj42o
UF7y6DESK2PZfGfZP+pIU/0nxeowXraOv5V+CBbF1IJ0WO6ta14o31XMlq5Z7LHQEJRiuj5IvvuO
DYV0DlmoNrCOKcPA4MViGppq63v8Tdl+nFDOO5pIqS1oAKQl7tmZJu8NFR/Td4iWRqKktayCEU4R
4sv8e7hu2gGX/Ss++/E6iHn/NSCA5zcmAzVLIR9NXUuudkHUMrtVTxSPimOpqCQYYwL5FF1QYCkG
BQz/rjDqU8MfAUyJMDZ1rfUma3GFu2hKlH2u4DjsNwn84+qgPNHuBRHHZcMLImCBkORTMcOlNF4H
PpNtFNMjKGikAOreF03v0a4nIPTejxrc14kHSVcMfFFuPQVArrq+2NPbgpFAOVuze87wnz4AyD1+
YrQLdhKfBy/gt7bEGTlEAEzWU+F7YXOLa/GGyNgeZDo8BPnT37rsBPPkwaieESsYm1FqvKT2Pwd4
f28QRuNby8FnpkBhzHW1mnOSoq0AKJ7Q0Wp0nuMxzf0f2Q3D5Jts/l9ts/JyIdBJv0sg+rxhBdch
HRN6ISxllypXHyExIuglGaP2wDwfC5nf3NW/Yj7b8xDtx1/vucerNVsLW+R73iLd9t2oUUXiidxR
RjzZx2HQjathUb0HisyCbkc7A/GoQckwwt30mrY+CvQ7KHHrGvmVaM2N9ewhE9yWffKuB5vrb+qr
oyGCxt+h5sEKjdKsSfe4RooWGMDwkcxOf2PetKfX5PWv5CrNiHZacL2+JWgZw1FxQBFNDPe+iGJ4
9HufPH6gBYAjPSl+5o4jLfUSVSq+27B+cbS2eER+UlujurULEplKnLlIrSyGJ2WrH2w7oze4EB8c
KOSo1NRizhNNC7WFqU89UWw0EloMRDzwevruIiwaZBemwS6lNgtf05Y2dYwB1SMy9fwYvTt190vu
UgLJ0+7wbpXyhKr/AziQTxcKi7EpZ4PuWrmweysBCWYJzn4wZVv6A0FvAC/Gn8j9gGRmHMG9We55
CsbK2j4v78fq7/9yywfhKYTP4sfbzArn9+7cwpBXHNzlIwyT5AD9Q2s5jUPkmstnFnWhiPyNQrIM
GtGhMu3ES76Hq6R8jYHSvB+dCyDFqGaa873675GxR9z+pOcDo6h6nqBN8aMg4ajachS+BxQCvCar
+GrTBE5aP8Ymht1g9FX8d3qnKbna9fKBqBcddhB1rFyVSy/Ud5O0FwnvmKBQBGM8/Oz9EcxIfAxQ
CK9L777WMWTYEOo8pUlS1+mJfJv2fziMT4TvZKjgY6ENpV3PrAzG+qS83NEf1ml85QXLMLDWwZar
kIy7wiatBbiCS4yOWRtfz6S94HFQw1bIvs0kpcoT264A1G/Bui+/0LSLUjQ9QCZvRJUSEf+s6zFM
tWGDbVV1d9WDlnfF48wD4gyeTAAf7V90QurbJLPcondZ2s/vq6XM+GVUM9Y8XoJe2nuB5JpU1t4k
vWnyQDc1z1/HIS0v6SXiSE2kL98Yikp9gI1K1ICJNBkWbahVlaJoZiFKPB4ZGMBPD7vjtH83vlhh
elA2aaKkTxMBxskkW/DclKlOJVnJPjzPXHp/ZCjb54mwtcrnoJd8rkVtwazR7n2NkqbYW7AkR8Nu
x2Dk9faRC1QNnmzm6tb7uszExdujV0lZbv8Mhjcc+dG1Dup0DfYNwIfGCdIu1qHSb6l1qm82sBlr
uH+juv8R6aIzoILaBmWuEUChUswMU7sFl3M8O8so76poT5tRNpUvQTuuHyipcQL7bF1MeMe/Eov+
y7EudqTkEmcIH1sjBKs0Ig5fB78VW5OoyXf3ijUsdJQjUx4+xk//vfzfm/jErs4H2WB3aNocgOca
6hkiQy4WgUrH0/M0bRUZHoMYDojXrrhW75rjrFDppBbtAzGYeFgHpur+baspoE5HBQDW081PUaGg
qXtHT4xoIv5mtDXyW9nEUBn90j8l7zCOHBMgIccB2JjHLoM8y4/VaxP4ghRBb6/zs2n7/bhLb/h+
xxNHie1g0V5N4ovYkRBqA9Pse2AgPVA6eSeZ/xIqPojJrsVsh71XfdTHEcWAoq45xMtfk7fkq5Gg
wfieHS2vzSbCOOd21ei4Pouh5f/VYthT+XLTyx3H2Ejy+M9M5nf+glQdhtaRxuzjNDYMQ+x8b50+
AcOd+7uV0qlcqstuHjFtcgCbokZ7MQuU2WGi2dqAKWdZGeoFnWvr/9tqXJ6mGBzoy+Lz+YhhpWhO
R9wjrWYOvxHI6fWN5A8iGoIn/en752A48zgg78wx5DqnpoOLEFbctmDi5/dlarPm5dkxrt7FDb9j
NQpEWwCr/9p2gMpKNokCW1Ok3c8dSc4fB1HJ34wLVfXofifkPXEes8gQa2zOMsrV9ra3+dvb4k+r
2PRYMgpaccyRvousHcUEfn8KroyOBt9UAkywvb/PEyw258Eb4J/lVvXjpvJ5EkcYCkKWe2Qv4NQz
h5tSE0zO6mZWwZ0WulHmyB0M+IB5uMPtKgwTm/4fnmwcbMbeXk1JwTBa1THm1/NtSX8LwOz/u04T
qImLeOy6J20OEblq4a4Lt5yHQhlELAFfH09nTVAiI0db7+CtrZsTd0oBjUzHoY3uYJn1KJijR6DU
1n9+Uh42C4LoS23s954vmxDJ3J5ms8WgNa9sNX6e2lasB3VQ+vq1rPXuNEUJu2CFKlOa7c+OCsmJ
cUYWOktCYxAF0f353IG8XWXbMDCs9LpBHPYVq/xwK34zU6pnmMcWvn8yAvRBlTAeS3SEKBm/LHPR
8cMvWCnASlr3M/X5aw1KDV+xqzHvYTJk77KDFs4rQFkPme8pZSRAtHMJxd7MGtwcZ21ezblUiwOW
lS5jSJ1Rn0om3GCcsEIq7kDftwFwAs8nuu0T4e8DRrWnsPNjm4G4ERaLCMEEDu3LN2xtPf6pS4nP
zcqMlr3L80Qf5ygL1CzEbqJ5QDNbpqY7ox3YF4YzkF90aF/gtYTb0FVoz3IqHkipF/4kBdF9fYgx
EUl2xVsOtQaIAMRwmRDNloX3jSW8Zpq2B+AdPo1ydM0UhyzYkdLawHXheWrO6OdOULBbibvX3+FT
IIDurJDuX3m41F2Oybnja0sbi2q+xmHur3i4IOUEf8QzU9gI/lXkbBHuW7MK9eViMa8f8qIHJvrk
grssn5w42sYJWita2A4SmIT/7GwtxdZKmLno2SpKITbIJlBWVthPSQUx1hk5xKlUwbqGbTuFFIbv
3ySupw/vfp34kXbgPQ4n6MN73cB9Jqp9SuRdfPh/pDIOKLOmXgHkJPkuLYKrLk47dg+3BnGX5hkx
ZBew/e6dslhdNlnM97hIyM0jJZ0lnczAKmsV4pB0VjAe8E7aRSV72J7Qlc6xQs1BHOxc3ah6/Gzl
5aOrxnINMTMB3sPBbeNOssV95Lh+hq8VMyQZVog64g1MKDqvw4OUCGI9jf3XdOzE1oBkA3jw73lG
kxymFnp3t5CXAUl6GySIaPF3r7JmBo5Kbf10ZzWHh/f115id6dVJErj8pRQa7z3GzdFT2Ad1XoE7
go1EGkoasmq4d4sS2gSyncJqlZxCNL7y/tz57ZvJl9j+8lT/SvEJJr3ODTYYNh3QpKd55PdQaHjC
0QjJ3R+1ca6ISiMvkWqvmHiqGaUYSNgFCUXSdNlIAI6HZxINlT5s7AhallvdPQwRD6S4Wr2lJK8A
BlFmEDIyRTj+rnm2TWQyNtanGcs0WDnbOrgm6a278l1JjSTToiydXCxD/VqIR4OR5k+HK4xv/Ohe
WCNbyfbALgYQICPxIn6MP4skYreSZ8IBILtt0TQ0hSZCDcGoQ4Gmsz4YYkGUrzUVj5L0FatdFEIf
aJQtrvhcMxkmMY/+pgcpoXUSoP6yc4TD90zHLnG84h6EmbOTGT2IKoq5XN28uam//PnjInoUBsGB
Kj+7QFW3l2amSzyNSqAQHsDWPG/BYRMEg3HSZPMAhOaiMBCxsRiCCL79uXOPTjvg085bl3IlUssR
ubqzwPtjRRGJWR4Nxq3IqgdeObuQmS/mgxLv9BAKquJljJnLYCZvri22EH6rBuaKg73vKb9IRLf5
Wb4lC1UfgKm7Y2lHMRar0IE32WJjmXBYJBWAs3pMMViSX0yElUXcoJr3xD91IrZIrLkwlIkDb/kK
tXKhNyyXVHG8DbMwdAdWhq16UeHwjdUWxInvLpFyqX61CbJGu84d1foC2PNKtf6jpWcjtC14x7XU
bpOdXvdw6L36NI7vnN/RmzSWmXiBTSY3zFlHaQG72rDnqcH7iy15aoeJui8oLNRLsh/LMJ5Rv9ng
hcj1UKTx0Sq28FhEFt1i5B5q19UaqrfilhVp6Ap5O0gmL6qMTqfETn0XRa7hdJ0Ln/SwqqSpYMMI
jAkZ4GqHs3oloc2yaI6WG4MutukaEff4AIoK0m5dPV2YLoE3ORG+uLUEteqg2Ct12NhzdwRkYij3
LRABsbL7oyxzQon+vVvs4x2+TCjKHo3hYsFc05Ms4R5N8Uk9uJQTj4QL291dL3YCW4GWQc3FAdKv
HBv6C92ptpW1P8rHw/hZqwDQui9gLOqXWDnMQ3mrmcpQlO2hZZfaFfWAjhKP3yZYB9I6coux/0w6
tpURfWaBlfy2ZWwCtoivSmHfrC+2BYnGA2pmPSdraqiiwxtt+yi5nqfO3z7m5iEQjqCCoQBFRiph
QPrtdiKUY99ZXse68vrXFaINCDGBLEVyoFzwKsbu3DLBVdu0AhPv4UAbfVsb+CuQ0Yd7Hw4LIgq4
7aS490a4PdRZl0KArdgyC/PIfv+xrX9LgnxDKO/5pSCVK3vd8J4hNLmE2+CdGTfx9RZBuc8xevHF
uga0wcKiOoUwyw4PewSAUJNxFFBRJ0RH4zqgWfVO1p5Ccb3R3LyOF+3MFd2FpWmC64ZJoaIEddUg
f51SHjyxlrJZJ+Vr1ekfgMU4q3K0WShK/z/hKRZ+UFim3kWpMUV++bFIohPHTeo0sQodz6l6t3wP
xtTXOqZ1/JojS/UhgfvTrE8sU4URVyHr9f0Qi0TxUY1TYJR4NOva8vKu9ZJI1RDbOEvSiZWX1y2k
mFw/r3S5hQk8nbHO2zigDeeSLUuZye1mMLA58G/YwSmG9FaV2dQt54vD1jeh3bu1fwjNUI2FNLOa
jAr3WNedrvj39qb8+vk5jWmdvAJHIo9bhtMugDbnNJ+JCmexvDGTbK/PS+fEJ4sUocY2m7+nUHRU
cHsHpz2MFYTfLA0x1xeHchNWFe5cqmb4SK34OjCp5C39vFTEPuRRDp8EA9BJvkeZyl4VBndlfj1O
riMLnRDUaGTyuubU3+H5ONyauj0W/ooSBYyBjUFHP55ivKiwhZGnKzE0TGWTGktRrZU+lH1FjBpT
vGGuh3JnZzDi+kfpUDq9DSoRP8ZEMBJXk7kUIbIcFISsIY2ktCt2K2s7awUY8YNeg9j5PpV2wXG4
pikw068SFL9bA0Wo8E42+D+oIvEOSkLlW00wOaGe+yhXtlmWjwc2rYO+fKSoKSwaYovJJWQDsIE6
kIU8WzD/TnZOR4K93SJpxe30ffcD6UeKqbm2lq9euei/zsHdRe4nmdAyFMSi7I46lq8piO9sOTgT
dtk1dreROFFYiF9B7zMJ0jCoS3exkDFNf2pz1tZ8SIliiEPeWc8QDGVnLsdcklvsi52PSrBm7PvY
sjVb+8PSxq1h0MHH5fqMo5+W0Yvuc8/L+G+FWpqVaUwxyhIZO2ts7sPc20aarDgyXILyIiTEfpQM
L+Xn7YDf71LOJg2qsPVkJTwbGceR7X/MtXCFf/TP8eCzR3y3zWlab9i2N2PCHX5A/IwJzSRpXv1J
NDCYPPLdJdQH72ZUjFpBwOhBaoDVm0eSs5SlwOnZRvdm9NV8b4SS8gTVpo+rqa6pC6TRjlEPkMw0
zdo3SDjaupk08RBYFgvtrpWwKo5bZ30WUhRM8QNRDzQ0HWLMZwBLV/W3P6soDPEyf/fB+VOvxJ3+
6r8sxSwVmkrnlOV28yBXfizBeGDXsgjtuTck1QTeivpJZ9o3GS9T2OJDORNgJ+k+V2AnsCRN1i0g
iiEfdXzIoWXn6o1RP89TlHEUdLEeTCNfs+SSGyLxHPHdn8lNmuYN49j0u7xCYeoLZhzN+IVXIjyO
2E7fwhEhNw6AvaDAhC0QVUXuSqooS72DG78DAZV7zFTrAasw+16IP/4ClmIX+AjKpkaMzKefaTAc
K9xX1cLKen4GkUKCTdLXqAcIMg3C9ayNRnEIIaqsnBT1RzeSKGJZY2fKyNVvCC0dT8s0OVYM8YpB
W5wYZMd/lAE2t+UCwgWkPblfOWZz0j7yNmLPDDTPXruOtCT/A6gTIYOJFhOi9wa1LcrlkHWT0PmE
Du8PlUNcLB0JnG9jf8eySJippE+ZhI8a0Pof90CmlopiocVkNVZVCRfRwxpm11pf2ssXZSbYmQmJ
P42D/lg6Q+t+DYZDQrSwOan5VFC8ncHtuu1n1ZrCFOcqFrd56KshSgD7ALkZasieOXTWWwT70rN9
+/pA6mGLPmjDF9vxydw1CCuTvDLBrf2VeJ2O3rA694LdoKKObIgU+0xtBdwYtgLTRyqDP1U5MJ3j
QPp6V7JF895x54xOK96czRKhIXOqxZzBDJmDI9rz6EYJcL5EfVhfksddhxnmvJO4Dapr1QHU31YL
f2eXkLplL/Ce+NxBfV10fC3dH5tyqmcv7seoe1y1fwc0/RzzrwltgDASYBrMyajl1q4Q7WRWIL5F
XyqmPL9BLoq4MqJuO/Ta36qNtUMH3l3Xks2cWwPBJvVrDzuHaijZvtD3q3YulBLGD006yBfnzo7g
dvx0tmUOYcdk0KR1yy3xIgOsuLeW4nrNh805RM+RupwMAo9oAanNVAIpU0Csqd4JlshdEB/s0IvT
8iZJdzR7y3tak6hSgQ5MC88PA3qxwP4mns32xAWrBAvovTkJIJ121uR2iE34P9tjmBP5StDa5S5+
Ly5AyCRhQpi/BhMqprheqdsuof+gA/1zNnNLrgRFDZUAE3DxQ2Wx9iUutNBZamnJ8jkVwzuqFctC
2U7aorRLd+WKbCobgFuthpoh2GBkrOzyxD3AzP+pKS3OGlXMINf88iOZd334CTJCLrbJfeIpTFO3
qN1vFc/6Dhy1VVdPU228n4nh1DJxUDu5Ol7OF20uTdgzje4qJvqxpb07MyDGB7K8NclAHzJQzzBc
32/Zrjk+7Y2fmCQZX8jacDsssd9GX8OSeor8zkgrcZ6TgtiwNNMudfdzuBw2qpcxNV/EJZDbIL9b
cPbTxKJG0aoYwDlV13fQSjjWqleYVD+lUsqVdrKsGLLtQK3TJFCay6mcYHYzuZI7Rj/Xbqpepmvu
gDLYuiA7QgNIKL7RPZOUAsV4hrnb+8AUk1qjuEjiJtfSpc4HCkyf32SGZmC3WilXIFcJy1ERqSu/
GI0izDAkHchqQd2YRCyA4CiCKWw+aVfFiLP3WN2t08GP4DH0He44naFl8jO7hVetdSBVzYLdwKg/
0KzEDVs/FZOKYkf3IZ9fnS8ps6Va1jL9r8/yPg2vjN2SdZGCkB/7Fv9JIVo6UFTIP1f3n4GHcrQE
1J4m/2CkWizIJ61LTbsbJ1MgpIdtC2/7NRbmbkRF3/blcZU8mGvNNDrqyK+Ym5D8lmt9z16XfBA3
AGIIqLp4pMp+QKfNuDKfhwcJLxjpoIzUaTzl2l73NXsdQoK60XBL23Aw7WQocxHL02u+CYwozm9j
EB+W7zzLe9PHhqsTh7JPstGPmyffnbJ6XVf1zBzYLvCCyvXinHtVaRLxxVpwlpydfr6AGcmwhDXH
qlt08hIuRvom3gLYLJ/7rlywbiCCQRfHALmfMehPlWFbLKbQt7FyiaoCsaZzsDnlwLe6VfYjrR4C
AtgC1w9RYbbw6X6QXd6TTFUtIlszpK6cj0XWIhcGufE8nMOCv3rXD1uN+IRoHD0HHDkDKpIZTY4p
0LgPp0q07ZrZ/LeOBZ8yYRefAu6Pmo3jr+8Oy+YyO04hHWjrR3g7H66QpcXRCCIVuhBZvCfTUVwV
iTrNbnasiKDJs/BwgGo3CA6s2vuxKYN24H82MIJKF4rFN7KwuuEatyqbFDFkYqju4LsV0Qkv0Exh
YQyV6qlirb5gP8HeA5ecUPXzfph2X/pZKR/XMPVIYiFFNdpAH+/JqSeDEeW1lJ8b/68MuJGRRxyO
z3caQAR0qsy40OgZ2bnDuZF4Pww1Kc+FdGDvwFV27RhmGOsg+ueKaMKp8hQT+MGwNpOVecoV7xYb
IxlNyQ2ECRIJbLAfFkpwWB5vAeFwDEbx4WzSEqFGhPJHvPg2kP97PJbmnml4m4OGxPYeehTrys8G
hxgfaSDOQfFKa+kOYUZ/RqqS65SMUSDyb9IrumsdJp030Ww2yO1wtA9QeJwMEbErCnLmau231w5N
9ca13z8gs3eikexb0S19PGYi7JSflxPjA+QOWBKYy5j9sgLifxfbiXUgM66RQc79WL0AQ5iq3/MX
8gK2fUxE6io27tjaOl/xJ8UCWUrUGrVQIdszbNRMc9MJ/FJ+zq5AFXnkbg+nQ1v8gqA90da8JvO/
+0ppOH7FktlxB+luGNcWPGYB5Upr42mzWZR1GAbL9VwCDP2W38N6h16RqJq3Suoy71wT09HguSsZ
slOevrmxu9HYRC6jHnlPi5DFp3QJ3x4C76x8MRBz6cvDERMx6RhUGCbu2dyAIU5QlD8Uny7KkXMT
5h7TC0Jfa6T9Uc1ww05upzg8GNx8ZcHmYnrAK/A4uNQ0PsjMBO39liKreeRjRV5fTo9IuwNUFz8k
n5+hwSEMarD6JStl44yChiAoz6YpMedOcq0Nq6Vn+K6Fzn8LsUbAGt0G8xy4f0a8QLeLz0lPFpgi
FqbL9ELrDxMWzmq87Fff7L+LC69V+zFlebvmAW7oKHVmZyQsmm8M9HHofQmPCLPqeWDd2I6L5/J4
Y3F+kbFSFibgmPDzhzXKY/Ebxn7AXXH1Psah8EE6qxJyf0BzS85lNF4fQLn7C70L88VNmUlcguUG
ORE+qaclQvZzPpoWvJw1j61djXi+rKAJzOAIXUXOCXNShI18AVYs7CwLrE27S5Hn+Amp0BNGouKl
4Yv5pdD9inVzV79hg8htmI0raLQZQOhYu9iYPDBtfYBnaMB8AzmslvNXs3r2pr5yozVJ9DoXpYaw
rzS2yfQHxNAOarHrZAeg460F7/G4OQcsYiBULYn7+3Rwh4eQ5OjQ/28aVuU12nxV93/8Q2/Ig3Nw
M25LS6pIKW5IrQO0u+eZf+QJmAorx3NYLk1NPYy98QsLzcP1PRBG2q/M6iwmL+eWpDenq5ipTQpQ
/+xK3UJh1W3RHu98XR3CELkJZCGcP4E/vFn2i8XnV81Kko0qUGAE6qM6LCA+7h4GDn8k/1kKMn3+
dBWtBCmkopzT/jCs+V7ehLZdo1ZDyG33zPD0uojLD8XgKrervmgo0ucCsYrSZpN6QIYEhGxOp4OZ
++7JmgZZHddwg8Zy0EDe5Prmg5KM6H0plnoHQrMCf1ihslGZlBloSBCF6GS1peRlCsA0LApozo1v
/kFAEFMHUZmwFX7phDZlZavuyDNFaYANTlrfgnh87bLlJWidrc9scflPJMvHATmlYAgr3sm0DSwC
IjNcis1diVDkPXyFOxBM8iB0gIuUVczsvBlN6jOMxIL415XLHlg7XICtaW3Gw53pypkob9Sd9NrX
d7elREXSFUsXsv/A5+7XXPjPfxrmaS0oMFxSHwV8L6UDwVKD8pu5KwLGesIYt03By5ISK0heGtjU
Z1dAkLNtRS9sITEd6yx5yno6V+VoJHnkdpA3/HVR7yhJLDzK71xtDMZXyXdAu1JkAdEJ2HtWFN2S
4P1wEfSNRN1LORoHG5Cc3RQ3VuAOCH/2uCPkSpV/v2Q5KaX9kOblN7M0NFjF7XRvf+yZbCDYxgkC
bgx+cCCZ6ECOb7kDOQGsR1DBxQ1XuXTvbch9eBijAqp7pi4YqUqW5bwjOXMzIfcqJI764+Le/oJw
PZBJphQuqluunzwO9wCJ42IJJY5J9Q/DmKFLJ2bTeNIug1PCzOt4r2/XqCYCCWzc4IJwJfVL36Dv
ge1aI7a9XglCyowuyAVjRCjID/r7FFRkH8eoklJwJyusbnwWTpYb871yxEL3QtzURTpSdjtrFSH0
f+cqjyAMAcFR5iWMTfXLz2OnpuS4gyLp+A2AVed5WmHb/ALqJIOKO/B2EQwPe5nmjxs4joFys1DR
Wgg0CWH3DYV/e5T+MSTuLWjrVvt0JNZ9KWk1rqjnhdZFP4RRuSmFlLV7u9JVTrIGxF/4QQGTeJGA
H7aZJWzCyNVJ/qOlGrDSCRWuVnDS0NAaPhTNNa8NSyuYcmA0KQ3yYhSbY5yH0orNzt+yyBn533IG
DyelqRtC2BfnbLk7BNitTCm0XWrgJppeKNraqSW9tQG6+KhTHdL2/TnuCOOOdCc+xPqNr1ZtYsON
eUXeHSdNfh7H8hcnY3qkThurwcs+lsyH7Vs00de0MSlLf0gJXWUrZ0t1O8IcnkSOxLAUeP7OH/mB
A3qQ+JENlbt/cgkVlMvc9lFtYWtCWIQm1jNkzAI7vyKuvyMBSmw3GABxwHV3mu6w+l3QMMdjqIWN
rd+HcRhwfdg3ZRWV+L9/0ks2MJ93W4no2NKhxXd/RuSDsw555YQHMfBsNEY5oGRkPBxKQhROjS76
yFL8+0uDbFzKKGNfEZ3NmaPplNJVYkVZ2xtt6MF0AVmEWen4dicKOHVh/yaJiafv1tQoPwEXtloM
2XC3YEWsZa6LyuDMBjte4jRc3bsgmm+tLTW55P9Xqo5lDYoCJu9BV6Ghw68xZnR8oEzsQu8RTSPn
kKbQSPd/B4lpy5mpf8LRmH0KZWeTa+HFCp8QGebtzYEXDl7me3o9NWKbn9q0IxhleVzEyAK+jiGr
gED7ig1FFo9ms+pBu9okGHH0z36WUxHXbTC4ebgYPI1LH4PTL07m3OLxqpBhs0Ef5FXD3hqLknQ/
wOv10Gsy8xOe2t0D6WyGowDRtTzvPf2wIpocckX/U3jOenNtn+qpPXKKaZIcQzGGZNlxqRAi9n7w
ENXKfr6ijcwxfk3Zo71nYnG1REpRrnMFn0tcGSjDh87L+dn7LhiLt65dN8CumItxe1yrHXrIR3FJ
3nlt/a6slrJRShP6cml3xYZPhw5lTW/e4Sd4tnNUGTSeH2iBr1gdg51I2nLm/YtGjd9pPrtxiSuy
vpqqMtCHh5M1+0+hnb5jYF9Xwlkag5NhvOdL9C3O/IAsUTRrb5vxP6uQCAvbIy7wfzxcRHf3TBWz
0dRQ6AtyPDgypr3iabHVXTwSY9pu8YJ8f/gB3Y5RkX2vHDHgbLNbikXaLdxEihayMJjN259fNqCx
9+2K8lq86ep7LKi3tvmYjTEq7fiwDHDy0cMFA0CgYZIdx5C5gZVbOW+etMJPQCVQgEpTZ2+Eg9Y2
PmTyBT62inAe7uYlUXDD+9ZuAc0P9/gHhz37Pd9j4LhaFHbu+Qi/G8vAGyq0oPL0FENoYc2++C24
V/smyyeqYro2yMzaHuJdGMWH8svh5JO5J6G5iPgrJeUTkvBiHWPtn4od7WAesOpe7YCm4Y7FIBfB
0xKWMTkKR9emEBwaJCgO8wY81KVFVx+0a+rhuzeZ7a8bjsrLpPeQUNNShwgsEpxsbbAMezqz8fnx
FIf8TbzUl4MfZhxVOuFcTzS8BHVWV2cSntN31Sg6GkAEf2HYANHaXnQLCRzVQMbA4M9Bo8VsZ9EI
F/EUW1FWKOZFf+HuhqhVNzZmdtek1BGZap+r08VhyUYn5Ufk1E4w2M6KHzNwj9JQwCCSP0LAosHY
Eu/WtNBuBgTdY1vzoBjpD91m3f1jFOJS2cKUMiDla59lS9BtftdyKhY90WtScURzEQGPZZko+Nfk
NB1VRY0p2GCHv1J+auge2JDKRTCDWYG8CeyXGRMKrchcn58FLcugdWhJxjZkJLsTHdmeuWuPMvVl
8o3BxJNnwQ5PvUSN3EaCLzXJGW1g1ZpRuuKKyhxYMpmB/deWHjJfCG1Lr1U4aSSApx73bjzlQy1W
c6Ok1VyODQYmu7WIG9hHsQ1nSR62bQngStalkquIBWDhuHlMpurkkzJX7QzQc6rv6FNqYObV4vEU
y4xkGWgLaP1qpheYaqLhBwQHBauXqqsnTCqTjvFEG0pG7R1FJIBKm6H6qXz1oIjD0PhnhRjZ5Jhn
ZDB7xDHxNczfDMA7yrCl0MxaFzLME1EgbuxGt4gxyH/rXYlUG/0+4IjfCG+WIsD/Ff/1TZKykdWJ
wa2mJRCd1KrY7Kw/XvaDcT1ysGRTyc/OwlgOi5FSN/d08jnurufiBtNW/CqD0NkMc8aukSV+vZGh
qe0KZJrRg5HuiuIPw+ez3SdrpfRnA5+YU8AshiBNNbFjxDLgOpTs5aGt/LV2SP3qGXLIBkVrOQk/
qA57xqXTgUs2wcUW9N+6c4vo4FzLZGnjMd5JT7G0CtrEQ7j/SFb8w5O3ZgabO4FhFWEWUZa09TLe
h8yhYq4jL7Q8wRjEaTOkS0B76Bc7TKimWKIT/Z1JtPW3HJIk5n/y6uYYnBRn6OPryDLAOFzjfXGQ
6Dk5caINnSjdCWwt8eGwgZYVYZCcabKzSx8BLOwJ6YSk0pc6Fb134o78ROC4lTpbu+0ATLgeQlzA
G8hv3SFfy2TUiH7xMue/+pa48mp8DzGuJxn3mZA7vyQOn8i4knmd8LXiO2pnKgDNEyZgunssYrQ+
IzqqiB21+7zjCI22qDK4qY9Nrofv0S1HyYQcLfpZ5ZiF+b7toAV2MtMFs7+ijiV4QzjMxiwKWUbm
hJCltRFaZZVnICx2t09bnsKpv21gTeqsXGi53mGOg3ZxeAL5feUKovjPz5POt8oIRgSPHjAf5l/A
8X+FwTBG7UWuCKl1BiyUtrlf5qpQ+krAojXQkQKeXsTg0gAwE7TfMAS7I70Ntoi0V8+HIZsn4iC0
bS60/uRRymO7DJxK27fCguHJr9jWH198UaI89BM+N9XucvRlCjK2mxsizNZAu8vHeBGsqoshKhd/
rTNB7L6B5LisFIsJ8NpNCDz5tlTdfmlNV2K99rrui/3dHm1ESMtMtAWYpK975BENbJ77FdwYNKcN
Ww9NINXDH3c+zi8mB1r3NZPphpQ9qIVMnZzvwsR2AyyyEt+a7msFg7awU3kTC8p+vFjVsM5Rybnn
IyqLp8hvX9bz3MgdN+ks+LaKiYYNI2g6+0On/ngpYQbKTyXXEJ01jQ0aIGfRR59P+LSzuihsKLhX
X+xL/c0IjbN8G2ncImqrJ+SURqqpOZ5Tl+DqQcrkoZdKJQcDrd2J1j7FM//HH3zLa9+Kz9KhYzcN
Whv9VxnMfM5gGMfgNmC9eJ3mV0C9e3a9dbbVBs3KbN35fpHdRkP3axS7m8wEsa1gQy4c0jl3Whvi
5ZjdvPzMMUiPbZ14eUS55v962Hx5Xffvzo/S1eCZ7k5cVHIpqbUF/Iwxtw/akIv+c5Vm1aB/gdEz
fowIRe1OJPZ6N/8BLAcwV2BxCTmuGR8VYzSqdOBMq3LsGfXKkjG1y5GmZRE02sNcpa8vyL5XIGAS
NoI5JfuGrkXOz9KPCSlXWqOsnj1f+v3AirewwcnZT1yNH63w3IWW0t35c8P0p5wv5ZwpOJJE19cn
2Q5YhiFn+eQR7Lh5CCmwcMajVs8RC0AqeJjC0CuuSiUY2yy4sWxNY5veaNCDRueEwCKHsgA4dbNs
d8q0+W4QmI/gKXkXHvEVPHgBwR+RyomFsyjJ/bkQf1F0gOjtnJIJiuf2meppQANGLIu/SNmkB0tl
FqUzU325klN4DKqYgkYpMuwt2x2jvQaGKVjoiwhsiYcVHkJjFAFBk0xY6z+zDuLEyIvb9z4FeBv/
EidbYtkT8PV9CwlcPe9vC2mdHo0mM4SS8He2cgeBuW1M8ejK1YffteHD4MLbm8cWAKekB2JwSLr9
Jgoq1NovCqZNUc+XozE0sCLjsbzkPCODbsODeT5+XAHDHrkJOULybv1CnfHVNdmsMO8Jn+vN2dAh
WNRsm50XomcVjwi9d7ZzLaEamLaFl5X6rN3GOp/b/Td5N8bHeSAG5X7s8aAwJo/GOrMUFXEZvbgY
YOQkuJhKFoumdaRjRxL7MN+mG4XZzgbv27lAK7TcXF99bqJliYsFruhLS+NDcxvkI8VQ72leMjoj
w+F3s6DlGiXHwFxEQJxkyUYBc9oZ0b1TePfYsjApXo/73Hq5TIdVJ+VrpwPsjRjA8gC6xfAnF2+C
ojFpeRkSLsWMhY0JsXKdDHHPHcG5CRG5RYyWmAL0BhmXl9KCmG+MNqf7wUwSqjZUxmJlg5jvorK0
efwjR/WL6huuoKzvq6WfWr4w85VVkx8ayc0ILL6bgkH7JhU9HkTRNfjjn9gSinAkNCPutUHWn7kr
IWmQIrz08s3Pi4gwJJ3eFCb40FgpqLbtAW+B3sLZemqZmIlBtCU0Uzb5CBvpMzsH8mQEosvOKi0X
kWH3ceWBsDCmWSUcY2QKEePU6UHtUG1vRAN/w8wFw3ivU8TCxoUu7qxtnCyQquwgau8d9wJVR1u8
sPnzBOH+zps+vOIUe+XElit8HGdnFQpkDgnaJ/qWCpXRk8hE7I8n1lkCJKozICv3fDWQ4Wb9wGUx
Vx7COTpatbpjqRhSV8L6i4uDHyBuNp0zfnc4S20887+peUzORp1Qx7zVlRu1lH6TboOOl9MFzapA
NgZvMhDYp7JIY4GdeFpyZpcmp06T+/thpwALan8JqVjPx2WbM8heQbpf8QhwxXn1mw8yzivgnfG6
iTbAcDsyLF2ZBnlkROBeFkVsRmwJ65Fur4RBJqLP9/Nx5GM3rB0DR/6gtQo4NnqyaY6MkuwFwUWp
D8BDoDENp7//HiqyoforSR+PkaAyQpLDqM21i99+G1vqtlbo2prHZ7A28+WgDnVeaXPopclY5/U3
svtQh7k2QR+JmtSeiQSip8/760WtVM3rSuAfg/6+r8bKBXU7qXdjiGArp/V+LDZuBeSEP+ZqBwRe
/pjvahVQ3hNTKWDfArPX6e/E2IzVYSYu5ZidBacU62yMoGpa88Oipkq1pxXJnFNrJSFTq7ezLIFo
vJHPIA9f/jntfh/j8IfPIrOU0GmzV8EzikfZ5qXdakWkCq+6YP6imHqQIfgLa5wNOkp5juTLLBQQ
O8rrOJ13ispPuFgwOwd0Ia5GAoWG/GItXiKrH8h/ZBLvgCiXyP7byttQsMsV7+oOHAGc37DKySJU
2qznTZgO4/z09RMHcUHsbVq0pvZeP21sfy7zKHZcEefoeaeqEaceaqrT/A8NK1Ugk8UAGJR2Uhw5
bBl8pSDdHoEMRcgmlOAzVejD9GFsFyMc2K6k09oAYfWbXKd3dKKbgu7H5uTVAcykkhDZoHrcQ7cM
klKHG/b35VTX79RO7UQ4DvLsL67gs30hrIbf9IMCDoRFSqlLR3sma3jXMY0KaAlR44Hol8foHxh7
M3/m/dvOz+SthK9ohdDz2bKZjIQ0V48cZkgTyorhjf/WxP+TsQk+vo/60maYae57Lry3dgjQV4ES
Ting8YOksKtmFVuFJvHMAB+AkyIonR9eYYnwGlAGEYSATzNt7AIV60kk1T1YxOeyaqH2VcWtYWH0
vds3mHw5nMr77hWf09wm/FA79iiwfmV6IgwdTAOPJnnQJlfmiaFUzMTuikWI/7lQzWXLYh7SLiN+
T9NmTkAgnds/8w8sxvwqXeTAigcXBv37Nh0zZVSJ0vII0K1S5Ohg1R+8ydkPWzedHQLcvQ9gFU08
Y/Uh5cycs0iZD/t6pefmvn8KohmCO3UtNHpOXqP73DrSn45zgPwbOaDWD+575MrkjhEhAV//hbWD
UllekxDKWuDK8X1qf5bOoLuMhkrFRSjy0gFUU02JUP3u9ayeat9lvRe3gvheTQl+JmW9wHCRl6np
0xi7EN4DGIxwMd9dBD+HpthMQsOLrwJcrPAhN8Ej7EUvXDKK6BUTJGu6qr3DqE2afpD55inx62G4
WEvtuBhDHcjJngIQ4LcuJcWkI6P0zc3puc8TP4g60cw5xKVm7rZdmA3z/q8pMhluz9g2wgu4bQ5E
AF612kGGlMUHv2vfcXzQ7KAspgFU+leIWAz9x+JHxHvN0rKAxLDzUOlbVYC6Nw4NHZIMLJKCiSKZ
qUBimlwlfe4m6egiRO0J7m+wo/GRsUmkouhnDI/1BoLHqtCkc7xZrI2al5HLGDCWm3KAkn7Mx5bi
0Hp7fRKVVwZfO2m1BFoffELVAAmE69/UHtp1jcZZqvVzjvhVCSPecittrT4iO026ACCNmTFjmqlt
7TPME+cwBS5iywVDq69dqwybpq63iFlW6oJdSLagF3k1bj8DZAMayFHyK1hfDd87V7oMux16gsde
rWPu+vU1Jds3vovWB/ibPcMx1HpsPSGHPErAG4h+AbkjNBwtmmJvzHADS8vkl+apw3ijlDpAy3Ig
9NFvk3T7J+CIfBS5uNxCzhhInzyHsebCUtRUP55gaKKedyhMaZfX8MFQtMmsQglAYA+WLQc89oop
tz72tp8yOxsGJeRpJyfQR9EQouYiVbT8VGKtOR/aIaJL5EMvHHQnfmTVzK5WGjDNpfYKduiqn3/Y
MUW2vcOGK+ulrtps+u//hPeaTor0+pAXk59Pw0Oc6dLj2a6KY8gt0ZqnmXqixed/VqlqDVKPWgHh
+vBdl/vdBfj+de9+agKOR6UvLDGWrY0aX02PyDy3JOcSCcMJiaK646K7lmLmaNFsYYO5ciSzG3HR
2mTbukwuXnEcfAMOKGLyihuwvCy2cWnOFbqgTSaVboL317uHfzWQdYKtY82Ao0MWOhEbUPiWLt1r
XnbCVh/TLlMW6WPJBCdmIS9nOI8MYGbWTxyrIe/HCY5zmAFxKcHECR+Lud9EcKetOIV32sKl+dLz
4jG18TsFts5tPdWqWcMGxYl92IIEArXn0ziuQS9v/A0D6sbmq09Jo1IDOsFkdvCMhBO7Hyk9CyUb
rHGRYPmyf1aZNh4/qmCmlRaqPGkHQaQiYgRPM5Lm5TTjE7tIKDA4JnkFWKJYevbPlVZVWUAFEu+d
JNMYcbAYGyAWrvWylZoIw91dYuorE9YLOPIAEDAQNGKVeJ9ZKZr0CuiRiaM85E7byNw3xItX3nHM
UJPRS4fL6DATdBu5YrE97h12QN3X0gob8dgWYYyuqsejiUml7by4UkBm2e6MGegbeVNH4vyLHu1D
+XWaa8NuYi4TlTi9DLaBrOhR7nmkz1bYGXzKDMhZhp0IHls/IIXcbY3VQDIcpJnQkoDg8luCRByt
RINgg/9eTnlh7ZvSXQ65KgSIo0fMyZGAoHL3nyvAORP4wGtfab56gLmDJmshiPY2YIjlOHE1t8jO
dxkgJDZGubUrfKy+Jxu/8zF8Xf/3yzyBYrZTI05u/IDKftO8G8T7L8+++TxvJXTIQyhdSCCUvPnH
i6h0OlSHnFQEMrT+gFoW5xudnLr/6lKb/N/zgEJoIVxAae3QdMWT23+IpdJ2SftgNp78Upbdv6Cc
vwzIy/hJvEp0rdRtBf9HjU3KEi/z1V9bt5cnL09QNU5uyj8PqSwfjViG4Od2gNFsgDikcA0nN/O8
1869w1jW/DDKj0YW/y6Zq/Smuc7CTlqePOaITvfKOvBHFq1qO4/evR4PF9gws8kY7a/5jRlPFaAM
dg2brDBIiIB2qx0r4kc28M7nYGV5z4PrOLHpJ+vXtJr9aDZTqlkx29QB6V/1QWc3EQgVgwAZEd98
9IK2G9GmVu3T+GHNraXBU7fe8r7Rm7sqB4mSPAzDJFdEN1bKakTANr2w5/IALBwJKHXBbS6EfdNp
Fx9SJxqQlmlMwzntt1jH4gmn75Aes9BuN2acHykwrDW11qCaBZKKSX+wkZzM5bA5YUrvB4kl34uI
PHTwcL5DIiAACNvEruStFy7VPE/gJ+32pX3ZpBJ7EYynBzpiX5uP4THthfVcAbbSZ83GkF4MvLS+
GO1996KQBGPESTYxgBAddZjvs0viniNnrnfpzI/uhbCHWmRcKGFEXVNq1MAUiBcDkzMuZiaoKf6i
WFqG+vslctVGAcqYqcKbYlgnutSZd0ev8u1K+YiEaXvH71b+WtU69RFjYy333WgNIAsPYmfi+4rQ
ViSnu7Xtl2pe5uNuWsb7eJFgUjNRS4/aE4rJzOWvwIdqcPQpOxgNT/UwdsI7NAxcxxddf6nfbjfn
wMtYWXwgo2Lmn249eLDpqTcjDOXU96IXJ/RbzHRvXqvQTBLKDQShP7EsTaUNMJaPoaiWcx3yKpqQ
Ds2XGJDJWpttCjgCGgXmraBHMaKZNCbRBdEt0S9q77NWeShGOnjiYMND2bJxnM7Rv9ZfVuBNCBiI
JwQO7HLRGKZSYfjSMm1GxRgLQQDUjmYAso3VAyMSlklyXHQa6WLuYN8jkzcghADQEu2JsUC7B7ky
7hFWWqKukYCkAk0xaU0eJ6G0vCeJg93ihmzrl/02hNJKpc43K/aXlqkREf4ec+OT7ywxMDIplHaG
MzwFm9mHlDYsjPHstdraZ7fJJzjQ+JOZ79Cu0FQt4/ORhtpXYXVj0+2f8SdBXA3LshDt09Q4ZOTy
gKVrOK1yxvRHXsWO7BElDlpm7UENrpptI+Od/BaeGjdBax1sonSLvYjPBgfyzn4263dtUSBpwQxI
gmD5IEtuqZdBt0VaiQGpNQFUbHBwQAQUzhahy7aBmUwa3oB7rWbivNQHAaam5S7yYzqpcZNTd0+C
zvtB3qtIzkRsUu/V1712x4Xa7cM0FLGnD8mtlihKusUKFrBwJhxPJ35VhPA6EPvbN/AvGDzryEdR
2lFc4pPq0WV+rl8EVEGoziCSKYuEFqSwkx9BgNkd89c6Mzi1y745Gbi1eivkbNzJMFbxnJXR0KFg
irw9LXwEw1mvX6//L+68lpdGhRLFLEC3sQHSScXBSoVojQD34QabAjaZWQU52PqI2iTvgw+4r6t5
BnrnrlehPnEVxbIpI2nPNYR/RTUd4bTieXErW1c+SFbwVocmwzy1B6VBPkVs3x2uJHWnqnnFQ9WN
CP57ZbMeAzT/dCZYioShFxQDVEv9hUTFKvcPLQgXc1pqVK/Tv56wyHgMyuvCvwt3qNkuak9zIiBP
KNJ6nOaCseJ4OwLleFBuka4ojfFkqTwgszIkZODBR8GL9Uj0tNqC4ylgYyUpbfheZshvE4G2JK9K
kEtPo8i0b/kowbwg5cPFLA4R+zTMYOiyraHDYm7njRp6g8n+wHnfaZDpKAB8Tn+CGlWXJq0L1rYW
BPjHbFKMztHPmcuo0x9e3/ciP6Rx3foW7lnz7aQ3c1DDSUI2pPL4cyVUHCa6tOJP/NUVkTOhMMpq
gt2uSuUfvnRrEaQtcSH3WaeROP2h3VSZq2fr65Y2p/0La5x7cL2I9uvnIxlBMwD7MaQjiuWjZJFP
hBiPLIeD92rck6TbosxOUY0gTFVPIxR/boAIgDaVYO+uGQRQ3NVJGy/s0uFiTpo9TwJOa6JCsZHW
R1/ilDGH9XqVLOJcp4bd2Z4EULlra4STKAG9qTVB1Knlv/EKek8WZIZf5wsDZkGDQS+hN6NIt8e1
VhJmtoXrXGGi6wPI+HWmCzdV5vIM/IuCVBhpdOGzN/5RVT9lDLC34WdZphK0T2PkpCpII2hiF5xS
SpJfFvWSCUqI3gKroHd/ipe14dNxGgtXUgJNX4KLgKBFdWPW29JhU/cCpbaxuVyVFMb+dTAIPfvr
aPFjMLLViGrgcsgnbul/MCM9LSRtsHkyX6OfVUK9+PA25OgYutmVDvrpCM6s+id/8h+eUaRbAVFl
3drcPqJh5KOaUN2Dbv3GrOtmxralr+3mQVar4fttvAlGQFsotJrB1mv2VoHFJBkgZh1rKssntK/Z
QhgMmTlvvGE/y0DnqQR9ZbIou8NWgZpF9iv/yYgqjqgnE9DAC4tztMzLvGL771YUeTQ64P4q6ZQO
h0FiwQdKFUuGK6aMA7Hrx2TACO33X1/6rKWQoD1md+z5ad6p6FQeuJ8QqWzcJPC79jFqQxApUhmD
oEXgY1AKJP1mJxUqYjgAX5fo25JRuWKpsqmtzXQvb5AOfEj0pyYQjD5dPBYzNDl+0S6dD6wJYuUS
KBdBKsRa/KG8di731RbCMKZ1rCRUigkP/6plwjs72PMND4lYcgqsRdfsJ4idnaqDNAIIApAh+iiO
wbyre6voDQQcfOolC3CvU/3kcIaTENql5C/sg+JGtT1y4sfmAcT7DDHijrngFWsTvP4X0GDTXdic
IRdQJb3K8wnCcJS2RlFHukNhM7WXfGNgd/KKptcO0Gva3VXPj/zTpjmcPgeGajTzB5qgJPmRe9n+
Pf7Pikfm8gX4uhor2LEsWVSoI+0zT7ggAsxedmWFhoaojTc81ekZGaV4+QbZ8Bb3jj3h+4sjyQkA
Y+9D3McEYLuXqF2tcbNOWccBNhtZ3+ytncgLt/3oVoEoSrbCOrS6tfRvwYt0E01PFlE2c/6ILLld
IbldLUf8tz026PLGFaehsnDm7OSq8gR2agPqGfe8L2tKbZPH/h9CHPQcRz0hkmBD/ZGGjG+69I4w
1Km8ODzSIukxaH7Kh4nZ6F21V3je2pm8kXkD9W6ElYXJQwRavle2wkOKHYmPZ8WykV2jONsaJkgU
HJ61fx+6SVYUTB4LQHLuwhTokPGdV3ZJjLRiv8Py5pgsU/WlfNYCcojQkdyy5yoqVaQi8K1es421
oV3bjmOvkbBaGtOROJWexoZ0QxY9j2j7xf0PBCyJv+sEq2Q7bNHwj7Te1npsA8N84SI9WBOQKGkM
OoTcKmJb2zhcXiKy44CXTgTT4FVoMG4yzC/MB0s8uNpC3+FqjwqKk9YwmrzVe4jJcPt7VvWlpe/K
SFKRz7gh7WQyObX9adZ8/3llVFFuu7rbuAeY0P5TEHjsYaItk4RkOnos2duSzYfU76/ejH+g/zLl
IVenDlQpX/khAXll4hS2WD9d/Pu2PHSnK+06YFRIUsbDhQS2ienj/ZHyO5l1rkiZ9dJoAUy3AWwb
ZWlKV8NPWIpIJgG6r9W7OSlTs5XuELUhvBnoC3A42Jcn+mWWIzyllINe0rM081MhdJkODLdvlPYX
9S0C3wqUU3fOhQ5XFCUff7YVKjvzxcDWoyoILQIgJQ+NrcXw+dZ9W+PwL6U8i/RfKDujOV7vujMY
T8c/Dxi7821bPa/9/Dw7nEMFSSHLOmqJ4yk4aJ3S1LKp3bHkt4CtxEFcU0AxvKYRDWZjpLPKEAqv
MNF2JE43GDjofATlXCKDwdcraU6gpFG6qSaMuJjg1OJnC3OK0XIBvNp+1Cz30HQ36IBePwiK4OmR
RiiLp1kIU/Cx6NCbnkqNgAGLE4enf5VBpFEpNhpDu4L4g6FqhmBJ0HDz2WjNPKxMgi2z+aIGhMQe
8KR4SbWZ8De2w2uxixcSkjJHf45kP5FM6oHxVYWurIN47Z6SB4kQwQ9lvpI5UMOrQ1AUO5LvPKJM
94ZCxx9n4YKTgP/nsFd6+hKjt4LkgT4aif1ODy0VhlKHv0bIoqBwcWBIHwR76cnEvo1Gbezem0Hw
KIY+Lika57AhJaCkbQJF/jl6hy2vsZOCGHHDXtro3DlIdweBH0Dd6Cvo3G4HeJdlE8muTFs56r+7
hxwAv9QTCc3kM1hxqbb8IJitvXhg4y+R3eIzvOjpjKn1ggbNcB6ROUCt3kdhuaEzBMN8LWacSuUO
dtPFiht0vJmwcrXUq+uOO7zPsIsOplQoNmLiTCuJhDBb+3Pt0si89HLXg67o7GeuP99zrFxN6MQJ
otg7cVmE6zGXJq2kcPtCT4qtHR3cBc6T/igx2SE6qtexxFaqfcw1mz/J+HJaD371y4/OJM1/Iz4V
kGstuCOscBzPufufyhTcmjQwgewRyumB9EGDgz4gb2i7I7r/altwjvoXxmFWj29qn9+hY5CWgwu6
biV7OMskZzfSUeaBEAOjEwSFrGc1HMBHch4GZdSw2Q7otXXk3Xx7vUH2CdZk2AUb6B2B01IZj1fc
1tccYEN6hK5q8JTqwClXX0dXf/r7Yu5EmW4ha29lFZ94PKmcOEU2+jDeLwei+KspaG6ZUse6oqo/
hstqcVILbRXQ40LeTI2iXz/WgRs8mLlFXKTSh5JZLFi7LyawvuLN6gWaI3TN059BNbdW2+zvfI6p
OQ/41NBx56iCRaRcztbFqVjZ8Pd94311wFXybAvpKUL+arKpoQkNJz4tjzuwZlZIQpOl6dTLJJjY
e4I4ZgkzDQpeYEYqhwIRSdIuEZ77Qd8gRl6HlLNWhX2N/3yV5P4IT4ubG4a1Xk+dTBD6OMAM9WfL
HVLJ1s7JCDcyLQ97822wCRDIuX/4o3O7vCzEYA9t9dcTo/m7mVYyoTgMYJvUSrrFOTX/97aQIbB8
nnV2pYu6cTuNNlDsoY/8DND8Z7F60SHIpnMQf7dAGnmZQo5nqiyrAIoa42lXoubm/1X3vZURdi7d
NQ5xiQEZPupABh4KnzNfbYDFfeJy8kqgRrvDKmVaKe1usUCT3faJ65fvcKPCt9tfCjaNZ+0NLKrj
6eHnaqzwcDTjqKcbdG4oS5ChjRTE9Szy81yFVXxuUrOf91ay2uCZ2pMrFunDkHGN9wUlEzotJY1b
wSpWGfMYmkvg9DxRRZc7Ha17B/b6lNdQvJ9L4GhA8TmcqrsNXp9ZOanZ5X7+oaryL+H9AMya3IBP
ycixhiVUeNhE+J4H6DscweUiRzKakebh4s2VBeJamcRq65uxNJsazbOGtyMYm72ObwRYJvIxsjAK
0Qtyx/0XM89lwGg666SQIbosHZN2y6kdVEd3m2KJpUPDd8dvn9h1jCUhWSCZJZrvf64dlq7RSai4
LjeGGOsIigTKJwPQNEajUf3wnTeiDPOY1lrkbb98xMpqQg44godobgFcpq/ZffW8WueS/jaFAfKp
9vYsQAITP9skJ8ScaXHdxITg0B2lQPiPy/tGUAQi/dsBExfHJvOvDtQJaMoyvJ1bgo6gUp9oEM6M
Ml0rHVqgM4f4mJ4wNFbHjpdfGjTl3p6Jgpdjy9vjFmEHavMtJShAw7MD8asVKl3Xre+buDJIATIB
FWMpqckJRlMJwSqj2FfM94uNQKfZ/1fb1AD8UhR2Wm9OxyI2DHKCApor1yMg53kyt2MX1k48hbGI
vHusF1g1GMDwtdJoIjpMgHgCEDb8RSXfggPek0URJWmXEaMJnlHFMJVVwtfMmV+nJNF2iSa6Vg0s
Uib2h+B8VmywfnKAxXuPLksfUcxG8wjMfQWZP8p28T9W5gPl7p+6bLF3mjHEJYA2C3VKLhnGIZVQ
rB9Gmo29I3BiPeIG7StzL8OLpQ1FFEKyH4smy4sbQ0rnJmOgF90RWnJ5brYMMv+3mNWnui+brwZ4
bzcq4c83eI0rUksK1wF5RmZG9g0Gp0CwBLxoDrXyPgLoXImomHWRfY3sA0rvDcWJA+89LgQQr7FG
Tsr227LkIKw+KWubYrE/hM6/jbCpe8jQyhJFvYhn8sHkBt7Si/eidAWMgWneOQM6LiMU2GRokkze
NGHrds0cudv/LUrEqLy5ON3G5jGY3WUdvQJMIH5CL4X4PS/LDgm0bOCb8QNi8iyVk/JbSKjChu+m
5mzsCbS6U+dRBq28Rlcvru2g27/57OIsY3ku2rrhdo+N9AkvhQGK9NLq8vCWSas8s7XT3XQRFIT4
81YdafT46casTXPpXITv9uZtDfzjpBhuNCTQ0fpIT67f2S77UW0rwUdNBcdMmKV8viOCTuHODghY
SvkYeSH3GrRLZq/MRW6vBzf4DYz6/psj02uA9jz9ES9FTmdFj4EPcUfBNk27IF+7rIf41qRbdYaC
OuZwMR0YEIlfjDRQ0EFGsP+BkrOli9ocd1LSh7dcL+GGXTN5UXudfhg2ZR7Y25/4tZqU1gKmlZn5
a2V5A5AehqnpcSGB00QTlBdiztfav51+lwdHADmIPZ7cq3r76DI4kigYPcEQ8SAOwAAt2b2DAbbt
AnJDLCuLrqj99Fv5wT0IC7M3/+S3/8wmkffKhWL38vwfw7El/2SX55H0rEHpJiaD+U2t+RVtoD3U
gZrlhB3ps79sAUPbBvezitTsScqQ3wKPeERQoCOVZ9l5Fmo+JrzyPVM7cp6jIQanD7Ddy4nXFIM5
mp4V4l8c6MAQE8Ar9wPDoYBXQnntu6AYlxzvqrvH6UP8I2tF6Pji0brRAyQiVM8rYTjXx5jgLqsa
KPdY/P5slstaS0MddSZGzk2bz0CvOcDVKaDrX7Oxf7Mq1W5vtGAaf9LL1ETC5BiH9sVz9nPUJg0U
8Gi2mHQyq9ttyvr+rvT02CGq25gDP1ciAJSUxNmJC6VnF6W+1EbbCtMQOe1Zu1W3YUQiI9ZzJezX
qzyReQOkSQhXqvUSgO3xCZId5GYKJPSHPEA3KN9N63p5xABIYqThYYMypoZn4wWO2o/C8Fnbmsn3
SwocbSH002hHW2dAamrwBjx3m+N187XA4axf7G8mB1RGWkN3R171kGDm/CoZYXnZtNNWZwnj+aBX
c1zmXCZhGcTWDUmQhR96chE8qiQyy8Y9CMhGHuQaftig/oSC4qUVg1NDwkWCEz5+9WrUF4rIe+CR
nJ+ATWxyJxINwAZF208kFG7bY8tnTaDcsm/SmWJI5YV2D+OxjdFQHI8PKwK51nKD0DnMGTpbsts+
A9WymGCrDctdFd0G259ht391D4tM7C+K+Z5xwZKIq1D7v3M7kG6Og6yBnS81hINT3dvNnWUWhGbw
qbFaJQmdazAdgyMWUGuSQBdLSyyeQ0d0DxP+3DjzaB4ZaM5tuKRWVKYLP5msh2+AMsZmZdg+nkki
9gtlPXk1zyQGi/vuEEmxLBnydHwERuW24s8xS4bj4KAFjEwZr/mR/IOz7IsnRWMPR9onVHyR8C/p
Joku7NyDsS4RPFx3DaWY9WaiXA8pXwcHYoNSmufN8pZrtZ9BQnPFuWMfKCEfl2XEQLG6RThaBF81
VHetbG24dijWqvzk5Tz6YdmnZPaww+KngsMwtUS41HEqO8I8tjtZ567r6i3/pN/N81XzujZpmEub
uppcuiQMY1nkuyF6+8YZiazjlGYXSj+eVAsE3qefXdYEbd/XT1QxZpoE9x6WeKNanXwK8qwafkIv
A5QvCsuBao61U27SDMqmG6qVrK7UhptuCAxa6ch9MWQc/2pZRhi/AGV8GjN8i/ejCKgqrmadFi3b
1ZU8LfDJr8Hwa5AH3YW2a7bX/65JhdYFPXxXznz4KQaxZd16sSDx0OPDtarQN0q2mTw86XVdB1fx
SDepZSxRd3lJMII5ZLseskPs6D2Lzw8M37+mE+V4xy91UdOOScoEn+Z2eqleLreV34dTDYel1+0z
V+Zc+4I5legZErFmr8lOOocE4b3ZsuP2a28Sk5U9LbT60riCDQFmqmLA4n2wujSKgWzXagKfsNVm
PKrOl/IMO6Ll2trXy1IF0MF+DXRQLKQ/wzQlNOJdqwA7mhXi7nuT0BUFGTrmgKyoCbfpH4/nJSIh
AdsQxXw5v42f+ltxdYDBpgvhRO4PSwGAMM0GgasvuLTDL744/75SdsqPwQRPgu7wSlopg6GVww86
i9clo8T3uzFRP1WTrtocpTLW1EteT6Headbfb0yh+3VrRRrDY7kJnbwK3N2zDkJy8vaKyKAvYriR
tpoYx0M1cOdv9dwCcqK/Qz3BK7BeBUmh9wpO2O9oeVbFzQJf/tIp0dMwCLaeYRQ54v0DdPeokWCU
y9JRB6ycEn0b/AqF31j6oBBCnEX4+TzAyM+VCz3zKizO332DAlB808Uytfs7QIianLiBF2vB0Bbl
XQ+hlW1JnjJP4b5mv82BiZVMU6/u4N4xGw65MqZQHtyidxqDrlxUGXh/XFP+Nc2urkI2YGoPA5K7
M3IUM34+dWlO/x5KOprLHvC6aAQ4gy8CBJvSj2uEs5nMsu68szTndbndt4xlXX1mo8LW7qCM8TUI
OA11M+sIq5lsw8wlIuJSXs94OVXze3xnofbn/ZoIK4sNlQkN79aK++lXl4QWO+gZYlZ8Z8xeDEuc
4I3pTRLsW0XZDZbgil0XJ1rueF9CFHsa7eEfFLgN95oQa+OfnymjyP11jyODsCEz90DKihQi0oaF
YZr1Nay5lIR0tr7MOfouTzTpcsCI0GpXzzRlVSSuQmfu9hWKUKdNtYvEDnqTK+L2bs15YV41C2cf
cSm+shBygw63gOYmxXciFZvlR9JqBbujXbjSHivGoSiOBU6w4d7Vp0jBDD5Kc3QK0mBsbAgJYSl5
5m78vaIYyPirzAuUuA1bhSy0bbYDJ4hJ7BfvgR7xPkSID3RtOaJqUJ4vYrLdb6TiuxmG92scylUY
NkiarR6FrlRVZkECPX+OLCWiCFKN0f98t8F+cH0uYugwAfsLH9UXYoKIDyYelsgd8HHalZMVV9wO
3H4YMLc1p1T96NIT5vcnMUHpx0aH1a9zSSl/Iqq47ZFx2VWTgX5bg9XxxrPM8MqUh0l2GF8WQHLS
oWE8IpetT1CaaxmSjxNn3BStJefdrN0ZnbQyUgpEdWap+ai1K45MvUrJVk7PixI7ZluYXEWyJGPf
ZK64+Bul7I2bMpvtVaRKW+pCfB2gHpivudABRs/TuBeFWEm8I/7LdTCV01TyiBTSSuYcEOzIqC2o
lN1r/VUxlOhf/z8vP2c/9X08WSBqdrEqH/N5s8A882vKcr7wBV81JEyu3yM5lTXsd/6O+5eFOcag
sdT+439YtQgqKIcOIdTeZfQsRnzLi3HmMRboRjXka2zyRj35yiBm40Uy7M82xekSpKQlFBBEWQEH
pUeXf5xKBb5IcJ8A+UAa39VtoA4mBxYKRl+p5/cyuHGHqCykLeZXVrFR8+9iA3GNUAqlguJ1dIZe
i9gjpcIuxIs+vGVHSlNCICOqllUVMX3vugl3COS6JSP89VEa6+Xna+OSDuL+/jZUYH/CMserVNEW
oWJ+vU/KXOormQ5smveMc+yVmpSLrgA07IcV6pPP9Nw22kuRV0LpMLHkaXmw0D9BWAGoduQhQTeh
FvMr/XwM+n6ABcJKFpt8S+T4+4rOsWno88cOe+ZwY7T/+sTIRg/5FDP9D0dcs6bkndenSEBK5OxO
6O+lxxGk2TsHMHZ8056OL4RzrFmOKCtqxSGShvagsFtXDS0V/GfYIoEm9GU+oNJzi/m1c2F/1FCD
AItrobiqNQTJHC/qYw9OR7ETCBkIW5EKRIOLdgMvNQubou1u0w32G+Z8731b4C7MhcZZIOFUaYQo
m95KDScsi2GF2VvvV2Plc4W7L4wbEX4N7MugHjBsjS42ZbuJ0o2Y4v8k9H+c0XtipBvdexx/V9cP
1X+6xNlBursQDknFC/I1kmo6kMJX1rsK5OTGaxVzEg0k1fZ/uxgLgpt3jiBVCBNuzqb1VRTcDKwr
3gV2K95OzVrVsrPR+M6qBi4LVAiWFLzGNBACPPGtPMxmhaAc4LiKFNhu1wLwInYyN9cUOI9RS+K8
DH1S1xh4gAQQte3eywaYTohzqhye3O/2xZY+9vz+5AoOGo0QRRDiJAltmOkk6Vi4Opzm2EZQ8DZX
ZUpmaQ9LRUICrjWDZU2JiXFal3Io1+7sCWGVL/yGJuc5Y9CXr9DrTubUiIhfzgPt0qp60CKlK8hm
uiivXwJrT61Vjd/6oH+zHWEQK1m/tCvPktPWPrbn0fzI3ZS2xCRWIVNXZb112tE7upASDa86y50x
DfhaTtnO/Z1QidgvMY+fCIYcQNo3Edi86KwwF4qDcTTYwe0XddxY+NXHzVmztQt6W49mkr4uG9p5
YFMP2O4MCBoYLnfTxQbLnWydA/y/vHyJAPbHOU02+PO3DY4bd7LS5TWZqFSV21wXNgACdg90yhSa
Nu7XN/XFoNz9HOJhsT+4cXS5dY9qanEP+NDpdJ38khiwVey4ikeYvgUV+p1FfuQUekPj8/PInewZ
c6hLMzhLvbVwjNFxHvJlglmmkpE0blRY+YiDIQZu5fAKsccFjSO11jphxgYTIcEw2g4/hRIo9SPO
7GSNXeZaaUIH4toAB67tQhI8qPZfXNfxH3Zg+mdHEQ/XQgNVAgejzfnpkHrNhpJhGJ5ZLpvAWKji
i9B/D4ZRB6hQsrW8oaXg5dKLcNH4p8hqKR4V+kVcmnSRZ3O+hjMU0FprGn3BrjOJH3RWwKXaV0i+
YVR03C+XJI+z9WcH1KWPvFTUf8rx3GV4TnPVq9rRf/HbSjqJH+epXE1jp0UjcC8bGEoOk6SDIv5J
87mGZ+2BFp3/x914hc4rr2VQr7hP7Pyh03KpA3gEXYi5n0mLm/YhuUzevIoK7cbaXQHy8bYpoS7/
QTEUjtl6JqzwpcsCPJ7o2htgZ/Zq2+nqPwP9Ms4K8E3OInJbq2qfRtKtO9qFy5aFJmx4EKFE1oqP
7/zU0LnYjWPIHbOB1dftlnmtBNSo1jzs4mPSof5sOikntN9CKRhuA0vZb05tC1ucbIeOqIWm6Jyt
nhWgcL6rcRasYNYlbhtFsQixpfyH0mwkTEiI90RE5qx0JsOB9Bg9IFZNacd37U2GBCGUyrs5Y/1r
HCYWG22z8wXDAZb+GjXySaal3EqthYGk2GRVhZWW1RnHOkV7UqzhvlV+LynKiBkFF2CD14tBg2wf
+3r1T3/bMcrwyY9soEifcdRniFkbiRKgGfO58+/h3IJePg9EWD00ti0zgWz8d6PgqsPsBzMbcIhI
9lOmGX7dSoP9b7SxxD+a80prSbokMxlDY36n/7u6SLVq0p4UJS5cpeW1/TUoaiJk1hoT9FJxmq9M
YV3FABu/rpJLSSHDNU2dF6MmD3OJx/RQKoo5nowaujD4MGkwXAMe78J/K9pu9wvV83tJZJKcf+L5
W7jCMea77zRYa/YjFhYHHXLkY+rLPuRVDGonYhuN7HJpkTLC7WlWtlTNa+OsMd3xHrE5gfFK1ZOb
Fsab5NJbRVpqae4D+U4ye6APwks5aMbShNeV5tZPxCtZQUEyzJFhxpq3t79fxzig2ndJcAf0dF4f
oyRDz5tX3dYAFbfOTTYCNCY9KglCpc6pNeSsZVcFrwF2SHw7yeSRmCZA4KXCkgvDIVa5OOo0JNo0
NShcWXfGUTNzEUPhsjpf4ESXGm5q8ASR36oH4Y3/CCOgKl5dHS4KPpw7s3VOfJR8NYxR4TlVsQ1l
GppxfcFwCs3Q0M/Zcjsk21Lc9bb1vNwnqgOrVA8cDjIiwctDH5ShU9n2d+HfoZUX78FEWL5GKbXX
ovo0w0oEG10+M2eGhWygo80v4OhE4GzVoBD2hlNwok2cObF1UEIV2l4rCGKfjL9JrwrFfUhpd1GQ
8SuxW70u8L7aC0InfgKUMmF6ITANnKjDgkXblxXKjgTA2vWuQSReAzpBVx6/oHxGBChkavW0B00f
RLQJ3jnBj1f7JCmM8BtKCTw4441Tbd0ZLiXCXzvztR04tv7TNYYZNkDeGvwHcodFfYnUMg9BxFz9
zQIRj/k4n+EzKU1IKtLMeQuY5lJ6mGzwF9I85KXadMuCs6CzBb9zyKtRB2yeSBkTQBOXdZeVyhc/
sFI9hgpifwE+mfn0q+Sdo/LRf5BV2UC95k74tWoVd9kSL9yQzXq2aBuDYUtyJCgsQKmbEaQtqmOk
XQRAYP0jznzwd3pfxHYtnAwL8jSR3VeQDE1Myuv7T5+vbmd4VVmrVqlUN10mjaEKFD3DGPqZxKEf
L8oqckl2efpe2zmKjvdz7jXFebf6CCceDOMNjB/3CpSaVmlTNBYSfnFCJ4AgIWmyixEHqWsq6wDw
6Ngpaqa7NWqXu5lOZlPVt+VtMfk7Kw3QjNZpF2HOtXjAtQ1ylnKyVuutQ8X+7EPWtl3Ppt1670eI
3fpXoQz7/syvnIQsbmpBYvdSxe6wPaVfBC9s3TBnugWx6HnY7YaGSiLGsiZuDPFQP8Bp7HmFMLft
42TeG54bCz5jM6HyjErhO8L1ZzPniyaz6q8WERONmWoqPGXCrmjehpo3lQwqc76NmF5mocMmryWY
xAo+vq2j9RTR9XchACA/+FHHpkSruJDMfvxd/rQTIEd1iLXDXV4BXDyOhK0tevC/in3WMIiQiv6B
VfckqF/3c6sYIId/fsYZi5C8z8NwYoDTO6Klu0GRRwrigWBHiDagJdoxtrIQXOW4jWFh7Fjeo45a
Y8Ls8WFP+MkdAu41hKsv8p2yTnls0/Y8FxJLm5OlcJ7iXKipaHjzt+wrZXELz07x8HYNwJ+Noi0V
rXUdDq0rg+TGJDEy4k61V9DryoC4UXC9WDLgCGDT4lSSbQCba8G7NEebQn7TSqLHxwKwjQBteYrM
jPIW4A2zDXiiMFYR/KhcVbRHiHAn2tPSlKuajmcNKXQmnGKoLj+ztiO30hAqBaHW/MVOwa77eNCH
4GKNG3nXuDSBNYh5JXdBja8sHiZ025n0Ofzz9eNCTMVzfH3SzoxZhUJ3QGNMgGT/3qO88s8rj+Og
8lqSNQ8BFnOUEDeG9rHN5ejfe2yxydK6ClRCOCPvsps2HL6yPWCim4Zth2JZ2t4C2Xxquv8FiDPG
rS4HAUwlfyGlz2VBQdDLfzaueL3KVUtPBV972trNi7PoPMIgyHavllBF3RudSY2yGyVPAB8ZvnfM
3jZXQHRrPSG9k0zoudVYCx6vw/lNBRda574lFtgIdJkM3qOoxTHToAINZHgCQdmoCVnFyjZBVeLA
MJ53NeqmwcBUiLfM+DR9cuBRLKASC0E7HU2iCKE/NgdQtAmNGpH2Rc2UoLPmJfgyDeldlyZeDl6i
RtytDpTtH2T6cuf9DPXx4KWtb8IekkdB6XM1CKborL1aP/rHdjmU6krtmrnrAYRKv5zNim5pO/JC
/KevKm4v0S3m4kv3VFI3DyfrUxmcYMXOwPnZZ17g1vJTOPqJvNWfwwJRZt64qbJPypemsj3abrtm
tTB2H0/UI1PCTPzhHTY+HQM7/1tnBcrcTmetCAA/HkvDgFCa8MFuicS4pcvy+bkDuaz2aX3nGEG1
oZ9IcJb9FPH/5W+ja/85Hoq7N9CHW7auX9BQo94BknxYzpqXRX7fNO1K1cAg5NZsO38v/ZUWUwXG
NhZa6Nh8WflVJduZ9Rfjr/R3FP5wbJloAIaKtk7BOTi8rOoi+u3KwvULXc4jpySsQMajs+s1q3Yc
b4L6Mak9NOZhEx1OVzNgcReAjJGlBmy4l6I+3/TAOQpK0ru/mBrTDIHI/MNZDkqzCEbW78V4WIwU
cq5fdf3+SyTG3kwb6W4b9+n4oO1+hRZ86Hje8fqxeXu3OWx1ZKUCXYrQCET2JEG60EPKntJeelOO
kaTmQOkfOD52ywEC15rRegTJLzOL3LI8z4TzDg74AFrdDeC4PF6euotpULMy1M+2n2CR+qS1JoOQ
O0v+4UVgPAe+q4jFLuivKUWwbL8jL99TReCiI5Wf95B47o5PIYmAJn0Jza7eREinN6A8UTnKNcZX
mHjxAus3yUv5sqgBkiVTw9DeOhh9sGCgSmlWvJgIA2WVOzdQLEedcJFeUb7guZGnkzptAooMDRJX
S9PzxU1WUOzfodq7ZdLHL/VqfrK9MgLLkXNtS3BGmqdQhJHYAbIDRXjOulml6AD+q7Vuj1ZslUkz
0Rlk73nwdImPrR10ekVL7HEPX5mwkHlkgyOVwgssxWImYoblGDP2IsLrEDysDnL41TJiFP1OZa3D
t+zdq5MBDkJGFe4c/iXuKf8zQj5YDkSMPtNbJ8eh2ZRmxQTml5qKK9WDG88ZKuuSRsnS6RLxtn0J
BapVtNIWe43DyA+9bvWoZ7c6y2H8fC9bnkAD/x/tHpB4rmTIedz6afE3uNs/fb9Q5byNUAZQEA+v
ghBNyEZFxkJStnwm2TYliTY835Ut8/aHA8uIddtp/P5GBRtHiALUf71FalsC78Qo+iK21bTSIzsT
SyMzp6G2O7cWwmieV9QuO5l0dNZBGhIbn61O69iJb0GigNAbq3kCqys+cIkc629yiD6V8cjYYF2u
IU1JJxRk6BsOnzUAVVQmVMCj9PNq/NF/dm9FILuXkW34mNAgOwo3779DW9U9Q8V3ow4uSinxtlKy
dG3JjtzUEjT+T7uBCn4TI4UKrGpMcLEtlPzM4wJLZB1B2Ypew/yWEurrbHm1YtsE5NMQUJP7hB1t
gUbre+Ie9WZw0z2GZZZXye+TGLGzM8XzrHBBwg+ppPtFeTYtNb48f4cm3ihdVYbGD0n+hsCTZz7c
foi+YZ7lIi4t3JgANaCXyvvwro/oLDlci3xLIq8vQjLpjxVmAHE2AS7VDMAxFvwXp/z8HoDXSx68
hl4P01M6uX0Yaf/4TT1kN4p3S/0ETaJJM9SWkqa05qKpjUVUJ2X1QJIgcDnkIKOBpTvqHBM2o7xz
Q3n+DSpK0TbFfVI8atjVAHpEvPqmeHxf144xm5EWPECskc6UHQz4tY+4RyCvKIcWZZTUdtAZ2aYI
zQgukqRCi7wl+WRZgMKGITjozn1B2x5F8H2WtGJxYyU7sFkHx5CGnHSG35D9CKGNfUTlBJvsb+b8
OAUGXqV3Dv7jTLrXKxJud2mhT17yWmw8MNC6NRumhQAoQ6qkyqbnu/UXafcreMqSQ+jMuKe7hsUM
IXv2BAxknC+BYGpkt0F8QqS1P0z0t6iMialEUxeYgebtpGwh2kf5RekeD32SpW6x8BWbyZhOSC5h
EIGxK4AlJmvNKlc7TD+Qpon257HdjGqh2tKm1x4btimN1HGT+pdLPOVQwa1ZZG9PH6klA4QRzoGc
aEWQ1kbE/qDE2u+bp9ssD00d4h7cdAqSiZB5DxW0WdIr07WEZhS1cyJjyFTnZV9VIQvJxJpy9V2m
jOxBk/i5+fHQNlwe+tb4Jn/3577k2aqx9N+TR6v2DiJidiAr0NLdxfAKenNutJ4kPiWUMdbg1cHG
vIkxKmQ2KZo3mbW8vDsYC/5Emkf1tB3NSe9QWANEqLWlM181T9dq2KovV5QFSZmH7LAoxoUrJOGe
9zDSqOx8m/wFN9wrEiOzjPWADmfXLdatS8LRvlvj9NAGzh8Q1QDNk5b35RoZMdp7aD61nELZNL15
C3Gzd1bGRgWmcC3EQdLMZzQZw+Ok3Kn3ald8YZ2ZdKqKSa1rAs0pvEGcb6DVf616oXOTXMdRThQe
HHAUqvUegfgNLvW/uMZ9bknrjQJXkN5568k0ttG0Wr84jgu1Y/fIMSZJdokdz0AjO0g3u3yuYuY9
ycj4FjiLtZE9HRb3idaL74bCcNIgVrq2jkK3mau40l6j30uPMvQs52XiyN84Bj2GcNTgXDV6Hz5g
cYFfD6jjzKIhiweDH0rNkC00V2YSHVW1b06YEmAGVLkhVTUrhN8Zhv0FNOv63dLrollG9F/19U/J
5DFrBCCJ5vGEI2pExTWywJSTRqb6zxnXtG3I7GY6TfqztL9PD2cZJxmgUndzgBXEBboU7vMPCK+L
DLotGWzxOGU2P3JsNklOWduOJWmT9c3ncYdroAms35bJTriVx5sbQ8qKsHCJDlveXOZWDvP1s+v0
3DFes/f4htC9c7vpLuT7fZjAel0NXvovQwF37p1Zj4guDXD+kYsaEYaSvVof6aOaJX1rzF7tMch2
Xi+cRmbRpWlWOllEmZL0hvpXbboP305PjMmZFW+CUL5NA+nDwosGKFaoKnINaJq+eoY8/SbyMBCy
zdB02oaUWDRm6AA1oVUgd3YN1WKhPUXqLWOd/vFEnYXQcq8DmKviNGS4dQUkIrsJvGFHIVgLgkGg
bt5U/aHtldIy1+9MjCxBTX6favx8R4rM0xC2GsMQLHyYAV8E9cVQlzUGIERBkEffiLOfu7Y2JS0L
8JnBL1VHmAg5isYU91VKPDDUDDuC6rxkU8Nj8O5yasG6xICAgPojwe/cDFCoYh3phUW7dwX5q1kK
ThS8xpGiGWWr06sCpt+YzsuXZ2Jj4iyvMyUz4NQWbVZceq81pchVC9bKRuvjU57OWMKGwN4hddYQ
172X/EeP5V3TLsP45l7SFxJs1v5a0SOq2TETvd0LoOcxMFJShv9vyeXMCy9ow5lczXqeLjqFVy6P
hdqhx+VmzBqqO1TsEsOGnzGS2OdBto8DMMYHly6+tqrZQT1n+6n3Nd/o5W0RBCoFKS1BI9J2Az7G
nt4wJypgzzk2MQAzimqcYu37RZXsqOfeQa9TPUDWc7cCw+LFS5X5N1F8DRbX7M4fbKgn/cA7gs9Y
0C4mgXJ11NLGOGLdAIQugEMrn0AM8w5j+NItiqNf/mydDZ9agt97STQmZCo4OOV98gDofIysPLLN
4R+7TSUH+SgNR3DExwyz7YQfzWOSK6aMVfhGJj88xrxsgIBjoz/yCS1xwWesUGkXwZg4F1vRSiTr
jXl3wtcwMIsJIG0TvvsxbhNxpt7uEOGAnPigvKfweMNjYXVltX98SIyq9Pkiqm2X7enwlQ3ogH9y
xUcFCbL2lTbvkVotZckgTrkaYjJWHZdWSHkMR3qJyz4m0TmB/fmo0myjHEtUsywCOx48PCQDKq8F
YQJJZlFMpWa9VgFGkx5pK1C7nbRg3dtgIz6bwCKG2A1XXWphUK5XJ5kwTIS01ZimIGF9x2y3W5mj
rYIGBOl7BuHbk+b+rXwl+iOc++074UDPUcJcxhwrCJ4viXyJgCgbpPrzBf0P9Kecf5/kRZhai2Lf
HMtTzQucOdbPqhJtlftAax1B0ZP9A894+T0l0J4feULhBBVt+RnwMrRtrNTMH8Ff3gifTnnvgEHy
lskIhUIyojMC/6AM1HW37Jlax0cO7pEcc7jXzSfvkqxa84L0rWlxEwggGhigVl4VOp8OgKoYWQvC
LUdMFlBxCQIiAUu9pOao7Bn6XIA19n1YZq804LTwY/1bLOlczRxRbEftf2LKk4vNEs1fG4qezxuJ
7RjzXbWaIWWHfYfCV0CefQA4NCCQ3uoL35M+v8yhNw0Jjo0sBhagkJa4bA700oUlHr7+RItsTIw1
VK/4Zy/KekkWEksbcobyp/EGR3jyD70wX2tCJm0T8WDGScnCa6Fn4R6vUBYS0s63/pg1RJXWKqzr
N9qhwBNua3v9Z9UU/xdTbmuROgznvIhMVx5DvGJJV0+/s5jZGzxJ5khTtAO6YPm59ybT5Fr/D+Hr
VrYhenF3rXl7edspYX8WWQ5M25zDWFmhXR0VExKc8CTyBSCq6IybSWHjlnTVNU0luSHqnPBrkewF
K4XaH7GdoBRqDnRZhvDuCgFcTOqubIA6kcP1kefda7eaAQZOYtZPSqB7NnAUMVGbPXsqT4y2Fy0M
s67FERZ1Y/PA00y0Yl+EVcXfLFsRvcksZk0+Dp8HDpsn8zTO8kwNWZT/mAUCFe0GqApywr6bpGQp
Hy3kjRUoMUxg7w/JnulT9QjfARan79albi6fxN3SE+3isX1JujcCptvhqobX6RqKvUZhji0NOUul
L/U865YriOs9xh0kHeGKPNbAaTN6NnX69fCRtPtyeRsuFcNje/FPl1JvgdWh8PnngvS9E6qALMty
tvDy+6eGCsZJ8Gh4ZY9Lj664fZrPLiB0gfrgzrQZqI3WwG9CVJq6+ZY47k33K3FpHh5NWTO75oDv
YIlvN1g+Fe8zR+m1ujz1sZOVj/fqORixCa2mVrOzuKB4YgAnRiixMTye/qKugfqDIcpog1PB49Ck
po0+XP//aYZwlfHjiJ3vrau6W1VFIGuSNlB3f0ornpQt7c5UcMSjUphXDmnU2UKomursJT6/BXOE
V3LxvpNgkmPziTB8+U8KabsL97dPCLkMrcCy5Mrk1zO8xubWGxqhWXKaX29o4y/VmoVO4jqMfIST
ivixpzzL9t30kdI7exznVqAW9MZGi/TkJfV+xoCwTDPeGrwVdwwilF8CHc5p+MvA8pTfoFJ5/kGf
u3hP39S1Kd+q+yOjl5Mios53SnMazg3XkRSwSxdke2p4NP71X+cvRiGpW0twRzbFrc+ux7pWuA5U
0AylSA8GYpnm0gXDeaR67DxZfW9wBWXbRH/WVI6q1IBhYpo+5DQebvCc4khmCp5Q6u6bmJm9vTCi
Z8yCI21Vpeq7/BDwBU1XKx2hcLBCOAuUI0+/6cXONg7AZ0fDWf5z1/vVRLbkVIsFFju5wWDOljM/
nGCV7ck5ICQwmhDvA2fCxItbJUveipgDp682dvN6ObGnHN2rHlxcgGCt27M2uHSvEo334Ywu1Y0v
fDuhjBAbUZpv2T2bd3PlRU1r7YTAg6103pneEWsdAFHHvfRssymlmUvzM+oTnpaWZH6ilrL2EffD
HMRcnH+TjHDzee4FbqyBFGdfPg/N5SiwjY1BdtbhSw2a27hWbbwZGsYJVmlINIWIOqU1xToV8qy/
Y8/U78a7g9eDYIt+3tGJ2MkvvMi09AE4AsAArLmlGo4yID6bIi+w/7b6eCDJSwg1gY1goB+u9jKg
9S3Mywo+2G9oIa2IWjVfW2XXvV77IZUeZzxtPkTD80SFXbhWiV9T21fM0SilsTlPKPxenR7w2S0H
/9xppZxZWKxNYlByjRTCK4qzywc5oBxhKsNMPwVERqXg1hdJxnkO2UjZhXISgXSYJX2Ik0Vs82/e
m5IT0LnEtcg/xBUbJanf6cUu4sOcHPXXLPRlOYIZjG92rB4Ddi6sI7W65GrDFDBRUyKgIMf+2ljM
Y5Dz+jbHAxmxlCfb03jN+X5D0xVR1abJjTkXhl9z4Z3zPfR8OBxFQNTf+icYG048Wtt1zikzAOeP
gBpa26zMWT+bbI0Jlw92OVkZQzOcJZ7SC03DgcOQXuQcU502LkOV4WA2/RFm7bBChOBKAoiGZQQR
HRrDbk03wz0rvfYHLQakZHjA54WcWeDLTGjKDtpHiYCxTWLhu34MzP5D04k2IRqFZ3vKYpT6hVfP
1FIzSqzyOU4PdWs+VOCEnpDl5/K3+UxVRupYiUYmdxC+3NgiH/j/dxKKshgGdM/fqUUBWTKbyR7L
MdbI8yoiWf+dhoOw95v5hLFxCWXkjfv4LUMlR/B5dBTiNaZw+LTKr1mwJx7jZpVMAXogZUPfRPEb
HMY2w5T+RfYW/fLrOSpSHK/qQ6pxgxOtr1wE+IqWPLy376rEuV1lslQK9g2TM87SquVTlQ/ag9sO
WimK8WPqg1pt0+T+WpSnrKNw5dYWLwimGXZ5Bf1o0lSNZ/VyW9k6Ta/7mtSeMjHiHiNYWWuS7vJk
mKOumbjPpVR4DMoHIgX5F4lfKjHU0yHmXiGEYQMjHBOiu6jk+zHF185yS9XCCihwhACI7akk7gNL
M6WaNmTUb07Dsony5f8Szh2w5OoQRidnXZ+rHEs5PHdClSepaGtLQQxTJoVKqTtUHpmxti4T8urB
SzWL9R3MwuG7mhVmJOdW43+Y8/ogE4pLGalgVJi6Xp0fPFSzcBoywPe98ohIu+GfGF8sSRq3Y/ON
E+RMFp4TsTklhY6/e2KmKPoTRaGTTVnniZO7VSDwgYNrpcj1uDyUT5FF1lH1KudBENqbjmq3O2uC
d3Sm0tD9Zzmm8hQhq4Ad3U8U1Suc0z67kNkRZoMh2PraCyBvrg3TK+Zkwyw6gCJd6sP8TtgPGCJ/
OKHvkPQ5GNCd/YSdAptMp18CwnCItujJ+d9TmNvT9ZO9CDP2wwARrHet9ZkoRaqGplsOWKu4xa68
yE0kYNte0/bwXCP8IJjzJH56UDWpNZGaSXwac9rS9RK20TxGfzBANgLxkfBgo4FBqRTBqR8TDjZu
xiXipAY1NlzWadHhV0TgjlBHd6wIogyV2hy3DwoCWMgFLMvZVDxoec45Q9ye70PJSEO1STK/G5iX
86HVnW4/u5sx9nLbJM6wR5PcnKyOD8EKPYlw1QcRlu48EdwLjFUfE7bCyoNtvjfbs1XNPYD+3N5K
444CZGxO2bhQ+JUrzpj0OGA/Oov2+7duZRlFKZvTc/gMd+L5ZUdMTuqaKtgc6vyhd64nCxvYSf+A
vzDh3xymDcBOfF10XxPhgM5Lcg0Yh3PMnz6LAZGr9PnBgu1IjNKAr98R+Pklelc4j5GSAkpaQxTL
IwxB57m7zvxFXC/OlCl/XgpXXn55jG7J+AoEig2Dli86iUnUIpgCO63OMvKczeI9KgVhOZTTZIV5
2prbUQ8xRuxDLHx4BZHL2XYKpz59nSKKiFpc2Lr5t68/6FeOG9ynYoLXMZMAW9NE0F4O2QNvJEV6
yi1bJSJcfHb06xNZ10X18sw0vH6N9ijawcJfXfy2QL+EUJq8WH4OMtNrRf/KilYaJ7wistkoBH6x
yY/VJlpadf7gzkUs6PCduHhDxqUcd+zE261yu8l55RHEMAARYKHIyNZHtQURDFeFj2n8kEAS7isI
hfeWwLZSzHziQRRph32CYQpeks3NzfSwPA6cpt3cC39lssz8GG3sQREZRMKjdn2T9ct16hnbbWeZ
PWo2lVy0r2cHB29fYdAgR9jFcvSqI6eypbG9VcAAIsVgl60weqUw7nlX2zBAsfqY6mhN5sufm8vv
xvF2QoWZOB4rfUOFWdEGF07Y/u0+k9i7wENXxHGk8wviXuQwaQpdoNsNJ2C+hm0Lx7iCQ9KmMrHJ
d/YUjP7Ct9n1E+zIrMhmdaPpGCV7it43iEGpdALD53tD21pNfYdL7LSnpISiAdMlFYQ3vg0hQv5x
GPtZFHDHyyaZ43wB2KCjycSKnLa7KPhcjHSP92DY0zX4x4GpGSwlWOG2EdhDkONmiHCId1uZQpSR
JSs7hEsOoL1HsDJ1+cN+tUmIwm3tUycSeANytw9ze7lV7UUop0g9R0CPqb+/WzXEFAGpUruM7/PF
v4naq9XE1nIGlaAxrAlIuJYOuGh+GnIgN/gg0hnfN/X83/h80jcYDhnpp3DhBZdD/5ssfNqdkUiv
ty7H+JaH629eK+iJxGdED63n/cHz96dsSIc225GzWycNpLnKCVUQOiZ5mZjKHTRLO3zo2hSZS041
TMOogMkx0q5DZ8bD3Dm/DlliBev84GiwXQZcFcPqKYFsO3EDFqZIpmkGT5LVA59Kbab2AASrU+jK
rj16EhVbVfnE8ESQ4IwuujyUu9Hh5ZTccGk8brx7V1+EK7ljzHZN1Tq25iyeMy/f+AqTLw7IaOHd
h5UMpgIWp338hyu4bv7C8aJ7HLduxxHF/OUPM4f30lIb+6ifJlX5lilAxECx+F9pf2Fv2qY6hWwG
PAmCZTFVJO6zfcAePxLsax8PLgz2m0JvATOSH+pG2YrY+QUeUdSI4GfxR9hoCZOV5NYJuVAMSUFj
3/UeNJUxmr6nIoNybO6DNv2GUYnApNPcQdtwxIV5BA7qeNoPE4XnmOv2lVZnXz3CkVMtP7SbZxue
8tvCo7vmFA31aEoN5f3jaICLTTcrjqFCv/SDGfx7EQvRw/STild5ePYWph18Mux65f8RO0Q94wfi
WDvj/sgBNt/TR7u4/kACXg5vUTqEi4T1xC4mdm5jbT38o9rJwnGqYVHQtMvyHoFcVoZhWspw2/sL
eOjAaqttHf/NLZ/yVelUXnMQh7tfTQRuO3vBGuFvMfR+ieJrgg/ODFH/zcTNRuDVXAm9ATcjhu1b
A0ZQymGzx4K8L8h6XwXLazzP9eNpEHI3m8nWgNRwVmDQi92QaWeFINqcl+ejZgBwPTjKz2ZIFcs9
JjAOUxMtk8M1ylwc92hfiZGL52cjKfl2JEhZfayHDnWI1pJBJqhF490X6bRcFvWV7tzxVHMclisP
xhFDTR4BuEUl1XrStl0/m/my6m2l9i9Xar6sdTba4hB0XxEVSQBDQ+4GkXmsUQNIGL+pGlfkzh/i
bE9bio5BZHnWpPVk4UCk8BVLU8p0YwnCKeXAEoNEXSOx1+yQ7MgZWNJIPRLc/uIIbT4gIwVMSJxc
TbzNPdU1rcLW9cri1mLC6cJEEcU5NplzER6vP0MhsNIcva403taWa94+qMwk3AilYnqIeSBpear2
mdEaR1YZ3ybEaU5sq93m8OO+CqmlMlfmB7uZhzNpbj/rB4xCHBBuVorMsvAM7NWaQIX2311MWx6U
0M5HULoZqomO8USUWo06y+hRr2HA4qEP9MD3eb/wPuPnK+tSOAgqlVvADEjWKGjvqXZhr3uqsjgj
HC4WHdS8c0eCX96ZfQMFRq2tpjvp9r98/GX0xKIm+EHLHssRSCN9InskPq8aE4ZXYELZ3MwtciEh
l09d4IWtGQ3ws9/jCtw0YJ9sigbhYofkOKMuwb6qQEz1HUcXhj3HK9LmCzdVrY7oN5F1L5JUDqWh
NsNBPkJQtm/6kpBg07+w+MFJV4dJa4cb8OUWzUgkUsYKhCvLFaDzPwpnqpaDzr1GGDsZP5q94ExL
X9eB/DM04Q2USP3G3z/aMjvb3QeDKoSuAWeNPVLWY5Os+rNsUS5tHl3K6uAz2XiLzrAldNfXl1/B
6usDrx6Earhcz1KiJB87BU2giQk4HGtujujiqYI6cSjRlUacdcOt9uxao2mD67YBQYol2Jcf+yo7
RnAWlOGIZXdgAg975U5OdjQLd8JdsrxyjhOuurqAj2VWFYXHOMktCKz+li7Io968q7fpfHMv19p+
7Ju7zw03dLs6luq3thqFf64Ju8gY2YXvB9tTcHJlfxcKwGRAIn+3Rvong8w80IgEpeduA0P59LY7
aKrAVM77VpUnOLJs8AyFfPmjQGW23n3raShJe9cSyDmsDXXPCvMMdOdDxrAWhKIF5sgUw7Y7dv+Q
G+kLjJCGhJeDjpTf1fHuan1PQYgGwOWhuY6NTWs3kUn+4iyWiHNX9p1TpOzZ+b3Tj5CqDb4V/eUC
LoKoGUgG4TdBqi1Tj8bPhcQCgYZ2nX/qndI4DOI6LhdkKVMdenc6ECODc0gCNl5pE9O02YYcpKc3
dKq7F+bVUshmcO/FBcb3oKM4eki0V/8ASkdigD6fvp+nUDtrWCRheEPFSjpN3Ephjja1uI0KUf+T
2wiF+pYG+yZeq9rUvlbDG7/Auf06DaPxR5p8EwRQfrK3P5kadHUxpeasGDMaqtDfsP1U9DlAuevG
XM2zEzSxy/VXXBVkBbZrPxVTyxDlMEHyFAGPtTZTYiPxQyoktS/q9oNSDOTvfSGOxWisj9a305Er
vZXFRlJmHIF+EWoShb8d6NV0/RxxMzIhLwLivOdU7Iw00wYzqFCnUCtxHCqLsM0LdWZ7zOzoI3aK
1ak77d/hmOCfdveOAk03wR0vy9J7qHU1Q+DCvuUo0S2YYcMLQq1y48RVeEFh+ggOcg3ts00ULhTC
cU+MuttJvCDnVDT4WtGGTGgRefZVxNTcbSfsBhARdbQ8mFynGFoUG45CJiBAA69DO2/O1DoBmNfY
fRloeyzaKlXVZqfxGcCYoKkGsKpmKZEmBgQWz9UKNSVI9fRJx0Rwt0K7gmi7s5wpptnaWoGGobiy
XqTuNUsiUolDhLj+yiXYnpV8XCHwMa4vfynFJsJI9Qi0gH9YC3Unq9f/2GqhUH5jrNqQGIHuDfx7
VnzSq1lFIf8Ri/PKVhOe1o1CZzF8yiRaseZW8B0XOXU6RcxoXAoS8sJAi1qG4lxQZzh7VsZY0jDF
K0IpoQ47jb3cuA4eCorWJp8PNvTeGEKWy968Bqitpj7o3TrDswPjIlLhj2h1c9qqQqRGnrquMUew
oeksojV+VCp+awICMjWiXNG5r/ajH0/8AfqxanzFamBxCvdH3r2seM4uvOSnyK2/MpZbPMTT/fjL
IKWdYhld9mHTaXfF+V0wygNKKcy509f767/qG0fxRnp28A06kGyc+unm2k/GmxtERDBWuSi+t/yS
SYZXAdnOpM6dWLppenQzb7wQpINAAmQjtwaFtmT7GQ/3OgklvUNmIj1/bVgnkYIdC00CcBze7Jd5
J1/cj58oqEWAVFaSCKrJDdDtrhx1sjmYH3CiHtrf3gQ2HWvRe5X6+TMX1Xpvg17iwX877HA2ReXY
kMNho+R3e49SH8Z/tM7wx6lopfK2YD65OL335pCulFfhkbK8aKDhsHLhBWM9VRmFIUPgg2Mx/O3L
WwNChGnyfyuH0CPlNl7k2Yd8OaByehTL0XZu3x9pn8rOi3K6VsRWD7MdvPyEgBaWoS/5P8DBmulX
1eSk2P+j7RP5o3LlYOARpUQuiu54eJpuK4h9BC90ygxNF2zABKJDwdZxqfJ8KZAYpxpDcBDRspx5
LpD0o6niN2sxCz/pebaK7fptI3eW9GXatVlgSRebTx8NtcV3MT2L61r1bWpfCcKAMDTpJCeub+aP
SqK7NzcvcmccHhRM0PWAe7o2h1pDeAPn3kIxohEE/6PZiGPSm2L1mPp2BK4Mtb9jr7BhZEu2Klt6
sS8Y18sIn3QpF8Y+CRn3tXaG0mIjGzjCcnUKnGYs5Q+HZd0VcXitbIdUULX57+9f6yEpD1rMZyan
X9t3g7D79uh99z4PgPsS7WwqY4VVEf9hayCcjNT5f4Begckx45dxuozk0yEytqe2IAks1B1XkY5I
IsFMnon7cTyTmBCYBKh0xbmu8n5JzLepqmuw1ct+7702NJUx52/rTj7vY/AGBUUHltEUCS5e3LKV
eMjRlktRYB7sNg1j/M+2dS2EBVPKlEebaQbB+rt9nkd3VNE2meuelLWWAOSKEpPzple5L1+PWqIk
vv0QxMSDJsNE7afQ0iwTwUb/zbhAaNSyIIRFVRYRkw0Z8oseed0oGuO1XkA86U9Pp1rUCFwQMds8
6DKG4JiPR/4UBL6Q4Pll4J0Vvo16fa88gxTVwHVi1uzwtkCO4ej+DhxboG4xoTWEz/hLLeiE4nOT
VqEqLrM9SYhswZMw2MDaOJDzCWpSgqFwfCLKtRvjtz9pGQpTxjb5cwYt0LvNQfadcOMiVuSzwlgq
44M3etShIps466dpkIOKCMdgrMkLHlK4xgrvQDjKSXQnxXBpQxC0MzmM5TTFXAi7PUhUuHEvLxkK
MZIPOEqHk4ZFH5Zk1MJrj56m0MEeJuuPFRxvqGrbw3o1gq5+VcVc/6+BwamK2NJJ0d6LNaUbg+sJ
HpvT+rMfnWmCXOoxGjOplHOjJKlCnZu/bN7hMj+LJPYUAL67Dcz6qwzysZYDC8mS+w8umWhLebWS
F3FiYqk4SRFxKLkX1FuSJCXyEEmXJFAp/FLPK2KuGa6bAZZCO+J9c1rTNc+FsoP53KON4D8yLSly
vTOh7xxDJlNjlhOZTfDWizeHNA6ZmoUd+FeXaIeJYCfI1dBTUfxFFkPhTsHoE5e47ZR4MfNKHLb6
Y5Y7G23j/wflMwGd3WQjn0WT79v5K6Jg9ad9vISOcChpFV+Fv2iwo18QsFGNma3Kz8QdT8Sk/YXH
ueZtJSfHpHkvueWGk4PQXErQL8MbkJGm351TEgounAU7L9y2nVIlnXxboCvPWelKCIzcEzwB0Tbn
n+O65y88/JLWEN3UfV1y9s+96khL4NzwX3B+1GgIPRMFyn+wMjh2iEbvCMefYnulQGMJ1PWn4ubg
ZKWU2ro+UW5tiM9v9yFVTiKP37aCGGxZ/ADKTgzWdGFtZDxSqqXbTjsn2CxFHGloexXKyNcZX/5R
RDFFZZ1HydcGBsHB6tI/s5Ldizav09pgKl/DN+D0ZfwZLAjMsmb4l/WqOn3cxyy+/LCwHTBeLQBs
EJ+Gp7eW3xrAOGVOSLcds04fI47tAd6k3RQWlkHshPaSmlAm6pDs/Es4VXQcMaAbqjiX+QiXSysj
wlEsNqeFh1DKbCmA8jeVL6UT50LfgzuaOuAjqMqK01kdAmD9vlBB/Z9Hi7qNRqZYu7itRjq+BHZL
WCwRk8mPaYjPWklqeeKxe0JA8xBksQrKw2tTEUr2ZdIMFBC9zv08ymaRIJ+nhjjL7H9iQSw/5Cmd
B9sKlSP6frwlI7vFVP0yyZkPXGRiSL80l4ipZz5gXsJ5zP5Xb/6Xz6/I0UJcHEcXMpqv72atZQZm
/u4gRGObqf0ACL/gVPWSfO3oKDlni+/lMG5unYQMiIlix7Q5lFs87tAh000NEiBePoRcXoMVztOc
4bmHefYJqR6h0LFWNCDTw+z5nFDoXLN0AXMsJI+efvSPogEGNeBDc/ZvvU372BcjZ7EsFj8P1MaZ
4dm/JldftN8iCkcLyiCQqsj0HS0pv8qAM7kono1wFAVYjyT9l1SPbDhyKfN+ag0P+Bf52Fo5aB4u
MdT5I94lPnXybaKi0dUrHXG1k83p1in5gFaAc7MnMp12tM8b0hi7pDCNGnPGhmpaRzpFhHTSF8Ls
EjjNbzwZmoiV70GDoFn3jMuQGOyPjMqOjxol+PjUn4tnl2wamhorNaH0WyEKgEj7y4z/yJdfypmY
GV2NOswYfP1dXKqQjlARXxw4gAzSYgLeGmfrW9DteIIrjTgvhMqfrlp0caXlqOEWtyr0aHe5lVub
Z8vLf7BzvazMbRMmx6Yc0RsicRQa0/rvmaQC8wYZlKBf90Eym0QRm71zmtFHYf9Jhd7Av+n5SQZH
jLAGToKyqWlvov/fEV75J5WYWEXRj0gUwDwsBceA8WpHMc3iDdYV9AFpYbDplxDiiPVtXLsCcku7
PwkrFrF+i8iEIU+BITxHJAqcoW2Cnq7WBmAjMvEb95gU2SZ9WOrVTgwW3OqerYbZ2hYlRO4csFKc
uKwukeAlHWqc2iJ+lAzgFd8BknBT43RNXY9yl+1DQN/U5Y+x9DPR4Z7BBQAmbcVhlKGl3j1CzcOq
9PoUztybhOT7k6aJIkjjKqct3egbaRLQOtL+US7IE0n783zq8Xnlt3n/pTCJzH7DJnkh0wM7Drp5
Sa8bTp61bLIo947zI4fBXU8IdstpAmDXAKYt4Hinp/MmqNMFLmHmBrjbrGwXlZjJwPMnDX23Mwpw
hl8oL0y88jnv2uQl3/KXnhUU8KEZNE2xtp9Gy8Mi4WEwzGIc4+RgodN+UOqRDbeh+8P7fNLQZQ9i
dCJ0t8ecmZUHGukBAi4QVVhg3Ls+STSUzM4/jPXrOrG/6Rhu2g4+4Wa4FevaSJ8UlzQQFeI2GI4n
a5/TpNgUwZrZ07jElR9zvRqVAPxq/Gu8nVYg+dP6JlnbnrH7CY/Ch4z3GIQFZlbF1sNXQothdYre
IBNxFuf/iVqjakvOrRU6q6KPC8Lrouv7E2XXfx8MkVwykQ4Ml+qw+5vO1+lNKa1sEAlkkRPkjILA
x6ns45KweWJG94JdHgPyhXcM9Y0WPiov4zm1peAKgMbq19gsJX9ekh9VKwMRzIKNsIri0cye0Pme
mWlF/zUcijqkmJu9SFFnxsMIRufYMrZMuAags+2l0EF3hfvExlw5Yv8WaaJr758N5xKySl9h3ldy
pB+Xd6kejA0nivvk2S7UwXa1KGRMRLRVJ3TQ+1BIlA1WpJTDvJVzMG1NIKcjrQq+j4+BESczYnFH
/+GTt0bKENQ0MU+Ow2VygXoZDmUn+gIG5AAvdwZ9H21Rpszem2IH4mm9yH2n53PkzZW+WHW8XlzF
3/zkC0tuVrUrFKrZzEdx7X2Nayo+55MX5MwJttvKd/TrKeS0Nu/QCWm9na8hAOllESNS5q+CoaY9
x/lQiPpmhCYpbgTyCWMQp9OW8xunLkc653eMJLIoelG0FpKXSmiRpxtUbK9wp9Gs7xJ8h5L91935
ty6ScLiOrJP16HzHp5XOzwt5jNzrcalgaIUshroNFfhdD/9WnjePxIsPQjAp4HFdNBFbwFS8lYwY
+UkyVSxLcWcLvfVN50c5zEW0sgOJFCeAxsug37oW9qR4PVKLHXS9GZyLHpnGwBL9QFgzatbmB6aQ
RVj9WrgiRyKT02t4DOsnrZckZwSoFQcQn5Gvr1VrvszRBboRk9MRAzBLnA057ZtN2m1dt5IwNpiA
b47SIUdHoeGf0hlJJkKOLWhzieSXPitFKDXVfhlvaCJUuvWbp9eMQX9LhLQGrnltuKQPzgBoJG4g
XxtS8cb8VFbndJbzexkdClKk5uUYRfhf3OWUDLhi9uH33jTKbdvY9v6qAGoklAyqenXu20oRG0mj
Tmo0y75PL1R+SzqZ3jR5VaWJn3g0jDO+THLxgvH68lpkuh3ISaHRwfz5bziiANj5dTbeQKkdJOs7
07UA1aUQh07RnqtJ3MvkiBROTG5t5cDZFtDrXWsz3ssM0SGnXxKE2OgY+Q7jTo0fQ3JCVO9C2KwO
onxbCsFWcoSIkQs3uH0VOu85sI8pDRAYzmJrhIV438hxJYZfOHSZtIUQ6UIfxYIFHjnSfSq4WI4c
UerLumem9CFloS2acSTs+S5+aTzXUjA4jmnb91W+5mOXL3OBDP7a1hrC3u4TCab+ZtsZGOUUJIyD
XfYvM3BGbK69MrPzgmWz63tdpIwq3+7ehPlhMNhlYSZPL857uBhCHpBYFmDM5zJE2tx7OrquNhcA
MjaveKtoVYa2ct66IGetFC3PjyiyDQO13XA+nZDRsXB05S+/8xEyvRwLuGOEdvYVoTQ7R3hicGW0
M29hIxmLIp4cj/NQ4slyWJSeccWG4LYagrxS92MjExuAScy/PEkLnYaemKGxrDJNluCakXp+Htt5
8qam8U3alxkfUkv5EeoO7HmiOOt4D1Yna5NMuj1X9iit5ny/s7rUjw/BmPw/APankLmwrwhV/v3i
6JNKAMYDf4b1005Im0XbDkoLX8sE0Xb7ohFtToxY8+SCJkDMZZWdhs4YgUcRHkIWGRc6ccIiiyRL
LRxLwwpZLdfx4gog7SWl+pL+hjRA246RS+PsgQKyIqnou1Lgk5eVqTk+q7SnokbtnRWJX/LAr68c
Z9DqVcENvONjHFjSoN2BormdkmenQM2JPD4wTwrZwgNfo4FjfGe57CWKwwkKnW7kQcFJG5nLm6NX
PlAw4P6HX6fgAKh1Dx/ZctoUAcEXSVxAjv374jc61gvPNEq7I/7Ge4dlTGHe9+GOMtbxR9TflelC
Z7hpuGDR78YfBP8w3SGzM7dc5Vwjvm5rQdKLkZHqfXDCHKTxIZAZS2yr3tzRt/Nl5CzwdQhZsfJR
K05/cXQNcM7Wf5W/ahA4oON+6moy1mBf3zxRr7jERwDnQqcMmZW3KhPGmKR0oZddiXmBhVbZJvrE
6yG3pXGk7WXfqzFDcKp8r94Z1xXN95O8+SWfnQglyZwwX19y3wRaqVU5heYUpPo0hfHb0hqSXT1B
CKxmb6oRTAv09fDxuwsfAqqKPUz4sU0ruy4uPvhxv2Rs2tqtfNsFfc4P1/KjhHIs//uFfhTq7eyt
naw7CQCslN80Qdu6CdwWZ6guG6Vt8k9RLiUGDrtT9koGZruXVw+jlJyQ9gl91M/wxhguh0BRD8po
yz74cZdzsAiNq6JIclPRzSLbUvmdqwaznxejnBPz1SA4PLz3VlDk0wHQXM0j9gWIdO3PO8cLbjmR
OJVKoHfdy/DtzlZBJyNVA17kvG71NEGlYsIo2FlOZ06YopcuXThaQeuGd6aUPx19wx4TyqPXMBFV
Fk85esib9izejy5OhtuwUWIf7er+7sXc2B4aR+AIxKgk8xJUc6eF/yNSZo3Rzg+fB4SaKFiDwcZk
j0r+WGD4jU+FmNtgiHF9FkBpk7UCcOZVc14Ku3cCjcmi+5MTjgW80RPyHYt6dEDBjqlsFc9NINAU
MGsWJ6aHfHMqWABRsZDoJhpgLhPYZQneMAqjtSIImH+0t2+GJ0NB6TktoipQofvRDgHEfwx3AHGG
HxW9I2pOIg8OQgji1jhdaRHxjI6J8zDV7MFWdP1vB/57iXJtdxDaqOUkYqQ0At5ZC1405lVGWtbz
7njVZMGVjDf/8snxCcbjTiLJf3fUjtQDr6ev4P7xLQ6wUl4FjrWfnij09mmWYKz0hoDDilzj92HG
31kEODYpwAuYvvUdtBQfGi+N3cg1poFn5mB8eddCX2H/KvBPMQSyBMI8F3m1BpKUnlpihF4YXzuq
750yGiW/fLRby445gFqmOtdwAFfsKCy4bWm97PUBmPOD+YmyeIBb/UYTO9vrOI+8ch5uHgs3F/8b
IyH4NIUHLWUY1AwsC00XXcTNs+GbcTg7f4xHUh3rxB2DtuTYKRMtFB5rXXRHK/JYrHSQQvksSAYK
wpPwW8c/czqdjhSQxle/YMrUi34ETtGKB5HzNuwweXwKlgd2Kqqg8KMUIjy4M+KnQ/bvE3bYbVrs
64366gMUHgUeUnwUWc1DQ3pc0kji0m/HECyDqWq5fp5leup17CU2bCpG+C14Y55tNIIVKX3dio1o
bkbCBaOzlo9iZsVRpdt+1+OhJPOKp/Jc1gv3JPDhzq90bIeYcayGXpW+iTwBk4AoDXhrGKYjP8iw
83FnPIZn2c0AfJ9pJi+w23OihUUhSX5Ez6Chm7p8U7W31bqG3vMwEGLZQOCWn3f3iUdMhfKJJSBC
V4rpeLZwkq9MmVDCu2v06BxQOow1+Yr7hn14u6yCj1EBtHTwwKmuxeU+IBY6jwXJfUidfm+SE9XW
CegrMHe7szuXU9k/r5DSjed7vrtT4WZSoJOHm4vTiFZ0PsICEpacg/knWP6TLppNdKlqVBShS5Jt
Hah37+bPTNKKyOZMNlaCo1X1fr6tu2Z8s5ME3oqJs/EOWToE83xGEvk03rl+UCHXxcB2N0/ng+4k
ZqH9Y4fTZcbIgqzAuxGGwgfdbs9p/URxrJgdoOolZN1A2mPOb+LyJtmH1NJ9HWk2mdb5jXwE0ySe
694bkkrF/9sOr4/KNucQ/54dD/F3IHa1zeVAI9DjV5JsV6oe8e8mjU9QrGWz3BPqqjo4SylUOFLA
0MmRmqYqGpxdnIqq3UsHa7VE3nhRofsq+UcwhR1OQ0Wg7RRHrM55Bfwdu/GgNmSEswoNoIfSjrN9
zZBfPOsEKYrK5Yld4C7DRDAnhfYm/eZXmcBnIgu5R1PBoY51lBq5tE6yY83aCMBvzcSfdendKyvC
6VHZO5Nu2jKBr5YJaueCVVw25vRT685mB6O128CBla+w36tWzpi5zYPVk4GYAq6wP5Nrf1AQ9YUA
UEM1c5E8lMSnPiMzs8FTDX2IJ5cTDem78nBb4r5/tx+rPHn0M42CNJ7JqKzj6o/Rl/a26JU7/uAV
m7SzpE+cpbT26XKemcrR2ZEVrXZ/rpVU/++xzLmCFraXE2FsblxwN9D6eB0mGnQVxqCKTjq8rWL2
MIgz0Cz1fjsuXi40nhbBh/yIAj5m4tNMJ9f/gHeZxKob4lZCBV0ghAa9+smi+pZcsS5e6IVt8P9s
nZ/Vf21svJ1RFqXNQ40HFJ/UE9NebRdOv8PHmvlveh3Z1orPkLTfZyt7jbQ6D9WYQayGYrAoe1JO
s+5ud6UGVFlI7ITS4O2zjR88d2KIvg78N+pui6eHRF57uowCndJ8PbwvIfRDnzTNLv4FSDGXijbI
xFsovr+vrSuBBucK/U4LLtu+maRqkrRGLQ1QgoPRjNrswiZaW1uzxgCIcrcZYOdzHaEPgWrB5670
pIyIskHUGDoQ1KGe2fqqST4hSOAiMlal55mlGd/kmSCp+e/UnqPDpeYIvyPRm7VpdEtFcC+8HU0M
3a5yu7JFdrQTbl7K90yf2MCuYjD0FaKpyiKNrqvCblyViPF2y3RMyMMlSlSrE8yxoEjhWylwoXd3
IbkVGm6SIvThVImEF/1wkbWOBPg8D3nz7GgvnMoVPAHTwtpoGf/F2nbR9Ia3vnB6QTYdhloWwHrN
JJo3CxMc873ZFQr3Ltbh7FBJ1IB3KcNrprLZPrkrB7exqcuxqkt22RgmA/J5bFRJa8vcLLXLE4kP
AAeSZRAmcbiaG1xz/X7NZMXvnW8KxA1rYJI4C2T5EyGvg3CA4xJt0OY4N0iiNBLYM1YXjKmgs4yb
MnNVgpdm8gr/Eg9GCPkJHuUr7JkpJBz5voB+E9G9N3URBgd7i2LaMe2KOBnJ2M5GTFUX7Wqf2neI
Xa35gmrWeGUL9JTtQZ2q0JBgC9t3oOogePTi3f56A9T8J/usxSuAVAVG11z5pc/ZbfeVcViY3NRG
rB6SApkgkU410wxfD/eSPWZpF8/mnYJu7lqLxVtYNeJsAuXPr874LUxNa8nar8b4MDq7u/81UjKK
/rBvP8IMkDBYSQJ4hLQO+sAhMyxNkSHC1tCtpdnFzVGSL05xclTpu+006AdXqRPdz+PLIjagj3yN
1KYqCgsvVa7vT+vVJu/Zp+NZIZvSb+VVsMFuKChloBtRLaMupMmWT+E9vfand6r7F+LOp6t6jZGq
GlJppRDij1oqqp6WLfNDG5xmvAOYKERtL0M0EsojgKXBaH0g7IseOCMYtK4s2A7sryMdVBLGFcyi
jGf+mErkSjsLE/SRVsoum64FzcPyPuhmt4yyc3gOSXX/Uex1c051h+8J6yFClfkYoXJBL6prHADn
TM+yOKwM/89uHwVl+PFH5qqEdXCe3E9sOhfIRUevlhkhtjS2FLU/ImMwaEeIsPuyVfAPxl4PZsAs
/qRpLLfM1THzo+Qn7nttQ4M+pz0lN/1DigTTTWSA9TtQOhGocXP688sHhSnaWARaEJtmfnsZbU4P
oOPrRoGEL9YGIM+vwMVpVfTCUtZZtU58O2w8JMmWsmbARoEvAXNx5W14o6PQkydp7pkVoLDYnKPW
Fgf8B2JoNWgyQ9TZF9ouh8rCY+E3zhkU3m1fPY/vcf2BjSK8cE8US5Ahe9xwjiB0RQneiTXIXFtB
AEEt9PwDIUc3Ke0tlnBqbIG2x0OgcLSOEsI4iG8UXPGupk0+FL6+nOB65KrhZ1kWoBHKkwWIbjYX
vDzdVFXKv0/PJN8JJUzKAfPy/adzAx70zBXA/NQifwFaxzdAjJFkUh0O4v0LWNR6+gj4eOfC8bZ+
WB21/yAsnqmMm7V6YyLHZIdnhnXjbC69apwxcqayRQ2wqzQ9HBGgm1RV+dJSGEPu/syVhPQzRVyW
B5Diiad+SAZm0XOJ0xXoFjSUEdZx+bCXRfgD2HbhynsLUkXJonsbaJpm0gu80fsCfe8cFJoJIQ9j
5YQtUf3au9D5tFFXP4yGghFU8QqFNT/SIKLqUHC1QCa+cjuDz6UlN4a50PWGdNGtT1B2gVgsg1q1
TdlyPgNAre0Zu8gi0O+8nXnGkBqMhMaH2qpesBp2uzcvA7PphjW5w87KU/jzq1Qt1qB9nsV9Htj3
lUigmGz1YD7rh01UEipPxMIBdnEY6uQ54gzAmPhvweZdC9+ZtGqJcm6sPdhGgxC9DgX+JpW9F3l5
CCCYqosQ31qUQh1KSNOG55yf0tC9kDO8tnid8itqE/JJV3Ca3ZJRl+UwgSp5xc94wicgFSXwuC3Q
azD6pSY4/NyiMwBlP4WCnfoAwkl98CSwpp2dUOfsEjmABUQHRf2Wb2fw6qv4Sdu63PCZBbt7+1t2
nF21/XMd6QlYnttIJPCaJmES53nrup3cpzgzQQXR9Nl+E92EryzRFKkyE7EdTqlPj/b3ro+wsE1r
AXb0JTejQVBXvvap4GbdmJAlJeMZpX4nrpfHtRrKfhkTHw3lUb88YeLgKi/IHXbsK6/X58Tnvv1R
j2gPtwBlhvGSguvJj0Kz7VKq4JN/zYWyiD3MPrR98tkiEp7oJuDIGsanmZXK5JUiEmEISW/B3N0e
G7YrUXyKk9Bmfoi3p21T3kTp3mlx6Vl7iMAQ94CxE+l4KDNt763G6BSLju0LbZakRCNj0GpQ2bWc
fLw58tAYc29ZZ3f61xvN1NJlHDVn3Jra8Fsbr1bponhm5OhH1kej04sqoVDaTvRQGSd2+AEDpkqf
jUERyzaozN9YgudKByYEoEvVrjFpOabW767KmnfEdE9xQMnya44UoX2RXMAT5x1cLHz1iFElcqTi
ExAF7dq8XZ9yoPE1dhtiBwtlm3cbKMDE0zDRyLIPUm3WSwmL2zvtzmY3e4LZ+aVX+4BH+XhN19EY
Sc/f8YaHJAaVultamB2CAsz7PMEiqyxhrwt+4WWC7Htxrw1TSPwNyGUkUgl3QX2ez2dlS/AFlUl7
o82yNuXfNOknDR1pESV84iwECyameujw8kxk0vFYajGsG0GX7DZJtUVf0Ir3LWupLML9kKCcO9jQ
bUIqyIuLrKdZqvlQP/5qz0JjOS877p27syQkmReDABe9xiKrTT0Ggc9tNvjrKh+DSD+NYYNMDIGt
4aFM5A8F6kT8sq0zpNjskOsBVr2abxO8I74ODA/MvREFPKqVBCe8DHirBpi9/YTIyRDrrVuHt0gQ
sfFtILVpFFYh9m3cZ/GAPgv1JFBDU0F/yZhL+uqhQm3X7yw/h6wYUdxE/zb+LfSm6uqCGDz5T4GN
fJ1YW3Okf7npedlejIC7J3HTV0tUEsEo/2cWrmVklZ2Ov4KhoxblFJqsi2kkCwdn8QrHMXYPN1ZN
vsRSROrdGzjSeKpoywDOiDUtEb6wl2ZZpsKf2XsxBy2D9hIMTbgCpDsgDOy+4BbbdzBoizFTN5C1
SyAq+nEk7EjvJaYoFxg++B6O9inRTAjFN3DzCI8jXF2M5ZZqKmMp2j9ig5qOnXzjqVXSqfMoJtzd
QuwhEGSWHbbbV8zwDJ8WpxnzXOdRBMYpXnNEEcxBXdhk4riBcdRg5kXDLL92UP53IrR3yKzU8jv5
GImR3gOMvKHIsBras5s4IFWdWjdlaQMWU2m1OO8r4aSWIKMjGJslqY+GhPrBUbRZKfEps/cyumym
8BggUEpvSQ53PsaFVvjCDOlGLF87FNC7/UxXAnAoTZG5Fg48uZSZrZLa2iS2ICYlVcbdkvlZJJmS
tIltXqa3n26QrkGCdUDwKM4zqwQvprZR8YM5bNZcg9UKZEH8PJ5wH/fLwoF/FRE1ckZJ6M78mz1c
MDvIAdPwX+ZAcPyRKKvUnr5TtGNx78H/9X+Szodlv77+BwY9COuytwf/WRfPUmbrYHXwpVA/7YVI
pY/IqQ8IFAUz0nGyIjHihkflMV0L9cRt6QhgipO1L49LLeogL0VerMGW06a9nsYGSGv2e/N5JeT6
nAuHx1JhEx9hCNpPUB/Ng0J+eeI3e9zX3tio51za7YhI827b1hpPxAFVju4R+N1FCdeS4FkDUeen
p5AcgCaxIAw3kq7f2TB1BlpaX1N5xzsk0BJcFmjAjet7wYig+s+2OEZFBpm+zUGqfsbDdCyhH6G9
oOFDVAt5zbig1vXjVh371GB9ut7ZK2MEHzAUVcJnMHnAk5kbeWPDSNjorZ95nFpv1M38nbvDBMhF
TeUNTTC9oFYJukrTZrFtNSWjpeJ+c5aMdxhdxLhm/CL7mQtd8Kf1toq2QU2AMjiD9Q22U8ByaxTg
mPzTYSD6p9TLQHCKHXoAJsAQtCw/sM3asjx4wih6MGyy9+Vg6/QUZfTlkpaDpAcXjgInQQSex4zJ
EowrE/jc6E/Bpp8lakN+yNEDEm8fRrVB5Hs6Y2l4O1qDI55b9jyObyWsNt+GUfqnskWVE0BcNGX1
w4GaGf6XXCTkjuC1Afa971w4ujNUQPucusGKoEtx1lk83E+aiu7eWGqqhNF62JlSExWgUXNAlthh
DtUIA0cp6v559W8/kBihbIIKQy6P24YsHrz0oL7qAROBscIM3QNlwhsdaHyXSUlOuWSANf/xuvir
T52F0mlxL99IuleylWwyVX8/C7b0i145ch3H6SZQ+mkPkRxv1+pdgVPrNRf/ojrfRT2kM4ejdmSp
W9D+TCmSCD4KtrA4hl/b+XDFZfodw4gzfjXlfwt+MQ5a1Og7jbp8XxqooKVqN39XckmFkVCUkWRW
vX9b6icy1MOTgje7IB0vs3JBrf9CQ0lRW/usF/fxsYiey8t7DEL6Ghrp6GAYnx7mINVd3byENJ1t
EaO3U8/DI0sobK7a+JX/U99wQPwJyMIrAewJBW90lRQ/4YbiOc5t/tO19ehzQReZ2VGWH9GTn7Xl
s2sxWS1CZ3njl2L9EOToB7aOcpT1NlE/ba2IPIlDBix5qaeiqa1zanYQUrAVGQ9UzWlhDFPAVSDP
WUvjtQb6YCnnRpJ8jgvLsWzls4U2ThkoxPkoewvooKQ/2Mb8LfdO8x8YkuzvPbFaKmBMKLrjBOmx
HKFyboJmuukBTqOFf06Nh7JmScj/7BQZsSUSNiSzHXNngsnBlW3eqKRP4V14R0NrsjyzJ3F81c1q
3W/gRMKtld3N/k14IntTsdwK5V4JrjImaMzScL5/ZRf+xGOdEsxRxSFxoWiF79ZdpVNAnRnQUhuv
tUBm/nY/8L7MoRiYilBqa3jn6uwNgiDNiCI5ksv+FuNtwucBXphgJFWwlPpi4YHacUwn3/Jey/+A
qO1C2JT6pYVpd/ZsG8f2L8fKJF19ptxDu8i60Sj93/m6hAnfEj0oBtXcRG4D5e5MnOYOq7OffDj/
bvcwlqQM+Tu1tMafjRPzdIFMNU5O97fsi/+aLRcnVyFaswCDg6GnUg5AuglnBx5naeGNTYhizZmo
mWEe1fTe+XEe2zjD/5RtpbjPa7Om8emCFpcDEe0RQ2KTEvGw13kXRCZLaToqPIEKzKvSS+kzDp1C
exkdqxkOrhW4gMgPjYuOh7UTthAye2zhJCMYz2raJYXhCD2EhYNTxK7HH0+r4bvwSHxLbbkiv3WL
Mi4wR4Y6GUikXByEkQlFbifGBDXKBzPKYi2az0GFTAhuVRw38DEi4QxO51yGkLnr3mFTU3N0aJ3L
RtHpUDEV5TKo63+ZUg+zIx2uJ3kvy0JvaAo5tknQuIPCqCwycVeQkGjxPu/SCyF4V40e+XkcQp/p
zRMYWb1TY3OdpSt7xXsiQC7vnABiNy7PH6gXaGvzavF38zuTVLq9p35ynFQuHpzcztSBoZ1JbD92
FfMqbyKNvSzzey3av5ypeOPSpPAzoz5fT4M7TEiBvfNJsUatWfafdb51KCgRt6GM9HjLzhhVYFA1
kCut7wACMLRJPclih69eSeo98j0hqnuhLyFC1nfmLfxmAjeqhPs+wTz5iFXZh0irFnxGCSbEHwm1
XaBrm/+Mgbu9K6CnW42SPBpVW8EjoxYrpDldiau0Xizv+YUmbXPUHleO4MAtVBkh2nMjaeFFkWob
cOtYirxXL9vsp4Yjy/LTp27Yb+H8M30tXhPeFEBxQ/8J/AVll+ocOQrT3EBKF4ZZD9kYlkDbDidt
JGAEas8OwCnrACt3nqeaBR2SwqpKzTFulpCbIg0npBlMV3ybN07rdZtxkNSXFHPSp0hPaU2Vhhrd
gSBQ5EWLf1ALdR+jrb8L6RuB91GIYVzjPzBObAo001uqCK+2Lp80QPwdZ4Kf1ER+w1pTlJzzLxkP
UWWm+ZK0KVwWFsA0Uy20XFh4XX6nulqc9yOhIKosW+09Qoj4b11PLbQ9A/vTpt6YIiSZsPbQDRIG
G3fsUqlKbNdhNx3Zh0ePtSckEykRWMpyY07f9zVNpOg8VOLKF0gVS2ZpIVEF/BFhISfhHj5EhgWV
cIOwRNLbQ/wXz0mYG+FU6t+cLhMUxfCTQlh1b0Euj7pSQSyji5+e+GK+/xtriPzalz3CtuNSaJdz
uG6EPrLWUXSntn9eQGjiDGB67LXE/PTjUR25+Ss1ALWC24bS8ZlsRkdzczk40hOofh3CRpmjotc/
SHWTJFNp6QCgIVSDOifb0NDHs9PueDxdyNs81Wlf8VqHOm1iAKGG8j9ytLNOsS5qKY+LJ+usw4qQ
opuNUnxOmajwUFPw5GbYFS7ZDR3kNpgkgfgkjsEDRsZt/hAU2o+ZVTtGdusWToD+uRtr0kjMOUCP
x7xoAJpWu2qDui7tOZvSqog4PYKiItPc9ueLIQOhToUSBwMShhzllZlpuR6h2NEwThxhML1+LLZR
pyOLqMgRCjTDhOSkoeIzjI3C85lL1unm/go44pRzGzjfmEpFpK4GWh0XTm7+AdH8bDT+wGbpYBS0
0RYTLPTSbp7rZJULL0C0VM+TZ4AOgSvzs0HJ+N1Y1AYaxkQNhamC5pmwi7FHI2+g6UPYR3S3DEdr
JvsaxWuevI1BEdaiKQ6qzLqlzauLlrRIE3TWVKDK/ZtgzuvwCVSDUpY/rgSKv11ZXWfaU3taekNO
/aR2fw4ntHFB/E9pm8rXOXAENXHbQEixgplOhf64PmlHLVSb345XfoVUDe1dTjcaCR1f0Wly8sC1
WaXV8h9eUWt7Dj8e7qk3KPZmcMlcE4nb/g8xe8mrbFCuRRBe91PgH9iPPyVqKxWlqzRxgMVOFVu5
IsY5puX0Wc9JMgPVJhIQXJvyK91FebESPvmo4asHFnP1J43NijZVHTvchm0KbjQFlUaNW2sIP3TL
0Y3GdUPSMgxeXjcScwzLFx+Eeh831vvOIA7mnVsqWjbabZjheHX/G4h1iMgeYLnAFPBh9P5B3jmW
fuXunjXwDIGbLDD7IaXY24ZyBxRfamEPm86tHmKh96Unkss4ofmI+fgArV474KQ17rXWk+lwlL8M
J3btoxM68PdiLhMfbCcrgcEJuS6WDY4cFPxsKGkEp3AAYh6QudObuVUpy7OZCUbOe6VYwYutKyik
zeYpX1cnREYNDWTWRNSBWQ5874OTsu6A6iddYxFh9ujWyTLXJ4TUSWQVcpKCVTlZXAT24qsBgQMe
/8wQ0ZNfnIMRaEtef24oSwVUXn7nnsLspYSwqHxevZxfA0FD5V3LuqSGxYm93P480MPF7YTKTEez
KuRwmDlK7VhTRZvG34b2Ouram+mP0rnLTEOe+jhv9W7O9ghxFclfzzWLWdo7r0NLD9mw+3saH5Rb
Wbs5uXQI74wp0FuolHFE92nJRIKbiZlW2r3W0t0uhkhqNIq+y2lstPUwH5AnWYpBKWQzKi6HZKPX
eaoAJvYc9FuUReGbhkHwksAYL7Xtxv3flFG1yR2TcpQMdrUU6/selWuVNz6mVJTxW98eQ4IdB1Ef
NDgoviVP7ahi7FzAXf6qNANclAWVai4pHVoOZefYcmjWs3DVjOsLzk1j/0lfyf62sc2lxOaZKPSp
C6n/Vn6EO4EAU4SmyTv1fXQ0hKTUT4WIEpaSBoVo9Eb55agJq0dK729jcnTuuflo4z8Uzsxo7wol
Lsim5F9FVHNmZIbs/UZI+CRQG0fyypW4qrDZCLAr70PQxSxnHs5B1LXn97cBGTpdheu45xl/mGvr
353Y/7jjJPPDMzn7vLdtBrtTzTuJo/bbIVkQNp2SHMYooIbbkKun/YkXTfc/bTtPKEJdm51Cil8f
7Nvk0NhUwKb+iwePlXwMYVs6OiwZK6/HE63pat90kfHaoNM+JLx9SbM29tOdmK0UkotbuBj3/32J
m+LF/EUNzbWHFcKTE74U6yWHft+sQdyn2Dd/a++2N6D4/RdFXIYjBgQ6bLGkcGyA8mjDWRtpGNIw
93MgsdWLGYZeW1i7pawUQGoDXkSj/ySbEdnjgFu5Ic//n+4lHzifFHayIPmlLW6fZA+3UnG2faqk
KbsDMyGhzM4yOotHQTXH6ugHYJTh3zNnFpvr2Iuh52uyv1iiPl6/sSERVd/m6H+qY/LX1QCr4GHc
QB5vpnr9nZTHyyVLdYtvmyGvfRuwB+lRV/JXguOfgE8bChiYq9dKFdDZBnBYfaisHlMQGpX6lXiP
vhzoZh0+Lsf46Uw8g83VjVyNXQ3MHf7EfJg3tCtvUM3CT5bAAWE3YJYlO9TosWguPMDKrsG/F89D
oQpa3UICusBMi/mO55JeY+JcZTh4Q3k9sAEU78oql1H2dkc+IpS//EVIq+ToX3VxPyyWCN3Bfdwt
t1d7fh8q+VIuB+VixRinvxplzFj+od6scdAZ+fEsx7mRhlSZ8t41Y7iD6nmAoDaTouKsyRe59DfB
zJGIPPutcdN5rka462/jFhEjSEu5KzlU4WlDbmGZ7ikt/Mswa6sP14hHztzBjHLI/b6SWQXuzqkE
O+w4rpDsm4jpPVWExfe0McXLWdAGlBrF5G0qioJ5QuH9xzDlHJd+T4rpb35t047+ajpl+obhUMyp
LO4AVNdUteWzvwJRZ7p6eR0U103+ugIdSwcI7nIQF/+p7BIoi5jDoEX+WhOutRP7QccgG/KvatuC
4D2oYIktyf42oWW9hJDbNysboyw107Ls8igBMXEUyrM5gAhPoLQ5D+0kddTgJ+XTDPBK1Fu8Sm+d
57DYCHruk9tKr+1iSQMCnf9nEH9l+a8+buG6E8Wefpk7lQSTFTB3C0ybSi1VjdtGS/FXsyYtIm8p
Zn0Yh8Y8kFrqKz+tqXE0CbynB4ypD5ezpgy2J661dh42dBof8Fjd5lyL5c+XWXHMbgdmIdmLw04I
xq3BVH+18F+uxFWEmCW1wB8Svzhc2UdFndiMBg1bf443VgFmxAEDEOaIwxz76K1qib+uWFvc3HLo
20HD2iezypgWL+p16KOzDWYy/MTuEI8NUAJA0LZy369Z2iZOVnRc14Um64/d8nxJWCiC4FHGqLer
4RG565EWs6N8f1BHGiz9b25ObP21zD1oDXdbZRvLLs/mkkvDTuCxTIpm8SIieLyAOUGgsDmiLRkw
mAzDlbtXuOhEP2XLP9Sc7SlcNhyo0YOnFzDKzl8LCgBzujPRkMHB9FgfHPssmHRZWyeaH3Cvo/N7
hEmiKsVmLKYyFPkt8nuYrQXZi76j3x1wK4cVOIRvCACM9z6x0CnYOVHLGclZRV8hnulqalSqAK9s
3md1MtYX8DcCgs4W8HkigNIA5/rRMeqTOYOanD1I5ZCQKsdCnkzxueXIRbvEpYxdVOUinS3ssQLU
O5gXQwqJLV3tB/QfoJ3U/r4KKyvqJbmcMHDvPteeniolbbqmQ6rjWXE5GdeWj+6OQYqXygNFTsxo
Tgs8azq9XHMjq1w1K6ilUFABaFxYLvaEbMnhbPi+VeQ6lESHJSarcIu2SzvcrNg5ct9fwcOmZKoo
aJxgYmUPC7BmelgJO7opiy9VJ5Ow9eqkkWj0eG7Mta7vGIIObB/UC4wYcD7US798UxEegq1CnYxc
vF+rkbOPlFyFymFVh2BGXPl29GaviazMTyfZ6jT5l0l5ake6b6KykiufluOy6QQrgnvvsJBdWCm/
PS3vIRvzy6DfMsiOJMtWSIdBiCt923EMpUnu5P7m0AhR3fqYYrxMlcZEqCbK2WBvmoxAI7h1VhYo
OyEcSstJ9I8q/SgOeeWaBSAZyKVdCuMdq/FaUXwgea8Kcoixd8DXmIQpfSrl9KT7ounb+nMxYwPW
aNDZ0WgHpJjARIIopNr4OyiorI5TMD4LdZzoaDdl37U652ACQ1BbBH8TkM8yQPWi4AjZSBWqA0zD
XI/LbwRoFrHLXPdTJLz+rsFcjEHXax9qgsk4pu8QZwhjX/67GvFivs+QqdtNxnRCgolD0kOU1TGS
oh76BZS0Ay4YRGROLVLr+mrMvItrTD6IrQvPSwN3l5ME7VIOOInTm21NHzDxU2c+GeWxOhlsjTdk
jiEpN9jDPyg4mokEoFdKJ+Egelr0n+6dQqidQHKZ8T7aeYDQ/LYJgLCiP595lL5vOvHKR1oN2mQo
4tsicQPS3PiUPTsjZ20ISS82yUBiATzA5SRmIJn9lJuYmvuOFqM4HqdLdMZ7pn9+q7NoqsIRTTWp
zOD2mGrR7CeUvtvsvzIbwdsFNvFZ5HJqGXXu1GpEPiGU+QW2OE8MWr5o7XP12P3B34cPsWq7kzbh
OXjCMZYd0yjl3M0hUmyTwBk0I6BLNMzp4cJYMA3Mv5u7WU6HpDxzLo70prQcqKJ0qiJsQoF0Ky/l
sgzqeP9gWvbelSfYdxaT9RV52/jV6qRVLGOMkyNcGBg0U95SQTGcTxE9I5uPHVGYYJiK0u5Kau4u
QB9sOTjmcYpE0H9hrJbPFCLu4aV5Edsu0ygO8NnJduakoLD4RBhEdwvNpztaxWT4yF/swVXXWR2K
gfJdB22z/IsZy5Bqe9XEJbGtu+B2RWG68qx1kfmw210MqtHuW9/W4Bufxm3FlN1ZZPL4b62P7em/
IK+cRdY5y0o87d0F6CNeV/7RQO+l/wsfwTG+JZ52YfNxsfCQPvOjc/Zp0A5d5wsu2QPIi/Me2gNp
Qkq9JUxqFNUJZmIjfuzduYGnJY4oC94V/UmuUY0JXdHs9ErgJGLhOgSkQqpeKGunCd2OCPreEDvS
RKAkkgz0BxOhU5eYyjCTKlQAqoCoKArJHCsbTqmDjzTws95lPozGBEFj9dAanUhxVEhQXDc6a6JN
2VoMQQ0OCu/EgugO9e0RoKufspbtkjSBNK3EjTzeiwwreMAWSvu2aJt+mziBlf6/A+VGcTtGtOHo
1jFV5FqQ/pOOJ6wuTkt4kVj2sAPEGJxTgAIOsyF9+0O9FmNeibOyZFUR4OdPhAoJQPr/XFh1IOZT
kTbuWwVaVClD+a7V22Y83mf0OMM2Y1GDDoUXaMmZA3AvHsRQPLXzvbban92vQJ4u6qi2JiISAiTR
jLsosytjMTWWOcrPkLJOEkvS8TUV/kVCw/GDKt2603jGBbRJkamtDJGGwcX/wTCHRnpqb+zW1Jho
0+W/0yVndeMtSnJIl9trVPmRb/CCuM1AMqQwyVSZCVtfOCULo8LjKJ7wu8X5eqeJHKfaoGwBMpZ0
i5ROctg5pySY04kkcWRqPLYvFLVIYHHPv5cn/VQFMkE+yDDQgIlo9chz0V62sYcwY5twr3craWe6
ZCm5n0K77U/a9B9tRs0yw4xdJQJ4rRQ5xHUW7F7iTCYUG8Demvd1kaHzmXDMn+wyzLH37KT4CJCm
k0fsFuXQ0qn6OPvzHAhsC7JUaGVoJF70pr+nqZ6YALJiULgENFWsSVLN14OwxvjxPr3K3Zq4lg7O
vPRtHyKYGfBmqvg/vXxlAgpxivxM7lvGTMwYGyceZc+JBbA4FSFUPRBjVsQi+zzRccXmVFprhHlq
McKBl/f2bqJOeJu+crLQIg+/0d5HxYwUOi4x5MkJy6P/eqEBkRqeEesd5XohiX02PsG8GcdjGaLW
ZOk4HEeyElKz6as4bwsvRhLo0PNSmF18yA3JH+5XutN/WyLMRFObb3+yhn7VCQtMe8zujz68oaht
46BR1CdIX01DOvP1NN9V8cdu4dFKZwQEMcAfMfCYNZo1kqBttIh+W3Ftm7sQkqOXUHRqDpp/pSlP
CiIOVEwDRbTk7A26o974Qwi0lQ7kW0SLx9zKtbqBkBP9H6vEMb5Ssty0C6T0Ykb1ocywANU9SuB5
pOPl7dNcidj/MD8MqOSE9Y59FCGWP4akTHqMnuf4BBBYFnQv7Y3VMVvXXDx2ZcrAFZqKXe9RymMG
XuMTcPbWFD4Rl/coXCKjDmoxVOxPgud7kXk/nWgeY2R6bG3fGanB9m9A6feFpF/UvWzhNGD37KBx
qznT3DflICxh9EYvINzkQPG0PghO3PvzbQb86PyYx+twpy4koBOohHgUweaBdOzqSDUReqT7QR2/
w2Fidn9cYhoBbDrum8H93SamaSTsURNKNEqzoaSp2eNpy47ujUN4sheAE8BTpF2+EB80KDnyRbkW
Kdzdq68og7o01wjKuD4oXL4d+qi6wN45m27eQ/WJAaDlyAyVGUR6I5l5hnFEu5af8f3gMnugUbxn
v3IaHN9nyjqDVmAR9v6LoFWrtvORv71zRzxTTjbmlJEfiaPIT1wD0OF9coE2kPKRaaoCmdDZ1i8k
/YfHG7EGFCCJz33//YIu37JMoMhx4iGaR/uRLyqZvXWo5hS4zFBGggc6/nP/JEa3BIVGhBovR75R
x5gMuYVk9FpxvqdI1iS/LwGgUF50SBcypldQI3DuNR+SdttvJ0R/AFWsH+w5+FVUeovZghVQMbuq
CfJ0aAv5JVF8M8WXOTU5pLbJ6su/D2yoXRpjBOpMTmoviPUSkJtXOGpsR/SAtwseReEVv3vZuDq+
qacxaV/Dkal2DQrrkqfAbsfRAnOwzlGIUjfvftg0Jiz719a011TlrYi5rn1v6epL/QMFxl1w7Y9P
Lwi+2WRVDMf68yKuVF3aS6GH9vCa66iokeqPvGUF/Mkt8Y1i0aL8J7bmXqLdVnbnNAELzRSqh/PQ
Izxcm7OJR7q/MjveH2gk1MPZJVNZKgcJyGstCxb0MEUPrDzD8B8rnKXaGlwY/pJUb7NXGZAo3y0S
rYXrpwQYxiL+fnZGH6oZwJ/AsZsGD9RLho5MY5B8SpYUw2UKT8gRJ3AC53e0Kl7zE+EFZuIQZFzs
Wawp6xlWQ55opwmZFkOPjZPwRrQFWPnEI26+VubZDIbCPtG4L6y37vToaUDPPjfbgrEuEJ8p9HCv
X4V3sY5DnPaTwTh9w/IRfv6WiBtWQuEQ3OQt6EEEt0gjktI9FJdyT6h7/YtECwIzuGnQVvQ49ss9
16rNUq3RgEflPxaxqQEzzqAuIYOehoDFUerKWehvAo40QbQArE2qJfuqa/4QgAayquDLJFOrQF7m
8sHo0PIM9bXm5bEhloE2AfbwRC3ifIXM5ZiiTTy2QCjGqzSaaUw5mTj6G68+bYshKdVc0YtNfLhD
HpHyBgHGISIvH2TlEWQkpwzuM04GN12I1u2L7yRIr/QXnuNbdfUgHDUBzZpDDqzZinuUAK1TJEYm
g9y4lxtFxtEEiNx83bRWYwbAzeZAUTVw9BUhqx3VgoVArB0pj7KKhL/v0lJKlmDYJVLHq0dSJltr
RUOwrdfvdbw7nGcgqzoFX5OuWoFYwkYixr8HwXpvJL4Er5aNQSiW4KpzOO3jVJVK5ir1ENTgnO1s
9wgLrWod5nYIuMD22hKwXQFSp1oNphUO3vNyXLJBG/qn6VakAgghpIKStah6od0eaehR+TZ9pKpH
E8i2MHD9Ccu7T6cIC0FH9SMejb0n86QFldunBWHnjzfhnp0VkxCEjEnNR3+EBH7gGq7GF+1S1S8e
0b9/CVAA+O4ZtpLcWMQNJ0jfVZie/lQiWThXJR9kccrRTjtxBx5h+x+qH7HgwuoOaGo+TWKtaQaI
WGajIMxw1znjxDdFuxL49CEjVl6sabx5xQquuXyd2c4o5gyRDL+N/DNWdTAzheLo8for2OA4fur5
wBILYVzgELTmd75ojWuH17NKiim3MYqT21ByUL/i6xB2m1fnA+AUH2/+lURId5nkdq7qllYNLbc9
/nroeBe0O8pYZ827c3lE10g2BcaJPNU8EP8QyvY85GFcK+w13qamqlu4gr2QONDvdGjCzmPaz7Bo
0fP7zOjOGzsdj/DXj1PRYZJEPDmNvxc9ilv8246dq5E1PAjA22Z2ATnbyybxbFt84RLJCzf3lido
t9XOas7amost6A2kTyQrEn0Ln+CxoANhgzqHI5aXKeu4KXak61mfF/W1zTKlVGu655t12VjPFYmC
8cOgIh99RpOuiCyHxQmW8odihH0O1oBs/+Bi21zjohDrvltEGkjjs6aYiGwtR9NdCarunNq5a8e9
L69vnj2vLvdA2z5pbZDkjYk8twXo0uRuiLatOX0hbO7KTvbdyZmup+baBf7rvU1O35QlTjO4hdkA
2SbZutYrnxdK6j/OvMjVZHqX8RGBglayQNKjaZkT3aC6yKWPImqtXABM+ALcMJzW+K3/4VWvf4jI
78TA1zhnip2BRylxvzMWE+qmYgvVZd7jy9gASjq4R5Jnb9059CQtWqzCpQnsh6sdVikBoJFf8c5E
di0g9lR38TIRJ7K6qXS9NK6T6HtffeqzgYNHrsFV/RqFDcWMJl4AbWl87i0nyZU+0KwEjDWqVbH5
3rAvAGUfIsM07hNmzE4TSwTDOt4Q+jG2WI3JX9v3uuBBmKRgTSBhv81R4EKiqTknLOlQpZmt9OW2
zC31/gWY0VJsUCU3m6k86WkdcyuezrD3qrfXwVWQktDljybnFiK24YKGRfyN3RIWiKPGcsNKhcJB
FOCwJgYLx7whwpiY1/kKn2YB9q50dIpykwcJlBz9tjtpwyllwPzT/lmwLonMfXMTLldpCgqQ02U+
fOf0X/lsjaptAvq4Ks27nmLcETuvIUo1AWOtuHaSae27cFt3JPxF1QNoVp63ste7KP4jyKuLC3GW
/Do3WTSLNdky2ukX8by10s0FvbzCHz5XJJY0jPNWsuqyuxlMbHOq+/mL0agq4WH+1Lu2HxkT6G/3
HNNeOqfmVfIweRSUYQqMAbLvLO5R+TN6M+U8ITK5txILBH4blUG0QFEP9nomMnzeH9nHd8gBQeGT
7IeaUQ0Yc2rIEuQ4rXEE3P68SqPoiYy1P7Hd9E3oNl/nnioQEkPI6lmJ9UrEQFEGOLnhaDeNySnY
US03CP7fa0PNOclvgb9ebBqgCModMMdv6ChPMeP0Q7b0GsLxGZkD+or0GprrOPsFRmeT1YSipS8o
iQ7+aQ4DPBwgSsIepJ04s/TIYJgqy7j+Q/ntwAKIPOMf7kJOz3gQlpO65MlOqQdEbhoAHWcPUqq3
zm93rogTuW99I7i1GNcwjn6NSvaoTCjXXHGvPjq3CTzyfOL8klYzUlXiU5xb3bn6QeEJQY15ZWEi
gwTncyglJKBtQ9Mh3pHkOZpKynyRfAGG0SJeFNu37FZ7VlSjfkBCk3OcaqeQfWyegNMedrRzNSyC
KVDQylz0Y8ON6XgFUcDWxul5R5g712yt3DxG1+w4nfR/cjfdTe6W8Pi9BGXR3YcczedA4VYX18OS
N5Ke6V8WzLeNAkMVEGZ5oRpzlNqlZK79BbzUBwXemSqXUxRopMckNtqG48buriD3AQ2tRfG61BV4
9uH03Xl+9R+wdJ3PIR9OMvsKVckW0eKUO6kQL814/KZWofIC+5QpDgKcXWNWFPjShgxG0pVrAlBe
zfJDd4E1LT6zZe77tt3YmNlWWTah4x+XWCSsyP+hhGr7QRps00BQRXP5mPgRJlygnfsbwiTNSOE9
iLA3DoR2DGKJUyzZ1gXXCPD5t4xlAXClVoMe6iQAZubpcqVP+4YXOUS6VHvOYtukmTiwhhm8jz3S
ESYB/oMD3WrdkbHeOgeXjM1W2Vnlkmu5lXADED/ZUPLSh5nijioMO432jf/mL61gAHILW+KzJ2Bh
zFVYIbS1Bbjf9nVNy2+ZtgAwJgT0FIYY4hGI/D/ayBPtplt/QgJ3UFTw+VL91jQOBWzLTQKbeeyS
8wvi9mo/SQPXBKu1MsWKaMNahZD1HhWD6OZVVMmgLbj2ybf5ef05ldD8RfYeawYtLb7zao9ItkI1
vlxARJWRJnydshbqyWycTES7pDbhXf+j6hQ9D0tONjwiBpOOVRsMnwlFmSFIuV9ZtNJiWmIFs+xT
EgLgwA3mvUVa2mXoDdze+tNyrNIDK6L/ohbtYBRsA7VZq6m+b8hEZ6GswO9Zo1TdahZt0DfUdMFI
zasDYmmrfmvcEOJO3AZS5f4UfXZeNyJr2gq7cRfzCaii9BThyNLQb4lb+p9dnDiodgs2Yj7dSCAD
P45ZdwL0mZP6eSET/eKRwiP+Xc7P0wE1fXejqJOCYXeyRU4u7URB4ylhVzwlQe/MM7kGBYPtqWon
C3ahSIYzsYXiFGpzDcdW3i/RsDhNNu59YRw4wN4JQnVKhrk+LG98CGxmDqqBpFwwkR2ie+2byteI
eo0JSIkFeIlsUXkyS7R5cL1Fqp0Y9xmzq6H7tpaAA+d1Zb2N1hhdvMBZqAe8X0OzMsXKyKmm0YAF
fWwYkh5Yk3w47eAg9AkawRCrrgmQWAeaZxc5vrphAYFLDL35V/L6K3+QjfKkOU8vOkS01TX0gDSj
bVQoO3n5TY6TC6Fu02wn6UZehWp6CJ8OykAayesmTU3DcIYAieXARxw7ZJW1QUNgYv8D+eavW1CZ
QbJTXlF1XpLEirDcNlh96+z20dIWmpecB3IjaxEq/WC8/Vt2R6jun8oczfliZb59t+uxE2DDQeJo
T8j4g0KmAQmxgLMyFytDC2YvO4GK1k/gfK9TxC8DLuQHfZTFjT4uZFRe9gO4qAZQi5oc7glKRjch
0u2W9XASI1cAxfQKfx/+xj3YLAv1B6U8/jy0F7CfxBaCtJvl85lOBrxJq7vuYKIpxSNO+K7dA9i7
ZCvtLFoA7CyXgEtn7tc94EeWP41Kf6+jDKJx9ktZ7saanpPvCUqIcb2+bwdKshLo6yi0xwge3PCz
hZ8TsRLHe6HsNkxgRHz15ZasdSJgJLPlv4dwWZ4mLlz5WHrRh1sJWMNqsP/ANQHGoMgFuIoTyji8
ns9djsAenW2jX/m+avHWgh7xkNXk2cqoevC4iYthaheHsczY/rScRMrMpo+YjFf4gZsChlL0pfku
D3SYvfNJ1xQgR/WERAglguZB1DLg6cnDwPLIsL86YDv/ozcdONgtRPwCjlk7N+XGxDTMKW6DCR0C
iNpKzjNwAC6IirKf7t1JOdIrEQPyyS3TM62V8qdeaTVCuV/1XSqQSURTKdWXDVqjuihDWxb4UnmG
TH06rrTnDLNEHtV5nlQ9dkeyaXnxe6+7iugrMkvYzsIGPaQwsmpisGSEQ9p6/dP78fYoUpJ6gWvr
/fcQnfk8d06ZaG86s3hnogHmEgL0xol29VXZLyhbRacmzzxb6cNwRzSdzj/vSvFyfFT8IjbGiv2l
S8RFUyG4Si/9+vrBh+2HNKbU/1zSvc0CleRvmQZysrou+bRgFIHwO7V24ttpyozOQuOA83SHccmS
/jCsI1y9XQt8RMlSNJyRzneFp47lg+WqiIwmHanqQXYzG1km46J2mdGLSAOGIs2SB+TMUrllNH+P
7A3mepei07oimzBWoMty+dVlqEaLGUWLMBTH0D5eU5wmOs5qgVJXxOlLfUHRLlcbYyZ8t4n1p+R6
Ba3mBVPaKwfmJCUpNB62HPb2WU1kzyvrayVPwIu24TmwdU1P/90DB12UzJTvo9/o+/Zgh3VfCO+l
/8m4Y99AmQDVMQAN3a9yZctPByWW9Vtuhywi12gvAOgeXhPT0k0sBKh9qBe5sPFfUBKXoN9MFBl3
+neHSlmGBi/DU1NvKXCOqlegloU/vHQt6h+eZ7uouDzo09zNHOTnODQRTQDKmUDDy/Bf/hA7DSjj
Aqaj4UBew8vGDTk1ej+8Q/L3yE35pgn6iJzMGwvPrRpD7oaGmYVNcuWHxS5QIaqQVRZtpwVEa87F
wGocd02TBYsIPPs6xZJKLGyQoapmlWA/Kw5RQoTTqBFxJSwPPcTjidn8csk9h0yLiobo1AtLRDoW
HJV/dk6dm0jYskq3ePKPaeRkCZOllUAz0H0bIM+RARMli7Q1eNJcwvbPW948Ad/0LzMMOwaTdWJI
UEzPx5YumeXWzrrt+2nPD0kIlPFxh5bzrzAM7W7reWzPWaz4DkGLIr8u0miMgAARWApWI8YScHrz
q21uL3v1qPbU0wDN7/ywNNsXIomsrWY0mMTnPHz1Sgux4JmXAS18gucja8GYrshkltvCjksRbemB
ABhF7MhBz5zNzCAlGEcEW8r9syiISeRWO0tF7owLjIOJWAIhHGzsUYKfRdrD+hG/IcbMkV8nfqxB
Ru3e3C92OcVdMmgfKdRUAW5p0BdAhg9vssp718aq83wpVyf9hFk4qbNdIedz9RIhsZt+6fjEOBAw
7RU45Uopq7WNdGVyM1xh8pMtpcfdmU19LfslGTKRZVYvYJufptMxt9IPjXLlvgnv8hefgxwrYV+a
KGIV/LaXlM3Ppy5+jDs8kOHHRgwGOLMo3yNwbG/MertZRet22LbMOtG+TdE4O6Mjd4OW4WldDkCv
Maj/YzGrgtO2hgXaOhU8gAtiILr75WN4QmIrrV7McXuEhTlqg9pNjR2xQmdOCLUMWgELPNGMKSrW
uTZtNk33z9s9R3XuQb9e8C0u37YqAjp3XzqLh52omyMbOJyLoGaRxx8hpn+nwwcN7WsY6w4SLoSR
ZbJsaIo7xpEttxPamrTKoGYnWiHfHAZgu0cAKXFEUMserIEmlKXSjx/jZiO/H0nZ830h8lMN2QSz
MA23FYZuSW5ashFLOSX7rLN6R2b4FTAaZm6pKPbmTEaBHMb2OjvqAiDmX/Q85Sh+GgbnqUWJQ11g
wdoiYkSmLnfAbCZSqYQMGAJqkGItz4G4rbtYyLJnXhyRV4B5RO5qUlQYsKtOgqEqUpz0PUqom1CV
/aq6wLxHJG9UtXPQvbgvvkJb/WOsvGQa18HrImMGV9Jkn+l/921TcpV+aukBcFcZn+x29V7Wr8qc
bgT5IdgrmzGuuE9OFjmEuIxVwxMyEIKd2O4O3qW3aR47zY247fB9M3U5MuCSZw0ZtUIUdwWZIXN+
VTUCAJhHMvdOAKwZhaDm9Dan1BBiZpmMvFIomCib3dZVCKfu4JUbW2ByHI3GA0xI3mphmSlySh79
2MdAjMkhPlJKZbUgsbUzE0cZuae61y0yFRUKjrzSf87nRA/Ko0ziy+MtzJLYl3XxmQbG17VYOvpu
oCnWo53GLp9C0y94T/AkF9zGnPG/X4G9P9ghl8EhKmHhsCAUlme2/rDkNEoNkaUys/kk9SoLUYpE
kDwWbQlMBxcNWOZHup9ptGfrw7bKr4Y9limeXa7jCYnonY2TupIDBl38bQe+Iu6iakNb7Sb9iLwx
oUEQRYzDgT/WHfRj16j8CUGdAl7VxVNKc36jXi2Ie/70epis74GcUrkJvRTx5I7N9A6703xbLZ2h
xdb6bSdN80SK7KXiDjI6Zy+x1mLohiVLvUZIa1o1dqbicclALKLCr6goAdiobfwLTROigUjaC6XJ
uK2vc2qzO7xzgCL/8EWKZKtOO8z7fqpB3v34xQh+gQNeQ5Qmty0tX+XsHGrzOJoa22QOADoZ9xwZ
7yIGgUGX+Xv8b41IFoi87ujq4SKFAGfb+vlfmxcCGNTfbxJQb6mhC6f5U08MjxGK8oYy+8vQvc8s
0rJdo9QlnyvJc0vgjNK4oCUoMR3nMpolxjujhcDvnyc6MmX+cVvNZdf9/uJnNwvVhrBq63irTmrl
B+bWywmpIOtYBRyns/vcSuRvA5+7BuoRAFeb3cxkvqqE55XtWGDbVNBF+lEmaAmu7K0bburQldXr
Z6IYr+HHAVB6GDzKT0X0bw4W9GxsOrosrODwnL3vyYOxBfZ8dRWdwStFFnP5O3HecUxoVryUNCTo
XkB848TmvwnlF7L3fbZRFe9tTvtWqARxgXHBR/3oOuKdb2LBaTOPrBBifsG5p+lfCnsLbRsxadYC
lIRH9ZVKqRrZD85ajidyWSgWGHZQShbsgyL5V/PaYcE/e8oH5nFBDhfHdnXHlQaWdraxdr3uFRJm
kapVEpIPatIOcJospwVcFTyW7PoHjk3Q6SoyNqVqU42GfbN5e6rfUcxfOk6loa0YouKLJ4XP4wLF
rRMACjpuW7iFjwBg38p/AeJ/vYHls4sEt3UqRck6lDIumRern7V4waMtTqepPYpP9hTEC6Uwo6zG
kw512QWFOd0IsTOFFyMjpM87l248x4n7WdSMh7aU9Yjm+fnlowh+q0SdZImh9S9YcBh6/ICYRy8d
uQGqJBGiZTSolUiQwJ7l8S0ax63KjBWSzNMxKGwG6bHL9qbwNl2X/88JGNAabk5NXHMVTHa6avaL
TjxpyJUrIMaWDpgOcMqvzfNWtvrvz6Gxp3XzeH/9CZPSJWD4acio/u4JkMLbAQecw7iKhSmJoAkx
yRUdahzpsI52mfX7HkENs5JBKQ0o3UE6lnZvXMX6MvShF0nb1/SeWHdo6mw7XbkOlv/KlsWZqbsL
X0l9pfXJk1TWeTXJnbx0ytTUxeeocrINzq6v/YIuRL6MyrNm9WfjsqbAOM41dlgS9/WciTtW3JLQ
NN6FIypl3dWvZdG0C8ikX2ayK+d0tqCM0ooROyDR/P34fT+J/jWijV0oEDFFrQ5zCs3R7Y9F8+UP
L6h+iehAJRhew0zv8ahw9smC9axzIDvLBUUpfAkl+zJjXmKGTIJE7bMoWNeRaWa0Ej8iylDPJPNa
VlleTj7zjNFiaQxRCodR3eFNCLfBKNwPOA2qwCVzhhmcFtdj+4nxKT1D0TjH0IHQaamAYGFqGloy
VsPC4rSl9kVDtzLV2Dn6YMIp4PwelphGikiFQrAnNmI1tw/cbNlGmP+3NqprTyPUdig/zzHNaNaL
LhMIpHbKB0OBWvC89CofQsDn6voDpiiJMtq1n4fgldg06JS89jsBSX3UJUbUfK/k3Os4UgU1ZfT6
pWOAR9UxfO/hMx3JoBNhqfx1I8I32vtmNQQSeUs9ZmSub0KCsI0I5eqsWKqC0r5LFaxBMCLUou8q
Jzt5L4Y7G7zBEFGaCf6uQ68ylNvikCqQ/jGa0JO1fBdTrBk8qCqm6gQS36gHbhPIj8kOMfcATwpn
XMPz7gLQT/Rb4nyNrJQM931F94vh6G0xbIVctR67oCC4ot5W2xzuc0rg0GJrNvAHS+HiNsXLg2Wv
p/nWNSfmDs9mP3cqlro5s9IJP+AIokTLnHPne12vnXLjIltQy2bmmiGrfLSYcEC9izeYb2WS1k+r
zEkRufKmAFPVpw1QvDreayf8k1IzlzCllZHnLWUjyWg8ZwUBdTXaloplO114tbzwtPf0zFdr2nin
jZJ4l6PQ8FQp6c4iLEsNcahJskNNw1CkS0ZJgVA8//ZQRib6yt0GQveTHSsMrpGDD6f5UiQECXDZ
r4uECV/CoGie9C4x80ImX/C5GuZl/GxPBGpE7kfSD+457U/XvKH/XzQG3+Ksx6Lop25oKqVyVakY
MEvoZCuMQ3VLK2OVP6hZ033uPmN5l44KmDvRUimYwRe81pzgDWrQhzlOkH6ZyqlecoiugBpXXLse
85latyagsGqsjTeGWpvz74jSe/U7B3JaQYQCEoB1MEuBW9Fvw55X4Yrl9fvvmrFOV2Jm4n/kVCLX
ikvOm43rdwujYLzM7kdUwH2WbSYgSDCUxoIl+Okf28ZCJUroclQbkDNmeKYm0o4HbhOi9jT6Z1Id
mviNbIbmpSufc54uauE0thsslbt9sDoMBCUDk9tDjaFzoEnENxZYybtI7XUohznhXe1MimNPg5wY
GEt7lUy/tRnrfb2Y63vnTYHpzJjgpHD2/pI/ZWYLhEDycBk5y0V3VtMoBSIBbOQtlXKmffINXS/0
NniBz4qKN6boJPjxY/AJj53S2/NAXaqZX3w/AiueF/i0tEx+zNoH17sxjxJguyezz/69OFt7LY10
/kOLf7iPkSid3DxVsV0AV0osmRV+Gl2odq0LtAvMCAcN0OnMS33E3BkaGlC4J2coR+6q/UNdCQng
39kZfQCZwcdanSBIEu62SJUFIUU2Co+uBZytEcLcJOcY/aw8SPVB73dxmYSF2WJcxm8pkJpI7vAF
VDt3H2g+l0VnskM8NMcOuGi8ImdxLCOzgyci4n0+6GADS4gjDEzSKR2XZjxtr82AJTbKppHR1cdv
L7nOEED54h3hBAFE5yTSZTDvYyzelTMwWYPmkRQ8DIpAm738lRPD7Cov+2dQ5UMy+GrDF+RJLISi
A3RiJ1Gjx+85OFJZd22CkHiC3gMl9+DE95lrGNhTo46klEfi9qBZ7wAxN6+YPQHcBWCJnxht9hRi
oODyEue7qsZBP2KPZMR7PgJ93jSjONwbA61jQ4D1dYTQV6+FnVTWo6NzH3L6fg/y1uSywSdFjaRz
0RkCTrNLwcq5Rjw69N76iw4c/30kVHfBOcXdW6o5lW4R3mpXtdBl8dr3vehBD8eWzDPInBURDXlc
jlZ0qZFRpZx+sshqv2NapPEjml55UHBEwBziGN3cK/ZE6d+oZuRIfE5yEfz4BqXh64/OAJEwK01W
4kGS/+Spqq8AEXJ6SOJBxoop15SKQFuAMwvroypEJ7rrcRRErrcR5OAcCrt9bcPIKLiCqWSOO/dE
ea8NSklFv0cQgvN0bZRGDzn3MAmoWJr0GJKEcBYtrwD5hSg2AD23MyGKdqqki2SnQ9pTtSD/UFZu
YRIfKJAbPJNX0uy1pDfmbDrY40t1j2xWTqR7yFgpLRLmlrPVY3fMIe36WNUdpBInfbWRXOMS4VXd
3glwJZTDHiG6Nz3PLpExsVH3oaCiiOHMH50BxhOtMHrYP7XlsFwjowQDWDhOu8TV53a+BpdrpD8j
u+izkMUtYGgb0BX95KtAfdeFMnKBWaV0KWv9AbTN917589AJ4t1mqICS6y4kKea04ILKWM1+/bgH
eXiEIEaclWdSTULZiuoKJIG4crpPcZGt7j9JGVaINd/pp1xitbZhWJ16T3bHnTudZlKEZWgm5GlP
EMkglvK6712fxneRyELUNpOlWInCeL+lQKwWdMZagGl5lhUdla5yO22dqi4whfPkkFRLlEL+82dQ
VEKrRlyrYL9vXJDYubMIyBljK86SzOem6ehdyH9L3pwMyKO3Yfc+0R7DF/0TKSrqly0WP1zG8InJ
JmujzfeYKYYWs9wArO5f0m2CHQFxx3nauPQtdlhVNRjphrwF2srEyew7e1kQXyZGIQmT2rbbvbDZ
8tXHWKpdIyWQ/Dr81ta/rjHOrjjCY4EgnXgJ4OcWDA1aqsk5pr4CR6E16+R53ZbI4zr/cw7hFkv2
G8C0YkDQzqNLt0w6ZNmDwtIRJXitO65/8l6eHAULtUtaZnbrHRVMjggUjZSq99m2EiUhwIHvdXgq
RuOmtWC7ZL94YtwRgboMtDoemAaplmKWtAIUlFi2DcsHVAnl5gFRSem07xg1yBCiRteuujYOeRFR
IyQ3UtFM/TYQJ0gU/W3Twd/+D7OmVustVGBSQwU80IdhP2ZAliFKa9ixLFIrxP6aI/H+DpWBaH5k
/tyofNJsWqo42kThp+qN69WhU/LIUCj7jO3ivuxsEHq0gWdMJqvHgq9Ta2hNYrLXjxyCL1EYTrJ+
/VqL8WJ3p4+h6FC2q4AoEMObTSfsHy2T6Nwh5OYeliU51SY34T0m1qMNE90hGuRIalTtJ9ltHM7Y
RzSSen0oFZHNXlCejr5aq6rXXzWXwIWeC53xMYCCM6vsQhzWSnwrLgDBEt9ioIjfx0QX3ZoquOuy
OjfRolKeGZA0q3Xq2SvFIGLOy//W676nf0lS0vEKHNN66vmHVh2Tjs7+fzBHTKa67CoIM6/zeVVl
0S+ilgK4yAF+ZwXWAEPlL2BjLxWavG4AodY0uIcDZ/k+RcCvq1dnh39iYojjHW/NmA8dkt1BF694
jywfwvEqGDMUeGNpsW5eq8SIzRT8BI9WsOiSl8CYVHiyZqFpQUTAqm0KB6GXs0bXAEez2Lr2f0fu
CgiI6sVAsyS2Q6gMKbnVJD6SudauoqtkyYJzJ8t2wjvtNPCDMqhLLyUhM0s2cQHjrgO2u5ZxoEcN
VWezqRurEQuda9PJlmfxSOLFI8chyx7EzZKp4BNF+KJlKAJDg1LiYxjHC6JeQqtVV6DZgtKLvQbn
zX71b8T79MLVHQBwo3DkG5kZnyb1uf2UL4I3QfY+PmF21bFkQKcn3R3/FI2khKeFk3cYrfVcjFdW
B/p0wm2IQUiJ6wPb14YJI2GNzYw+7fxb39g4HeQRBQD6Qh1s/tePxvJ1KNrUF9UswCQ58ytgfJ2K
snBzOtME5BMYJ1XqkH9xm2UiEWGBEux4qp28b/UNGPe7MJTTzLmzBPJz1mU+kZ6flOgCUK+PQfbE
TX9Ab9CBSylHtHVbmP4x4fgaVXvJMkWAD/3PZJgh3rk04Hrjt8C2ZiXLYIJubMq1yYhFi6q6+ksW
7B+mmy9bllUWVwvyMDpEOHZgLT1aM+gblZ7CmWjFV12H+bW6d9B1Ebu7mHrglgn4SpwSe20t/krQ
d13duU1r6qj2JNUAculHdf3tow0PqtcsDkdWcULPSllLlrzmLXxj31UITsPWW8ohfYNzLh/Vo/5W
/YkofiGvRSnC+mPYe+AbB0RzEhYm8XPXc87nJhFFeDPIJ2WWS6Pj4wYdvONTvI2n/mw5cMS5LsLM
uo+ef5GMYQliMU0xReSvSGM5Yggwlk9Y5ILPoRLRa3ahUg0tyRKarmuLWW9eXDS10en6I/mnRNdT
59tJJGIqjbVSUzzh60hASWOvqxDUwCS06/Uh+pMgKVecjcxuMJQU/Cj7lOGtWIGf3Fvc9liEza2O
n0KiE1mfXiRFXUtljoqr0+JrRJQObRZGiAidUaJ03KmJQz1zNXBCDcOO2EgN7+VrHod4+tMsOcGr
XOBSbPQVBdYvQe1QFofLqJhBoe1FylH7duxB++eqhoqx/Nvdhjuu3WVLG+vOAuLYUMooh/b5+xUz
IA07QoOdMFxj/7d230TZu5lTNjal4wrYESgZ7oPteZJ44lWy6sO4Bl+uskTPLzQfVjoLdhFjKV7R
5aaSmxQr3Dh8oD9gW6ty+key/F01/5YileyyivhB8s4c/RCwLtm/hQWGEE9VuG/e/QPr9exzqxcx
gYhBBx5znpxM6nZKVZBpo/u0mjqQrQ6BwghxFpCts49sOEuy6VGJ8YibCn95ax/W2yTYCLpVm9me
XH1m1mLxihVL/ldL88CzTs6/0UgpNJNnjAWnc2Y8Xb5yabFszCR6LkxxPWt6jPJPp1pngJEdO0a5
08zxWrscimLVq2YtiDJUYawGu+uvl/9oHNfWLGrO+2TjbokWshgm2tMjHho/gegDpuFw5O+6YPXq
VqSEV6BJNHbhfi3MOxe8jYatAuud1BWkIshAMPV0EiUIU7J738my/1X4P4rFqbF2hsbv8QbICM9h
7D8pW0R5AZYPWzHIKZCVmuu1TY9cdrrCSdKEQS17QDQBM+hEzJx7ZF1Nco8vxPnXs/4nWKbgM8Dt
gDKQ4VpD/XueV54I0Zc/FP4ZcpeCkpl8xFbeS5yLT+vtdrWnrA86WpfuQEjFb85V8xVA6bfunoaf
eIkb4O3jOyd6rPcnu3WX3XPokEMMaoUozzxvr742/TBMWZE+WeivSypuG7aH49U8V5LLRqxcznvK
Lj/RvI+OPndrEkhraoXR1KtaPY26Fy6XkELAyL+OnJZVKucAN+se9AXI4tlL+/4bHe+mQaWDmJuw
kUB8hHDFsPobLvVl/PsL3+tSbshAyKRMGEdHc5i8SDitCcjEyY5V7AM1A5mNf49l544E6tzJjkxi
QVi0CjKEApJ2e1jV6KTL+1tbS/H46LRU+U2uaBwtse7z5Sknl7SGnb3XKY06g8nRYnoQfq/TTARI
7x8wsdKLNyhoZb/z8galDroPvPDt9CjbVVFbM7aBm1NkUlNQcIjnGxPS8zOY2BRwEEWBedQTY0ey
WxKxR3XeFToHqIg1IWk+Q6eOZ8SSJWOKdmwpHa03tGXuih2eGMUi73kYQW35yWybmYAr5FzUIYyK
j7WhYRICc+mM+N1DSRrS7/gKc8uXd30IqPw1zyUhI8br7B7oJfK7b4es0aids1KEoUi+Cvq1T2wj
9ythoRKkkDE0z6mITMd7mEeL6mjOCKqH+pl+ZzweP5sMW6SW5Dk6SrTUglbT16g0dDDzKzIIHKLE
6i4dURGEozYhYBnrqrvkYxngPajM2cv2BM/Ge7dfvv9w6pcvSDzfe4uUiJD5yB7E1uu9MxryyXE7
gGe3GWFaEev8ALkaC0Nf1L4WvJiPPAyuxmqPfrDgg5QjfZ1BWGHK+Bvez2cxN9uF+um6YnLLb3mo
3KHDUfWAt3PobNA5b8Unv3Mpe4pO5OVJDSZkKxPWQ/w3U8iMX07W+j7yjzUigb/tPsrxeWpjAnpf
5KPDFie1Kf4E8f4qhVJSnVyHJ+aUqtWwJhRtg/JHOwgqYY+SAuDCBP/DGHgkVxXt6rquxOjIhdyf
lL57FWOrKl6U7s0sb86yhxNDB4mFOBY09TQbRDbmpX560OfdryRdCXtEGZlflgSr8w8LYJycWQyl
Pti+udtZ1qcjUbBoYHSyk4V2f7y4B5gx/NDyRgERX69+aOnJ6gAbJTzIqtd8jlc2lYrT361KE7Mq
HzN9vT/uIvvhE8Nj4O/Nu9dgh4e9XccOPBXRbraRr1cGfwA85cSjiVJtCi/G62u8l/Ap8NB7qnXu
CPH0tezmPqjLCghgGt8HmBhuBE95wbScH1xdBQI1uoZZ4ZC+7Ad6P23fQBLnQYMR4qZ+lcIq3Hgx
ufeLQLNgg/rbRaTHGR4ZR/xtsnJ+v4plbHWV9zim6xkzVgX9Ya6BIYRZHY7iX5T2MDf0PmxoAJZL
4OJ/q6BjL34XT0oMJSCklkSowNkI9ew3hqn3PtlXI01h7O6/riUlVP3+YP4BaKs0IaXgFaZo9vFz
UgyNelCXr2J0G15q/ykt/T9Ekb/iOD5rC3Q3fNEslg59bnYw3uth8B/lDmPeB5f1M1tAzC63K8wl
5WhQBXlzNdnnUPobFcTcDdCwqbem4u4Y1AuUbRO3S9ian/XKk53O1sA3CzExftLXR5p6dcWLTDzV
Klr5Tf0wa0bAD4aIyCq8ic1fUUjTdb6kPjVkgfw82aMLNSnkmsOv248qMdo0Y1/ZA8Nkg2jQ3G+5
5BGzKvOpIXekPvLFsmTYRsB74uFBQO6LIAnabxKwzhRbQdcnC54ZvSP8DhQ1bAlH6TSk1rW1aXPg
Wo5Nvm5tZNVh/SuH7GMh5eOecOZ1SQMhoxgpWLuNaMxVC0MNlnFXwYU9tzG3UI+5qe79CzE+cDHE
8llJwE0uEQ4l1QM6lJpTA8ecBIAC6aZ2sCpKZqW7sjLXykP6mtOyBVnEI57KyoS2w3042nxD9ghH
EtAZsCKB4jOZh9x+UYrd2zSatBWJ2at8RCKqq/eYLTtMQgBS54g0UCbMR1QzUgC0cPH/w1svWh7o
UHvBOLuqQXtPtiWAJoJGeA7T77L0SnJiwDhbagQpVYN3lTokz+WA2wtg60IqmtlYiqH4FR9EgUZu
vr1ChU5y38P96gS3fuVCkTLeHD7gZXA/h9ElWFG/ZgfEs2+bVgdra2+oXSRwoF1eze0p8G3tlAIT
BgGr3xMI5UMRLLUVQCdGlnppNXASajh4d+1WU8DRdd8iGhTbCo/3F5k0Qj92ZXpR143zC+UR4o7c
4lqAmN3rRuaMR7Xuf7U95szzfLPSSOe1FlM4N8fh8GVYWr6YuN4HTwLS39IUUkqx74M1uY963p5e
piU9NGsVq4jEYVUw/bW1Gx9dxjsQNfq1qCjJA691V+xWtUas9XeIcTVD2Z1KcM2Jew47V1tkbfXp
a/dhnxijHiKN/F41XF5WBKj4nxOzBposfIR4Snod8aOgIyW+Eikrw909J8e3OvnDee4VJX8ubhkr
3P9wOPDwv6R3j1xMgpKetQ8XBhiNT3Y5mtfE0h6uZZhQws9MdP/yspFUx7KXXP2JAQIvv6oZYFPB
cb89Gpotvow0uR311dHjzBeGovSXSJWmtk10iOu2sWJKlsggg88iAK8iesRrfZEvnAwdJ6E3FVT2
64mbaVXAV3rWXCMIpTeJSdt2yOedi76CFvcM3eonSK2fNK2CPeNY1KpoU2+QzYlQJsyrGgvy50iz
RGGfpIRsmn9DjhEA5vsCcMsoorvruhXWDtZQhkAU7IzXJQJwrEXlCQTe8ZzerMq3nVGxyIM9jP9V
GvKkRERZ5lJJs+5Hc5f+X+SjkfR51ZB2s47YWTZNQqTAbIrzP12Pas2AjM0d3wz7F128GxPhJW1S
B1zp+ZHR+5jjbA6FhdvLcZfdM2ZrUXOhfwArdrB12I6WBILKphFkw6jir2eV4Q8hu8+ofrC5d3qi
TmQE8RuscRZxZDUYn7x++mUf/OyurEdulu/fTCruNv/ssj+J0AzzpH9xBRXKL7o9n+LuuK/Fh3z0
PPacpqjYLnSl10E/NgLvriz9LfgIhmEOvSiy8o56iLwRXXs7IwYNZX4nE8YtaAHIorK0b6PgPPHb
zSho/d6ln+WKb/pWuqkR1OqHHE+Rzi5s0pQ9TcMjCeNnQQdm7ZnXp1sydzqHfNxf4uDGawBWUNbZ
Gh9BBHkHj17h+gHdFdYJowa8fwAGPg+4XRR0pjxLR8QVasnbR2JWQdYuMMnMmc+WBo/JycEUswt7
u65edkr1zX11ZJ5kMTowoddFl7eACDEREr1Fi8SixPBdP84chIyytT+jY+AN7rJmmUC3OmJrsHL0
lZ2tGR0MFJPp/uinLT4DsRNNfHcWJL3HTieuFTEhUMeM4KhOI7rM0xNDVJIoyyo5xn6WewTMdWzV
JhMXNawvDvH7LT4o2q3lPze/IRjr+CQNWOEuAWlYcjga+wq8Lm0Tg0xg7VI3DybwH8ZS4QGE0u6U
N5MAgktrzZlf8veusSmI/fOTW7ES1UUd1rajFOA4zwi1ceuzDPTgF5XdXrvodbv+IKQBiR6aUy9Q
Itha+n4aKehTWCca/wvBL/UFybdZ3p9VygDPdcLTstVBfKgJnkfaq45bVyLVGAbeh2KQMLvJLIks
8RT7e1Og1U/Wge0J9ckuva/IfQWPWgcTN1cCp9nBojkunMld8FsygK7s/+mym/mfNAChSpcI3RBx
BIw+juLCH8n7eD4yd+pTgSTZOHBatB9LSRy+ydZetGALM1h6SwnHlhUUgD1DfmR5pCA8H9q6pMta
yC/oIe2wsap0qph5dcgmmk5qxbgC1vYDsLf95s4u0I5OfcoPbQtPa/r1vnKOOg2HtFasYdvTQ0br
CLNPFQqd0+OsDrXympiT+oi0T06zO6/WQbVDzzXBAmAfva5b27hJvElKKfrxpATSKfKa56DS3tyb
vMjmhfUMaJeFbQ75awjru5BQEw8JHCCLYUxlsJzlQASQBgQw8ef9FETi3LYZb5jzdkUhnC/wJ9q+
6MGhnvNxIOiCf5EZQSl/ghxwZWbpD8ABsi8d8LMcygZMqoG6MULKe2FzDHmBJdWCnumNZtTsqw3l
KkE0CJEQoAagVDvvyU+ipfFThHStI/Bg3BTOHlLaH4lZbWHzcs+iXOlJNJQui71g2CkXtngp4df+
01DFM1HHQXABqlLib/oc9VnJHpRen71g9eKHBOYJ9FLRX3jajO7XjQYkN982vGhZa7OlIUi+fyGM
2ykUpPfkjMpPfd52SFSuholYipeG2GfM9nZFRnFNIrTB1d7QmlKMovXMqgcN7SWs4IB4G5157NqM
jNAexuNOphXdkVilgInN+8Lk4Ee0gjYLFZbdwd8rIT9P8LrzZFHo0cCFm79j0Ai0oiufkMuSTy5f
5O8vU78hd9OB6LHmEfixhh77hiPzWd3VT2ZjakpYoKYh/mbUCAPPQ7pKCNi9vTwAIK106kA4ePfl
55ad07bSGHP6L5bcGNlc5CCYd+nyTAxk9soLKVa9yNkKEpdGb684YOmqxGkwT5nVbmvtnbUgyQOx
IS486/hzh2QFlMXa8H7RJlgQ1+LJE6IgQhqLKziAFwtjP3XYNgeqPFLYaMnMTgJCeR6vb0dxZXKG
lOwArHKss/Zy6KTCZfx6gmhKeEIqeVJbZ1oIHXSWw2t4u/PisCjURn0GxVFLW7tqr213IgcLh8dW
qWFHSRU27mReXcE4QKuCiHAp+3BX1CvvE6lOyYJgn2wXoltiTBpc2MVOIdbKUaGspOJ/hFf0DiE8
vAJdSCFFpIpxRxeHiAvgpmijIuak4jxnGcWJpclXRSE7HhvCormWEgXOkyRLrP37jepPdj90x1gH
OXye3vyns71X/XnA4XEq/vN7o3IM4GEajaBGXRsDroKWTEkaYmfQDPKJbIpQTsSqkQ3XzVGpUqj9
Pc7aU8a2VIArjH+hKWYhJty6hpEmn+CAq7bklVMJ7qW/U8R77hTDT991CbffOoqGJ3VH+oIxq8dp
oyk22gp93MOQh5zBcpCCkf/GkbHq+aNYDrc78/4xo2PN+udJHO0ginRwnojMWNAbel1r+VHz+xsj
YKkBodtwtEsKQ2WNJGJoM7l5E9kKvlT80HAfISt5Csvxr4A6QlYhktDyCgus5nbudNYw7PNQWt4/
IrEDei6IrELtPIxjoj7MQWUAHOa4mBFaGxA2a6M+nqqNDfBgEgS3R5/X5RBQShNVcWfpbrG9ENx7
NvZWQpp/LIXRc1UkZND45fuSWKgU++pBFdgz+XuGqJqElYvBHvWW2tzoCChh0l0yOHcZ59u4MHA9
v+InygpY3WwwFqLzSIrKNFpDvkzhW66KBuKrZxMUqgnrYn6ZBkoKC3p2EcYu6D/8PMgqzGNiPT3R
v8GkM8QBTCpjS9hEFBtt+4n1m6b/g19/OLlNBqjiHBGu7f3DGJ42gj5Mjx/LgfVuk684JTV77Nkf
ldYNrEhuvgaRUCiOsInYC/bYxkQIqkrjOuqqZC5htKClXR4NDda5VN5M6VO0ZlIHzez7lJ3rk8rd
M3LzOjCSILLyVVfAwAHPGAR+OvwKTFc997yI6NvnlQQ6M+lvV9VsDrjQwUVMSjN5ewIBMlOuqukD
YVL74OWSe+uENFduOeizPgbzzeQ1bxRwMSLSlKVv9llwtCxwX62DQMqJ6Ve4MVHa4i2LjBIDGo1Z
pvwJvvEgfEncF8GGx8RpeIAMCI4AULWmksFqvrbzlv4OjlCwwBTGqm8zFvjlRIyM5MOZkUzI0OW3
VrV7RE2JdnTzLQumZtpXsO1/BdcvVvgMGQNwty8XLbu8xeAatzkRNtN1bRbGu45IX9dC+JfRFTSj
Gszn0PSEtoSqN2GqxlAO2TFJ3cBywneMqKj/y92MQ2srNoEXzmtlHnOmAT8KWtBXBilO34V+wOer
uc2tzaYbV3m/XBKcEQDior5t8OOLBlc9NyQ5+1zxPtHBV+N+LJ5MxHke/X2UUkgsRF2yRo1AJG9n
cp8hawyHmj738JJipV8IiDioYiwU6BY2otaG+TLJlYDeIXNbNgpjWw4FAqm4jsJVfOyKMrLrWre/
d7fcXl6AO80ntcwt05Zddb4waHyus6E/Bls1zVc1rBl10Pl6mkhxDcF/p5LwV1KZJOKT7qRZk117
UolddvoLOqF+fbupZYzqxfLb9S7hhtlkU6TcxopgloZ4UiT+1HCprl96CBQlVqjs3+XXLDsFDe9v
92RbjJnavmUbYZBTVZWe0gl33ANEpXRaZnzkflcXlbpq1lLpBfwk+WTxroQIT+6swURWVJYKp2g0
u1h6fQGwBb3TOvacJY6A9kV9703it9HpIvwA4Y184fWPp/opBU8vgX5L0OQSwV4ZMBuk7stE93NR
UOgyefZON0xOuANT4Hpwk8zj82HCfJ+ByAokhK4nO36JV0p+SeOsE3fCUjSYnckgDAH2+V9Jxl40
S3UWpF+C9J88p3puCCimptcVEDHF1U01TmpQyDIbR3/BXI63RhNeLi2qYjs1J8Z/xlYDGcURGbsP
SH7H405t8+LNwAqw1WiyD87o1LR3o5zW3kAxCVI44HD/uzbJKmoCgO1mNkdPApLXL9doymMRpVPb
mTjskGvC1DnsVeFeZneunUNfLi//kgpf7xxH21SFsuByymEIq9dVIh4dsIxzM7DO6I9wH2bd8FK/
YBdIF0rMG3Rj6WLNmpDe225O6xRAOMJLATtb5Eg5wmdyNFKi2hyxiDHOwwBjfG40LQqU1MYC7KOn
pJdiXZfZNMXMEYxCUfVhqEdg/w2wDnbrMqftdKpD36+i0EvtJ7qo668ty/3Rbk0d+w3YJ1wf27d9
D2tAdv1Yzkycr/lOVt24rce7UoFY8Okir+AB5MDzYMf8r8ZANfVrn08MkK7tqPyU9yOBNBtQFjaa
dKF6tvaqIExLMeG7dQ/TLlIGdqMjknsZmkGXBzSM7VvBohCTQFF2ZqkU+eVQxvmcdy0aL7sFJgP/
NaSp9PnfBsl/HCwUOfADp0cZrJIGLi6WRC+lhuI6pfEyX3WI2B0FKgYMUJvny+Y/DHEnYlJ9Cm9d
Le16G8DwX+ytSdtWeCrGF4D/9jEWX64pbKqv14yzpbJwwa3Xm5wvygW+95Pm9Il11S66H2UCgxvJ
JAbUqc3a9zv7rieVPvmNbE23bYe0cv5pfwBY/b7ovJyyt2TTa/4brQU/xBZJ8JRoO9L/hoxVVpx8
/wDo3tWguisS2VJ+w/j+I9PdxpmNHMtPrSGEXdvtr0xwAT0hhenrJh+/5hbtBdWioQo89oHrV3hc
h6Yjqiauc0j1fbeQ/T4Y9PmSQG+pqRH4mwTAgpHDHkGDueSLo9kebC5Btm8WsuPRFwdQHXP7cv5f
y4bwsqpMeoFTNZr469HZrbvr2euCuZdIdQNpBJ748zKDaOZaFJzXjSptZL1u/Yk3msOaasnKn5mR
731X8cSGymnEeTxt3Db36Cto/sXwv16IVngJQ02aXwSVbC+WzGsJKW+zT8QVcIQNT8JHYSEoBubh
6EBQRQnmG5LbICopXxkG3J1Jt39ajH3wYqUioXaivpJAg+92o6lVvDwnj3RPWC21j9LWXkno7VeV
nDKwMBVxG7uWfky0Kc36L6NETVuv/c0SoineUdmZp+OR6frGHvpQK7MojaXgwbke4NQYdZYroVIZ
NtxKgfoH81Z2iQ2iYp7wdxuvLQgfg1J9zXACjJdYC+U6lqgBogQYH6GTqSAU1Tp6ro7iYL8Z7EzE
Tt53V+F29amudIP4Ar62h6RnhiNPcSrz75DtRoySVNTSGJIqCFVXhR20wk0pubaMvF5PVwOUscUv
S/KRXzIft7qJDSO+osLG+eHX/RnulVd8TnhH3tHBzphv0JKWQs7ExWSppvXgLNQ6qMmBPvQIGKj1
d0lgN0PHdXC858QOlQQ+mO9Z/8ZztVX5eiTXT7qo93uuknLBj3nrrUAC939e/tUQvwGYi2jh7/E+
1DmODkatvHxRiyTIzC+2Mol7kVvICYLUxlRXsXttk7qdP2yPnMDa2QdskedOBeFdf/wzbx7SjXB1
IgnEeeutGFS1wNC0C/+EB+A9Wr5bHkE68gLA00dZYra4ugn1IZnRMg5z77QSCvj/v5XtF+4WBWEv
O8PLaOkyO4jhjXVgXI2kWhR1NqcPK6nUMwyLx7Kr9AyMJ0A8GUtOMpq71SLxMplRSlZ8aEIHPGxw
zcjVRf0hjfSougFd6Pa+J5CONOzNH5X9KXai7tR2oOAKJoo2B4yDAp0TCv7cUht7Y9OKo8N4Vk05
ssGycU+Eqx8TIiljsnV03DpSDEmNxEOrO7olnjB5jI1U6frUwiKaUbgNWLvkI4JQeKdv8aznMCg4
9OxtGs9Vt6Xb9HfJAi0LgbYbH7TpzrcryK18mWOcF6ljr7Q84u1WtNhMtQy0JQuBpvBWjenOQt4M
JRryyWTKwTjZhHWIL+AxZejEuiVJyPNI1uqrWuKnuM1luaYRBX5PABLrR3WMSaBDxIdTJ6/doqVA
lNJV0H0BTkZYNnMGnSOxAOp6eO+SF7SAow3joxZ4UHyTIqa1Rs2L6Pzk/KiHzVBxEzZJwknEnABx
/U0agAzYRRPuJaolsrLbKKa6sbESatR24sZy1gqjeoos+KpUU1oQ9FXtqy2DteQgb4sGfzc86HPh
yQH+CUrn3/+SiF3JkS1LOQZt3QEKrQHSRh1PkU+Xi9WVPqis0YjbfspeM4vaqmOdXIVlfH/iacL1
qvzykyBmquQZmqa+IsunJrGdBAOMYIaFQAnie13PxXSzjPk5Anx0UvhJ5va0B2ySg5M4J8ce2iUC
yD5THIAojcPOKzZv0vQTlPyuPf57XYmvUTbicFhcI0O/kWX8IOOBSGijy+QcHLqcxOjpqxwj728O
HjLemDFxPo14I+2zb0MmPm3HH2DzVIaO8wcmnqWBgKUeseFPUf9XoR9wbLmTOWm1ab33AL66Q7OS
rEPN8MW4dx0IuF1uRiPDcVrweEXI8UZgNdxV+6D/iIXASK2DOOCYkF6snkUOvOMa/rP9aYE9m/YC
Uvm/GufjwJ/gvkRPz1jJeLhArHnuCjQftIQ/vSIX3aRw5BGuw9Ro79XH6PnWiPeSaUb5ieDBNlcu
n2xAGsuM9dnE4R0huakHK6MQUFGt7GQ14z3nkhRfYTZkWTxIE8QbuO6uQY4FGPVNWR8MxRXsn/13
f1XjW/tuTmhKk5M7jhgWv6i5IrSQwskcRAZvz2SroRr8pYaCyVSHZFkY0VpGUB7o9uiVPAOrNQ+4
cr70Z0c4C3mhlTOos0l7cXMa49ZmRvsCrp9ZGhWIflhBpiIibAjo7Tbf++X/rHUNqIgcXxqMadhs
lpBYQMLPpYkycRR363vNr6kji6GdmdqYWX8BN9rB07NKyUL3XrX0Izv/kSEZedAurQb5h0cClLIF
Ccm0X6tcQl3tPY8xo3X6e0/1Ghgvsy7h+/h0Ijwqb6xJHSTmvxVtGIKdFASxPXS5FNWveqqQVeKT
2YVTktVUZCHCYQ7cOMIgT7cC2Vm2XaALZO/FiAZO0ekN8a+6aJV0f73FzoLhZcVJmMgVcy8DxNdy
qg1I7x1Ai1ZYiBKmdmaz/ZEAe77R8pLAzMqcKNWEs6Lk1v/BMWf66ENY4usYE3EaWK0jD52zjzfE
dCt/uLMlUsNIhAqJQ10yMIO5zT5spdua13GKddXVuzJ1n2UYvGaH7GS3Lw/Ndjl35noDaQ1UjKxI
EdzuuyD6FablGx5qh664OTSgkkUxwQkKphdUkYuswFkajC+gG8FWUlEH+8hdDlg7mgTBj8A7z4JP
omrj6JNI1UWbUdfy6hkFupAQzWUajbeL052h3nA2RVgB9mXZtMlpO07KfzGMgqbs0qykvlpqnkcI
9BPqDUtmUAJZu1KP+NVDPgAdB9dsvp3e8h44uFl0GIB5rtvtHJJrbIyI6z+ti5sGh/e6n6/18vnW
akjIqVwpyhzLVEg7Nc+JbdRBfoHuGM1h9JtPEosrRJrcghjwi7OUaDCuzQP+eS9n+uymhk03uD81
4r27uZj3wuFHNYpUiSaO0NTzv/Md9mDfI7SO5/qQIgCVtpcGafXiBHbtaO+b8oWsGDjoEpEhINWS
2YKZJDFu3B5Fz4cDe0QhzgrR6xmuY2JndOY48JcKpw67mNwXd7GbuR/8tqFSyjOkVgw2xuY1JGqZ
ZWeTc7Ri5KiaMd/fbfTt4f0KSbk/Cg7D4NFeVPXh4CW9XwLTq/Tj/Xfl5K5snpWUVQ7b3WnkjHuS
2Wwp30tCgZymfaE2lT0rqF/6ZGVNZpO1wJX3N0KR1o4cBwIgQDOfSm2x3CYV1B7oWJIlTsW1a281
wfnmBh1F/2C7jPJuBK75q0Vdp1K63cE+swTiZlk4/bI7Oxj/PJfCzvMyMHxFszCJVqpokf2nFX2u
0Xfhy+HEou1FRJrJ9amKSACD3O/cGPwE/WNIerhmpxcUk7Fah1MGHMyhtxxpxUHLralCjARBlCYF
ATfXpTBo00cgJWMhCQJn1meUfC7buXfilmUF/ZOF3VozEaRn/evR4MXbC9dUC3RKFhKIljSHrdqq
pFbgzaV/e2Xtg4MmxS88rFU6VKwNKhXnvx7y3J9UK0YtOdU3wZctdvEAlApomHkqQaW6Hdf997Tv
5wQODgwFnQoZx8JrKOGSroixL5M/3nnntce8xeCEzIcybSo1HG7wI7lHBeN2MNnhn1gnEM/f4AuY
cd+yI430KmekIsFey9fdbOdmChWV904AGjNAC2KzIZ02AXG9JelXt8Fkcg4iHxfVboi5NJ1tnP5J
azXLC0KZZuWGXsCdFQefdNdukKkpoOVGjc2+oR6KQ3v7dbR65LaIsijYD8ClbTeyv5aHM9VlObF8
BbDXwajMFL7vaM5OWkpXdg5ftGhqlIKkXhHy1afLSGMJrFdatXMULzClXTK2ptwZXQw1Nfg+/JWP
BkraSfLy2rF0YzTNm/2BfpPHgOywLRo4Y3RL32H15rrpN25MMbsnMOlfVIc2jRtLFhkXWkr/Tvxm
+vF4T6b93gmAM0okKc/AZjGZtpKEoamkLXjyi/UhvOPC7t9Mv28L1WDVD7oHGyROLHSTrlGJydW1
RYZJozWD98V4/VBlF2/0K5hYC61plm7/PwGVDOHqpIXTeJ+OXssnEW+eUiKZXANA0BmMtj31Nz3i
YK1Nuh7PtOXB0bpqIiQPbn6xSW6Z3cgP3+uRlZcvW7IWI24DtbZCNHqm/4nFUyb9yBMPtJLOTQXe
+DpFeqy9t+ksCkDh1c5mPKYi54PL6DPeDeSLzYu+67CRWT3VjmNnekEFzfPnn15XuI5QMnExPklH
FtAaaJTZCjBIIbT/IHXOawvswwZCWAw8pXQdJ/wNZQ44aj+mbMEGdZdxaCfqwtA7NdhBdp424aap
LWVdv8TaZuiQ39mlZNx5viow12n7mLW0gtMie6RHViXCrzKA2f/8DPdad0Ib0qjjfFrMzHiEGHRW
yJXn0FR7f2H7MIU7I6XOmYYEmxRp18Pjvjg2Y4PCxLj1CeeVqdPa/PZwKNhduAl1Ue70NeKjq/C6
MgCDNteR0iQJFWjmWZyGo48QTRZT/z696FSKoUKbRO3M6d+hPszEdA2dNf2l0/AliFG4QTAjmUJc
aIQKYj5sdoWEbW6MQq78doxb/x7s7m2awO1izkX9mOdhfZsBzUEdtr2le6/5Hj6Y33zGai2+ogBP
+9UIBzJOjfCwQ0kq+dMVpjuPPzSLwsOcZxjjoMseePih6gPAPNROeooWQr37bGiokBm4XwSYeiAs
YnDztSi2zH7FblOQxDRU5N4nhAoPqZnn38KrqJdae2gR9VjZ5C92Xrf8rX/ENFosMB4tdGtTE0eg
8PjjWRPXYkLi6gqZJFeHW8/v0hJtPJri4hhWPi18iYO1VMWib/yDaSFh5unq4S0T5HwUqENUZRZS
A1dh68sj+nlZ4Wr59gO62ey/rRv66Ly3mBHBXpCH6Rbt4zL8dPkJbA1KzoNsxhbZE+voCKUpVLV6
LTlNikIPcqzfYEVvw36Sir+YXpxZ+kqZeY1NwMSMtR2GloKKe+/1vsI1I4xXg3Sa0rdjf4jDlY7I
jZu/vqh2UFreH+VGwKoBd3JcchNIRIwEpZh7do8M4AHdwk4Fwgy2OAOUB5paFlsgjher8P5WPqBa
/KXJyr+sYfVNV4xliEqHLkF46ls2gR+2PiPZ3Pm0hQsuVJaVwTz/q5gZTigpw98W4ZZlIuikZJRZ
RVepHSD6PXQmqyKVF8zIq4r438ufW6MN4bTDfrchlR8ktC6T8eOe1S0jZ0dRhNSMwYILA7hrUvYA
wCUeVP9YKcN/BIuFwuVUrVK8L5E40kz5Ki1WGHXmz7bhMPiv9fAFBiPSpixWg0n4RHNYjq0iZezj
RaZNAMKaW1zOEty5iiYRfqq/8l1m2aWN5dL0Ge0kkOYWKoRDtCZPQm4OFcDSWiNFuY6+JD17w7IX
Defq47SEOAhkAKmnvcMiDGtXkDHQRG4a80YM0JmaiVlLHf8Pl/dyJcyvkArxISYqWv7O9tO133iI
HUlNeg6SYC4QS/1spjQlmlQ2W75nqBBL+kzmDfPPvOZDiZbnHWq+KiJPUvYR6UeJY3G/crIglRmX
JT49z8bIBjgQRh0XQB3om/CEj+PbwqFKCglSjPhD/Ly2w06PPXuC37JwsOvz6NBajLe5/22j0EBj
4CEJSJDFqCXi5ETIbVLIi2pO34LoUL08x6Tck9J/5YKzfXraySW0AVAO4gjuV5sgDlIaOEVgXkUP
7VBmQPBvbFeFCfqXNj4kKSWQjxQIG6ugZ75xTnY0i7i2e6QZ38hZM9gOQTGCV1wdcygGFhPzv3DB
CPcJ70/Sn41em+9rbIapxuDBzDZaujk0vaS1PYUEyfZpDNaqj/UUiEwElaRiAEK6pSxDstqkQRcl
mY/9uru1SRNDRXAB49mAcnayjWZN9h4XUrhNt2cXaQhj9/kshGLTKosGJESX33yrsjHVHXIQ38lf
yDU7xEeki5aS/6bcbJf+IG5RgimblPRhxdblymyAF+1LFLzjugSdiqTU0lNw1oUJp81G+KPuzE+G
xZ6yGcoxGK8eLq+xjM0z90qdVVWvuN91EvkdKnn0BGGE6TEcgUDu7cIoGHNnlaQaEempjcqhq8SB
v3GB7lVTQZC5mSlUw/fRAbshgaZOre4LmFB3TcPko5S6ExB2GGIJBBqshF4vfqu7wFuy8Kbbr+l6
Dx4AE3DKu7ckY9+4K32vGXYLMQWenmq1dThOhnwPej6LkbR1lc1ftvQboTmS//N1lDnYLmaZP/xK
OqjAFxmdwJ1B5zqmS2pPJrjZ+FQ1gdB0cmWttEmMdMTecC97TlKzgZdczi+OIqjFu51viwIywuFM
0K8LWxlvOQlhPlYvV6p9/LavhZnx0e0clcRDiiTD/o6ZYVENBviceisu0KQTWa2VnltsoH6OVe4H
eRRqOdAT/N5rrK9jzHEEBNUBmYCnZPNfmw5MEcFkNhg1pzuNgahsEYSeqfAE6iTcFIeGfhtauoap
he+L33XlRvMbiIyZ3XGdagqspicNrqWttBWcxlVqBo5jIiyOc9c+rIHKWq8SBuL+mwFEoXtJCJiJ
5Vm2XqmeXl5g4/7SU4sftn/aDIXpYnBLhdAuMCpY2RGc5VQQkr7TfabLwCG1wUV5o4NSn7NmnZar
IVuBfks6fe6bjRcViUZgJW6/rtHevzzPnc9ASUbzHs6agTJrA7Dht+2BvxgO+EilYFJ9nJPP6HLL
BI903j10BQznjBTv89WOMaDPJBeLDsJdM9QlAqLieHLhhJPLmrEiCZqRQ2rZ13CXUY3QOTgWBfY3
jeTtYC/qElMkaIn4FvvwUWCtwd80RDanKHHaymKv1GlHBNAutgNOJ9OyvjIKQnTBSpRymsX8OtpR
q9RceCCBtcG8yccDaWV/YXwvFr8BdhQ6bh0Av0LWz7YAK+JIC7VPecOdj/Mec0Hal7rkVb2mPIDo
aqI4nxxF0E+uxUOnYbbbDR8NhfOgV6sIRERIFeyAE6xHDKUEcBYIUc7mBDR05HpYfvAOXOHggg0d
3VmYXKPLZVQCvOFbaXYj3WKcHHbmVnK7ESyW3vIEaOR1C/4ZrThexPscShyfo9n+Rr8Sz3t0LjRD
n+l4rfjY9ijMzmdl9K6eLzSA0Bbhlb1DIjxmrMjBX43SoTscQifVaSL7WiN/VAMcIyHmi96g8bTL
7su4Xa22TCt6qrTVsjImSCkG13mix5ZQKJfOqQN94/nk57SgEHC2nbQM49pBs8WCO/h80Y+ro322
CwvbniGGoqlg83GDKRac7o+4iBV1N0pDgIYmw9Zc6xRj+rRvJA+228dQp/cAdlWLLI7gVLMjKYVm
SSS3yrY0FuPNIdfkaZEYXqgHNldgzaLDlOfql3mer0h8z3+hON2iy5Z+0EHFmOoSPqsm/RebJVMn
tzUiP1csMkTi6F4zp/kPTXthIC/Wglkd9gRdJ924H6H3/uhYZAeMPWX7FU9lSqtJinqoNz/2vwIY
N7fDGaqZNNsV5MjnruB7cV7jd1P0IEupheIWBg1raKWBR4UVB8Te2EdRbBUloP/DqAMUN5qKVazL
OCr9YRnb/6dZbRaKggm0uiEeb5AhOFxe35VVeinAJPbUsZHKlzr/XLJwjvYtmPMInj5SCfSb7JF3
fPLF8XciMA4QdeA6DpPfdAhvElLD3+IbKheqYkkiAGBnzRgSYzWiDulZmS3eXTZTCZrhl0OyJXZo
BX8RXI+LcwzTMHpZUnVUc4rcDLvZZhbKU+XxuUTHtykQiQk/myGu45H6COC1k46f7QPzfh+fd/g0
LTTRB23IGv4hCWc/WdGKPHvpO1ruz/3bDsl2Fvjakqp0RTwlv3ao+WWL7BodlZKJYDb84HlyHsD1
Vqh0K16nNdAfgG4ENXQFSon8PFnG5jBuAe8OP4EBpczALjVc/VJjeEW6fDxeoZgDl8SoT2YIacZr
wfpPf8ycXGDjNY2i2XAql1GAY9ZMu+YH6a9RLceaPu3ds/yIxlnAtNGko5HSZWFHAOLjp2w/K9cn
EjBzRJnhF0p0VxoTPd3Yisr8uKXySqM07SbuA3JGH28PcWbfLZ8aGqlY+lLiyfID4q3L0oy2qwqA
8xXxu7iqCWd/H1KmJgW2YOMHeQJ8yE5vHC6FogGUzuPw8gJxX2Fa5MkjmvuSydgOK6bsE9YcCKIF
A+IFcavyB2kYHF9sJOAsuiDOH3viMzGMg68D0J+WdHGP0dwNR/NldXS+cA5+F7CCqyVUIn8qONIw
xyo/2VYSDOASsNSwNu8qr+imZkjKfR2UKjiMW6Z6VpO342GfizjyKZDVu40CYsKG5eq6hdiw8QRf
nLsq+jzWv5gSCQkY9CHZO71JSfQn19pVThpLELVqphtuHDmzURHyOXDTznuBXae8HUnROEh6Ke3b
BDqppcQoi9lHV7SujsSo6MiQxAJ9R9UAr7k31i7uGkeuLUqV85Fx1KKRz1GaWh94KA/OamaiT3Lg
VGlPhAWSWXZ6IvuneyR8b1UmF/Am2h2lnUCTIc7xDkgHPCHfIp/r2NDeoYk24IRX5GrKU/GRs7RM
4ihDQgB8sO8erYjM+FfdSKJj77eAVeowVB3W7WYG5a8n4MDd8epYg4GRl/LXWJvXKcFDDvDlICCn
wVMS0bY/slGF6cZw1KCnxTky8YlIgX00mK0jS+w+T5fCWKXmB9dN89g/qfnrWvsM+Te3g5X1oEnO
8ZUq2KPN/bpVbVdNWdbadeLR8KmuzSE/+msmMv57f2hVAO5PneKKHBdE3a169jrhFDEAKLlIrq0z
4MSD36VhzEdEqWMpiZ4PKQhPMpmHBGmQjLO9B/Y0iY+DimfuSh7diVaxFuhDW855+2VNEysFMPWH
azjZEQiJrhWi1yPdv5vEKrzj6pwpbFbn2FTzSQw2l//GYLHmVmXrZK2SkBoO9BnQje/Sqswavg/f
6Uw/YBdPxBfigW76v7Op02BCr7V0b76roeqMMQpcF+dd2uMrQ/BOIOEerumCZ36XwYvhXALtibP9
EK7UMgqiZhtRjPOMcJvuPH7JcdhpCLyepomHcCvsT2xllulfAC70Y++gI1XMt+h1yBDL7cTg3lA0
W4uAarW8P6HdsYXvVrisC7tEElokyi+qqMCfl3JzdUscMMqH1TLqyUtnKG5P46cp2T+Btqc9s/OC
qdagWQZD26IJ70oS4fYeCSbCNwb56ThFb36eTh5WqNTZZdVv3S899YyeGxyrH1j7RqydEk3HVIWe
wSP0tblT+9stH3PyWLjz7shTP2fZUYF/dHNjYUmJjVk5Itdb8Nr5LYp9c3U5t80yKG6OTTmLL7Yf
1aCrfpa/2N1Ahdz5L8C0UM44/iuJu0f4E3Beqhkfsqn0+8TJ0Q2DmZ64MzNoT83gIdiAuMIXmGef
oi0gOZv5dQrZQAaNGx2ObRy+O0HYwhtaaSksOQLad24zJobDriBTQFd5c7ws1tilZ7KVtwBUKQ9c
C3FMQQj9zwO5EbR3h5G6kPT0K+1sKdIXO8W/tDAqerQkjQ9xvgp/uNKccn2/WoJW89gzjeyT9nTz
OWYJRo7fIbZAz+mQ93d/2uEuON5AETRiti0Apr3TS9HwjUx/EolfVIdCsN/nSFD9wjarAiVTQws8
eQHY7zBwRMAv1gEXmNhXezKJceTgHpViHK5peM0fPiF5urXzyo2k+p+endzuRajemQLq7F7t5DKJ
joKcDfJF8YhcbP5OHqlLZoK15tTFX5GUf1xuxmBveS/Ky+aqs5vRh+iEtO0OtU7KYgjHoPrNv1DV
U0WRR0HdZTTFDVxKBd/SJW6Zz2pmFtThh5PIkFzWifYZElXR125p2wgj4Q1cOJKhH/Vy7Aepm8nR
k4ZORXOG8YFIjJI9JOZEWutz2HZduHqs5yie5l8rV/SytkfCPOAYSVKfDDO0hrq7BPxdlEXzj47z
OwLJuLUzkBMTGm+yDEw5VwcjfkHYd9gd8Scuitoc+1DyyGgTxrz1mHi/NNcT8/EiHhZZ7FovSYq+
xpxKT9oCJ3B4AMPtsuM1R6rFygCr7JDZFYm+Bn1qjOzHADqFP3t+YYGH5DU+McUELTB3KWxz8qNl
8LWK7NnBf1OkpC+it1nLfhmqoARohzLUyutVTr9OhFZgnxUZLh95ozQwxQjvown82Hkgrc6V4ze/
LOvG9kRlCr+NFduUq7Vjo3+YQ+oRnoHVTihPAnJxUuc2PqexxwDxelE1lEOTffCnMbA6CTh5wzwX
VKdtt5E0efUoBIADUDlXHSG6RYX9zi0KjGlBJeK2g0iY0Xf59TCa+N3Cv6E9WAXxec7OAHTNf/W4
MsqAwiOTvpRm3SEjIYbkO+ZmL4BxoNQQgXhhvX4h5cOkFBbkbHiTVyKFdeSczkVJoj7S0WDwzosh
9f+9wYcHgoGcn7G+34wGAUL6IDxWbAFpVDSQYSyLSQaftjo0ddtj0ihUpvygQoiHJBUPSyFOL2Dl
1FEScvFOvY6oEfl1e7dY9TNB1XIGbCFPfp8kRunRlUgym7DZFgLSJ8cRzKqeMFjWuJvKhXQQGGeX
XYQVjPFBtlKr8vecDKYfc7+UfKrylyOi+0l77P6fh50skuMcuLMwKad9A95GgyNNU+dToKoUUmvx
tiZxUq/9tekQIvrOuzPbYd5MA30BhNXiiBsPgDD+TmnNeQUa+yHIVZ0tSLT7YEMO3TK+QYXa5H6S
8Qgds7ao4kWmRAc0qvT3H6USiy0qRo9LxTB6/bs1uKC0j1C6mf2eP0KItyGFSHNfgRV+YbJeXaAO
m1/UNuuOdaeHD2Jtybc4cuvUOeZBlXucZ0fFaSx1uSdgTRjQ8p9DDnVaSVsSGaAwlV3bZW+nel6s
ezfjvZTxBPsQgcz2hfvr5SAdvR88lmumIquuizxrOTReDs9R1H1oJXcnMvbAenSPQadrHqWOmuFq
piPtEh8rtYh8ClQQlU+nznguw9ZgPjulCp+D/6LpTfO2UPmtz4r1Rwk30MuKJp6aUj6/z69dAjl/
W46w42f22OqSPt2t8X6E0p2fxIwbLLkR31VrEt5irqxgn/k+LQ7gP7wJwYzOr6T4JhHIq3WpIILa
pRuUAROztTS6ERjQ9xoede/M0+gBESwxCeLtoTbsGxARNq7Vr04fHEOR/cw4wPYcBjtc8Rj8+dEA
vpGldsXTwXLocWP4r43OgdliQRKL/ykVE+LUtcXJ0lr/6h34/8UcDiK2g9UR8oQOnUWrJh6qP+0I
JpSo6Hfoje2A7Int7igwtZMaMEQHbcU5jxI+X/c1AwT5LZrAr0d1II1NlNV1DabE0s5s0dw4joPd
woEfjYEH9yZjjw3sEWBTMXEDqDyr0EGN0re6wG6+4aoLYUFydD4wtepJsbiRM8uCtHBxfD19FrWs
PIWgnT8+COKXNnSK3OzfEnm++KSoLoScwTr3dkxsGoB7PpDmCUnLTHoD2HEwQoaCGxmzYi1Amifp
4VQUNmnjXorOPa88JVGeaKa6+HuB6B1CJTPYCbOklq6cqMPvU6gzMslBbtp4+hI/+/8HUwVlsk4H
Yl4DHiH942kzRen9X4uo+l2P2YQt4gqfZKqAzb6TYJiuDg2DG7r7+Gv980YqQ+uyaVAzG/bVtOZG
P4Y1MCPdsNA5uZ7CClymAvR0Fu5ifv/X9UXDKmDUHxSVRk6OoqPOXbcQ58bmHpSQHGyi75C9RdRw
09hR/1SqmfHIeTJATUfRQwUnwi9r6uu4xCzJfXG9b8NiXNCVCOrJu3cINkdq2MiUc+04V00otNNN
axzf2SgdldVqkQhsOV49r+g8auEKsjv1z9nn50RuCSDClOBJgMhoU3OZ/r3BS+Kv6/rpbsrS6S6C
eLTZRqttt+Z0t+suiCWVTy5qoCxmpj8Ft3I9lFpX7XeeXxcr8m3t17DymfvGSHKnx95vfGDJPhSi
Tyqh2yHLreiKY/rGXp2bEDbwPGFXZ81QN2HAGDOmHGh2zWENlRTsPvLCSAPQ8/x3FtdqI8oyZCN6
v2KnIEr/4TYLSsIhLfboSSoPr+e36gGNCWpTO0RQZoqSjfzR0V5TkpId6+pT5dDK2rZ+JmKF7LqS
gPGVg31+fOW+mmcGpxGFr5u30SM2gpGaBtpkkxhH9V1+3pnETXGFGQHGdGknnjfseEKAsZsAvd/O
8qa6WsDIsaVtMsg4yzGnlT3+vkPrnuo+b3uA5knMaMz75snbK9CmvCYqn1DyuS+TeIizC/d5/7Wj
m0SfIWFC8LL67etaLx49UODXSNPjS1wn06Zg+TjMsbN4vnVFRKfRdPftbY+OHfITf8W/ISgbYesG
iLUnCLqaldTkeQGVrqzalJ08buaT5M3Dmrb/xpG87TQh6PMITyR0h7piFRHte5whhtDKVTQa6zef
cohrkqssy2uSqohteT9BOksf5yjXDTqIVoTgiCMrQdmdAZGXaerHAMvNTfMFfkjOMXmm3qHLS/r7
wx1NVEZmqv07HAQeyuURasX09momKVTTnTfcVzwHQUan/6kUowQUdtz8P00OPdAlw4rh14qsXpFo
jdC8zt8IcK3Yo8xrFalyf6kdsR0dno7XIxE3+FtcUXsCDAbG1JWlmc+FbVLZSpl0X1Wf/wM8VY3P
iIRm721UhmzpcxWqBylsUrHaQkYcSXBeg2oU09+iDec9n67kiSkC0l9xKjX0gPyCcU1ycu4lFivx
b58QylXm6u3qQJfJSCsaytTRt/1YLp7zpZ2uZy/sMgvzQ70OAudw5UtVABc87uxQpoReNey3MJtD
qsQyG4LgXMRN5HC6lEBdU4MwNCkC6Usu3r6GdbgsOU1qlv61UGquHkTvFN4IhuRtULlsbc6fBoaT
8Dgp48OPVMKvjM1u00dnDKPwGnHPVZm7vKqxYxluhxdKcbstxt2HZYysP+IUIidSDizS9ziS8fXr
CnUjeaxIHpDtOrY4jta+NVB1/kpqPgpIg3TJ45JmETPRLvZ2xjRg1ed+OoOQhWiR99gckPDSZ3TJ
6Zc7kH4a2K2w1LfAMXgJZj+0oHcTE4x4yJLIC8v/SH8+lqqH/Xp+X8EN5rH+cMLEMdEZEjNw0ayu
AsMO9sQVLjiQNNGb5R2IW5mvMV4WK17LCKlLg5KkBLbnV9FStMsgcZEsSPBs8oSJll9i/RjgIxAM
/YHy+mwbe9ZUNBDIlK74B30ZszHZxpLZd7Z0wts4BddsvY6pWBR1BnyvSEkRGe43keYFVW6V4IaG
8EeH8m/Nzt/r/hBhwLMSMcdFF9d8PGEJVOa0zgKXXLqw28kpoHF9uTof6s2wYhy/xIzbRAPq2xz9
+bu/V45hhU+OHZblIX0XAxbemCK7XDVEchm2vhEeeuz1QXK4fNUOzELx006qkod57G9LVHoOsSVr
A3VLXpQmbVr/J7AzTy6juoeGL87kCdUlVZGpznibnXPvOocoppMCnf9WDKk6kSyKdfw32NXHsNc7
8nYbvtG6ncPAkuqSq1QOi2E4Zg9LnlDii7TMy3K6zfoOWRyuU5cuLlrsTqKvX666A5/o7bGoUIly
BaHdH/0+XPeKezTeY1TO21WP/lY/CJaMkwnqLtJSuvWRluvACxYceFD0EGuWEPPz2IZ2+NQZjMwM
Dr9UI5eW+Iwr/j0Q8Wa7zQav0pC0CIAthPi0WT7oZkVLEIcfuXzRSd3JbPU6equ9SgIcFIzYiQla
SVfNrprMpu2/MqCPrj3nD3Shl1kC+3/oWsQsRqtadaSfDNRMmg6CO6pjQqBTKJd7jQM7KOGBIGUI
RKJIw59Msk0Brpwnv76ZUXZdGLRQH1EHwMSJ707Ahh+HviAyyPtDjT72LeZmZ60Xm/kyjgnCs+SA
yrsds4NOIMwj4VqQGqGNh9KAbvL+A8ArDwbuhkKvtM2TlpE3ZI7iEpUkDEUFeWhiyCDZhM82yM0K
xN6YAY3GfT//6jOEdOIeOhqqEZo9rHKL+ZwiStxt83+qbB/jYC8pz6TUWu/kzjtfDuuh///Sjdwf
9wMIlTojeMixQvegzuHL0/H8mxXdfjbM2rDGYTiWfsR5xP7vqKHUCBAutQamgpAa5CQLppquH2pd
eW8TJyi/z/0mvoYFpawFcJal8aHHKh6h4/MXc+NoGYkWQIoMHvDV8Y05LQk61CaUU3ZV+GOn/x29
WQhcK/RjIBtnaNCjMwNbKjKyM0HOTXPT78YkNPOub/O9a6scTCsrhYHkBV2Q/GWlsSlfPYK9YkaS
MRwP1Cr4xucc48pt9cRcZpGaf0L2ikOsEpap+lwolSyXlXuaQ0l5Vw/hof4B0mctNKezVxA225zv
EKM6rQPBYUQhsgZyCRztLx7Mz8ywFUi91qHf6+KzlXzBDCngdrCLWTEypq7/MpUxt/B0Li1aw9y+
++pKZ7PYSSD352aK+7FrZ3ZBwoc+S/DpaXiC4v31DRilV09MjG2Dj4pQEr+yFOLusJXR8O5mg+xN
Z+wK+cSdywsqfGjyYLnlZfiMhRbkn7X2d9kiarXbcfvU9T9BzK1jrqZfkqQX5G3ApjTvcvTgRRWg
PT3qBv+cDhcCVVPLn9PURj/Y/+AMyNNFHap/GZuWr8hqgNasbnDDH3tq9qxUlOiFperieASlfzT4
j9D9+j1uQZR1uEiERq5aIo2izeGZZ1+TpFwTknTYAoZ6UzOF3M4Y/aZRDXydMhXI+gbqZuEFBF1h
F0A+1Dthr9h1PWXz83TrJjs1OD4n/vk0iPrDwdr21uwLGOqjJFKh1fcTT7zfkWGsyKfJPgB3Me7C
BBpGqtYFiFGKMQI2xMQSpQPUaFEMuhg+TLnpyyfdK9DZVZ9vWcZ4SS0u+Cp4rVqxVDo3hwNitbHp
oKkNE7CvlAYYduL4I+albHPx5EkX6DKuQtobihGHbZYiP6ZiYmpbggBZvEtc9wa15wZkUNRVCqUj
wcbgFlw0WjHAto4wjxf3aHHHLDphIR6K11UVVsyFuLAFA9Pqmc+R9E5+C8yNw+c95tOC6dwiZdRO
g/88imnNIS0Kp+FM8VF+u6h1/LyZOemo7xrz4JPfx/An7blNOtKcoR6lVZjn1K6e/lBDc1r0BY6d
SNqeXeoFZLKQ/o9wr3lJIbSgT+1FK9pd9KWuPBVnFL3lhIXIg8h/G2U79s0RIVXH2fBxYTO7p3qq
DB/oId242TZJQ0mFrt+v183Nqv/5YE/S4bMzWAjh2E/D554hpxgkQjtjuIUh3Stri6ku1f7leCnK
8uT1TTwCm5PwyX1Jt/itVGfYqk0YUDFm0wT3wzYrjGRmIdbZHjVp9cPUSWc+1mW+1byb+gnS+1xv
40NvWmRVqqv1RV+QAdRu8A2CHWTfCRYYc2C1+bXjhAYLsPelK2lg2BNVKTTAgpdTUkRIwlXqj9RO
fjl/o4HAkvHVDYIE2oDfmft8t14sxYwUeT8diaj6VnaGX+aeekD/Ihn2SHWY4g6PGYNmID9D+EC3
S2unT+zi4kHC6lM1hjlKz8Pwk2V07YxbBjGWhZdavvWr4wJIfveWgHLNvDx3O0CxVuG8u/sPikiC
HN3QiHIo3oJZH+NJFwIAzLei0WN5PFM0aRtyBNo9OdNt2X/10K0NzZVa0/LqIADba/nAt8v1ankS
DolmdNwtx4nMl/NxE6dQUWApzkgS7x6rgXF88gE2Sg31zvjwvik4Oe/3QwZVyQ1rDI4baAv6c8sj
tn+IM/dtcZFqTVKknCsPiCgrSPhW7DXNU40smcIa6tru6Mc6mRJvqaMEd4RM1HQU+i0rpMFWi+6b
Tzly46aI4hU8ECz6IKqYREi+n2ZmjjglYIxjWvuiVD/ZGrsudC/75GhUYtfiPIOvjmWFUVhc0lAb
q/f5UXU0C7j84nedgOeSJwbBuqAECjlooZaBZLl6Eq5vmiy78Xh1Vv+hwD9gIz9EzbNIiktOnpNT
GM3NIbxvoflNiqGU2zNeI5sRfvwrSCkOBvG9wCk9+uZxpuL6aHApD7Ng4fE6jwALQoh8v2K/tLD6
eU0fr9wnrh6npienefT45c1Q4p7rEK621dh3Vj7IEZviH1tDmrRoDl3ujNyyQzrGqn2iJyq/6/Qv
c91uPe267o8YviZURltqJK8U/nnSdJj38jWEOFu7cPWBMFlgzod5XNrDwb2dky/Q75Xd2T9TicAT
H0IKN43TUV1N1Je8D2cIFcls5M4FSaTmSKOcLJQ7YzfoAcWC3e65HaZWmk+SOnI8IHZcVm6MhC5K
j6YvRmvHrzh14wDP/qPMFaI59zi+nI5+bl2OkEaDllrDqOXP6D3CNKIakW6R7YGCzmpHRp7CJx2m
CZUYJfwbFhDmblWAmzLrRq6hrkeJZUHVfN1Djr/GI97stONJTLeuajXh4FkVUDXTQQqFBHydbWYq
aw0b04CZF0i8Zt0E0YBU0N0kIB2fwk1EK4EfPvGBAZTuYrX3U92fUzMZv7ygrrstK4kOyXKx0zYA
P50AJ+tUPVxqTfQkSEGQD6eR04uCEyrQtvyNk96PGBZcHck4bXUQfX7JQvCK1JCC66xERS3Bks9H
4CAepzbiboR0xibcWcgD2bhdb7kEt7O4ZRWg8EO6KYlCWThQWq/BHZtkMNlC34O5l5nwiQtLX3ms
UJlO44uIXzHzfy/VUSOIWQSRO7GL2zXSkABgSN++mMfJxASDE7E+4wFqZ/dRededsUCsvG8CMv+/
upELxwSUxLa4LT2UiU9jI0SZTxdxievFL8x/EJQX+RWFP8ZRbig08vHDOVhq1QqwdG40R5a/EjmK
AzAI7Hp8z1ua3uCaHbJxtC7mB9uKOUVaSASwJ4wa2gaICBMx5UJe6vs94lY7HhQyp3CBqauXy2fZ
eCDWR2JclYLR1IB4KvIhc+mRD67dAF/8eU+ZNdQv9fMu1JxnHVsCQFaIUdfpONqWpyIENjaWF2WS
dB4OAbi6gw4M+vcxoqz20lU1qt0NVv0f12O04Fw4a89ill4mrHz8ILKF4h5woNhFTsQw34uXfxSP
1PC+IIFyJv6EpT2WVX4Y8gZH1s7tO+RVOlCMzRSyz0XzrOzXQiX7W46l+UMK6SENWNDJlrbq67EB
bKD5kz8+gyl02cK2xxk8TvzJihzpf8sNwl+0Z5nlBebnrRcs9leUjx6eNz9dej558F1bvqtWKZTQ
72DrNSPEh7Y8zxW3ER5sgrmC1VWRku1wDUwFA0jSh7TG4hSZT06GFznvaa4pMi7noNnZRHTFWshq
pbKcit9qKgcNtTvmIz1uGB04nFHZDeLy9F7KA0pLjWxYLE2V+hNZYrDbjY8NjsZ1CIOiohOHULSN
Zc/eQre+2xJs7GhW3aqzGKcgDZiU7Sy+dvmDhzNYu6F2XnF8iuxt/9TxJeBH4tq4r/JPlmn4m3X8
j9Qg/tKIqvySrDstSK4blswK9LOZzRHS8lVwAdMcguvouhJES+NQWqtRFxzIp/WuWx5icq4ChRs+
xumssuetmnf2LVlVpRsWLWNGOOLbjKsKUkzrff1oxh+fVzk5p0NSEpIAaO3Q0/rHqhYrraZ9cb1c
b6FYniE4UKzrZ4jOsV06MlDz2TeMXpEj5cIrVOHvAZMNMIcmLy4+ThRkydHPO3sIsRRnRoRAczuS
rdJbxOW4IDXez530/428M/PJG3yqG8zTiIwu3Yk6wrJ6wPSEQJ+mxNJ6dr3WBbeBYfhq+UdkoBlp
644qpKwGGKXOa3ULQXHiG4iF5DdSTGZy/PF+JI/ZJFTKutYxvJa4k183r9H7WM3v0lpP+8FVis3F
IsGe7FUGjVRJhlUSjesyUbzVzLtFJoVNI1s6IxG2ZZ/c6VrfklqXY9XhHaMMTmLLWAn/h1SB7MEZ
1gtGeAsKEaNen+L6wGWAL+H6nrkSy8Gu/FfLag9W+SIX8q9DTTq/GUBoxOP9xbFxvouH5cbfQhT1
04OcYHrnNPpDCB8gx0u0zmCV+jJzosYANiS5ludwtY8bj3zb/vvBUvjG2gYLHC12uucZAYA023GV
gNCd64JHjucMaZNp7ifQIZaLVtQz4A1UAt6xqhdfNf4S6osRR1vnvKCIq/HOIpKTsAMFaof2PRBq
rmihFx1qzqm2w1o4HwdID/4898kZujoXgDsZ/a7OmTBKMKx2yw8NqsIGnREgeUQyVE+UxtagN3uX
/AuWOho0otYNO/CKmr1S79N8Mqy114o6g/09ClxG67k5UN89YeVVsByWYSu9KVVQ6S8w1A+8RRcH
JMJVyN2vHRFbV4hxYSTUNZmP5vXIC0INvGyRuchkbV51gvA460e9SB700uLbUvs8ueWFz3qpq/Fe
8F6tU5LkwKQFKd4jJOn7O8NfgIJq0DF27siNIaqia/ZH4oJiaFOVYiTs8MJteDIiUjHtrlsevn12
xM+954TymvbgJUJ3ALGfpkYvCIVfwkn5O+Ffha5lv3TmEVg2LvvNhtXjixNOVbeB7v1lyFO+kj76
ockmFStBiGaPhgPi3HwbO7X+5PRN98QKU2KVz9pBIeV3graljAQqU0oHal7Gzg9BdJqUs32nnltU
Xlz171xZSPyydFmgtd52kq+ZogbSUisP2iG2oWF0/tBftU2+rJwcsRfFJbe68Rlp+ase73ArtIa5
8m9y0UGpDaQJhZiXFNDBPmgsGsbcSWR5PbasXucJ7AKLu9MvY0eGoLphtigrwidUI9RUbGMB3SAx
kJjKJz5snAJAbUVl4CQOBUeVNa8aEPOIADpQlBI04CQmqLTbc2cJXT5ijidOpbEWNB3ZWtqyxYdN
nKM4jwlcjB3sXDm9rIeuuCwi1yPT/ag8VksPEK7IQCc+z8okjwpZx5rR1EqRPR7fwlW5XPrtlZUi
RbAmjyYEI20LLSct7FEfyFitnn/Fcp7KgYsgUF/BkstMt7qYQVPIojPTewhXNx26fY8xHK5cbQ+3
eztrWv5Nn5DO4EeNCZd/FzQCx+90mbzVNbiKWSoVIsrnWPF7LKE62YidL/Np0mcd8n5TDl5UhU9d
HAR2+MGD9RX0oVueMRMdET7/4AeBkkOx7Fb5U5JTwQtXpWbRVSV2DMMaTRrEThRzq9NKMe6qb7/C
KhSx+1L8zLmGlqYVv1wn3VkE+GcLUdMpBuyD3UFf5UnRcAaYvctrEGsYCL7SCfBw7en9f6anAkZK
jc5oXm3diHU8SMg6BTEaX9sfe+Av4/T3Iu6ok0CC9wFa86iEOU+vePHbTZdErLGT7xyDGkAv8Mbe
6zgpVolCDx++FRaTcgPlP1vcEXb61y3vJheRQUD7Ng8vjY18U5urnuhq6ADKcdAITUyvBIz51uMU
bGgFd1g6mJvSWbiTMmVbY1wnm8/jkLchXFPq8XBTMVbfAspcvsvpWhTZ5CUaorIoyMq12aqEgNMd
0vBubHbqVIXseQ62FlCQBV11DCwDRe83boExD+IBmxeAvyxbT2dpZH0qPHQPq57sxUZcJ46S78Ys
swNHv9e5Y/NgG1e0D5wHUu8P6mbXx67dHmDjSLuSQymkOqmakeclTCO3T4SRK+cVxECGUnnEuBKB
irlL7W8WbjBmxeIaJdoqCFl54MhPMInvoh/NpZOCoV/uK+jlWDKG1MPHGxph3suHozN1npC5m0zu
X5aliX8IskASjqKhRpR3hP8RSSw3XHENwx/lV4OJG9BujPMgTnsikYIABjjF3XWFPn7tdYz7bazy
nyjmrG7+SLPrJjeBzZB+VWDduBCp8nrosD533/B6OhMWMxDq9RuEQfi6I93Ak208V250ijPI104R
PwDSD7asDe4rk0SsHKOMI7qgwiQw0S9URvdFsG1+fTP43Q9omAZ2xGBVzKiWiBdIG+IzRi8dtTdp
mHb5nJnzh14xjIqKjYNUB6YR8c1Hk6edmbb5lK/d4EG4XuDr+KTQ2lXUwP9TMODNIBWfn/wSrtai
sXuS4r7r2F7YoNtNEB07RvEXRRQaYX5G7CEwablOyKJZiKNK1qGp6pqeRhEoqi5ep7736YhRJNon
7iTwxNf+iXyYpQwdI8XhmP6dO1AcZ2D+f+RDp9gXmvuHe/lm32WEHjjkZWu9vOCVUevERLio5M1S
r5PP1jhrUcvtFRdlI07kdE9UTtS3pBgeiVLPxyWLH3udM1IINlYm4bqzZcN7kSZgE+cyol3199kd
RkrfkK5cv3NBZcsP3LRtI1Ne+JagC2y616f2CZ7Fh+QDNzCZKGESMJFeYEUeHZ7SyKd+YweIwSdT
dEQiDcZdU4cp0S/atHxaPV3UV9iEgcs8kiejuYRRrJCkZ3XUssiS5nvbvuU0KZgVox3L0390+uJy
8awOZXmg0W+Or7dT/XKudrJi/3HiETlTh0b9MHt7UzZIu4AnaNOwa1Q8ZN8qfgeSMEnfgEqGiJNr
+x/E57ZuD5xCGVotHLarOZ3zaPSC49MDnDQvnPiLlO7VYLs2YFAqptv5mB8eJ/rkI0mvzrD213+4
cOCXphDNbitDeg4Ox4OB+NWUkr7Hd/mpWmEYEz2vGXAzF+3WtRk6o5MFUkr9xPaNUc/w+jh6M73u
CLuYosuzFzab8Oe84QDhvFNsEZF+lbT32kmsdJZ98r/+PBrPRkXX4zVGaZdO4i7nxrEz0H/qvDMP
K4tYWAan1UgZH/QAt7AVvDcfMA6UXUXoTJKtdtrU08PN4t5oaq9STTDXgdrdMrB62Fs7gZ6RT0LQ
YmQsk+uWzMbZvrTLkBkVQ8GIhPbcycTVwFoTn3XijFjpblxJCkOP0CBIGUvtyGLRBywHXBbXC1Ez
W2z25goB7Wm6jcaUxV7IJi1Qy4JZ3RwUzurRuEzqF+l+XSLJYWu9EN5zbjxde7hgjfomV/p1ZnGM
ub3IBalxUuUsdjsEBzRGAIoGBYRl6W1zP992PVxrHkkjFUWztV9I8tuxzfs4/Xd6R+g89GmiZrs5
PWvD/qLwUNmBS1fTG5anHAVzZ/39tKaElMwLylErZggkoIhqA2w02a8tFlfEt6NbFiifBoJ9kfHk
lqbHbSDsOUksh/6d9Euddg84L1BkIxBQQES2ao6KnTBGpCXIij7jEI+97qbIwK3aV4Jm5BKbvtof
zuxn1a+3E1ypR5OXhMqqywHm8RLzGXeCZCMgCiQ0Ps5uAKDO99+qURyFT6W9F37J1oOF5qL7edDi
WFQ/Apeah9kY1xc6x4VQJ0Pa9UFfiiC69D7N/6JrcnABTqC+u37o/REab+hEPujhbxjnjx2tPAqf
1Rby34oNRTFsRV8/QL2L3KkLAOJrrgHE+fjxmxUyx+wWKBk/9SDWBujsxRdk2y3j5FsQilOA5xJz
7CFKearRD39aKRbU0uhCp1w0/Haxa94YwWebWHdIK5MF1ZHBO5Pq5FKGSdP97w6awHPCx+JjAUgx
3aWgeT2pnirlAObPhA/6cADAZTjkwXjWA02ejGk/uGAJTYM1VKlvQj2KAclXcTEdMJduuDF6e124
/IVIRw60YwVSNonaLiklX1EIakPUlYSGoF/Hghpsg+TgqPbLXv17Cmr/bF8D0GWZZNk7pWxc/oqi
Wu8CQUZClyf+pZIARcDtAISJ15p8NfIKwyjsXQSBZbpsNukUS7nUduDCL12762yZWWtIQyDj4cAp
wrk9YAzUAL0svKnyBJ+2XMUp/mFqI7jh13BoumFJfiKIimN8XEocoVfozBF3/y412m/4MzPRYddi
Qk0VrPVcaFKjJCOfLB3wqStQdctn+cCecfEg3AFOIFGt/F0vI3ReS12lJmzgIJSqcQ668Y4xxTo6
8+7JEQci64krpU/95DIurd0MC5CVHO+K1rQwWbaHJGEqM1m2ZGI9f5Fv7cauBrobyGwdrUMjgk6r
uUZPJb1y5Gp7W8LAcL5oeD/4/ylEYNxhNg6VzYB+paG50DJpb1f1DxFm6cUUBR7tV3oA4nanxSYV
Zpe3a5U6u1hweQI60gFPn/6EAgSrmIhePlPcda9Iyj0idccOxlLs6C/vrCYgXKs8maKKpJVbKmDv
sz6NvXt2nOOP6bDRy0QBO8XhoI1+KyJkM+iWaLeH7UDXu0+fzN78aPDNsEX4xX2hsiuXr53iJKES
H4k96ovPM7cskMXf8OXfo40mF+vgsEEegA5CKm9Zc3mg0ebs0QhPy1+1H7EAZVgD3rbU5gZuqnH5
oj28r8oAeCA71odVbdZH8XIuQmnu5UuH5SiQilqDy8xRr9aMe6toWu8hNJkiIUH13VXrJRtcQ5e3
QlFuHg7/0/lMSk9Xk8MhrQRl/Ct66xwrk8Uwl2fLZ/o2ejztTZVD+6gHY9xH5YFWp5/LJSGRnmLE
EO+JrSb2qGZgfKjciP6K2pNHEPwkvKy7YVLsHExhe4FzufoQroUUmDjHEkuQQvwjQmXIjkuPyZFg
J2ZogFfL8CCwhgPtEYSYfwaSxBqHAMOMCUoiNNOL1DLlFO3vBrRIT0l6qFt+ET/eMpAbyDt6MYQ4
KOEwA9qmZW8CJlIiYEDm8gS89U8gc/SBwDmtO3Zbnav0MKDEpsKdCy0qZNsWMemYwVts5lJqZfTh
bf5+NK/wqlo+r/KjWjzqqWxNkNoRl15x92sy31uq9Ja92E4XCPBfanhU2bbNoXHHjJ2E+THGxGns
HczDIrdrov3QNjtSQCXmLauEK+8iivdNcrZaRMnmQkrMwJShIr7zUOHWZseMa1O5W9slcGcXmAxw
j+f7oQ1/jI0fgzyqJDXLGasEQoQCFPYAU/vFElZTAHiJRhGFiEI+yq3RSkyosq3p1ikEccl/RkRQ
Xe/QXgZYrYgekPAxRXNr0u/bjaLnYnVg879r4sop9kRXl8T4nNSJxqw/MRRPaAl+ihLNM1OIUNsf
dLl/3+PyOfOHQQnM5wLC1I2HQX7BHMDo4SILVkFYox6mFkVHOxcn7aLSdCxiGjtBUSFcab6anJTC
WdD0jPeLjvZ5qpSk+7gM/SO/26LPvFdnQraQ7PzT8BSAIbwap9OnMZu8QnnUP9kRAa3W2prMzAId
yGwTZ9VZDBbuvATMoiwMJy72KgjpJznHbfB6PI49KLb6T+LXuofjPmkWAVKepmSLZBACa0AP4VVL
zEjpxIBBEF0jEkTAJHYSA1bcwn+gM9pONqDQo6djKsuhV3cq67r42zCjWCwQNsN/Oi+wSnhWPmLt
FMwv+76aL8wmD7CQ2HsEMKDBBp/TUa315iij69t4LVj+P7X+JC2NB9y2/k9EwCRWexRnbV51iFGm
ibH44YJj4/MyE96oLLZI/s2OztdSh1w8YMUP01ML7R9nxiaPLXTkhM4drUth77w337egqsTjSTf0
PFZfXE7vXUBbPTkISMnqtwv9+AKqUHSEcX/F+3k2huvQFS/AS5rkiLGWfT7FJZt/NxgpCu/lZbQC
l3/wobMl9rDJKn1KJhNBDxzlkes5abJYe1TNUTwOYZmbXg0xzQ5w9nY0/Ed9/fklb/wdlJDE6dLc
XfewMeRXww2OY5+AQInYGbobNKFJz9ie6H18p1Nlw+IYrvB3lHOgJ2aj0iMpU1o18kGZc+5Fx3dP
6eOiEce//qE8BtBSH5IyFZCSNRikHpXuon0kpDw6NVnZ5rhsPrB65bWoQtE+uqdErvP3KzDGq4gL
p/C/W43oA4q6ZbyxlVPVchSWnPuyIJ17NmgNHmpiaAbh3eLlvf8cfuSGnO1RhJiAwyMmODvciHm7
NmTunQyAzPi7aAB+xtIhVxktrmG34/80SGMD62Wy1YvVq1P4y8bSapLbBd/+ndAwrBdpBVr0iyMY
CUWUj7ceIMwEWqhHyugBbaE3dW99CfTD3X5wrJpp3eFz+Pg5f7sbdotcO2MbiNTtQdjOij7pV5pc
I6Ni8yj8tYUnQ/jlSFVAWmk37X3uNWIFhPVqUf9t0vLVLI8aN23/vdKVKj+5EwtL6xu8TwiKCZGa
Ja6EF18/S/riOlzekRksrLZT7JgMXHYb6eATLcGLJdqlCtzoVoVpcGxoh1YMuQmJ1vV3rNIl9i37
25FlSBwk3C85HMQ/JnLCMIyeH46ucMX3SdEfd2K9v2uU6X4lruiqtegXAFsCSDUw/4EWlyXUBxSQ
ucCtyVecHA35rwg3v2mjt08kA/Xbl0+8GOR/iWTUiw+vEa6vuvDWMqwssxrg7+ZJZJv0Mses0xGV
r/Iv6xPjzqIs5GptffA4IKi+IKqLqG4o51kV0nZ7u10Yw+ATKtAC9l7HzP1uo1HAyyzg8C/fcZxk
Rz5ZE7joIDdcsz1U6sb6vRNel9VpdPnLxg1c3KyjaOrd2hWyWYeEp0JNO+xaJmxaAQClKbcOmZ8U
lVkYrGNrk1vIdrVO6759N+svnbBhGzNXVFVECY6BYp7UMcRS7D2OgkqqSw7GVEZ3QUF/Gkn0aGHt
ckmCejw9GKWcxjstVmgRW8ljqTrfqxny7S2SUEOq8mNnzB+K0hAgMRUvpWFttsc48vToJ2FiNS4k
jlqIYJjbHkgNSQswnPUjtI7SPHnSdhqsaV/B+7qCa3Hfoeu1nKLBZGqTK9KaHp/qMCUqVY4AuaVS
X9jj0tpOLuH6VMM0bLKAQ62+H8hkt5lGPsEFKOTA4TiFURwFlXkgeQmM+ahW8SASDO037VaaGt3G
oRfVLGad2aP5Vu1Ce8TozASIXQsaTNpkDUZ9mcT7psCT6QOPXzWbV/Jg6GZWnqA4cL8mr3agoN3o
3Uy9L/LYtUZpyN+3z3napcqFnAKkZ5zBbjbJxrsIODXC13JwIx4HMCIU2Fy8rdw/cf4Tzr7bXqe1
DQXkf0jEkkZhi6dSeq77Xb88WVRzuX4ubVyQqSch+ys0d8o311X7Xg7H0jjVkvn4EGMmFTQ099IJ
ikVZZi48BzM7jtSEPA3f5ILL/zud0Fh2Z+jqP8KSYIahDG0npI/MNIlS+z+Yym3amlVdI/kjm+Al
Z91nTx8tvn58p6zkZs4FLX4VLfN8TjgUKNryy21yYmt9FwYrQ9Kk2GwxNzvYdLmLkG84idMXVKQu
RDF+3lTLNntdcR48r/u/H+BIHvaJEwtX+7EQVTz/IiNWYHCeaQJDDJJPgYealHkL6jLYOrURduLu
3zsGyi9XQNIe5sG/C5lhsn5zQ1+a9xdw1tr6sWD0QvEQr+bj7CVBjPaj5xP4uaOVGKhnAgm+/yvF
s9MMDxCzDbONiNyla01ceiQthRWvPmQg4UDkEW8ObqMJqk/+BW46lmr9UpLbuSx74zw/NXeU1AOq
81OJlpb2mJ5LNNqJcGWgcj3oG9i4exxvFS8IOWqEvEbYpcK5+/z+vb9UxnD4KUUdqZQ7HF8Se/sc
eWNHNdvMq+9SZC8u/AjC8EsUtDCqM71aUY9i/Q6DHbLrma/4IFvgBv+GZ4gwsOC1dd7QIKYAfX87
LkmSP9XZzrf8lZtJ4MpySi4uYdrQJ6XnkXNqjgATJLOFfaxED/PGaG0QK1drY4AgV8MViKN2FxSd
Wy7Ue9tw+A4HiAKiWJXU9Hr2x6Sbqryqk+IgqypKmdOrUX0nelko5vJz05S5xfSegHge1nKRrpkQ
RVOgfAXuyhNOK3JbfZfwqSRXTILVvykcvC3yeI9pfjxG4cDKAonR2STLySZjEO9C1q7CIe9dT5Vb
/teFmts3R+T3BFcJJZlIIS81V0ppFC7mi36ZE/6BeWDKSMGzg+gcn2w1nJzGKwyq99nZdi6mZDsi
DZriYHbH8DKx+8OE6kpMeRI4uBxaB5Tm1jtARBEguOvKU+z6AvPRD2xQBLRb7Lk+b0IcZOMHnw/y
SPWNIYZaglJT+UbXjaSznLPhEABigvri0mowHVmsBI4iCsDevwAEiQ0CchKEm4a6zW2EakKtwlvT
Gcp7oJ58mpIBCOI3HcVFfGu51zlznFfzx1wMRklrT3iJrQe6ipSdwBgBoIIsbsCGN3d945PRg2du
UVWhwU60aSPjiq/SUnPjYA3p6rR5WpcoZwri4xUaOob2lTdH5mSog3NiFc/oYrACJrjb9oiCKtLM
yofzYg7EPR5FLjEFzxDK27JoQPoRn7XkXlAX2ktSryqYJuLATjdQB4Et/zAbYc/zafMZQxjpuyyL
upApIZ/kuyq6hKamZ8JYX/pYaSPg3eBLb81UCNXJfo4Uf22sFFHEvfwJFChWLVV/cg2wYxU5JqHu
1Q/ZWBoM0yuxlSGUEE+L/CmRgR/kavdpT3/QZWT01svC996xZrgiN/8hW4DNvIrcKb4U6erMGFre
LMwp0SNorIfbLKXVa/j0Cjmc6dY/COle4uU/vi7Wrt8mYIfrkuyZLH2J8DYDBzgxQf70g+gym0RB
r0T9toKRigi9FPQsuPtGk3RSswJi9BR84k3EkkbFydlqvBeUvSoR4ClFPUzXeuSOLq1ktyWzvlit
bg+0ns4f+yJZh7lwXlvdxZDl49xhgct/39l4o5Z1nrKsey/jZ2OzrLxSvr8ETLDTecyoVbdkxJQ+
K9rh4sBc6VKtGgTy6mGM/yuNAUyjkI3X/5lTxlGGUSuwUV4W0LXCjT3MX94ppksCK7pLvMePINZ7
X5p6eiEnWKNe3YAGjPZpKli915iHfg1IWjbd9sHsiu2Ry6Q8GbqNLYHMcgUzZV1GqxYNGO6dvp0J
xLXUpLhrgrqmhvpQJRKJ3L+TMfi0ZHRS4ZNyCjwC0fSTy1r3rGcaCVYZZxrDNqBb0EVEAf5YnZ5/
aShGXaNQhNcC2p3e6YGE7wZlgDk3iaQLAvSAghItO4CjsVNJ5bEcQSv74lNToSjYKemudw5vIsqd
Cc+qGR5HtlWWKzaoErTkAN2terQZnAxGSbvETa3PPeVojnmSaP5BQTAU0mgMFEMb3dAgydhk5La8
l0qzuojyywleV9s/htoS426sSTul4cI1D7lzUWKptZJMjXOkT2VFZgn0VkWI+A18dGBzmuTtMg+Q
QC3me8rVaREcRwGftPyJkQ21nTH1R4iApqYvNmNgORX53bGZtJyrmHCKFRFlO4jXyLIZ99mFOWzs
quYl1B26YtI6KvIIalhsFPyl4/S4Qrz6g/wpXyzt88DU58zRLRJhIZyKTVfJIebRPK9SkN+48oWU
xsK0f5rxsgWMZQKKWIfwVIcKL+l1fugSY/KaPzCYOkdw3hcwZL3zXcjpxaoMTFSYoIG4iTcFm24m
M2k8a2+Ui4PedczGohfQ3luZ6FURszNAQtE4soQBniL/1LSc5ML3IiPDcaL/XxjWoGnE3DEXaqxu
D7N5WhNyODnw1RLNuiLlWL11ZUl0n5ZWCMMXpnI6vAfkO8VQxklxNERrR6NcRURp9PyTawCUCb5u
5wdOjDXD3hNeyFzbh86s0sAchAff/2t3EpojO3POjiK6MmV5po5dM4prDdcOiBY+7Px09797KiLn
jOALHaMEpo7/60hP7rn6OunPbmIT+SNIG8nP389obFpkIvOiTbkvkjVoq+iP6W0XqEYGrcIKUdjy
svB+0ZTmTEe3MmpTD6X/lpmizZHrEMKR1Fh6InYqqsGKaQuufOwMdFn8X/pbIBn0YkCbbIsB4WF9
y3k7xlwkAjkRsKk+DisPoCzDHPw4+fT4SecuLfQ0JQUVDBjn0Px9ts+QX1HfsMzSxaR3+fVp8s0h
T8LU4hIDZ0vL19TLZOXYmDMSGypbRveW3Xp8wyg0IXhAByF5+EeY90f4Vd9tZ5OW3xLXDySugk/O
Ak5kc1E55TbYjKiYG7jkyZWHkSz+qlE+L4S5ziFe7+xlFyugH4c4HNVrJIjVCJWHwQGCvgHTwPBu
N07MFxy73qKcHCJMN1KSc9KdgI/MmMeSedJnE1fbuxhDDxxzgIUvcx3JhwBMG+79Db0knH7hQwt8
+vbpYIQfW/s6TlCDkSFc6v5ZEkg56l7G0LlUguioJ27gMN9N3bwFI8r6klHxmm8OGfQLuYPbnHTA
tr4C5E23uLpf/X6tK6eE2Mq/RyCZEjepb3N77T6RXfN3NPaRhirt/2YVBR3mbaDY0+24kT+lgcB4
FReYy5CzaON0KCuKjS7EK8GklkMeVfTrq8SIhbDuuKHG7mqJ4APV8jDreIy1tnJlKi0iDEXLJyxb
oAWfynuv7yIKUc93SzKjtadW9hR2UDv5br4wSMFPWTxhdbapZNnmZnzKBoCqCLA3f0JId+NUOZGk
KKq9o28VutI2nkWvsfS4J6lKYebDwkuShO6hEhqgue8kyTnzT6Zf8gXhbigY/Aobr0EeUrsfZ0Vm
s3kpHMujzuU3r/QY0buYSxNUYKt1HqvYYRYUYOa0d7YVGIwRsnvxr+8jgYwz9Q76pPJzvbGm51iU
KTPAf6DC6Gfvlndp5uGpSOQvZFgb/mI2X4uJrD/dESw3qU+O+Tf0HGTGEg0l0DeFxUC20pusIVsX
1uwo8lPufaB3ObYxuURwRDGf+Sed0ZhWhXBawmIPfIjLl2tThSrdm0Bt3POvDjzvMCZbMhAP84Vw
DkF4be4hiWRq6bEJ8mv9FATB6Yb76dJduQomMSFX2VDqZApB6Dy2gP7bp34FHqyjxOmv8DDQi3q0
/pOcuYlNz50jA0P9ZCK8zLg58RvTWj46T2qUv3nrCfWvDV3WXGMY9QvuF8pigCUF3B7KWfVsJ2Ii
4lmfRPou1f3nUoS4LUPjRFCQCfEKywGOiPE3CreqwmoaAiT+OyCvhTutaXONRyikdYLxxfvI6Lor
wTacxvc/jXZUP7M+/dpW2YXjqwz+0lZrSi3gvjgzg8TPIYLABH1sGHGHEHDTmb9TvhJwoLPR2MWo
SA8xudjV98MedEdKvOv+ESXCaHldpHC3CKLYc4na1XkFQcmadedXL4Sbx1m0VIoA0BzHrfCPOtM+
hgtRQeFFVtTK2U6FfE7GkrNja9bzDP/kh2yoMuexue7k72ZDTuX6hiYhfiuBzDJ5k0vMUdVSfaii
PUvsUbNiFyo9q2+XosrlSgrn/aqedFfzS0YRXqQj0gKqAftdW3kvk1ix/QbAgzKf+2+O4UFzzTl5
qTkfBojYOJwery84M7pA9d3pwr3bIew20ykd8ihKvSIHuaM1ZqiK6Fpx635GWzQBBeCF5wYYsTBb
Vmh6maOi5kQazizgx7WIFKngIpX1x0fBZ3twAQS9wMjLaLTXxcxF87ISj/Y0csTL5hX7+gTGW/Jr
zb1xQdYSFlR139gTxw9AFcgUL0U+nAthJWdnkLeWHWtOOBPZgLtY+TdX2hLu65R8d/2XZnPe9ODm
fbh158+8vdQKpLlcUaKugscX0gaKmneMjBaqjwK22DmlDKdw/u0R+3nxnYelt/icMJvHUud8rFcK
f1tQETC8cFlqBhFjscDNrQzz3LZclFToHex2q+7UjNmu8V63BB2PUzCc+3SUHDXYEL+19DP2gYQq
EYh7TgNLOetqgW8zPie82LkFOitZY4Oq4QKG2Nbo1GDVNwbgYHnaZIQJ01ViqQaR8JnNWlxrdBlE
RK9NUI6/wE9vuAdtQ2aXxJi1Of5hDr2y1Ae6Z7BxbeXu5vH5nmZUFi0cJ/TvSgyzXocuF9LwjGjW
yzA3pV2HWS1xHW/AFow2Rw+ryDrMPpXMxZsDX70QCsLMSUN43MoSTQ6YmPP9uqv6MPwhuPzauiyY
SY++zd7P79v8Xl7Vh1mYvFqrGgren7Ec3oidsVCxvrmNjySp0LhgHw/ZTrF1ItLHcv6GsMVB6IZL
TyOpa73GmM1N83/D/SJ7Tr8G1MCe0o7Wa5iKr+yIjjLAzj6RxoR/oq8jYSuyI/XqLSzA3fbEV68O
OuoCG/viFQfjw6zU7xs4HYfoNbDXKo7Tn5soo7E5F9MkpjHMKydYw72DBEfoXNjAu3Hahlnaj8b2
bEgRtnhdk3u7ybLjq5Zg2EB4KxWzPScWHzePTa9LaYaVkNecrhP7d3iaMjljZESAtRpVhLUb29uq
598xQOcQWsBjs7Z9VqYfpNwm9oPS9CmnypSpchSG+Z0WP4KeAIxsjmLQPSktuUJjcyoGk2O+52Ya
jb0nJBJf7qpc2IIzYzjOKsV0agRaq/IH5iWm6ZIDfhNW++KWH12I2JnLbgT5U5nf50+H3dBTuZHa
+oXbCoOrXZCv8rQ8Myg42ymN/4iKOvkPfmwgN1UqzCjuQKW7hocH+D3KqwInDQ+utQpFkjZKs6+u
tRDNtoLc6hcN4LRXai0erdK2HkjISg6jU4QkmAeaYqJD6DVE+f5uxPeo4DGswSgQy2tbXP3I+JCA
VugjqESJayQ6hS227lng//lsGeHdzSMzvLVn1baN78SVmPl2ZVK9+pVqX7nN8WhPbkEiuK7pw+bb
A+TuP7oDpqlgxVksMvSjC63W+whvURCZzqkBFTX7FF1PkhyhaJdlB8PPp/YMS1a0VBOAGKpxnHQl
SKrcasf85SndyIEu7tE3Bmswgl6lg2Auxe4OFard0n3SvOrFi+QxDIn8rWhNw6L1XgDJ+P42Y9ug
PNGzKj1rseivYk8Xgi39vHPi2I3CFWAxREmAOjeTy6yLEhnmG6gN7wGg3Rh3FG24adGPFnVvW8WX
wBaUwBNjmizyaM6HzKdQ2U2j1ANkPmlUydcEUf0LO/9TeidrtxpL9sZYdCc66eYnH6X+5kiMWI0D
v4h4Qjf5ZKTsyK5gqplMIrzq/mX6toc+EVrEGMRIISUSLS88wTFUtOXp5B2DVMJPuN0N5kv6Xh8Q
fq2ln50sX0f2lFRTBFYl4ND8DJ+rrkSGqRh4B1lLUVc/14ggBOfRMp7NcwDIdLXMDKKWD738M4iZ
g5z/0pgckQOkJCDn17T5d53mqK7CvCJxgPQHBGK8kJwyC05J7dq+TrvBdDIU/7cC7SrtmRQSrgJS
v9tPD9py7Uh6vPMG4UvS/NcdOYLOXYcEKidMfOJXnzIc1AsJcnhoc58VcGFRs24EklbgBplF2jgr
M34k6w+hPrCElD8DGfbq8NVMDiRw75oxxgmDM6g9arnHNOdNV11CbZj0sJ9n21sv3W4VlzL5ivbR
bYLqxNQ6BgF5fc65Q+euyrgn5aqewyj/iKRaBm9k8QrQSU65126FPTwVhL9VAyrmlQqemjOhH5pS
fqzwVWu31xDOFE0Ws+m2prNiEWauO6vhJuXuTkiteelgjusNe+OsaHEfxqjgCwa1zYd420u9XSRD
WTG++wtnZkQi0p5EKqJQCiuoO84N3tUsTmO9VFeNnesJUS6FauauAdxQHJkpfrTe2vmfJpEZA/Aj
Ny19hTl9J6WEaQtJ1a2yjPC4bMD4rT0XC6jg8wwA+cSykCb/M2NW4hwmlnpfBdI6egmQU/KjBlMf
uCWoWlGb2l41DJ132j5Ds9sjZNb13/Ky6cOb83eUizIS97PfI1dJNs7fWufS3N61oWHk/lji0R6f
8dI1bOpU0UeRL0Z+v+ArFa8oHPWnfqqPbiEKe49f1upfnsVfMxrx7DSTgQRrSHL38eNQGGaRip6z
Aa1MIZct3s+pgQ6i2J1aW+sxm9UiS6X8nTVVD5Ft9YOvmMHkNSSICi7AxOJaGKYoXLL695GSnVMc
/bnXgrlovLHEYqlz+X/IWVyRBi0dwy0wwnIszzeXM8ADzANbThq6tzvEjlsHDJ/KarPK0VeYOZ9u
x4wdP9bc2AhijCY1sLi3Ye+Q8WnLeZ79ub+ouOKop5tMPLaV+WTuLtIkP70265l4kt7J5q4KZovv
GYZ+Dp4v4gxzb255Aa5SiShX9SD/XJp7c5SQC3WVqsRm8idWAr1S777d6SX+GkkLMdDYAAxD7G5C
Z/AI16cVJOelTw2+35Y88lc8P79EgpQXtw0wyyNaEvzG8qzuaYaTsSS9cUI3sZ3yWyMIGpFokvuf
hzK8fpsi4z7yofoAUVeOqEquJitGMINkEmiHZ0QpGQ0Z75tNBHxEtrQFNYrg4RNJImbYk4uEiaY7
82wTDbxiyrQLcJYnTrofA2ZyNX4u7F8vNXPHNkzftnK5szHQlqgJukmRWmkluxGxhq9GUsahZl57
09gZCMiOrZT/SDKvwSyHqzUPnEX6vLXgHc41wxeHSbcud2apy9nmFi7TuFScZnorsm2Zr32Qsnjz
5bYOsVyMGfnaVUrJPRbCVYpFRk5RvdK93Prvx3vTsOG+Rg88h2/2NWAztjVflWFQ6Hrcxuca+Xty
4ApmgN+KdugT4Mh/6SKcui3/YJVRl8NHCf53I7YvXQf0nWKAywc4vuGlA+meyWozTrjb+095YgpL
NlFOVZTuSawAbm2OwCacDlHf+ezZrCjk6gLViIHvpKMnlGH64FWKWjEI36844we3JM74Myqe2O62
EQs+m9y31skzx85Sr3vNMXVRe9Z/vgNrS9p01RIso2/qrjeToG/+9PvxQvv0opKJ+SZVzHM8j8b2
mDmZB+dL2Rtr1m3br0cWPd8BTrAEI/SiinzTnnN1jvjE2vxd+AHTmZD/lNYm5mWC+mcvf0jBhU18
OO0HoZ6p4kGx28yVQD/aA1y72eVS/Zf/8tSN6BQnMUdQxny6sjR2gxsmV/EcCkEuBNppVNN2eaHa
1rg9zcuFtalaSooY9rmunICyQEPsvpeJHcMHDw6Iq54HmQRSXBzhhUp15H5oH5enX/40jIoxddV9
fZd3NLalGNFUmCXIGYBWWGVMjH2T8M2bK5LmfEV6+aJ5+0xWVGyheu9uKX+keJma38kjV/BJlT2s
+fny8X3PaVdQEkThuBQzDp8gYvDfQJXm7K9KTrYZEBN175sPaIpW7C8Fhx6AxqB8blpgaem9jv5k
ODfOkxfIfVYmuma1kw6+Yw4/zP914mrk2lD9eipybqO4rMKPjRYPmfzRiOc/6v13BeuDnrw2mMg0
4/hjoRRkkHXvwWSMCtUvwmzOS7lj7KGGmqEkVxmel+luAdsznRwnKHGv67gOWbkaJ9N1UqSkQqy5
2six61Pav6cyqX9gk0r2OmTJELDP/T86hG72x3unW1reQd7MKOf1cAJDW7oRVxZ9kRSMqAz8drJT
PEaSUQyql1cephFbXKDGTFIhpziDxoGAbs+Ul7eOOeZpVhjyFbjx0iG7jQTAjEOgIQvQoRUz3OYx
Ewx2EFmOlAxkL/LG1lnQhzMRPGF8vI+szQ0tbR0K/9Wa5bhE3UVK0qnPLyaVMwR8oO+X6AzZeEY/
Xms6Dli9iOLiYwuF7CmOWrEpOLlePQcdZYHpUupis9R0g5+3GINJw0d/TglZxtQay/rVmjDQlv2i
PkErsSQ90BY8qPJJB7O2TULhMtxdQCcx2h09d4bRFrywc+MMHQ8fKFTIUxrQEP5iUZeTjiwpFfoP
CUESDe4okSYPnwkqi9T8O4QtoXxWm6syFuRerqNo2zIppnnrcrlnN8sxQ1y06xgm63S9uuDElwyM
4arqIu6CRGDFDd1eiziD/6LZNU634MexmSr2/28jkN7X2wctMeUmIJCK1EsoCvsc+c1LOCetEjyO
2ukuk6KJT0pFJstbAE+80zB+SFe4YibwGHbop6G+tivgz3lIT3Q+SJno7LxLlnzTwmRzH2Tj41ho
6Oxs9B3gW6FwuxKZLiK/j/m1qDGrtEyYQZmaMn5jehhTOaBC7yogJl1bNqnlPrQH4F+HGI0JtJc1
G3RDM5w9Ht03+4znZ2nv329DEtLlKEV5GUpkunpKw9JmgfMtw1AADLS0O55nMT+9gqOn6ES0zIqB
ULSw8opTqAE5fvTbXW+gRK2JZGmVpN5sxH+HsV8RAV0bglSYAn/am/T/7gobV7m8NTXcVyTLaGCp
mHGwG0t5f16TtcKqnlSLUCaD0YwwjvvYhljUMWtV5OxnmiaPEeUbqigkuaPNMg8hnVadFmzZDylc
mgo4CQ6ZNVsYmxYthdhzNzbTOvxus0V2BZt1bfGOLVccAU7tN7CzF11cPHkhA9cP2pmKcLJ4N1UZ
JdbG+DZo792jOdUMh+puRAcWcrlCr2sg8N6SgpgrYvNT4IkBFFU0wbNdSlimKOa3/wYTp5gQl7V/
iKgPZoPY1K2kbV1p9qJxCJhwCI/9RDGfPq+O8Vz1FiDWxFXBMV1kYwB2a/pH/gESzKw9n1h33tpo
efbaWjgN7rCgArU3T2o3vo1BaLagFiJkE9ZGsRw0hEF0uzxAxdA6xJ1svPIRvjdhTwSm0u/UVts+
CQLK616LZ5Hwp/2R3QVDjbJDVN+WFAVhgBDy+E2RGPWyIh72+b6/VtIjbrTQ4TcNT4YNmNZIJNVo
zrOm3e7RoM0tbXKfHetg6sGZO83/hpCM8w5S0VS8ZCpZp6v8wgls9aahoqlMuZgsLUyBGcI5pUX4
3JiTnusPO9TG88UMcU/m+1UecUATOLVdyoh1G9psC2rpNSoXiou0/qak7EXXoYTrt+Ek/RwTdxbZ
6Rdk86+nXYICtHvlbS9KGITr/IZ/dEMqYGTi+MbyfSs2/CpxLyOQyUGrOD9oT50XeEF1JXFsbOEW
gCi2iyqlwP9G2R14w48BqV4/ZutgffSNoBTMOj14iL1nPhdXHrhf9SeWvXjrS0tPoAeJmPPFWIYa
Imf5KIxr0tWXhm5oA3o1uRPLvV8vxggDex2Cbimw9GUTXHItwuWJ0js1Gnax903NqioiukdaaK+J
+1d8qNT808Y5WlXrcOtBLa6peSW5gRG1QeR0EWvwzjS6q+o5TijwSBTzxmoM//xobc0bAjEgE1Km
SVQZpFAWO72XeZCLN/dd0Jr1BtSgtX/ycHCE1jhVtybajyyAmwHprl3q16yjDh5fcSSjnXFnvqKF
p6hY+PLKgl96c2mNWAY04wtLmwaxR6kh2Z3SiG1Bt6xhBc15BDkeTAoCRvlMhFHH4TXAzPz1xox1
85ebJlPEqKkF+rmwMP6//L5BrHeLneTrV6oWiVdiKvTfyXjJAf9csoIsNUGsZyI5G0B4upBOn3TD
oWla/LTKNrS+7SQdgva2KTrycB3ai140c2g2KushpeLqd7XAggSFPtdSP3Ek+6icwTgTmjq4H055
MZsvxtXqf3POVgETI3qXgytrei1529+uEWTKZRt+ktbGh7AOJPf5Sx8vjaspdutDWXHxKX7Ezih5
18ChchYK79z7H2lkF1Gzf0KXL9d9L5HSaUmQu/seWnkcrXTuS7OD5ty+3aqAeY44fM0XYszP0nyL
zKOGaYspE2+HicHSWh/9VQDWUCFeI6gxySsPh/52uco7Xexm7pW45oBGQcEnx5v9cERcz1LfxfP6
zq/nuw+jk0jYUPQSGX8zNnnp5UqWHqvRHSLNf3nFjOoHaFiGDbnLdGRyP73RY+cKG52gGL1wzbQz
Z2f8JgWq3fLBV3BDAxceHAILplUK431e0opZhlrwRDStgoQCxA7mC5+ucnkBUkmvikR+pHcb3bgK
d6bSUeft2Glv8pDRK7qlI3mJgI+Y1rZ6pkG5kjuBQi4DWUuGsZTPbQMrtJoGuHPF8DjUhm90h9pu
LKemVo4OqbrmSJIjMSa0rPphRE7QnrvXdPuCBhxNaaErJzM03yRh5VYo+05SE8qQGvp5I28v9DRx
92EtSUQeVgM4VJ2XFIQDeB2OqP3uyhy/4rJnXagTY4DMkRi+Y81bSvaeahA7FlwT3lQw/Prnz8GN
0nPXtcOZw6+hbvPKpk+iIHV1y8r6R847d99Yiizc8g/4DZvtwl7lrNrbmGZfLT2hBRnBHjDdAguh
0WnKenj8ZCabvBP/ngNWRxUd6sWnJcozq7d4FjGLuthfrlZcNX4Q5cyxS+deoL7NctsHuUIwLHlo
qa4kZtHnECenT4T4L1DaQ8/gdMtCkDlM4TK+JXe7ulUc/ev6LtOCADKpSsC0Ua4z02VCz4d7EcWC
uyuNACtp8JQc+0HQ1pzMUaoNdcEQuF3bdc6SkQoY1qiS48/wfGA7t0p1iuhuMiZBFqSR/9cuKAn6
D2V68gDxM4uNQNmSbJt6ol0LjdOkGA4ZjPylW1ABHI2QlMa5lC7T+RvtaSRtCswyxAMbWThIRpTp
jxUjxCPyhN26DBp1F9CjULEpPC6ZvOTPXCjsQ043acRReBjpmIyZKQZ1Iydb4RTujV9i+HIxlLc2
Yh5JTJ0mMLvkwGn73l8Js8Sr6bZjsLTGIC+MuFni5FYpG4/n2fhqvPjKGhGrDJrDzjUvtdUsdyMj
STaMZhjLCqmPT2HvUewWRJZ3lp/7h6LghTSLFa+0EQ5NVnNboThonOs0goCXNnCTj8IT81kmRN9j
YQBEWkdPo0hsn4I6TOR/BaBptTBiTWFNbN/m+Q372rU+d+jtt1I69Xa3ClwR4jJ8ptaJzrTEYowH
zotzsfdqPTaQKhYjp6fica2/jYdK8icIAvWwhxHwsjD4XeshRAr5V5VBXYN/eOJJnoB/Oe5JjSWq
/iIVcCvr5Qw9EtFAAvJdXeVj7SjQoq4sPb/01KztAGvY0jCzTsNIUaoMqJmw8FUgetEMmkoU9Q/W
pTsG43NQGZMTIdYFZIALL5UVZTsjQ7JDD8LQ6w6grHYJEFLgwh5JNjnRX0HjY2HlQ+8MN/1YwyBc
8ZFdC/80Kn/7/46yNKYEUi153c16wP6nN5UmBy0Ai58tnaZFCpAekVXkFWUEImbbLLhL/aQaxNv1
l27EWpNhVIsM7djoduFzS0rbHqImSTweA+XIfItIy2i6vUmxoaLyhvT+kOG5TIN64H3G81mRhpDG
grF9ZsVgS0m+38sotnf5QJlOGjE+ghHP7A4rDR6jvcBj0ExikzbATUtqoezhFY11HtVtGft69ver
2JPONVGHj9lOwS0sRoeCpCSoz9Y1ev1+XNgKUn8sc5Et0f2FWbwNQYmlAtkZgkyIGu5sQbLrh97M
JcimCK1+ANEW0yX+HHBDGwIsPj+q+4rEPVSaAu9gdEw2bDwWXV3AgIuIlJJLB6t9C2njCNaOSE87
KzdFj2HW1X5sG0qYft4+skT1yHDuv/TX50WohX2uQDhpJFT0n8Tt38/0FGaL9aOOLaACiyXryV4x
fdb+3xXcBvRED/x0FGR6IELOLZjYSnTpkD2Ng7pAm2C0f2buSyXA//rurTXXeLD6bso7yZDOLF5f
0lJxKLOxLLQbe3g+8eXPIJ7IvXA7YOYFevyNRa+0SBaJCHAg7PL31TPRFvEbClsVGUCthjrL+Z4p
/I6ofFqi4wF/3xs9cJl7aHkdK/BorS318miC8Nre5dnXxX+FnG9/joZv1ge6dccX1mlNoZIMyhq+
2vKG2WqljSdRf1LbYRMtgIgfDlHPSjdpgUXYDnOskKsXGQSfKXUi8I1FXyQUP6fyXRCVK6wuR4bn
9fJt6kZ7Aa9hQGinNbnN8b8lJnkJZURSDnKEq4FS+WALPi0NK2IRiVdE4jfI2ga+LZjhdvtC+TRL
qoydPkCVVGxqTRfaU2QLdWzczZHWTRvE/tH5G7YFuoSDq44fm4keofZC6jdJfahEXXkXzMTbHsVw
+CY3ZBfhaFjMJoJG/SX5URH77feRJ2XgN+XYJM7EJHrR18xJzaQi1dl0CHfOLSC7CvO+3EvJrw/W
ybNYoGLJI9LFWhZeI7XLg/8hy5P9FGmE30r+yMewNgHD0yhP8GoF4GwoWuxUjD1KUYSUFjcAnBYJ
jTFIXkOXTIqr+1x1ofowyD+5FytoWoKow2B+wt15YQZK8SzeZ/Unr8kmXz1L2CrxlT4vC8vZFcsi
SerCGCxeKDlbmVo4UxWRqD9TpcPekTvmxfEjS1aL7PftST7OFuIsmj5eT3ZBFnxy2pUjYvvSU8Jj
iGBhaPQ8w2ptRxpL42kluoUMCLp44mLNP39+14GkyN8PHKiTvMr4EApItwaN1Cfjf4al9m7aUjFr
3e6WhlaGF2kP92FCO4O2x+O49NWRhkyZB7ks/omeiVTKpz9QxnngUcL6Wpa0MW+E/ueKEWeJAVZN
njQa5crkBazuFbco8IMFJiQcUR947TH/AqfphAYJz9eZphf0ZUON3Hda7VPA5Ov3G74mlNpNKTC9
tTs6tcX0VujiV+dGj3gNoR0SzAsh9w9NJtXTVtPzSQ0LzzehRUTWtD6ZviLOaI+J2jjMN+b0V+Jg
oN7HsfE4g0yXTAhY2BP9TcjgH/sRlbehMDQ0qq0iz/4Wb+verkkBJAODXZN7XIORBBrJLPNwZME9
vNbit7ddUSHRJU5OOGFNwRK6laEfvHTHnHKjBZ6HnplullTnuJISdiT5901E0F1nmxt9ucD3eeKk
PTZUt9PMflchFFdzMGjpbQPm+98H6dNyuc7k3wNFltFpION7lYxKHRo6sU5vvhFcju2PF2d4ceSe
D+Uwsq6esu/u/kOYv4J58friPy5dGqTB6avb9d6bXuKoUpX/j570McCk9+RT5+t4cAsqnWtH62wA
dqSm+N1Ejf4sdFfuaChsyW27I8AvrGilO3NXIOKYAUroN449lE61NhEQU15kMCZhKGd6Q7UNMKc3
Ew2bciguEkAWucZXHut9FVU798IqKhYWRwoxwuhYL3hdfKOEqa7cEy3Cxg5ao+PyZph8jxkRDB0c
DIeX6C0C5SC/SKPCrE3OovH2VwhcVkIp1WqxLb4BiHIGihBl5wwxZc/dk0SMu/an/46QqQ2gmC6w
7gFhl5xOYcYvFUWvf4r08GBrox5xLMIicPChwO1fbsao+av1NHpjQQQw/leuDese4duuGwjT8ZJS
A72gslt3hIvXoozwXTB1GQ0RawdOzKHYos5/QQVqVR6oGzBuL3PPhmwcH1Y2jHh4elDBv+pOG4AS
q3DemnSLg7rCPlshWQtbka+JHsh/mEzzE9cqYOVJzclL/Wvt7PslYnltSZAxnuHjlqWGMd+2pO4m
6DGF2ZGEHWZIMkxk8u5A+AP12AuHIaWSsezwOQOzIKHdCtRESThYHuxgoZziJkmSCsl08FMjDVH8
aDr2lJIm5LC4j+VYnpTtNawC50HbemViLr23VVNzsiNNDzJ4dpaMFI6PvWu+RlFWN0LqhKKy43/y
VYeMFDyhJ28Ecc7HJW1U3vtnHbF1NLL3geaCfv16kR0j5HBd+4ZCIW1r2rRZG9fjX5Wp1JOhbn1e
ciHl46x7UQryLVW7jWMul45AWYXkQuxDrFRUqFcU3JnT0pf/aWwG9/jvs+o8ZFkyt/ThS68NIMG0
ebLbbhASxM0D9CiDyTiRTpewS5yXP81hAnT8p3npUqFF2wmXdC8h+WQl79pSPj73jkjfksToIAz2
ey/1onmQOH5snfN8yO+b/oneZ+YyeFRkP6IoKaDURdvetMsozjDQNn/4KOMChD+ptnaDrYSOD26S
JZB2zeRN3CUPZVtMfhOF+4Plo5OJWEMPwAx9Tvl4JKATdG1TpKxcXQxUt3kAbURG9BE8jYTuuXeR
EJOivarptp5wAWrI1sYCnX/RpGLtPZVhOMh6nOzJGKDifHl7tgxEEmf+pIOjiGbG1NTh1c8wX9vH
9Xeicdni6WfSR3k923cAndjffAl5UmQRo3tE6KEOB7LRAjoASbgiWwSjbbSHgSDGtnxSL14qmgWb
ycEdTnkoH5r7N9qQZXbolsuc5uUDNqL+40KGcMIAywwawgPRQeaqHouWAdNBonVoi/RTvY76as9s
dNOIb9Nd480KkCUitGL5Qa8ZhtUZSTi3rm4x7rWY81T3FtahJCMfX+KEchoj4GiVe3vLjTfaK0iu
ItXMxV/c/Rnk3/3nfrIyMNd2UfLln3UrHEaDcKE4/87q4WHSJxKoJnQoI9ApVjy9bBD2NG5oynsb
w/TFJpR93BYnFi11jH0j8qsPvzEuaI8gSjmzVRm2CIG73x6XdmxDw7guKyO4QTCrCUBZP2dcprck
jiXaCY2O/m9e0YxnvXnc3HsCLflFZ81wPzDnYj1nb1AYXTh7IV36vzQljm8T8CtfL/xHQ5+gou7n
6JBfnPZWH8f52e4yschprVKjbOReR9V+//ceW+65zYNokboQklimO2tF46ppPVfLqlWy7Fg5DPob
DW1AZMjPvevWp5lbUpf/4/B0ycz0Yry6iE8/v0bBrNlPAhmWn9AKrVerVJ8RdjYB9KMA+/MV71Pj
5xXTrJPqvoTbqYw8dENW2Pe2oU20y1znR/JGKMG8uS2XxqXcjb3MwsjdmRTi4rMTM4sLcrDZ6/uz
+zJS4VYBEujE6KV9RmMjqF1W7lpr+o3GepjKN5LBJbbhLT9YNSWnq/VOgnvlierl0DCNMYdJsNZ5
Wgm+AHkgwn5SN/Cfy7rpWhrrCN5oU7uVxiNyXJ+j/8FKj6qVtxZGvs8IfVWLRb9quzl7q2nrhVDG
LnRa9HPEXT+3CTIc+OFWGtnlJz0aSdmadaB8VY2UfbCJUsJvk/oeU8Z6RdnsORLXe2q53M9GShw2
+Ouw/nShdBIvbnfvQ7U+3jr8oKzjSUbZs1nhB4JNQzzrgNFsgYrwdPcQBeWYmGFh5tGm/IQwaPqa
x+axmakOBM6fWOEoUbtYKlJ1mJbpguNeQZTkpsgekwYae1zpT7r7fiFCNI1pD/4/HAMRTtKszD1/
MkzvHDcw420XyjquV7ywk3hIGy9d5a+5Z/MsHK67vS149g4jaEj/LjW2gAOmz3h0ocLU0ncoyen4
dqO1njWeaLHmRMSD7LKWgnOOSVCin1jiGQVojgBIDMw6nF2KNBSX47jefhiz5etYtu/dTu7uBjc+
vKvVuKvMrA1IlkSo6i1LZSaSxxZJv9MZmt56AfLapvbQzcmRvsle8jIA+S5V7BZ74DSfuNfGnFee
dKSIz1j2eyT2IUf+/DEaRX3Vv/NsctFJK8cgHDs4w4CegSOB2tS5o2e39NcnOk6BTKHTbwk5oZDp
y1tkNV61fxDYYgKdwCYJEhiZhLirdniDpzDPk6H4xBvjCc2pII/mjl+eQsjdhNz8v1Pqx3xlCvJi
qdCxArrfB1bfvTb1QsfpsIygGOGEE5ux/p6z2RxmvgxXfGK9Pa0TFGyHLeULIQ1aUUh94o+zHb05
aSMsVKNXu03WwD2xvtZbT2xzSS5xSr1SyXGSJThNffPEuhSG2u7JhAumuSpkxsc+uxcgYl9dvCix
UJuhyYM/J0aVUipA6jQDMgoYjbLeBzt3FAhE+Dkq1W3mi39lAXnVQNKWUMtlbdhgWaOOs3tXODPi
eHWmJIicfhC04oU0SN1LcOsg6CfzxzanArCemU33nFHE+89qCs0C/I3Yj4+HrxLS7+oYkA3JO+UW
lg7b2GUmSmSZ3nREsXhALp4E7omjMgTO/0gYceO5h3HB02KafEWkMCoYd+NRSVa1h6h0C6foI3gd
4AEezkyeLybMyoLoWVanUlmyA2sRXw31A2LBNaLIYhqLGbKTxGgwugj8TRFZrD5eJJ8jMxb4e2/k
fryoYZ/pUOff/6YJHjC3RfTIh/UdPqniGa+enpqGNFG3eMZl99wWBtUzKArSeuvU1CF6efFP88q/
mMAksUPaznHIN1023isxoqa01R9lBKz7OSmXj2ihB45o2GQs2mI4oBdx3o5CoDPZKOmjiUxBl/Qd
fAdaNfIbqdhVTp5281CnnKQ7oevUw3vGzzHwKdaOsDXe26IBrqajZyOsqhYL64xkOe5zoEGD2K7T
kOzNFoCz6oU3xXzj1lIJqbfzLx20pjKPjKPNBWKgQtDVkVQgzRLXxIgRZiKVLtSRyy0gp/fSVYCY
E74zAe8LsrlQbjy3MWZ9/epYep7x3bZeo4+u22DaQUVy7SbtooIrfAnXOPauLL08Sm9TF13PheEN
MlmjR07fUKePuywP8h81w3jBmlLQ5/8HkfddXfsIwH1/Is7FpaLmG+XYmaJJ3gTZnJg+if6tIfAa
NNChBFgfFhzsesbS0VMk6xo1S3kTJ7eYhgKBujcJeTnYAcgxyAoJBixK+ASKqnA4OCmlF2q/JHQe
OoE6unQRaA5G24oF5B4uThCH9Ax83JaoEy+NSCwZYRCckdPKvYjTC6MLYLt0y7K/DrIGh41LCiAR
YdyHPzCORCuESNCylIvzK4SKH9CpKCWAA113xgWxFrbznAUAcwSYyqpPehapCM5b7LV76B4IFWt4
yFLfymqYZOP7YLQjAVVAjUycVmWqAufqxxrDCju9aHDJtWU2BwAGPFmqOMuRyguf4fGRZ6ZGmhjt
b+3CFzTWccNe1/m07SJ2xiuJFboM7tBos9Dlh16DBqh7C1ZEO50rMZdz9dytsjFCAin1ruoeOnNr
mSeIhsTdo9WXI17+DdB488Qf691aK6SxctK72/pseMfQ1BAHOEWu1/9xrrCvtn71CHWloRd4G/k9
NEhD61XDX5fduiAvdeWbbbI7yyCa5oVhmT4crn4iWpaer/5iWrtFI4HkoK4rKcu4AI0862uLnJw6
Oeud9NUqRsBpbOoua2IcqrIMBkZvQC93CNSf6dyXkwxokja3qhuAhw/KgBULfR2nysMql/NYgYjm
H8ACPIW7jQ/qmqe6a09VJ0nV1jPbRa3rgyOKwea5YPJXS1yFa8YniXQC96p2UcBr7wvYIahG0dvL
tH5MvJOvtWOjGWxL7t9ZP/GU98ttqeHuUqM+ba294iNac/hu/jM1KoOMF7kvd49QyU8PlQBnhXwl
miV4tYtfRvGPYXX0GVTNtJMnqYfWFu6CE7S3iwB9ukACqWxEekPCVENOPzr6Vp4xXMt/IkYqYXoK
Rs9r2bnyB6psetisLXlqKrKpYpPYijXJqOLrPF0EfclEAUOcbJzEGStXyPujj0e8SYozRRnfJ8AB
gJPeLrpk8F8/vmBaIM3ObHjl4MNwecJbgusp1yUZeAPufllDaTGmFa9QHjC8irDfwEtbry8ILpN+
L9Pn8Etjuu95dbpdq7rtjGS47ZjCgqmprGf14wGnxeHJv6tjZeB9eKlb12hIPpCKbTqbMdJMcdPD
G+Hx/W1F6AggSh5vYzhcmjkkuLglTCykVDUMQRcxam9DARB+NS5G4/hwbLXoLmWfrNU4/TcfcyQI
sLG9761PgT1fBOY/Mb/cYwyGzRbnDU9L1ct4p6RWXAyr0zraxFDUSgEBbRwgbVvxutcaoJxlEo5f
FlHmhgtsWYnpmHcM5NwsBU8laFLgJmakyh7afWh8ZpG5u/tnlfqk+CCoaIcDqFOZxY9aZNFexALJ
/vpvEJNGWxODO8Rwwj+Lhcbmt9K6HKm+8fvCqmpkVRhu9B13Oo6JoOK7SUqpPUsOTVtvjyeOf+7K
5gdPB397fSzFN/CYOgNpNt2K3+DrtRD+Vco/YVcVdk/mt1D56nZPusPBJI8fqGwME9RGvBA42/Qm
aa+URGxtIPmMGb7mYO0GjHZKJnCApg0En6yite0+B4Wbzc3m6c05YG0nOiZKlLVRdiN/m+xOfLi8
xqWHZGytjUwnPtBX2g/PNNsPNn1DdUlfVXB4cbYsIsludoqJALOdTCB7lIN/iPxWDn20DDqa1G5K
tIHLA7+35Zg384vNOWky+fKMuzKG6EXoBmpho/toRGLsUMmCoUTMWnIi/msvrgkjWIwer3CNLGIm
xw6GHCQOYhDCw4VGWXmX2BKR67vzXSjmujoeY442EIn6esMfsnH947eu9/z76/aWcWv4f/ANSR4Q
o/Ezg3PQIARIYs5WmmGM5bMBF9oiuIkAb0+4J32PMBQfFvxtFRr2eKdN2RsYQhj6SjxLWlujjsKD
Zivog+Kpj2DSXbQKKToj2df+9uK7xPoLnj8ZKA+24iPoyHc1EKArcljmLZTAZaG7V3Ra0HTeDnQ2
eBipsnWML+yZsmqlQc0xYuueOiRrYGj5r4bo5DPnILk9ZRnmRys/vC2O/otkgfYM7tT+F9SJpCB4
KWWYh62prWZyu0Qpel9cR+mQUeo/LGMHatcxtmmhx3KlZfqVkd2x0HGUthoNGjXgm3mzEEKGFr7r
Q6A2TcMrZrxHMY2LE3LWN5YT1cYfbI6/aYMrJAHXgXZ7yoq0fbSYAVHy+h+9o7914zKMvxo2yeTw
XqigCnbzD5q0QlKkvNj45Sgmj+WpeTdaUYmZsHuynV6PVZNVnVzXOQJnQ5hC7xI1wm9pGz5UIq9a
Ig44XTQqMPxTqSZT8hL0edn5n+6y2tSZaf8GhHrRtQg5Ys7zBLl2FqcM7sTM7YCqPBfUPZgd8y+w
IsId/1HqWkyAhOHs1vAerPr1idK+48VLElr+EBd/fVErk+dvt5ChxMYSJ8nzw561rm7OF8HJeuOa
Lc4UiQJv/8bWAYpsd5OuKnKN+sj3/WJ2usOAFgIlYaT7ky0OVaizHJMqcfWOmgU6w8XgnYfzo4ho
90FKL3JNDcxXBvNqazW+z6Ws33ImlOry/Gf4juX6s75IjO4gHUbb4rDQ2nrX76/A4NnycBvVoMEI
KpyYVu6ABxCKSDJaA9KTASJlFUAly1T2Y+uc3LRGkzkZiMLSg8qvyq4jOGFL4/6feEt+m2v4rpmc
8OvPP0DPqMwnAWIe3WXe/mB9pWGFtXM+faST62zxjurU3TkbTMDcRvqLfxgcXDxyrYq7LHl/nGzx
tZWusabkd4pjMBg2Yq8lddfJb1gWG2oyn+kNiNx9Ctp0vU8CJUwUYYlXLtZkbsXjyGwu33Chf5zR
RrKxDuazmLWz49qYogKkASf2LtSwvvP4710bVp8IEIzhTfKXv2f5TJs1yygjkCZOpezQyBeD24MD
hhIeEz55vjvQ94CPCjQVdSD1F1eAxqxTbhYVM0YcUXuYXEPtGe1iTiENZ+Ut6SyhPmMFbd8U3/+7
fcO2DAVLklKB2gocDdxmyItTRKxW2+Z7DQfjOw2mUoH0mWEOV8TqKoe0+UwGYR6/4VN/4+TNks59
qRL8/g62EoF8aTc0x7AeTHuH8Qc6yst7CGCCUUuMwTJvcmsocG+SrnHVZYICNCtNDQrA15lc90tU
HVHlIDjhuSZ7eNtbISn7kP4fVKqghkmGSNuRavswV1PrmDNol7Rqi9bp1Hbin2NVBlqSie/OwYTc
F4hMItE+Wn+dRkGtEdLs5sGtXLFzIjKTB3DBltLTIH3OBOl0w6AGRrw9NsSZyAXanMOFE3lTX9o5
LCUa6MEq7XlfI54pSpaArmuSKpa64w/WfJYaZwzKjqLLND/CcVJtP4nuB16v7JseMAUxtaMaEvD+
XwHWNGlFqSOYwu9O1A0Ci8im6JutLjncu0LnRlXDP+8HB9gK2O8w/BwwCeX/xJlf3xehO+/VL5GH
XXMYSaU40PFa7GpUtuwb8xtp2CXUgVGr4l9vHx1O4DSF0+pt96QJqhTKKa32tky113MdF8fG0Sv2
JAJoo3bu801bgfrpMGg4jOTW2mP0Rl2DuX/peOlYLWoVYMqGisxKveDEaKgnrwgEujBQSjtzw459
/7qrWa0fRy4hHXMPeaCw39Cls++F7XTp992gE0hlAbCpiHJsVSyDOPcmDTP7HYusDtmZpWV/rRJ1
GjYrJguHwBxFj3+XA4Jc52rmmVb0QxB7fAOSekhVJW+epabQKzEnUHmvA5SOJ7QWr+jwrBnNPKWR
WK8r5yuntKApApxW1GZEyh/m8xfcb+S1uKnRKoOdMTQc47nT/+J4slsLpbjNz5mHVu/ADOHNRn9I
1DF/bUB1P0cUfs1DNmIgM9ImdaFZz7DSJ3qdNVU/Cty0j0kzhHg4aZujSf/6g/tRljttKlwces3O
CfAhd2lP5v7/OyeYYJPrN8fhGDu9jhq5yE4Vu4twu8XwDwhe86sypy+rxNpbyq0FXC8Fc9J5i9ET
7xu3KpKe1jqgOFdV5DhKMk6hspfPuMk3GfjEqiqMThw1deVhsT1aP0ZuhmhyYt/gJn06k0maMJ7g
o08dP6o7qNXpw8vxyCZnNs52aSUIdZfS9fkHkGHImDpokNei1W3CeYBxOkTXH9r/K4sjsG7oLJJU
9aLBZRSk/NyxvE6AczM1MshHexy5vrKYQ0InpKJG2snCQQ4hUG8nND3LZrY3ciDbY7r2SPQ65stf
6xpz9hkP3DFpr5l6GGDoQv3h1TJxUeTXEtM4Lipby8LfaaltBdZe3wxiKIxg716/8vhDbBju5a8b
3oR1sxi43E3rJrxKmHBQr6mbo51JNpZHYr5JO7ooYzIo3UUnd0W8g7EZagi11FOke1wOk+HQLFhk
9DrWSVsAqgHZgZhHp9xOIsDPTQ1lgbVMLgYifvBKUYFFJdprkNzY7HN8k/MtsZjQDhSmpsZydCfE
fN2HUeka+GGugNz4zAsG8EKBsX1/+5JRW64CIn+K7caDrOjvb36od8AhSp8Rwu7WYyHSb800Ra+S
ZP6AEqoPgDhWD+glDUzIflIIzDy1RYbilFuh7vhrqs0bApj3fP3slRZSgHVIkHhNvy7+CYJstr2K
ONh72ONBArY5F6i8uwm3rOWew1OCGECniBxR+izQ170OA1OqQpCuBWyRnRlLrky8dsn2Quld3e1m
qqKjYJ5EMiOAsKQzUTZ7yRa6PKoiIvM7++2Vqz3QQ9L4WtQK3F7+zEuPfh7dtdiXhgQhl1VsbyeU
5VcYCjekzu7OW3QeaQOkpBsv0MvElIUG8DarMCiTrsZyrghD6S5On7o5wy5IEphur8o11g7x9M7j
2IhUq2Bwfc3W16amMpyHzXs0QDQpmJnOqzYbqmRTjH3Ml4tvqRWdsKOPnjoGJzf5JtrkaOARYcUP
A7Bg9gliGed6HLIOh40mwWEllTjRRDD6DV6Lxw1rlwcCKsq2Rq1XtPCJNJ1WCnpqNl4lHzuGybxs
Y34ZwMZy0ruw4tZe4gMx4Dn/AsFM0QKEag9+xG2eBREyUQfFP+2UhbCN9DmSXvxbWJjxk+gqrsLo
YC/6C2V5uVjqRwqM7c9Ux4p+4F+sarU0FnGWtTxubryReue0erWUNSeBx0VpvKnv2OjK+KWuBDkS
vPOfcHLxsIJy1vVRGY3VH4vUl/nip3wJfQnLtc8a4g2t8isNlWIJvo5lNu/GfFY1elXaLQSjYgAU
JIG49aGDx5mq9SU8PGZttq2cJxdTwDm64nOQFSRBQoKq+PMs2H7ktbIBGEMJTe/hSRjqteMXUgTq
BT+qmAuw+z/BI/741PEUifA6HdUkuMBsm1Ibi0DaCb/EAuEF6/OSd5Dx47o5V5DckuQfHsCYRwZN
Dl9YC4nVprruScisJcfv/q7btcjvsVe9qtzvPmDiXBfpLEb/fdvi2i7v3oQneW87bV8CikvQMD/q
WqibvpptwQ1M+Y1fH2fqKbOjcMiZIBg3rR3I78d2gTdVjqQP8cf2tX5ErjWnfW85J8VwCNf3yA8c
7jltBLWk+dQC1E3Uhy0vV7IsyZty5VaZqRA4i3ctia1U2XaxrIihw2Ytt2djqVtJrHkVHwR2pcYL
rWBk1QzS0cwx6v4VOYbERsG8mtNyfZiSoMIaZYQNPeYkI1bBKUpvGfaj55W+TBKwvRf9CN/lQjem
q8bjYOnNPeWk0du5VUYXF+W+qW5InfY8uDF+MzuG3C2oCYgVnO5aIgI8YPSh38l7BPtRDmG7hli/
uzYxgCalLrL4Cnv9In/SIX8TbV3ZmP252DvaMm+szKDoBWctv34eX/VM0LMt7u89PcV9dnZyAY/Y
hkhQZDjEoCKoG7O10Yx4Vrh4si/m9QWefrSf2zH8BTMqogu5XBXk18gJ3MkoIQo34g7m8HiAiv1d
8H8cfwBhF6slQYBN8iSKowOe2bWWPBFZdDjguYi+RmIlpC+ky2RtZRVImxFl6NTsXqg6UzMnKWxK
tVqTo8Rl4LofYFeLCC9aF1wBveog9x0wkfxs4Zpv1lOsT9lSEMuN8zOUrAfrpr7mW6KD28XSqLb/
F3Hu02jeftxs9JAReag44vU+b7f8hr8MI8AtaFerdK2o1YRIkITPjSrRRmHek5RTMy5sn9ZxaX3D
o5UnzQmVnYgpYdkqn+Uv9Ip77JNMow1whE74bUeWjayi6+cs79KLuw0b5dIghd04Ge9xXQVhvSAH
spodEItxKM1ytKsL6iV6Nzqmf6CgnAklfdFVpz+NyqqtFzILGlorQKCRuinC/ld2y3iaAoqGyIiE
OFfOqR/6Mq9GDvfyXyE9hdDfe+Jg46470NCnAKJO6gaeOcstAW54XogLDQkKcAVuOiJf15INTk60
HTwKRZewSeu2qO3JlzW+13vadZKLDdxYh7FJu6sUfapTptFsfKi9oho9xsEOzBGlCtiK7OjjuTSl
EcQH2bCbzLHVFIQQQDzlSFzXZkURfgMdb5HC9QwTp6DVQQtj1l3cG7rHHL2Mmvak3mFernQvQo4j
CZxPqqofC3IMKIEWYHBkB7Rq4H+VVOyL02t6QPfSs6iPpqnnIFCykyLeqptBvSrnKSySnabQFWWc
qLTgthaZRZ+42YoFKyClztNTUOOYnhaWuXbaZIt3H1N8GjyB6GX7oh5JGc+JjhMDrHM9HCcTWedK
am1c5qZq0HO5TzwZePyK8RWpJelGa92xRoI7lbCBRyrwCS4/QIOsf8AF4nLhxQl+StARmEGHyhIs
kkvtxvUSRLRhYf2P8jL5RWc8M3qvG0J6XMuhADopTG7zX8mwvh62JVmFZb7AueOKJzRk7KDldNVt
Kmal37CBjy+s1Q8NbScvf27VWhmF4Or3xsR+o9CQkPiR+a5VZztBS6RXxpgu+BBPzLCnP3ieCKAQ
GlNcaLZ9xzmvfuBgFg4tCBDtpuCwyVXKwNmGTGl7mFMXdkDVBj2aYwRkT6de1tLuWGu7y9x9jjnW
s9RTxr/8oY8ICOhutG5WN3U8aqAracmo26FNKWUJefW06oEuBwcXa8kI/rKDInHD2tG/O6xmXIrM
kX26c2tZuPZuVVaTd+Zp3ke1DgiuMi+6dfejwxm1sGBwHurYoGo34na0xyoqzCz1AvOOf+M5O1/0
bGINnnOMRpz/RGFCQhEI5x4JAtmm8uCVCS0+4Mq5EIl7f2mGOpm9X2R3tfuxQijeSvGllD9dvc89
EjzKmDAqgvcOM9iiusV+npZaT8pzd0w7t/fDWQL1XzFajxfTVHvghZohb8GJA4pcUgIk5MnfePIt
JQ3B1d1HRBeo7Uuv4eY7nD3FZs9by7o4nXflWUA4LGPEpzeF0fVDc19bT6rarrhwrqbzAV0CVBc2
SGncvUQ48tUUiBWlL9k5azY6M+Yirbzc7lB/gBSvm/pRxxReBpfYo9Z22NIiZfPLTUtgFBcZlF3y
eVzq+9mDbetDJtdk29zU2puv0ei17LSH1DG0qErJt19a8MT83ZcY+YPR7E9Jehyt+Uyal8RR4weV
DDkOqb/fNX7g/aJyuV/zDgwoBEjqWOfZrfHpX3YOtgKpUI0VGAWkZxNHW34uF/82ompL4GvVeuK9
2itb7Iq5i0jozzbVod1035QH1VC8Ian44wjLsT7G3pqNO1X1EP+952lsnTTun9XGR4mQxtKkprBd
CTJEBCJGVeWgDr9r8aIMgJOvbhNQpv8FLn8jBeltPNOdoI5Y/0xtjKwKcZv28acRowRObNOBqyEL
tQ193/tGVevHXnvvVo/XwZcd7WBwNyaChHUZmV72t/JgflA3B+TE7opoScThms2YaHxymTxxGdeY
Ya2clhsooKqkcDCNErv1V5bZZV7kwE9n4drPdPqe8QveE0XpmjOh5vSMRNshQpx5Vj+eDywItRfb
GV5/+kNOm5XH2OKDXILZzgrjsn2N7egB9W2eni28ubEJCM1sxI5mqUcLrvpC90rZgOe4Io8itpjP
cWjTAUzmjxpbp8lxejE+z++BRoQa8ROfKoabj/ip3Ga8y2iSaEs7VlrttypbOWf1cMUsojUVnq+S
+FDhRemUBdUgGrPo9O01WG1cCt5+MWsfDzdBZiEBfj19sUWHkfU3hXFvO1qBFdHPWSvfJmb7s7Ad
JXFCQy1NmDj1z+OBRPiPXndaEUDKC8tOAJ0x4IUBjvE5Qs7LqBYwVxkJVK4mnjMCTWEpi3AuuD7S
32xH1kS7JoaPV4decz17tAsPlnYRvDKTEmISdqnllgpy2aJeaoRDvi1MLuu8r/PmmBylp48M3Bev
1BYA0ASoJd6Fzy/nsC4K+E168NTxk0ENSvPKa61niE8yscJSQoHYnH7RHg4oBKcLubUtfaSauQXW
iKK93p3xhno9BzNutHgyawJRBlyI6oMq0pVRMLMset6ZjvEBxpMaOX6VuC6ERgDFSN5oB4fSS7Iz
amLpt8yryhUqkDjC2PKk2GOM08ILHpbAkNKwRG6AHbTSmDZjekWfRVB+ZHQzvtwSrYq4zxKKbM/0
oR4YJQnwT/+HLV4bUl7m6BUGeQNKNALTFynJbiky/pLZGRVvZXcUG5gnbRJyQYI32Al4+ljLCSFC
WkDEwXGPTHBSfDKSFZlljojgnH+npQ9/6LfHRI/xjuukny1g9LUYGW/00YvvwunulxPZ4yFnEFSa
DW/zYZgKVU3xMaefsJrvAjPXItrP8aksTEZJ0LZLBnTw7CkaU8ORfnAgHFLoeqDsYxV4GaenMkT6
kliTmdRykeuznoHR7QiwZzlKm6rE6yTxNBgM2cTcBoYMSfF0C4Mez3vnVA8fORasuDrWDfIdTFOS
CpWyFhyoz0mr1yijZx1VJhgX6QBYygD74iGT20ZHmdx34ZuyCxJmXG1ZO9vDXx0/tjov3AYnEh0w
uyuqeM5UPubfz3Ws5X6PpchfT/cDrj/jARcZBnmll5Gy008/Yh+cDeufMLB4fFNaYYwjTV9oaLW0
mkeKjtwc4Qw7KPnOOrZsar7KQGGUlUNS7LICRy6VD2yX6JfdD/d73oRTO8RwH1qVQFXpEyXZf9w7
BahpgKpNSbh3OsuG7lsnwDMMzRQdyB0+X6vubEg/2o35rhLuloaDuYgHkSjKUIp4RbXuNSJ8Q7zw
yYs9G4TO6UjiXxpYap/9kZ3lXkNgCfziB6BzHsyRmbwbVelhEFwHhtpVscd/4ap4tEdwu1Kf+S/5
NcNC4yD3NJ3CRrn6DIx6OTKtyXTWASG/bC3ZjL0E8AjuxMJ90i/KeLknsC9GGMpn86GLNr7EWwaq
GEemKO85FIDhV/fwxgxgqaKSPM3QsHZK6BO5BKLTeyc6RAtvUFrU60bb+kLreqxPRDFWzqnmSgqC
r8JwkZU4MYFSl+HyICmG4lRDjW4np5jbELp6kSV6jRlBGqXHs3f/PMBl1O9WBRicr5by6jsuZdW8
/2876gcuzg5YvN3qvnv8Skive8KxiwjB6HryPr2BYnOh2QzsieFsVHkz5WB6uoTJCfxcH4Uyd803
sfK4Y2o9B8UdaCyPzj4ffQgt1yLK0GQYp2hzlS3alxRLss+/fRPqOh/INb5dao3gT2+Ej4jf2SvI
TCvfTXnpDYVD0fZKiSb9ogMBfpkwORhi1pTA7F9f/INLFKOuOuwOs5FliVjU5JPNoW3ij9njsK85
C9bEQyuVws1FTHb3qt+aVEmP6QTq4WWJlbSYRe1RSoS2btQ3VZVBFYubsjJH5XMNsOUJ/qgX2s5O
B8JWQGZdq9gAE7WC/JHtuTnzmtwZei7HkUSAywTXSQgtjUHZqhiXcKvIet61/hus2aJG4JFzYCfa
u0TKbzIHdKuSUNlJw/f8BaHNjQrwLSolxMhyHyYaG7FzgAABOaANSs9tiQlY/WzZ+IvpkOSFZHt7
caGL/Z9NWuuw7xzw+AEavvXIMg4fKCi+Qr9CiXqE1ErVYvbaeqB6spq6s6dk3M4IDNYWj6Wzo8Zr
UW5IpDEgfZ0B4GUJyrT9txEQ7dL8NN0Z74m6jMNqJMEOfA8jP9dxILo0FtmXcEp0Crd1H9eDGrcd
XixHyFCbr3tDHnmO2ViogOqJvr+9YTP6dmoVxV+AkcLD8ZjnYOMy8FMx6UwKdbx8AAIvTyMvQzJd
zQMpXnVfI5bq4YqS/L92kRXbBWh15oGSoY7vJmHW8wmEIMfaupEQLu+mhwOXtzwMBADE3HaBpHWq
9HdqjLZ2F2M2NqWn2WKXcNAGVZzibE/mxUFD2aA8kfPW/ivlctal7IFUCTB9uf3aVvkqwRzKtVhy
wdhrcPRnD5UmHRo4EPW1tPuJI+cQ1W0tD7PRVnEc2lVRTs8kh6gir9sY91mpFm94GhHX4mpEUSgm
FVmDyjs90nXw+r/qPeCk2vglw9h0DNGo3HA//2ThkrLnxifydkw0w5Pe6BgnhSt+POIHQoekH3eM
4J6cej1ywv6Ho4jRPh0W2gFmk4RI3AqwFKd+8g+TgB2mUCv8L140DTFNGCmjrHqycyD8avUpxtAG
mFHtjeVyee1/4aUOPsdRL3ehEfmucFkUn7q7rCYirl7OyDLKF9TvLEsAHdkb7XgzuuAwPPpNMYrc
e6g3Hjf4e2cuXkthnLbnBvIyFFRCjizVrJM8p/yjwTePsEMACXErlMoOMRTaU7vXWMITLfKdroYo
IRfKZ2toRLccolTR6TBGPbgXBVEhJ3yK+No/X2CTaTS+h5kHYYgnabUspgkIpunrwGgyOD6ax4G5
H3DZCkIicOtdICJqTCiR4707k/lJ2C0S9bkVK7vezCte9yLvNc9hzgIm/4N723SuAsflERC1P/FE
LxlSIOxT0CAyBu6aozlFJ0oqlyPRV6Kd9WwzB49vanxyJeIbH4ymybyCqf7ov02WHNlXl+FZ6bxH
FwlDAxwqaIPckUh/z4AukYWLct5wS74jbnsyUQUsOurZZLaMvdCy5ggYS00PCed7S81GdLN9j4Sq
WXQweneKyvcZq0mm/hXN5gdn5rh8QAIE+vwO6DKu60T3aYx2JbusQ4jxR2IkMBXQl60hK/9co0dY
dgPGJ9PHW3CuBKzU/M/1JHsmx7vVwjUPqFMjqUWN54F/6NJ7YF13w4zynhGeExkKlBGE7R+Yp+el
2NhHk274qBXck7+U1EwWff0Q7ANXm8cIhfvFt6/HHVv6PDd38HfSf1WHxEKPSpN54wMsck3DIeTs
Op0NyqdaFyhCvTzQMu/y+iUHeOg/SXTLk1pxmelWuBLFgefWQ+T2CETPeLFGl3pgn4fA7okkjDE8
YV9S0sH94G8b11GorpuW3bsPAI77jubIWZoUIFoXr/IDL5nTmaVJVbQalONCzh9RLZ+I/xfDYA7y
euZjwFh5kvgpLXrUjDorHDovBGPqnGCoM+w9TWmJlUZOK2D1fwfZVyf5Tqe2NQc76/lw98yN7Fm3
CZUr6Xn78B4ax9jQPehsuRCHhlKV98YYJBPCa3s4YnQ0HDDZkR/oCFQSAVkSu0T2wJQwe3kM4aGC
/WRFBI1AO/s52R6K8Kbjb5uMUFFof/BiPtP4lv2fCLFZ72YZ3WbgFQfbz7snrxEoxe77Zv8yEXvM
qlCQOSLiyB+Acqc7stLyslA4o0TPrqwHmstavG1ddWBxk9ILDtANLP4R4EZVdZG8phKuyFf4OLjH
BYJVGs1rezxp8b/KwJLYpvd8szzUFjVq8FfRG2CoFTTymYXnINf9MPOT4kdbNAXOU/ShTeuFAC+N
zgs5rhSAREItzn0ompC8PBM947IahYG25iedAp5tTcDIwEoaDTTTGAn2kaPlxwEgv9ZxGyfe1XxO
899sPgEgfNCAhhOs/v1qXDJB3KlLYCq2f/ILyV+260Me3jgiCf/rAIS58xBCS2hIuziTJNlN5L78
UvPWBH9hqiHZ56u7gdz5z/0kIr7zm6vL4tnw0dHfPHqUYkE7HXy0uIJdb/s2swPgC8dicdmcEC0L
WTrpOQeo2mMvDfhGMi+5MG6A5XBFL0r+isKhVySBTEyYyX8MaW10Q7L3lLheR5YPI/QpcRUpcpMU
LUHAPHPH+GQlAT7oD4sYPoc4nApqyxvnrqMRFkU9rkYbZ1u9D1w/OxwZQKzC+1mpdpDMLMv9Z12a
KyG8pMyhHEVKPqJE3pfWBZwRQdD8vkREP/wR1PgIcWt8wKOKBXeaSjh4o2WFmHubA8JKRCske1bl
V3z83EMlVAXsXsJUo8/32WN9Ef0rKzj2tv7bngics2vgFeAOkJa9t+ySXpoSoGtaygIxXd5bGPOm
0IzTfTkHJYytk/Z1Qnor9gcSCmwLzXAKJOXLei368lW1L/vz1HMzLd4f2ZrMvPtBF0xzW0/K0K2T
PhWRAeFgcUckeVkVJv44m71W/EFf1OCyC9Xg0OhR6HgccjYtKaKX234raZ4MhIydpStTweynmdm+
+efLGhllhoHs9Forq7nOEy5yJ0vpjLWZRsMCiSY959z+ni0JYQI/iqeLPu6zXR9f9eBhl9CHqZV+
pRrtMHUC6jFFK6nahUt2spZZtIs5MD9x6PJYdBEjmkXq58439aKCeIKgT7vj5SuTomRBDzQTynlZ
zEwuvMSYp7kXwgSHNFkOjXN1oT9OZpdBGGWptQte58PbjXM42BQqYo59lsTt/N2DQt27Lkraps4J
XCkyUViRF2FDJXvgmziURLHeYY9qN9XhjfIbrqcmBwVRUbkJCNox0fBaQseWyv1N2VffLHuWorCb
qqbtsgt0PIJrHtSQ1q62ViIKGQKNj8oH0PJl2eIfXTHZnk2kBUieOyQU/1EgVtnXTkQl/TNcfqVw
3SFbUhy+Fo99MGNnaJ80u4ECiD1BjmIHR+fo048WOozjmhaJsIkIX/bxv3axAZGGHahSIHzk+vwN
QUvShCA6eeQQXnu1p4J/PK4NCIsxgHVrSRRbKAAysiARVWrlEO11Lt41wQ0RY5gHM4ROtGi1U72a
ct8sa69KOdJ0y5qmqWUa1PxAOISfiDO2B1EDQbWblnzpVnV136QqNV92hS0DxLKYbZYERpnceTcI
48KWvtDxV6Ua5D8IGOwdDh4fwqIVnDM9n2qPEAcv3dVqekkqkXRpb1zUYNjef7etDe9BO3WsY3Oo
oUBOCAGhjSPiaPvjWjCSybh5BBorYbKFGr1srZabmFij+T2/EOmrRndpQaHKgYsS+oTTjWcaqmIF
Y2q3kXcWIGv5EEnWIMh1G3cebetdGmCs+nlfhTXLNmqNvNl7xtSBu3bXzaiIa9LuQ1pIzaUfSWbD
cxNB63g3nktKAC87tJeszzO4N/xlsjSowdTGZXl4e8wgE8EbpVUIqK4wHIt5onzCD+ygoyYRdAiq
lb560Nm+t/PowFbo9ev7Fb+2wI/Mt2R4YSL9tj1VBzdbX3Cj4k/ZW5kkdcFAvovkRIhKsAeyCb5c
HVtUKCFU3f4fSsqh/iPMajLggS1pNgDuNsm0LFqAW1+N+O9/uCgid3kcRgDUA/05fEE0yHJqYhK8
Mcz6p4Tte6sQGIrdFEPvLuZ8IJGk/DvvsFFCBsaQP2V8fNhlT4JpB2PCrzsjgeA3iURI0TT+7RuC
dkGc6z5hgo8Yc3nPIRzxAu+tPxMDOfmPN73jZuYY7K0psHokjxLw4xi7Uu3/pzu3gK3gnR0xjk4O
wrqJhZUwaGY3vCsrkcohn/DgHHXyecvobR/J5HuhoUp1lvC1EJQsSo0CjypCu3t4uPrwdsacfaa+
dw8CN7fT6MJviO5Ky9OUs5J6jxwDTatqIaxUTfFMUiedOyw6KLinviZCl9lIXZ9BZLEgOibFhXKX
oPWPHKRIaB7HKVG+0w6haIzCmSVFxyKf1q+lRLYGwNaZ3iQQw4VQdkz5dJ7IIF8N5F9Hz6xhU2sQ
i32oU2ec5wR6xPd+0Uo3wNeE5PjlHK2DkUdWQdbjG/F8g5im314ztONSf1dm+LrmwtPds+YH4nFi
WL/DyXzFe9HLQ1SecvD4NkfxZXI8hrldDLIu9Adff37FBaaK1fr1m3VZJk/n7lJPh8ZrBDoTdMzX
H0MlGgiaxsOimdT7FnhNyagYoS041ehEGtpPqBB89G50r5zLwmanQ1R3SXqsaBmV94F3JnPUuQV1
RrIYiX/I5alnSeXPomalPm1vGNjwhqdam5kXNZ5Qw9K1k3/uP2h9YnsVuKRLTp44yklJWwsg4Ynn
BUZZ/vbcf40tD0kC/7phRKhMMhWaAcI579vUxVKvp0qZ+lK0jU+XFjMWa6LehlyMULRg0fa0OgCS
u7I9Uii2Ofo+YlwS0ldXgqdcwXhBfgHdTNq6NwWidfqQlzmo1+gVYFzUwVn2i3eqvOv97baVAoDt
ZVNKB0grJTkyjFdLpgiBtj16VL6xd77p5x4dXyGvoeeKeyK2MiSvw99n8JqbpVSfOZPrbjTxuXV0
LBIo30b7B3aeDl6oVh3c/wEX6pSOSdjVlOMiIteKUQiMQFHCOjM0ScF8E4sk7ZORU0K5QMxNJCj3
YnborYEZ04+My4ZitNApJHmrahVcwa1Te2LU5RVBgQq2hQ7dlFZ0bYa9hShsS/R4yH9nr3uvwuqj
gT9HQ1jrLb1GAAv7kOBY7Wo+yLahypButg/aZ70BiNLaXywRMeYNiLrZRgAssz7HgUL4R0kD4xcv
24BTz/FpdMv0B273pYnnz+ZWGgnWew8tdfJcncqNr3bItLYAcvvW4vXnFYBcmkILqauzBbSaxOce
yJUCg9NRcxKkT/slmFPzEOVlQqHdZlNUZJArUmclKZO1ethReowUv4MnOJTfUcDbC4gZSzI1PzTN
mG2ZQ9DgL8zotEOonM5/Ok4sEVwP+Jh9nrxpxOgBy94dtoTaoym8bhCMdtLEVthDgMjwvuY7NlHR
afgEDLg59rwQ/nX1FHXv/ES+vgH8zcI2oP1QECTGxBpqTUolAUE9QRbeiIGYDCqFzcs7NsU+grwv
A5BEiWBAVX93hfgjPKJzBQ/sV5BdORId19G7uQnCEbVOvYw0OnyDlu3MMysaGZeWEWGo3T6yaQFj
NfJhaHWWWVn5LUGvKLI71bP2l6aP14/SDpBxZdRWK0BMGcUKflUtY0pB3+LfE2KvGBHgzZ2zzez2
YPWtq1o4mpzvmEIm8mKlJ5kwb0JJ4sbSjAhIsPTx8aSggfz/yz69xiu7juJCNkQHVuV3cYLobVvC
uWHFRerohWTZTmuQqIkqdIFdPaqzY78jm+qcjTKrpL3j/4l9YJUagSIFtxgHc9lljc/+wSwNp2wL
Tz8OUS+62Cnr7w6HaxeqYMZgRVpCJfUjf9rxOcmhtYWJHENFNcj1vq6S+0GRYb72sa1UmO1WKy9g
pzJhKm9RyaD3zIycmr6QUiEX+lEa6qHDi4E5O7iMTEJtJKadhS7D03d+SlV5jPcLmC4ayy+9Yre/
amTIUD0nSzwRP798Op/O+FHEyj8Cx+zyO2zbhjhlVIP/9QRABhAlY0q8PYiJBgwyyHArOfewrCoE
aCO5rsCeuJ7q3azUrLtWGwC0vG0du5j4YJdyOPpr8rAy42mOdxbp6pjsVVozOt9DDz61t/264FX5
kOErirnyS/yl4bPf2bvFX5zykziTlSmdFquQe65RlL28Ouvi8TrB1kbVxblm9ADtS5jdLEVO9cJM
ppxBETl7ItmKMJd+4UEnJNJGXDUAE4RlHjr4+J5cwnN9DdE5w8AzDWhs1gJcLbAetUlFdBz2qDXP
DpPfqBhYJq6jqo+TSUms/vywpGdj8ID0r/qG2RjKwr1HcHbHcjTGG3Nd3UIfxomy7go2UdKo/RhK
yEgjBCCZNj7e5RaJsMsqmit3dEUSnuTOkuZ5Ji5rrdXW8VrFlUM2H8fUxNpSFXWhVtW0G7FWkEx9
dojKHxwzP0zg03c3ZFlNmXEG23d+Zk/ingmP6nVc8Ds1TkIMqNuN2Gi9DHhvAy7Lc2svxDAEMhSa
Tydy2calIr9AU0e3HgOE8qn71TO/EUv6SkzJAZo3jVD2Zlm0cMbR97M3AzMmtMdIq2z9FFurCihR
G3Vwe1JFggkvFiC0Ql601G0YQZmvCfuOZuYd8GShFd7ElYpBUGJPlYB+XTly/yVc5t7eq+Ax6O86
eS3Ln+DIs1qhUObwjBuZBnblKHBnCcNiaX8Jz1SDbjMBA//+9jVNiQp1omXsC9/6ZbRHhG/TiC4r
iJnr/f5+meHgo3epvGcJQ/LR//d41DIjTmFY1ZG4Ex5tt038H+A3jWzwEE+M0yG3iLVyyqhQessy
OMAbwr3oDbXD037rHsPSwPkkCEzpDui0iI6I2sc7x5C5uP0bbHAe19KrCvZ4g/xErX8JxdJYWggV
M4pfLMNaeANfeIl4KXaOK3Ej1d3X/vBGFJ6gwJnplhtEKamRphTVfClAgGtsVXDwkqeB3I/ft+Rd
SUBtyHRXVXKHQJLKGLAeU3J5QJdPYKgU7o45N5Ob2G4YgZ/L1LJK554SizK5HMlk9FuR06+3lJjS
+FJqxuiP9KbClSAE8KNWgNTyk5rGtji0llH6gekvsD3sS/OfMZdQ0PTuO+Prr4Z2QOtoPQh8HoKF
1wOCOTgywakwMqqaT4MStl6GyU9ShIiAQlIbq7gcJR0TNjc0HCi0BCYfRa+eLbLb2Q+4YI6GRYJL
INsXB+VWmMRfY9vOjoCHYcxEDovdppGeC9bpFYZGL+x/dbdHgTKc0P5hpHyVNm3DCpMFQEIevxpT
5c7GMa43NKecUTY6hwbZNYnRPdnuUm+ScKAbHHNONTthIZfY0BLbhJqds1uEFsA2YHFRIG7/w7Q5
Ru03SQ3i5O/p32mlAZQyv462YBwhd8To9NkdN11tg9Wb9lBaWP4NRSOPPcVVkpSiubweZtScw/D1
q+S9CUm1aW7t+h911+N8Nui9U88RZ91hgePCH25zTX0yTYtPX5Kr2lKZ0wuz3y5TzOm4mAeLud2g
9R3m30UBiTG5w2fTxRxDg5JwY7FKI+gXqGC0VJeFtLwBnqP33DVZmUm79w2OpLJQR+RUTXSYD2Nu
NQzkRsuNHjhEZZlUYaw7R8N55kNBNGoDDBYwEuhSqFr3vu5xr6wA/6oK6JW7R8WOPnZCTUOFX4Cd
ieW0OzpNsMM2ziElp36kOA0mCOxX7YPVva6m1UGhwYco5+OXtUB+kJAVlYAlVVswZRYpW62+ZnpH
7krXMfXhnce0veKf8CSDhz8+ihWgtAuRzVSBIy83nmgmEVc5SjVkBG1yEToEF0ndHp2cZiuBRgBp
3rMjkF8Mpvc3zE6ZdnTZcPMqd0xLKT64GKPmfBupWbRRb8mh3kHSTGadqyaQCLJQyyQqmRdStQZk
clGjjifmM5z90ImI18n/k4JhmQ2bRbz0ZUjpiwD4AiXnm//X6jaBR0k60cAh0WjRMBGUaAAqMFpb
Ka73mukYuuFSf7PF92L+tGiiCIcB7jcc/M6IQp5JQlDCKBOOD1D8IHQvMTTGEw2PHvX6AmX5XJ2u
13IEzLbovbVopPFGZwfmg66yXMF+wlmp75GHZJfr0rVPvbkg67/pAiNm/wU5btlYYqTUJau6so99
cm2RDgYimN6vs10Z6+hkz1f3hwL+fEbrEzEWriKODA/QzuIui60rMJgSGcg2+u3nbFkrs0+hG0S8
TgkmY+u5ECMNLWM/jxfMfJkxjNwaxULf5wWtmvleBiTEFYF6MJNfwC7ZqHVUS054tnTCVdMs5CAI
ztK8tE21QwuNFlK0Wc+srdxrAxDHrBB2zHXU048W2vUYrnQVwnWafZM6rkRsfrn96YtxzMZ4V0bH
g2sxBmH9Oy5bbonUcx3QaClvVcDtI88Z1tHIDZbJ6fBzg8dk6UKrp4m2rdHJSXKVojIC1SQrzShL
/v6P47zFn2nohORAMq3qAwnmWjPgN98vnwVDWa8A7EQ+fG1FyB985Te69tWf4FK6cgFec7FPN8Oj
AFh6rPNcEdkTDkpiaFOVNRlAtuRbaKsiabg/5TyHrE3sqT4/ab0FsNxIelQ4onbwyl5Uu25foF9r
P/616ju73J/Sll34HWufH4eGf3hAxWLNGG9Bu0XufdTimlORzTt2LtSD+Y6dXupfjpS2iZEaW0iJ
Q45S95XuW1tAgbUKqdBorUo0RcZxPWZl91A0Ql8vXAoH4TdNnLZaqVEXjeSEeN+uzlgoOH1bHEGW
sL19cz8PP2rLyHJu1bsnaDCxv9nEDt8apM0xl2GwIWYYhzRDOuKusGuu4mLB9DaG5IfZys5HqEgn
CRCjbN5BRNEzLceGJ5EuJuMI8wFxcqJDqemVMinTNgYd+k4G0C5X8zMBEdyoZYrb1fc4DsWknlY1
X4dzPLVx8ed8TVMJ2jU3gwM0/6ORrgCZLXfySXhl0gOCmZlgoGkOKVqTQI3FSNPZKdi9/Otb/Mly
ppZTt+5rjXLzMtaCtLCRNqkWWNlCja+vXNwF9BLSbrvScZlKtYZyIqeWmxUhXgRVWa+8Ru2ZjDOV
2Cjh7FaSundgepwB7V19gozuB+USDHmnfiVfaBW3nj238w5C4CN+BJ48dwJSorQLq2oxiZgwfkWu
JOu86fOk3wsFS0vXXZ8LJCkAQgHKDUfUFsvbTRZWbdS1Vk+2I/ziZYCRY/iyk3w2lHyuDRvhfUlx
33P/mg5hilL/Un1B+YZkDeFuOWeP5IQEDmjrt9tKueZosH4oAwGJ7EzSghyi1bLnz7Rjh0EZP4iI
SlimqaCKWg47ddgFYqSidloZPsskBo2gqfpq7+TDkig4iARuV+vie3bZCqH1prRNqeObi99XQcBv
23GV8PPG/faMtP214Pg/AcLXTksHjDN97LXjo3UqJSWXMT2Y0vw3isT4gx3ToXO9Kua6ff68QSn0
KaUqBWXP/0cMLmCqstuWWfm0kB+JcBhxLSyxywtxZ+hAM//RwVUK2pnN9b5i9rJDFr8U1C+5eOw3
lek9CogLoDBjTeeMcK294xImTjz/+z7nq5uyDA/SmzEKGSy64KSNG2ohZIGi/S4QjfZC4+sWf9L9
gb8roSkJVa2O2TW+2XYYA9LqDtVZjXNXAWPnOCtEldGjiMhN1V5qcfs/8XITglVz4hvSqzWvpJbk
aqu23zpgMwssl6itE3J5gG7DqgHGQi9uY2g8syEkoLEzR3goOd117wYPTAdpcW1biCKNmAQQPce9
K95e69omPN4J3iSyRSZWTFVz/uYP8iZ/2zf3GHiMVLqaW4q7uZa3wQjeAWeLdYcvCTuhnoE4DZaX
lSzW5ZPta3S+z6o/uQpcEeSEBd0Y51m1GK9ntU52IYs2xhUmN+A61pQ+MAGgQifNJj30l1zLuqP8
H7u9COBgIxycHrtdm5YtISvP0xTLIdxx4Z9GJB7py0c13lMZTGxJWbAjbmhNHmU5UFOwsi4rU/xq
F1ukc8VBYy/f4LdokPbh81lmaMH8iKyylZpLWFd5tBjLOKDTAgf7bdo6fRsP1TudC9rGrdVaxrr8
+chAkSzhmFGuaWI9cPqC+aJbtZdeb2ReFtRZ7jvSf4GOE6zNUBj8zh52u2UkgfauAmct+fTQuSM8
Law9MEY7RZ3iW04XrH3MicEWucZF6WaWAxUpv+1lVP2hkl9YMqW3onJkxrST+sGY0ujv7nkLGeKy
ReO9nmNu4lWzhWRnBhxAUKlIqgju2/uj4CDT4trF2kvPeT+z5ZpNeWrQZaJz2KhyW2stCLgHRgAc
EW/FoCm1uTeit3ZewGbgvnu9ZtOZK3Icyb0R7dxBuRKVjKsNC1D/YLd/tXrgP+17mPf/FZOhxChV
99gzlmxpQtYngHmlCd7WBn2mzkGwfgR63s9EK+Bstin+Z493+MqWbh1V9sY7cDvIxOc+an3LQYuJ
4+p13dCnooL35taec3ahfl1xZt5RPI7DWERJU9nLhvL9GMvC0KJBQb5rThzCcSOcXDiaZ/eG8UCn
ldLFFNAkYmMSsBHMeo+XRIRIqx7U5KxT3kJKAePjJ20DuNg0fbitNIe50uaiR8YRC9q5SjOsCzr1
dqZE79e9K4M5veLrHBFvIiDy0cZaUFt9XDBJ//Olot1VEbxNjQEiWz5+dqGIhJAF+hOxdmSA3UnN
39ZmH6AwNi3jKJZqpNEJjmLYeXrIofdDmEQd5qZx1Mh0fh0qTF2ZQMGGkznOs3uJbJTKvT0a+95g
9jUZPwfuugGNrttM5cejZ48qcdtl4uhms1X0RL2Atvg3VdYEncwAyyriWsKIRm4XuhaXLiKXIySb
L82I5gKOjyXtGxyyzve+NloKGiq/SzoJMdiwZtJxexRQHZYEbm2BHOxcoavzLRg5II0LDnVWpGVK
SPykbWXkDW1/OHA8/4S2ULQUOgIAyDNQMu8bCl42ufLJBhiuNvigs9/j+VCCun5d0OiRl/GMhZbq
61Xrcd+voPTvvY11GXA3p9tKvOGydQvA6X4X1lB8HElnn862FH7p14vT4QUTi+YgXeFkQDm+4W0A
mxZPBgZx1AWULl95uvi+wPjbcCtVfTcDO+AvQ9fqYMN+bjqRhdFutb+8DH60r+CuZsj9HwcYH+Ab
6jajjwwZUNP2mYb4aXUPWwED3KUDhc1P8Yh+Qs5WyQgvltWARqvtYTHIVKy7G6E6Sa8YYwu2auSZ
XbZScraZYntrR8IwInztipq0DcNtqC2jvwOt8DNNIYjk8R0P+zepem87btvRMClRuhSNS85Mv/0L
EkoFJBRspEiMBUI0lPiwMv5bZ7hmDMtDk3i0evg578tFl8qfl7hY5MrcgBBQb++fcFEYrZsnh4SM
eu3KmsMzg6aTMuUu8dD38XTuUs3D0RsrR/AZIqk1iuk9LhfEJ+groxQzODQpYW9ZXhkfBbPdiErf
UnX06cEldupBg/xlxpe5RJsC+RZGPjVpr0sz51X11e9JCpLHac2BLSmifq6KFhVJqyK6641L40Ne
vktch4H9LHax+P+e0ggdqw67dCu0JpCYrY5iOOIZ1xINIblUP9/wsrEcR2JinWkd2ihOF82x35nz
gwbtots9mY8VtTotbPP/XVQbq2EBSwxGCB0a+G7nqPYjzYycmqHH8H+tsawGzUkhK5VfErkZtp1I
eBQemRtw719y8SHmWuo2hS1V85XjXrk5tSNfLHNiaCGLiWb9Op4iH+nNn4cvblDOOnjWb+BpiiQg
Yus1yq/wxiMe5AP6yh2SKNtmItRRE3wx+5nYprWU/K86ez0F/EHPBCPDQnQYNXQ0eEeFqwSKlKFf
DwZU+z9EGMYIiwMGyb4PEL//5XYk48Y6MAjnwYk3KUZuvtGNUocqhePeNDuhx5rOf0S4sUu7NK5y
4si3M4r9CzhHlemXGVvfDKWHdJYKxCh7KUnI40Bbac9LiN7N2ECWglKJzTU3sudYxOmd8Nnn4ZIX
FTE2uaIi1J0nYDc5qUYWwj9QzOX+rCWZ/j40rCmpzh4kBX/q6rFqwM93mRsmyk3zkveoxv7VTzIR
tod+oiOEn9599TyYRPl9ScTtBD72srYqcUAnLRo/F+mNXiSQQIpiv/s/n5k/TNWv/v+ptptROLfm
trB8brMFswGTbslGje09wpaRtycloPcMaCWNwLaXJtOjr0Onw8U/ItOUICaxu0IJJR9TJnOolkuF
jBgITgEztTDjuzPFGupLDvN9P5Y218zSxqQOFH6PjUr3ns7YALS7Inwm5326wL8C/ArRDv96hNa+
kBm4U4XvThgGtbz2X7qa0XOnYExfGMhns5GDlXyv5NcwcQBo2LKhX1Z0L1VTWCURrmRjAmwSKTlI
qc2X66JTNsRUo8nBFaScX4q9uh+IxekSvi3hgbZj4+vc+NUPCrHDnlH5xngHVV/vhi1zRQ9b/9PD
sJpbAW67cf88ZQ7e0phe7pST88SK0+w46pGA02M9tEBEVBOLYA4yp1xCgL1PjwPB9l4qDyjdvi78
+n9g8MDI2tgaOqjeCYAFjnpPZpFUlTlQio1peSNM9xEH2HiOy/7jnPLAaFjvcepedH+fWMPjBwa8
9OP5bMCfIKghKQSOyk3SNQ6xA/xA3ER4eUAtZSJYe8XrZEkcr9WWs5puvVaSJW5y9HsQl7/t5B5H
I8EojvKSRMx4DGI7clKiBaLyFXwlKAi2WhXQPNEK54g1iFubMHAORQ/aojSEUye3beAAHnhXSHBd
3JfJkjsPnQtxg9T+ZoNwysxrocOu0YeLmVOLO0LwunZ1/dtgYFOdAwlIzHhscCFjLZQTEphJLH5y
mCDYs0kebkY2aPhbbOuizMtqIsf3vTsj7BQBKee2JoefSlGxqbLNL4H16GDPu7ti7U814C5Hd5pO
ctqxvZEHk/OWukGfxlHfwWTlfWJxIYhQ+ck64z4McAd4xiNGIM/Y0iJXQ3qCeHDkT8Kk45C411n2
1hrZQI4hv6paFNigpxl39u098W6aPUaL7oThcQMO6927GiAmhD7CvHN0q1BuT++dsrD9l24hhYva
+Mr1wlBCxRN+WARWKK2woNbW15A9/CaRgOF3yRMp+1ORs2moIu6zPTYoWaB1sczXzzd9Rycq2KEW
s/ImkoKJPzzuq6V78aGAclViqILr0e9i8B2uv2PgUf5LTFsFb7O+bcZgojtnJ5LlapZE4GpqoeLD
9Uf0FhngK6m/I6Audi2BCuO0TXqHwrFMOWY4wgyYEqHA+bhLOBGYq3D5S8fyJi76d+kPHZOHkYuB
79LVwETPe9iRp/K2M0zJdBjrgdhqwGFtE3cq5Pywn9QCvmPYhnqU0KHGkd1tEsdQO++8QsQ+aao6
KsqTKZv5wc/vUEJRa9IPMGH0Sfq2T1LXTkcLk2akull8PbllwcLWKhkqF0dYNYo2OJ9yTOb9pOSe
jGQ/xrl4RGiCq81Y00zc4nn9pzEeq5Ng+IRPPdpDOFVoVr7Yr2+OnM4aCA3lcIv+8+LYZV5dRHtJ
mKa69cwh0hwV9pvTzHlQCfhT5bpBLNNn/hyR+BI03E8Ze12RUXaKJov8wUBNB/QmGc4RkRr9WXyY
sWX5+L80mwzXLuW0WRs/1m9Je2Y5/snpPAekEjTn0vM++Y01bYJJe5QWBVPQmDB7/x03gclBXKOU
uROMUP5lz+WAldJO7ArSlnBRCCjaJ0l7m1FdWwvQ0am219jubihaAvPYuNVYjm7g8lxAInADEQ1r
M9CJDexnZ4dBFDPkZO457BDMTWwGN0dpzmQo8BtIf9s+Xa+MPYX0djop1+eXPB/4RsnvTWDLJSUe
dGeM7MRyYCIuJjuAaPuezhmdC0jR0sIsTSaKxuDgzUZ/tok6FCSsTneY34Uz5+Z2iYP8hqpBvFDX
tFkXb3PM/jCQdKwSjazy2E1Q/MBjgxL/COWigl85OcgUKVPG1rvapn0M6gc9H54jfFxEJo6wL72j
se1OZLtNKYVP4QhWWUVdrAK7DsqdCtvWgbeg3OR0OvDqTMSEwoS0v2NLPErYCOtr6Q4ZGYIXyPsr
1+Hjz/LH4SwwSQUREisqvnx9UzyUDTvIvzIYp7O3TTrz+UN/a1XDo1B/tjwpvCpbsu3veN4/wzk1
EJXn09JmqG7dXzJ8bO+/vqTa4F2B+0TbF1J1Jp03ji40GAK4tf407F7kW9irCTTjpduxWUKwVnY4
95M3nZVNBFWfdKqO88nClP3j464TYcK72VwPDiNLkooJL6cpdsmID2gelgc3DEAu9uBuBLwYYVoO
6LMJhL8sP2T/hNpGdNzdgx68vXt7NjK76Dn3JxMxj+H358FHZr6NzJ6vltwr1HrBJPy2ETknp0dE
kTW+1DYJ+Fw2KDl+9UwrRxZYQGOL0uhTiZzu5pIElQ+UO5Hbui8FmYGEfIsauTKEygC6Y/ERJx0V
mhv5QQ/Pwe8DaX/agfUOAP+lmsEe+9sMiXX2Kljs8iQMKaAQFq4tbkbKmf2xaCGFbCYOfQA6i6gc
+wbVX/eID5hO4H9XuV26xItIYfb1kQKYWfGzhlAVosEcTCjjnlhE5PiH+hLH0g4ApnKqnmY0PCk4
LHDrnyuv8oLDSDMdRjD/wEZEG59NXQrTkJtdKVgDbDxi5FigvIEWsnaJ7LEe08x/g2XOWOfGq6f8
OF3bPHArYZPDhuNf1QIWYQhjHTxKtRyy+EgRsm6US1StVw9SrI2Gedzc2LqAjmMsej1bbSYJprMN
I5OUuvptD8cvAOljhVtR6UEyJvdz0RyDJXaP0b0JhMWosecGQ/WUxYKN6yO7AQAcsVjQmjpNDxLe
oYCNADiw1pFHCMa/d1+m3Z7RF0Qdnsavp+dcU7E8k95lki1tRU+mkNEoITPbU2yNtsum3On0A+/7
BUWZJPnpgYyE4lHafP5pLZB5bBQ1K0zYMmMr3AbQFfsFlaNtLtgU+jWyF6D+mrkg/yqao96zLNx9
RcaZhla6pyVNGetP7pSMASDXwd8vZKfMNZBptbzdxN9J1QaJnnP6ak9j3L0EKlY4GbPTb6YqCp8a
UZRL8+GSpk6MJl6Tl4LsfNq/XPdpmzTDchzmYxL5b7wfjXGWm9Kw+sAJNNO6LQk+WcJic596cC/7
n8xyhZ8OCS2s4sDM6RkA9lFx2IjdD19/fp5+7EAs6FgHQGrrwQi1vty90CC948G/kyTYPA9zCtoC
g9WFYWYF86oSkyN7cS57RmOyP1Jq4fOGfgglOAMdOPyaBxL/t8lEZpttCo9JJWRcO5Btw862xRy9
SuvadXlMNLrAYBCUEDAgi901roqDrBtcvwkkMrBw1He0UKxD9mEdn6HhGwi4r/7pfiK10DdEQ0/I
3AvMr44VJAmmxcK1b03YcKjDknfJt1dd/Hy4ZhGP40SELAweaA5lxcOKPLeanH19i4IIbAT4vljG
at9Ohpk4p+Ib7GbBt5H7oa3o4BlFdPD6nndIE3SWyEvxDJsq8Vl9rgCQdfDc/uOl/6xdhHXxBldl
pTVV5UjPX5BVuVzuXuQ6lKJUOtrUtTHGcBywvhyx1rSPziT3p5qxMb+HahogGHFThykq1O3rz2wP
2sVwtt3zDhq9RsfkQ6MaXmdgmC+qz/S64rExylnjDVe+v9l4MUeqA4E/nidnmObR8T22PWcARFLC
kIYLx9LrLf4W2iFUupdXAhAqYYQwWhL+B/zAcDATD1awBy+l1NqoSzLONa1pC6xbFtpjTQfPLBu6
L79KWNAvdQ4BaxV6GA3dQWIouqsE94JPfeufTI5R6743DK1Igxfe0GlWYavGgUOQGDVEoOjdwVG0
BRr5xChgjPAczytLh5jEiBOKtnQABktNL9eEy5u9MM6tBXbmLKWriA8JD8ddgruGeUY4GzQ400Nc
S9czV4OgD5Gipl6rEGYQY1cWLnNGNqB6l1311bBmuorn6Vmgy3i+hJFE411wh4WvLjr1oW3hyf1W
9e+DyusSK9bcwBrb99K+I1vS2iqwD3aQVCGujTnAgUhECvXqklZ1V5XlmJvuT2BrnSfND7Y8qArG
+ybMbN1GA4UdvILnvAlE17oHQkygcMxVbW6gZhxTi5keZsuo4jRTySy4XPI+erbERqYfzIoV0enX
OW1wPVbifbK31Xfbd0f6Q7isPf1IjsWFVhTcDtLr0lJ/23tUlrUiGwdCdFrz4BSeb3tfRLOf8gyN
RTJq/r3JdsbzAIRO8LVsQNifMQSqk4jIENuiSo9DipRVE/8cqz7g2jabMu45g4YLTJhCKunOx46D
CQJSyWBApobW8ac0X7ah7pDvV+OJLaauor1KwyS6JnLpI2UUyZ0KJ3uFMIKKAKMMQ7OgBRaZOfnY
SX2A/nVeeCbHKZFfeM+f3hWoVdnP5v5Ax8kMlrT8IPn43g9D1HI1IVygcL/iHNmMpyhlEHkkqq78
bXzZsf1bnnCTPQiG4gB+UWmp1nMi6L/KQvl49klcLn/Apxx/fLP5Y9rw3uVwbAuvXadrSPEH8HxO
WfUeow4IFpfeB4SGiV0GX3X4Emz7rfqkMJJXJIWUlBPwXqg5hZL7JvD5E4j1SInZnEcyWE+L1zrC
5YrxcOJzghJO6fuVwN5x1rvzbHqPHP1/I9/VQ/biRfp0pwakGn6Xu4WJVYIVexlVWXmIRsz0HkyG
9y371EPQRWjyq0JCU4++HYchg08wDeHUD14NKoXOCLr0bMWSHeWZG/i2l9ktdedwAkZ19kwR14D6
vBFDEi6OILExWrVo3cI790J/3DNFR2yd285PVNHBFpySM/W4ReP/uq0oN0ZXgjxkqzDWzwl5fs4W
6t6S5skTYkV0vQxO1Pw6mre146tQ6doiFfIW2zwiJI5rnOxdZTOTRU0zjVfgujsS2QXxF+7VS/0l
kJwKyyR1Q2copQ4bt7IJiAXZq4Ii2kLuZzj/IEi+3QUqgrJkAM7KVakCTWZ7ucuN33jYkwZBq57g
TMNY8eU8x+cbQU9XufRkixoMKMmH644yHoUwxrbxopB2SmRXON0jboy0YThs7CTe3+5WewJehnzT
G5kYOxKrc749VDbGuqliyFtTIDMCBwVjBiY13pyh/Q/2TbMSSbidyEre368EvWXUmxaQuZekWqvL
Czw+xNCMR0TF90uHRAYFBoyt0VVuBoXB15oPxR+OOUe1at8Uab3QzgN2AqOH5VrIKRmVsZdqvXYA
ZCFEuXTfmJSA8MzJkt7YyJ3B0vAqleQgnzBz+W0vkKphhsxjnILhPk/12QHWXp32or0ttxmnEHI6
qVEGwgbNf2DeRp+9oF3wHK3/PkLOT1St0zg5nZAsJz65Q+Rt7FRMu0Th9zsfMNpb2PLil1mCPlAH
/pEyGUvhmiEJ7LyIGqoRv7I3YmxmjIIigJ25er90Mkh+lfm6x5LQ0EWJo513MRY2GG8Tzljsna5m
JjexaUGh9+C5nbOhi85l2mPYoRw1EOs4szBR7F0UvcIuRw/4lP7077+Sg8+PUDkgCLN8TCKPQZPp
k8wt1Fj2JQE+B9fyRjRRQmf7AroTVvHG8gd1U26M8sN9bQD0VUmON0pY5AWGTvG0uoz72RtcnKHg
Bw4r7fR9RASlrIAdXB0008XoO4s5hx4VlxlB8hcobk5d9WUkCGCn/EeoHIBONeBkBiaeg7bgg8uE
9xQ3rCBi1upJgZy6u+0e+bY4lZv2yBChh/WNRlCVtnatKT61+zmddHM5ZzvV1RPpM997KerxbC6n
iar4QHBTGW4rFiqxoRyVxU41EzOyCn9lKpslI4p855XiPidKtYXUW9YfK4qUaj13EJbD3h2n/R75
rGAZb1S/4y1AufCPRqpMMS+PnfGObbhPr8NYu+KUSu5ODsufqTyJzKHLCFIOdqGca0+FaAKRrJir
ztSxqnt0ehi+Wi4meAcDfBpc9RVahWtjW+1VzLgVwp5QOFApWQxQjR47ZXtNN91YP7vTWabpw/2D
J3QuK74J6q8i7FqL8oyzXhsoS3UYkCj9Rmw3V/JVrmxdTf7o/LefYt4ReSpCnQXOP+zHYFbkEHi+
nMTmdJ8VabfLBy4otJfCbBsWP+Hk42RBailnoGz0Ivay22DLRfsGfJI653WCV9HOsevQxjGD6Zha
Dd/JSEfOWe1TbVojXgUHy6X75LZ3ILWVuzyT3YSFE17C5HN/+FI+TPT/JKRXuha8hPTbdEKzz5Wu
xwSthk6dm7j6ntbZSqFTLqNw19LxB0n8YJru6+nE+ovLsGduuznj9h6/bxRc9todx3uvIe2cEwUX
IDrjys/dL+WNHkdWq2amhvxEeOA118FJb5Fe+5t4ceNAXtz7SqVKtubZBRTVPQK6NjPy9aoMb831
MUJmjqOGZFYS0seGMWMD4XJ1bNIeMPhRUYAax4jVgy6PVoVnRD94tuTecJpRMV1DcGYT6fPoDTdz
34hczXsMW4KSAy/2RCKlPaCssuG8qMgou+HbXMDWMNTra14M1YBKkK6sZuTRtYJ1d11I4OsQxRy5
SyrCFIwQ3yev4rfM7ZkyE5rbcK9zxjzD3xFKemzpg/PhNQmzGB4b/vgDbQ7zvMd+c0p26KXv2CzU
n5pXuC/nFdAY20J78jLbPTQzGWl4IeaL0/ONHPjvaSOYcakNgnqvxWUtKYy+V2EoPCHizsIDqMS+
gzpJFL/BE1YKrei7DXArk5kjIi5BWnvI5873TBarWN3TpppkcswsCnGGbrzaMdlDFUOHVRp9VCXk
uO9p59C/0AWQ7GxJorWksS5PvvhXpICeZMiMdjDMR5G+2YXx6ppVaivqH4hMwkRfjX7hU0Zus9R9
LNvUEIPynBfLrs5cddSY+Obx8uK95wCKACNDVvpiGOKMbpjJ6GOfzKkVQ/Rzc5zKgfH1rNYfkG+1
urCXg/w3rk0idCbg9XGjWRrSftfpGE40O84qBFZ/HIk5ZkUD2RmQ+kq2qUURroFnPEMAUDs+JNqs
P5A1CrgJljRCN3mJa/DX5hvAjWFDzRB5kTqdWHHfPyBl9Vc9Ukekk0e1TRUPlC9wFkuVpJCVCVXH
VCmKfyu171GNATAOpA9sDtE3pB9oh3hT6wKaPG6N0BgKs5P9ZIPcrs1za/X7kZoNjtzACUP1ZL4y
VxGkN1175F+3H5uQBJiqQbr9ipP6Ammny0x2s/vG2vzZomauO2xxZv2iShLBD70DwL8tdd2/n5bi
toQV2Dmv2ncB69WVsIZ8zkdykXwVg3AyFvqKltJfsdPTnInvucaSsxpKDcGanIRlv9L6ti2xjnz6
W29czmdV250ivSO8R2ax4p2kaum/67X0JVVFFWwN2lhIOl7cSku71cgsNTaQpAmVbP6mDSApzmWX
9b68jQVRvoVnwnvFTQorGEvqFjUXAbnlqySrSwK4LQo5Xdlaner9QxIeZsepdp9pTbFcRmABfVtC
yAxTimjqoocLz1v/GP56Y+ErIoPQbc29d+vWFFWqaPbobqOvZThJ4V8wJKSotCoo6O51VZxlW5mt
rKV0Q96dNfy2G3qbTRLrOOnFdiyBafMcFQJYdDIZpZOU0vvJaoV957o0Y2fyizM3fLrvp1IkL8RB
0ni/kvg7kv97/CO0oVYVy7oo1Kc5eaMAjZ5Wi8cSKCu1xSMCQoCYY+NDVo4/kZ//2RWit4BqbLur
L6svU/iNd0trFy1xN+qio4xeYcHhq3ezl0diYGfbj87k2c63kvQHnG3n/Cqf0w5jIr+2BdS2kM/d
G5wOrZ9Xi+ZqaeWa2iv3ziPhQpGQvgdT6ofz1V+VMqz0iVciCftI8HnuOarU89LIot6uOHGIt1Bo
7QjTnSxRfNZZsKihPRwtHMhPYJgt3qmW3R2TbktsvAryfr9KigmHShJzknwcmFRlhQNiCgwgjqgr
1ZfNn4oG+YBwaiE2VXXxjfrQovSl50IfFWjwK3BN++VChUgcOS1+p6aceDEFe15sJTV90WtmIGlf
vXXoksq3z5SSQtZQhTm2aq9izun+jsVqMAF2TqkAvEwU8ROMFXKgdcNxeAoHgqdggZcFTh2LaECl
hNaOVzMynCkK6ecg7HpvEsUx9KJ/TR27uNX8rJxv/LLlRtHnyrWUuoUfdFCc/491PWosS9y1GhUN
TLaP9yy+YEQJXku6RqVQNGhB7aD5nJAkS2tk3UAtQjwJXer76GcLuCIf+QRpZsATknNP7zmmtE7y
opKFipve7/PxqEg2SWH7UTF3JF9lrc/ByJL9/4sahI1kfOW9fojm+5lWkQ+6tyE7bxM5lu4hDbMS
VRGkdUIkV/SWfwmSYG2X6yxIMBPmDllwdOJxftbYH8Fs1Q8X16GuJOATJ92w2IOsCAj/eqAEO1/9
1H0gjtOnCGuhS864rjTB/P9k6zvCHMB7Z+Q0z3RE+rBt1QA+J9tlOR8ldZq7dlq/jIB8+X0zVk7c
hUfcdePjVfcGJssAI0/WWzLAXpVUxV8siLZ3UP+6cf7CJgGdm81gIGc0N0GgiE6x9DMqykutbuMi
oppMGGrdD1eVBI55pWwtoa5Ro4ZZolTwFNn3lUre12K3NmJby5NrNhE6lY05g3RODDT5ttXjpVft
pZnAp0623bH2dLMDcbL9epWw2Dn+d64GU83yj/btWO4L+oq/oF0842Pjt5MqMt+Jo6HhhSLpCGhR
d8J/OdLMWHniFtkzBTpdmDM096ngdAkkQJZQQ8ztS9u4Wn1NZG2D6jnNmuVKNwBNkIHkr+eOwtHG
GaIMJ2qDc/23mczyYA60GAdV7SbFKH4KQjdOh5pdAaZS7LFvDh+kg2OY1y+AWPZXGgthN8y4RsDx
oPPtGEBGRKbPAKYEOks9OHrtYFONi973VTC5aa4c4dF0EcXtlNba0d1MIBr+Pe/7BRKg1MWA7QdU
29hgyUI6N+IPlHKZZ8iScfJLpDRqWFNp5EuJB5P6xvKegkAP+H60HQa65EW9bF2CU298yjF10YqQ
EEnc/KBb6tG5fUVbVpg8nRYuxWc3E47kP/ojcrYcSLwYpovPUtPJNQkjIB5F6BSXglpEShSCPIvl
x0ENzS4TdnPBig9sV7NEUyus49YuKe1qoAYm4OSZtbDUKWS2bQLFYDNh5SGyLd5TGFy2eaKcJj04
HsrhSo9A2hjHhIiXCtJmvL1G6gB+UdaCGoOjQ8bGSRj8GQEi1P0bovvULl4d6PnT0Cq/2Ug4J3tx
6N7FWRCOgaawa98mmOuympgZJ4ZWzTDmzwSnTRvpUcqzyAK9bOZ/zsrli8bEXgcddlknWEVZKGF8
YJOPXk1M9pd3/INERCglCq1jA2Bs3TMchB841Ra5oI/c6xK6c4pbawPHEL5yaKbmrORJLt62aiQv
0UNuGutGKp+5b2xUbhDegg/v2C9CwpLvZXrYJXODcgahWOFlLnma7vC3F4koL21fTlQBaner9WwZ
BQxErbIGXMl4YbHlgkWbqsniktD3kKyRWbHJSmyeqicxolMlu2yP0uu7LgWsb4a9go2P+fpJksEM
u9RpJCwf9/rvU9L9BM32VypB5Q0VyGA4oZrFn6UcVU3eVAvQcSs5qabWbxweDCyf7ci9lccqIAn8
LErSel50t2TAvHAshvoPRt/cAFUxnULm40QPONSCmOsVu90w8LgBl4L+qUBNMcVtNnhvXcOt28HU
dE8OkaWMWavvbzjT74gTzTFcnB9q6xvKvJvoB72l5pBKyBB51Etoa81vAqNO3l4vpTVZfCzfnztx
1RhVa9daZLeyexeD4gniBL6JUORc6MCbgQK0qyv2FI5YSUOwAG2fP/btWA/a+f+RxAjlQ6w9/uHL
2yaP7dtKWTaszyyTGwXPDZD6y1qlLEz4bv3sf3rIc/oaT6UdBTB3LmiQCoo1azJQ21uiadZThmaF
Q4boQmYKMXccXb9q3S0gCy8O9apV/L7G9fMVGD4uczH1Ch7ELXFs/5W0US+nBEpmPMrLSlNC2qZg
Q6l7iDQKpQDNjrKExHeVDdDs8IJgA5J509Vm148PRY33MvioC8T3/mUmYUQmcuNoFfZ2bNXQZAJy
XlbVyeGnGVcSH7+SDKJ/cWs5YH0PsdP/vlK6fj2MtJDk+b9M7cfmSwUIdMtrfLC7i1Yzgh9qccVr
xp5Ed+J7zUdQr30V8NhnjPrX/YyVoNvhRrF4XVoN8kcOr74iWRBw1xECfaFY6UAE8aiEXhnAXb2f
qfI13m0CtdQv0EbpIFj7pE0Ori3rJDFFnubKo6mE/fqNY/dtttHJRheKB7IJ8JuN8jeVLAXNzIUK
JdQ6/bNCH3krayF38VL44PdgYJoEKKEJnuSLL4bsHCqY5V3m+mtKexcD52ua/+LU+lncaj0RB6is
1ov9lWxXVjc3TJFYDUQF5mMZlDB+YAlw/E3QIZ81BepfesObbCuvaQIKjboZ3BORj3698ldsDuNB
HFNrn6Ww7yhNjNBiPI5hpeNwUFfFal1Zrw2ZQkBkhNH55U/3OLLSslyayTyiDwclIMXajB95UGss
rvptQAwdxwsOLHcqzgtTzWgC259mgd1RrDLmtGAGpCjxyHwCICXcN0ujmpHCDV7qGPMegmENhFQ2
HlFBA5ECS20YrKB8FMIvLekwqg9EBpsAPTyByJnQe321wnjLKw63h2zE7mT1cRvkme1okZ9cggYR
x9l+V02HqmZrvahovYcoeAdNPx6UoWEv2jNVtQIQx84qd0bEGI1shiQERAOVoPCydxtWSt5iRKDP
69+Zidbk7Zccxoaxp8xd3eIwIPQt3t1oTvaX9nlze9KKDr2iiGA9uc7Vbbdyj89f8wgMTiFlCo3j
87J1LuLmtLpQicEYNLzAXd9QzXpIfMvBFmQzZhKiOjYGiDHhQ0J8PWxlAvVN3IaIX0fjameqOCHe
5d/hVRtlKVYgDeAA96NMrgcVkgHKEjMB8xpxIOvTk1Qwl3zMhaD8w2vvVo1zTjvjmZLZ0Svt8B8S
RVWzC4nbIYhlVOhaGi5Cihck5np+ltf+VjM1wWZ/ILQRXvlSPtZz6zO/T//BKGwb7Z7mO0X1xHIr
69wq/9AqvUSCI/L7tm/Ckep1kHWT/7tK0SswzHFyYdy0DJb1jumjGA+koBVB/uKIESYFgLjA2UcO
tCCrrv7nzNzxMEPPaY7WAlkHw92M7qDTo+v6UE4ZTOCz1fjVXpQE4gH0H6oaMrs+0t9KJcLpoL8z
FDpD5wiRNC3KZ5HbeV3YruJh2VSZ7tITbYAV4/wlaycpVwRjERIDK9B9xi1vx5P9Ukpxb4LXYK1T
u9HmZFqOaV1BfUOiqBYAphglboFwclrw5PQzrP+FmbkvdU7k/0ZXaSa/wRatmUzwBv5lhzOwoFu6
Ej5EjfxckVRl3U2WqUPn998ULdEo3NZG3vnqzhM8L7jKkZpXd2BCUkWbBZnZ9uKxKdko3yYPVLNf
tSQtkczySrAx4aJJz+ESj48JS9ESfT2/4mN2obFJG3jq0LK/JkgjyINwDPVNoTX6t8AoZO0+RMCl
ZHqHiq4KZLjZQBcQlx5Wr9z1qVotmUSaQlmfq+B9dypHHv0nsb8g+m98ItScu9qXWcHHgnHEcZnv
dde5aHrU/qiiKPBHzjK77J+ejasKB+ZpTVTVjXzty9j1USGm/TNC5TKpnH5RDiVBpSw5n+oN6mfa
mbfkpFL5QIp88w3G1fgW1VPQsLqHGqRg6TL9aDae6DuWFcHRO8ShQjjiZsLMUdqTfnCSw3uQiKnv
x3bE438e4GH6b/xjntQ6esgc04IT2SnoTW60boOG4E/gr8TKXA0TPc/ZFo0h2RUfrPFnzOR+GKgE
nJz1bc60WKvWZuG5DRLtWOIoaaW0i1w66I066MuHWpH4e1+FqVdQhWRNUKGqmsW5ccDw1G/uh2BZ
0EoWCUN5KGviz/oa3Jm97gpSjjtF6tCkOUabacZytAdJPmttqci/SoW+a9ZUElwcAdy9zm7ezxKr
1U/UxUYTpDOxkMss0kNYdTKDluR9ZKtfpSE9QkCtAAL8BXxmkpoIk+vybeQR3YEgpGydksRXuEkf
UdaOMIIRIMoieH1/qfGScG3tgaVq4anuXQ8fYYTKu5c0Anhrq56sWelTiSjDKcuHkta2jTiVCCsy
i+SoqtLd05+z4VjqpGkvEzMC2UUa9iOrxIqSuoae639W7Z83SZJP+6cgL/SDNcjZlB2qk7eb8r2O
yqDfD3a1zbQEhf+up1YrFC0Ukza0u0Y2xmI0znb/dFtSjnaJ5a7go8mcVdZ2Zj6Cg8toVLZ2gqHL
8e2wg/gPMuRCo7YYSIujTxIlgpZkRKJaUM9KV29oPyMM8wSCGNDJkI9QVN21Uc77L8tdkeEn0smt
JSDCsQaT3MSxOl8o+N9TE6nOZ5Y0OaZ74/5uRDvzqZU0oHO8AiqrjijCQFZmNXj1nctwAdfV/dXn
nOGBqifwPNzIT+1o/Td0Nrg3q9RmQB4ucOKaHBvUyVEZ2tkLbz2hzDOrlYVNMThedjaWjCRPOeZL
2TgKfORJoTxBtJiPwrgM6G8zh1m8yA1U69VanS6azu+70coFKcFMe7duH4FfrDeSbk27ZxIxXMQ8
Nj/03AZTGYUcpY/Zod2DwZTpwOQrTrynCCxtoht2lQy2buo+aN0YN2xjWH3veA2Hlbmh304d6Map
20mzMzlE4y+d9c6BxVLplsd61AcuArPYxStBXcKEeSI7jNmth3yJc/5r1P2PcvRRbtEtwN9WAdGx
QoPIBplkgQpDV1Yxm6RRhaOxJ7lCO5IQ1tY0gogyD4S3zCaBHcVojrG4aDy/3UXUk6ZnLpcgPy4L
Fa2K4ANMo4zb64aYAyt6rP8WV35TKQZtY32lCW2X0FGhdjpGRiiZmCaG+Zpx/c9Hzy+eRJV92H0/
xojs0PSmTE750s63V7tWU7iaX+Pps+v8to7AUzwEeg+g0vIJ6X2K2vT2+tKqM8jrV+OQVz7ieZ0f
8KUI9cLI1DhyYHK49q/dgAlHzNZM1NIr0Jy3/oomY+DaHb1wpScFMEZ1ZUNwt7cY6Fv0kqGGKdOm
pJOp5HCoS+JXpSqDnzgPoxHjnCWDEoL4hs/RfCze6dHJ80h0WOqzb3RcITnA0eYly4w2VQwDS141
tt72ixvg/4/FXui3WLIKCmREpx/omeIOHIxWTG83KaJp1/QH8UGDYDCCCrecY9znCNzYTsi2x8xX
FUUs+8OZwJnnE9Hte4WL/g1/ndU7+TT6u2GSau+KbJWE2MC5h7Nq80+CnpaMjfHhsCm77aU6CFpR
4bIoN70M06vE5xahCHcbvMvKObQIKgXhQrDXFF8245CDNmRLpXB4+EXWjmE8635nInbGxdtvwga9
aU7MYddl1RhLl6fzjkCEwaQfqQOhsR7Me8q80PSM8RHyeMwbriAJkE0CDiIkiXnCDzFPw1H4RxDB
B2+k4lPyRgG0dc8IvpjtZZzDpauqcYpBGPk9AIXQDz+4xFTJRgLMN2rKQ8TjO1n30l5Q78cOL2ra
RnFnfuvALN21VD7hlKmE0at8S0LHx+Lp2RVgbsxv0Mi4QQixyFqfOXfKsTOy4YDAffdDgxMkjjoJ
85hlggRPf8hqV7/KYc3vxz33gKUmfbSTTalqDxqG8L8jDqlsr3rZOSrRy8I/CyHcTb5Mly/rEYke
ZP+9/NpKGktJGxYX7KqFgqRMKz2E1F4Um2sCTXTET9BFxqOemv3ta9AEckkGH2Y1Z4vfcB6v3+8p
5v5Ah9nxIBUYibM95YbHQMi3qkdImTBhxCkdIndzaTZiF/0Dimv2EVu7MGPkbb5SGRp1Fl50aEFG
pjkSB0g7+0l1opNS9RZW03O75P2k+ldeQQ4rpV4p5Fq0F8mtHsDaDfpnBgKFnXXgustNKBUZMGFu
MgyeTgKsdohnteK0F5NhDN81O+XpzP8/MZd9DYquC9RvOfDpGZ9fxn8gBk7wItnF6kT6sS0XUINx
IfW7DtLg9+1hBPWoKMTNUb88xgbROVT269N2yb2d8Ty4My0dDUmm7ty+4b/9hMtLsWLuwAG1xA+F
vJoibCfpOptAA1frZkVErlLX66G7yrr4HZ6Mu7smalwgyZIkasXFGlQjA3T/MfsaeYOLY/cWc7hZ
5GflxtWTm5BgfdIa51NMM9zort8GNSUpPIrDtjjf/9A5gh8uK6xvxyPuFE9JiBttbddhQ1q1xgKm
TMAQ1UwbMQnlwAwVVUZsrwXSZ+oTOg/aXBwp69LXukMwZdeCg1sUdMyAQ8gHDh/4DlvXJQLJbasX
EJDuM4j0jf7TTUb5QP+RIT4TEbfy8i+I7hi4U7YGXuTjCA8BMiIJJ5fmRKjPRwZxF8DRTCkfgTpF
BTkOxCQ2Yh0I1ZGPX9oFFFLcNgLAAxWL+/Ue9EE4KFi0EifFguf+HX7nkx+Cc4i6qMWwwnObR8go
iYuaUdx1udHMVvg6Kb1fgIHYddlhTgVkPvcsDXtOymXzMtLv4/nfIcFL45Lx2c0K80Nb9HbeaJPq
hkWBj54+TCJ5QcVZt68vMdMlGZsFdssaSlI82klZsLTAj8gd63Hu4n4ZL/VIelFULuK1PCKNcV2H
ULlyhmSPG2Q/mfANujr8mRX3HKGDKR8/4cdHbXgrrqVpj26Eg8CUSFshHAbh/vUr6sbbwpnss4Kn
CUrOQuTSS/DJj5x0dunyfGjzT+JDERyxjyw8qn7WvuBj6UikSHYExMH/tK7kg2VLRNqqMQJ+QGqB
oH6MB49YJtYdFwdWYOXK3oGUeB6FnBJrEWeXhfcZ/2O50FLeYR9lwH/FYM16mg0eOrD7+ij3Zway
iLL4SGIQ3i5TQzBaqgTnlscdfN/QcOwXEOyBLjPhKYlbDMGY5rE1cD00Acx0kNgc+8QYyjcoWVki
MsIobzejLqQyA/wt6mG7AKc3FhQ0IQMZTtqTJmxO8bLiW7VFx6lMLahS4ScZikEOop24oFXWSPYI
qI+R7L/0Fp1bliDZupNjEbea6O7ehoLFH0t8sFEuhqYwQ8NI55LpBxuDb6nvSXj1nRYYzfSmhMBf
IUfmHc8rjfhoQAWu0HzXxoYe2Pgz1Exl9sTpAKMJk4PYNAzccfXhTnek/EgZyC380jl4EEeZED8y
yfhdq35v2wGSwGd2Ao1e0DvvUsaciNw4RbI2oYpd/BnbTGQ6/mN3ww+veBGGFC09LYs02m8zHB+f
AwCbenS58avnAQ3mgSacQwvLvlInA3PYkkGWvmbMbHDPEIjc7rKY3ADr++iPukiqq3LuLXpZvEaF
Btha74c00EXBi1RxqRMUUfwd5lvm0DQmkxPyNMJN8oMgkuE7ADfPY6YttlfBAVKcNLCi4xkqbgSz
wQt8hMrIW/L8+CUdrqkM+3Wq8kycnm2CE3ZlpBi+jk4953mQXh+Ay+oqM5C64V4o3KkQiTps7Hrp
9ZXsx3NLlsrRWIB4QhhnxhyLCxXjMZFKjdanhS1kYqbeyMsvfPVs6P0R6wUsxh9K04YF+zZLl67z
s91/8YadBEbjNsDGZZF9QJNGPJqFrH/ByK05yGNJGKax6tXxBH5tt0dJlHVsU/JiMGqAshgLY6kS
YXunMUjAGDAgR5Ile49VG94cYxdWLAfbWRfWACKqoXDYvSeSsuxZ3ZsdjDqZ2NeUsNRvrKGj0Nuj
A0kCfmLmz6gjiOApqik/l95IeryVtvcAkuRjTWZ3cIYep+/+n78v/xa7+ToLhe1aVpjpZ26JpBVA
NHr3dQQBr4mI3tz6ci+SdhvnBO9rUPKw+HO7jWFIPg8kjvXgfVJZ/WOMr53gMFiNMF0W6yyfnAlG
RezAIX9tHHnoSRmGp0IU7pqLE5Lp8U8S7Oa5OTxgAFiWUHbKtYnNwJpKpDg6Yt/5mNM8u2nDbz2v
VyxqpcxHnxUnFZBys2WHob+kgZUORACFhksNpUVe98NulMb1B3aGh9OfgZBEjsV8CTDAhqPPNjtA
VsdYPnlb579rI9ITzxQQ3K7+tt8lFiUe4viSMH/AZeJuS2CGprq3zEZpV7WulTaEfdE0pAnTE2MH
5QuedwzJIGi9UEQiK5Pm8RXqgmUq9DuMor5JVT9D+NVpQeYYucLGt3naZmmaUu7aTx6Pz/n8KfG0
4PXEV7PsjyJ3Xs+32o1yQlvUB1RdSFjqaIDWGzmAUCZRQhm+m/+Qt8OCWMBD8lkr9LTMWEXgEBM4
IAT4wIEvuYs4+Vj23D5puwnkIEJ3NcKKf3fdTfwqiS4xMLbbtJ2AK5+gTjiLfEoM1Dwd0Lc4xqxs
zjEkChqo++DQlToGjYOmRhYe8rPO+bq81NmvgfSmIILiv5qmYfx2oa/0y8a7zY43Uo3XsIxbB/MS
L4F8QeNevOs0097M1whoJLbRTp7/QlFkADYfprTUH/eNiYzGH8n182mZU/HTkpV65LkPkDWxvWUX
iUCMRjaoyPx+CHPNe/XCnHpHfRXl/yhEsdJN4+2twwpUhadaLhRagSPxinNU4IEjP2mkQKb7yJSa
6C4Eaua16F6ZVFFVkgmBxRCLLVNRbqwDh1DNK+c63a3W3SrKXdRxYoW4FI//kW+WUFFBtVrW9W1W
IN/zFf2ELWiO3mJBS4lpdsI/uBZqhSKbtroTRbTb+JUcz9AwVJC0kQF9N7UqZw5fzLHEuZeZD/6I
3Qp3r8XM3WZ0cCz7WT7d/Op9SuKlMMx2R0HosZq5sNU5XHurKCDDrkD1PZaybrAI0HMyX3JRC1Kg
VBAB8gK/8uA1Kou9YUZsfKB9LPZ8XGQppmCPNxGaAMGQGuW91jNbM9iA1QzhF3n3Cg3zOoS07z0K
OYFUIckvYva7NjlERmID5oABdpHtS0k3YufoKC4oxT5/nQDfAPlc/iv61EZfqaeLWwJuP82XMVQl
kTKdHDQUilcblOaGwpVo/HBHKBbOuY7N+bJZZbEyv3X80MF0xvnqh/k+r4EUTk3Zqg7egE27z9yA
03e1dbaenIchAAKdKFsyxjRFQ9wRLZwYW8mRXpU1XNPqPpKqmuG0kl08SX7uGwl2LbsbuheHHF5C
rlGRIenPmZKFt616JGOesk8w9S1qWHznkmlqiJTe+LPZBg5IPk68YDd3RLmOGTN0BR5BXIWmgXFS
GxjG30lazv+FEuKmL4sR4LNhf+J6Wv1Mizq/CigwbZ+gwAfjcKDkUy4yfVZAjhWVeb610iEvWOwb
sUVMci0UWS72aW5cRjIvLUSS/+ithCIutSMOCg1iWtDqqKACsXdcVHnlWX/FSkPvLeJDhIpVzLSf
IBurPnDsVAbUa+fv/2MvDDZ+8m/OtNcQ/Gd66s0kU0hT3JyGPwi0f4fBQNJznm5rcusbidVEoK9t
VYLrZbZiUzyxHkcLp4uX3FmhlvnI2UTY7WM+wm69fs9oQg+Zmeavb7EZyXwmtno8wFczOiyT1e1P
bqyS7lL+TRzp/az4zidC3ibilsUBFBxCOPe2m47wOkuP54pswb+a5l3W3LJL2j3fNsGBBtEtmV2j
H8TCMTCqUk65I/q+Y39pIrX8tMCiDphUs3FbwfGBKpDhdCCgyFdcG379Cx3GtPPFMI3G0j3rnt+s
pZhqXTZcXmyAGUyB4SHU2frch4Ps/poaR18seYmC8Eo2KKRP3nJt8lyxm7HpN2cHK5DFy5Y3wTic
jWVDZOe+faccrdKBrxVs+l5AAK+0oPOsz1PrxyMJbeeSknkQGchPbxM7NQ2vJy2mtrN1MxZOnu7v
Oo9h2w343SwzKN2M1rexV9msAiYgGGhwHPqeLDqx1gfbx6sq0VyDxTLHkIEJ8/LehCrHKbGWQ5ay
F9aP4lcS2M0maeVA+cFr8I5TD8i1+0OYQjOPwtmkjjUlNhf1Z3o70FcT09M9LISU/FiZI3Y4Bhzx
8c0+Tdq7fEITeQqYlULlLaDENEb0A85CrmwQcfaNXDA0/qLM7/koJM14tOok15Hnw1OCQLLylJ0u
qMq35I7J2fVK4o1ppG7A3e4A24AIn7Zu91xwCgnngu4cK59ppGpPxWv8nqpd9/5gcGoBiOMpOT6N
hCrKIVgHizZJ4M42G6QQbi+w9tsJVn3yememh8AoSuKJrUZtDowvr8L8p04+5byzrICfYcbFIiq7
7EL0+sVUusVVs1XTpRx4bIz76PnAJtY49SzyHrXZRxj3bDkfWGCerSQcJy8RrgypS8MBi4NPLTPW
zTUCmnkzczDvV6sWI1AutnyyTzYXezq89PgGL+us0hL8x8kU3nklTUrIbvM00vzomuKXtKvv6MGu
Ghl+QUx+5XkOUPdrTROobM/z4nLx4Mr1kHUckxKTjmjq6ZYeFKNILVqr3wnSXb6Cv4jVz5Abib6L
3MD15zjrmMDL80cyThqQG5/l6cxK3D2M0NI3faxrzt1TqdzNONMwyAqCSA+KEiWF9fd28qK/jszT
VyQh0S6M7x0eB5gSVFJGhf4oskggAAF55YmPdsNpRgS0QywbLSDzJn9FuLgInJG9lnrZhfCCP5k8
bMhrBbrZ7Gr38rzqxR/4N0v8q9/tzl+E4gZNNU1vm4xYLCLT7oQG5CdI2gK7Ol4l4PILh6GKuZ+W
jk/asCbhjJ3Kn+Y0aQlw9dhRBPl3xLE0QpqJUr6AGOwUj3VGGNVbE+wCULyY/AoQxhgnu8zcyhM+
Q8okFke7lGQQMVxTYFvmSUy85zZPk/b89WVUgQU76dltMiql1GCQVkOZE7uBymhOEKO1QJoylvrJ
Ct+5majAuXYzufihvA+2xyADvfE0uo+XjNMmc6GnWcbbBi8uV4YsbzXSzCeK/d6R5c63X5m8zPMz
cndWCa+fp1ZMyvEBcCm9mkCCRYnGz3DgrpyQBLO5S73tUMqcKGK7YR3oNl76z4hyArHqchY8wCdP
VmucMGY286tCccnXT0islAGRJ45tDPR+Xyc8NSiIW28uUlr7Uh1eJJSkv678NXQjG/Ag4z7Ic5r3
A6PR3TQP3N4sC5tQKuucqgkMm9hdSzH9aGtzlZPOoWFLQYT06c8bXSbv3ombJ/tPri6VYn/CiJq+
5nv9v2D3qzAN752h5tbzDh86c7MKcL3/oVD9lyhcrKJAqY6CSizRJxvyGEztMXD3kPI7w9rbzEFc
QBvlhsXh0p3BcujzaD2jBCVZOeQ3e5NKGYovEc9lVOXVbR0LRnh5Mfilre7qWDjqe1TEnpD2EYTm
1YLUBNWOO7VgkaRbLGqtij9KPkErr77XHUZzvGlC4Y98AjL5e13oiKyae9KtBOYWhlIBjH49JzGy
6xB2Xi8C29Z/OnYF31Q5xMxU8JFWn8hPhfJz6qo6EH/NlZvf24sm0xym0Sss3P1CY2D0xqgDE1zE
TnTZPOXDweL4I4CAcv6ofGvA+RSI3EqOb7VLf5pAMNpYVOIjeay0wIK5nGStRpxP3czHn9JwuOmH
T65bBIiTgSbx+vrXPLPiraZg77PTkn+9zPZbzcfhz/5R60mLe4dm6H6/vHQxuuIGesB/UeA6gqRf
xO+IJKqi5cJvuMNZgzf71FP4Snla/klGTNNUlPKAO6Uv52oKt7w3cyUCajUhe09NecjHaSao+/JV
M+eWMsrv9ofzdJ/X4QFw44mEtSZg1VhEa3eVtl5xVwVBCGlRzlfKsVMu7YH17EdDMwUZ37Dv4Kbg
kijKG00MhtnSctrVpVlKeQB9VYscuitHwNhdUKY8EQZEClKuwNCD1CWclTPdAlnLfBu4AekGnqr3
GmR42M2SZBkL78heMB8BOmXlLzK9/Oks4+slRHRLUOV6OnI5jyfQ/0fvkd3OEqhXAGhDkbIzamwM
Fpg8U8ogqEPcov+dTBQVQlhiDhRJp107QM4TNcS15bfwBkWKY5GuVU0NAyD9twrg19Lq4wd1YRJA
GnKewmvc/5btAT5bk7haEufF3L3PD9pCS2fVVHFBOmae3/EG4ZL31FhRfsZvZv2bnp7uKagSnAwM
TCsxdebJnZVfqjDewJ1WlCqyYlHC7uLE9CxaREtRWfxcVLZRa0TqwYy4noEfZlUX4SiUycLi2Sv9
xPnmlZRTWluj7ycPoBVQxf3NCmlZjappBc3LU2UIzUnF4/Hft85dN0j7lPtMy4z1Z6y9C/etQKHx
ffjoQFDg8tm8tmCd6VcFIivK+VlfSq8BwEoITQ99LYXg4Ga6C2dOjr1P4yXI4lAKXe3sOHKa4h+H
tWtPEAx2h+ihAzjQOYOYNz8Zr0PhUiRz34wfZxvcUnG1lWlknnopFJzCyH/1+K1NCReKwiABSHyX
DpAQCMLNx4l70qSdAZ6s/2vn6Oflhrh2wLKzZmqYXKv8yJgylnVh91D33yi53aaKmk0g6kiknTYv
brZcJ32GTbuwnIShEbn1Yudv4RkQwIBLnW3wTRi1WpZPNPhpUAr8WMjk3BaPuI5gy56OeGo5HfnX
627bPMzsCd8ZnxsOiG4XTHr8VjzRAmIQSBaXFaR9DU1vRi8RK9ph1Fkp5nvU2Vv2mp/xAc9l2uja
6bDFlBJvPCbIHdqmCMKhpEtuglCBeCVWrCiGNXcsM4eWFxwORbqpxoxgFh+l6H9Dsu3hcpypmvGN
Te3WvDdtzJeROEgy5EkdeokwBbY1j02YYrv3v8/wJBOUjaEEoG27i5m6C810SLeFilCFQq7HsbDE
2jevA8LqQb8ehb2Ggw6kRJViuWVykcdbkLHP9TOV2r0RU5A+iAPJK7vAOqM+oyA14ysvAiDBkVtq
LDfIg3sCubModUYq7RaZyDv7GX8aTDlfnFSSwDxT67pu/SmqRRsnnJEAh9pVUhLZyQkcWKyNRpbO
DLKTs9tNSQu3qV2hXntdJY6zx+a7d0oo4dVEqHsDvKzfzJTv+vqqsGCgcGMdncVhgWDa2u81eq1T
pIz3pZohNRLJurxmDoX1xuGnySckBn8f1IDc/cuYNjuiftHxb0QLiew+oGKkdPJ5wsB64xxhGPsX
w4O8a/1NMK4RMyJSo+iHCdEiWzKhfRHJT1cY994fzr6YDJHln5QsWEADNBOH/tZJpz0ZKDw/5E4B
4XUgdQ5XfAcaN4d6mKd0/LMJm98wBn/22uClwSQa7SI/oIobIp0/tON/6UrVb5OTIRr5z2Jo/m75
Kd1K+VvZky+mmda0B+vsnRafapLfbzYtPbM1uS3XHpCftAoTqtm12EqYtP9brwjvAJQrAiAeAdYn
l2Ip5OT+mf+BkoM6Rgm/ZVgiuNZCuMd8Gv5c3hJomZxzAcu7bVWYilQkslZBFfVjUavB5kVUllA2
wTgFIumhUTi0nMczoE1p3IJTNZkUjHdFw1/IPw7cljc0Ek7Pxi/zJDn3URPobE75GIL2n4oSN42e
Rf0GCdBlYdvoogjBDBT69PJlSzcsefs/BJ60Iqx0rHmdPMAw3g13wTS3tJ51hNZ/2LXee0pAB0EN
mgw4UB/A1vQ/Xv0WoQpn1TD/R+aZMfSugp3j3ZqtNGjM8s+PLuomAb2m26MA/A5Ryq4yJ6ttV5xs
LKcawMeyR+DPWyzBzoJa4C0c5DQJp0x7cltuuokHMaV1sNAEDfNmUHLec/debHdMJl9IT8GilJ4f
jY05a4tXN4ZjBJzc5B0ESgYwVHdc6IGB5hgtAIHVEnEwgElPqC9cfzuSTDunuussz5zw0UdbOS9G
hVZ2OjLsb8XxlnUYtKyJfkBuj+r3ri6xPsDcWilxgUaFrg1sDW8p1aOWR/GLzV1/VVuQkYVXIHjc
ErDk8LyO/KF/RLycGxoysU6QbMa1j7dhh6JrdrA98+PQvySKmzr2QqdAXex/YfUpkFyLJF0ikymO
bOAfDJHI4xbyXv8Q1qxWcgxDT0Hy1HFkCXTi/jk8iFDjS+XzOfvZfA1QavP32wtvYpHcTBpR39t8
j9XBqM66CIEeZ/jk+amxK52w/Dwe3Ael25ZMd7CpSc+Rr7tSJmVLdu4bOPWvIVqy6kM76I6A4B49
optSubqGAvLYez5MXt0DqlFlNML9P9ULAlkGOIHoYq0EtKuUgOEJD3pttdiAz9iuGd6xOsT3mPU3
Tl7YjxJN87uUoEOxPTKRXvYFzh4AsESYbSeVX+7D3xqBkufwOgNtCOEkr4XBgvyQvJWaLzzHrOPf
F0NPapso5u10dxMD7HnR/Y2mH9jzuJahDrusBTLqPa/Ckde4xM7GJl4SvHwY18niDQmrLOEugZnx
H7gngZcPxiWsWsjqxCwSqaiBPbQlr2ukjWvGA4GGPrEyzC0agrzx8+eX7c596dmAm6xtZASOEdw8
taRPBGhcXSQx9D4JVoR8pEBEEMeT08oqZGaT8SjXy34XAIDLDn480ZjOHEHjwQgWl2CAg3V6ivVF
1bQQuHN5ZBAIlRfvx7yiXRl48pvz5UYCAqJp23UDOKQ5LcnjtVQctot5xco9NIpQNXyjPNSceX1m
BZy+Q2053xWRlV6SM0hLyiLOsjvV6OkEjR5rk1aVyJ6+FhnjXcD4VmobSPzQbw3uVWy/dpH+3i4c
Nf0gyR6/e7BDZV+F0BNElzcHREZ3Mc1V+fhq+Xp4NfgjlqNACSXIq7kYQ3YNz95TsLgCFe79Pv6F
CgJuJqdJqAj08E6XU8weynEBmP2+zbeT9/dKFir88OM3XR1g5V4lz0NG8K26ISaHx1p1B6FB46JW
YQzv05Dpl4og1bxENPug6KjdRoXk4WJ26g/pOv6aO1G4mTOoC6V3FZCXgdSc1m65RG12ZrpzSjXi
AQ2B43oxNKKvsBjTeBVefEa41LqlB393zmxNcvxtQi7o76xRU5ctyqSKYSUNH4q3Q13gt5lvX/bO
QR4+QyLbDAIJ9CsAAiz5RhhBhw+HCBfvr2e6lsjfUcPOmH/KxAT6WTlNbT3GbCvO8HZjp1dW+tjQ
BHBKdgwT+gEp4tyqIRGgvtcnsoeRe2+0SKGH7UueiAEJh1rYaQ5/y5eAn3YOyQ2c+X02kXz7qL/j
hjGWN9IPVP/Zw0ph93mECECO2TgQFyQHKxYwA/AzTbqF+aSGVbrsGvYyQQAI/oXctYadHUhnxbzY
qjvGpDTptVkuPF0K8ZTYClAIuXB3DSgitv9dYQxsoc5Quj1LdxgB6VhTuxOKHVrRtTfFh/azbMLr
WdiCW/qpo6+d5aZ+vBwyoPorEayof5LjLVE6StkG1E6wckQtT8MqTtySE/tnELdXQ9b4DWw/HIYv
z6EfduT0Ty0ttszoNCKWJQyUftlYlMBr1QbXvm8pdnOc9RCGAWN/erIH6EhB5687avHfc8Y3TZvs
QQfieBEnE677qA2ZjLaHwQLvOigN8vId1xeeCOOEuiOcrBgwm/fhu7VdrylAVKfzpOpTJN+FCkQ5
c2LR/CUY+YvKbVG1uLRb+2d/JMz7sDaqQ4muPsAy7h+2cvDGF1XAfYqtppx0XvFFweUuZ8RjnSKN
WzoLHNMGfIGenCegIv5sc22NryiiF6vgII3bwc8ys1kKcMLStELSQAviwU/HOlxZGQAtjfX9tFUm
9s7HeGON3FbCNiTVXx3ah//bSJdQFSE0gCoUblrDorzrNJhNqzBJB5oBXckuoX+sS6CgfaKgmb91
eK20Ta5/y6vaz9jIxaLrJ0Bd3C+/dmCfFh8i+Z6JGzpg0+4guA8yzUwgE4Gapr3+Vi1RrgJmQmQO
Ools5IY32geqLhNz/BokEvnx6xa8vq3vrFkuMESReTKIesRsCK3G8Eeuhc8hRRf/536wm+TmD89Y
mrqq0ZP2YT7Xk8VKBBbLN40TW4KsJh5dL5Ewycmb8b+uwRRZsuLjrPV9eTwQvpe1LNG08pCuD9cI
jUZQhpj9vgs07S8UFQIC67W953EuSdQvTna/ciCWm39lkZhvXIfoqjJVPIc6bK0urHHr4GVD/OSZ
g7uTT+MKsFQwC90GL8xFq8B74zCeIVx1/OTogfBYUSNNNx63LubtbplyOq+57R3i6a5gFDL+zJJx
tJUr2uprU4L/TJ5f276vj1VTZl9YAjEqr+dv4WwVeqqnc7h2OvxYfKsAVpu6Bi2fPUsHQ4W1Ov4n
/PVbA3fSTH0b9TtaczeKGTMTPoZCIVEBlAWtJfeHqAHFZ2E0BWRdssqxgC6xp7R5F58iLTL9ACj0
lXgEN71n8CdElChG5nOXixeksI691NJwWV9aefND5bYRMIUwplcFQGT5BZHOBvAtzU0aA2WhZqrU
GuxkQusJh7ZFLNgupajaKx4Yk5wtVzG7U7xGbVchs1inxT/oAkcNDp2Vu8ixkuF35pNGb2Y8foKR
bd+QuCIHirLl7GUqzdnhCdaUeStcWR3r7I5PiQ2a9L0u5JIFvlLP588u0PUsyRq213dC0N3Mv7pj
T5d+f2Ym+0RbeNEAx2GwpBmBhF61bA9fH+nVWR8NzK7UB11oP15ymT/q571Y02MSDLv1rFSysrZO
HMXMffYTw/zhH4NfQ1LsSnruR5jZutNq7SMrrxDT8jVvtKGHykqWwgrc0xhfqTp7ZhAVZaWfSbEU
HXkfHU2Spz4Tjyl1PEUNIiGUg73/SFkhriFEg8usXVMCIyeMI+D2OomcuL7JSN4XmFb0SaUkhUFz
BtbpSWN00YWCju/YEJHH6SZlSDukrqyofQ6NMH3YpZyvU6XT7k/CRvDIfHpR0xSCUy6/PStUkcKL
Yx2zEPIAtTYU8Lf7TVhyEAhe0VesMJ0AuNK8UEAQZxVgUDDjQl/ashywoVa3J8Fv4JWQxMxEjs4G
HKs6CNmzlXkqvnVYxfXb5RzmFYpdUeuRgsgcngQnFLQZnbOeKieDlm1l+u0jI4GMW1nafdsQlZ9S
BjYfTScS+CpOAGNNLSlPjZWwp+WoagBN71jBP+M+stzsGygwgKz3/qLSLZy9Drbos5OI6fY2Lc52
CzmaQ5L8obaZHTYozTaGbSlB+hbmJcTu7RiTeWtBV/hOKS8tzMXB2OQzbGcV+p96R61jOqqxoxqG
Hmek8/4iauGm/anbqSpatlymsXWrZiWtlReWObvqply/h02Z5sodXyLL/0prajkiy4X2vjWGOs0V
DOms9cR8nY+EaIb+ExCbTO9B8uDUpEWgiMDStfxN7EogP9QTwooSjZsx5rBxRtqgDHoWX5OrjY2c
tjIwjWSWceLf+NOoY2Dgjqy81BVdyG9B9nxLwHWWWpXJgPMWm3p+/ZXuVxkxX5IMuwI8AvAvbNfp
BZ+VaSzxqnENuAeGnzK6eSH/NNV4dDOwEA9Bc7fCrl02muU3KF2bT0KiQhjmn/xa1M8Jl7ERz0Yv
yi9CaWrYRKLA1+T5IkrqKBXvBVRoY22Mpg95v46IyNPnZcZSvSlhrpyXEzu8Ct53Z7kEbbeFHej0
pw7i2qBwN5qyg9LJd7tFXAB/l14q2hR0SC0hp4D8B90VIbeMi3a5j1+KfLMlog3NcCA4btJKn/CY
U/ibMpo6DL1zwFlRlsau7/ai9j8QlcsaqpxtNYdwk+w3Xo1La8Bf/JYyEe/3E74V8WdxU0OZKdhS
y3NEr2FNEM4LCeY2DGIVPmInXflI0zWac1jqahXAjbS6NQS8Q4DJmCdFtLdyUfJ0wh5PKEcbG8Md
h/3cdQlCrZPBkU3BTrKVo3LT+7BjRqfE9UU6e3jJPMnTcpICOYNgrCbJAQpldVh4ZwjDs/B8Qu8+
qHG85VUDt+mCShdHOb3qjaaJsgJTRQnIDHk+mzLCI4L6SYnezVysHbmJFzBrxhBZOt49JwwKC4Ig
bG70m7uIBU5jBkcoieQpQHir5FPLy+Dbw10QUBxlNtxZPoF9R5gZDCL75aY0Wwz2eTurdBSWQRyI
bRuO5CasnC8hIzxJOgcEhlJL2F8XZAJUzEYYLO7NJzlQCQNW/hD4nvPKl5iMtVLgyJGt32On3SiC
xl5GRgj2u7UhH3zvCm9qEPTYnoSHC8dXAM268wlEsYyNzhafIzBaU+gjESIogZaCCSahC/yYkrpU
QQnEgxn8/upD/tQkPT6VKVqYMjlLFsF5J9GGr2AnbNk7S7pyS+Xpu9vyZtOY6nJaa7tOWPdsXscd
DrGcc9fv/G3aolVoRTbG/kaBU75klwvgaKMAe2sLShvLGtuzBoBxsv5G8dULh/nSAPr4gykadvlg
zO5h0AmLnryfbnnKd8asc34W/sD4CqDt8rcY8jXT7ZBDpNmAekS2RXUZgbjgg4bvSiTv1UY+Qaw7
Amq+5gUaHKxswkxWuq8ChczCzRtVcnywwvjLuyA1lBQvEP4Ps/9KUY+b/Ig1pvTaradvBmJnktWo
D4eLOkO4RWc/AXZn4kqUtd+Yx9vnfjOfEZMDuT5Viff+5tA0aPMlW7nxxF1y+nProXHl0ebPq4NO
zXS6TrOOu8tz8c1vOVkSVsCIhj2Uochrd+57ISE0yjTvr6Vu5aiTymdztQqSuu9SGE5lStohRQwC
qNwAVdgbTqm99Gm1zNKRF8E0cQ3Jo+/tVrwzomqck4PxlMI5dIntOHf2yLqmCtSv2/ixFmkIVLk/
9tgseH1dMdaY4N5ni41r5lqypLDGXCqV2qPvjgCIfN9plY6yrFWcpZfWWVU41qy84rD+H3O9sVAH
HuBhCBXN+bVdgC8BNoKKETYh6m9/2tVyybTiNJiRw6gI9+Ww1/2k9QeQz+ZbBnnddr4c8hRmKT9n
5oFYgtZT7mwRKdWDGB60vwS3i+E4OP5tWpfOM2LAyC3+1iFnDVpId0OKmYsnyYPxR0anIwXf3dJl
VGziiCsKjCZjTZwDOF1QxLqi4w6kxCaRNhaeV6m83q0X9BTVMj3L5MMCoPL7fnKqe8zsmBPPXulo
cprgr3QZzg3R9DJ+qMjcay88dO9AEVNXkLuT6ySY90js0bkSh6CC3M4kCax3G9eiK8JsuhtbvdKR
g990u4qQv5d9Fbq7e5vHAmc+DwOggMrzH2CZ5PUHfl4qH9jfWbFiht7s0fjiXyTAOAJBspAxTTeF
YhUn9lppNVxKGV9GBBFl/bQOXsvGxNO9mSbDJMUcIo54uo/IdYkMTwRXl99rYY+vsl08gWcYMx25
NH/NWY7or4LijfTAsGB/ueN9ylC5ybm9WRt0Dg0vnYCJ27la4ov/DN0mQE2kv8dzFIF2hzv4E2IN
yhqBNL8KMF6p/2UVRHB1IApbPYHgd0DjlK5RGWuT2ULuZxvA0ySwCZap/cATSi7iVPE2u5V0LU51
xu6m9kKjKYIvJIe2zXJ73866AFugW6av0cc21QdWzAjNif8ZQh0aNq4Gm18gZdZxWLOJwPfMg2WW
c9XtVFqDfQNZd0YhLpZAOB9acIEjdN3h7n679YtMDGSVGJA8jVG9mPXq4x+8yKTf1y94zNSjg931
hT4Le8QKMrL4tQ31BzZCORWpaqt12sAI5wx6Cy9c4EBVUKvhXxsEZ5dNNreF4Rc7iHyZTcZS8dPE
dmSdN1eE3heCqGudAhqRlZktfiLaYNb/2ZTD3AKFrIXLMWu2iFFN3CfhbWNo7zLS+5sz0r17LkpW
Jhc7JXV0xSVDtQ/xytKUSa/4n5wQOgUQ3vUyz5S48ZNaK8GQ2dwQPmhpUtWFU8geK6phVLkEsxo9
6ABALR3bQ9YEbPpWzmq+0eIBw4Wb4pAWgbshP6GAPLE5OiThKlONK92m53VUzbFXSslPN6T+Sxv9
ZAdry7LzhUoaYwh4xt40EDWd8ExnTtKIFou2u3rB32R0rhNaOjKO8PmpRwzzTsMyvfJ/4PijJIR5
6gjswk3KBp/Iisf+G8dCvGsxKsw5Vu4aUwxudD+BUuyw3XlpjFaYIe3dnIQ32lnBwtTq4xZFFO/7
CysUN4M0fpgE8HzZ07sojD/reg6D5zsU5ei4SX1uIpM1Nvk8bEMfaMkpkJTC9ZCGPqeGx8LjBEtC
HmIpw9h9KFBj2dxRwwWNNMF/+hjEk0+9thsFLttalaA7KSVrYL40d3B/v93lrjx3CDPWWdFx++xg
p6+BDiuhOXmFhNeJTfG/22mhYTSg8alFuWEQkl6zRr8lAlT8/BMAK1reaDdqKXfIEo8zZM330lvV
NoFPeiYvkrWgcsWaYhdIflT+k/iGmaV2cVH0gefBTqM9KWn9vrA/aJ1i695xk+jdWulw9sqtuby1
/KExYrJYf6Ifsfoi+JblW+bv575NXJaeOF67wT84MxIHCcOgEuU1ZPnGNBLcUwUUI2O3jt3JF6UI
KfmdixeyDKFEK+61eE6fnPTgrt6312YwdXszQF6eHMlucxDJazO0FQqgUdz2sYazhQlolM7Qltx+
i02/YK8y1cmC7ExHxSVX/kvpd50bLUPxa6k746G4adnrnsEVLYAkdvIhnjFDDx8Kqi55+wVcNCc6
5P3HZ9mVvzAPh1nxyh0AaKO6ryiTwF0RBLUdRT0+iX32HkRQmoG9aVe11BWAv1UPrJpM02FAlMKA
QaQG6mO7q7AM4IbxG5no1MqmF4/3ZN8skkRyuSQhTAsYRJVgQjvv9lJr/6T+wIBtcA1n/l5gbMCd
ZRdnGa7/cqCJ6yKJVyea5FCdzXz7T7EV62IEzMiiROSu6SgwuINzszDjExvCP8By0Vh9KYNM/rQP
jtc9MK4Ip5BVhPLz/sk4Y2HmVXpJNZXJjrMHEvhTLPC6kb/wmOLrod9KKsRvPqvzqsjatpr2D2oH
ILgG7mdWY/lvWcRsQsMUTY/Rlkpj62/ikcvvONF9aFOl3QdLeTxzdcbPoZIGFpOIWtKF+bPHWm1b
3ytXUxvMFsouizEQwXHwe8xJWi9UtwbndFTcW/vRu8AAfvK5tsyWh0CR2AQtxrLZBbRa3UONykn+
wYUlNuQUj0XYfFuhf/XbCJ6BKSaJ52ozlhErC9TDQ1956LUYw4OjJ1ylrY4olpROt2+WGKsCVOcm
bYrHYq9NM6nSSU3E2fX6vu1ef8ebbcvAXVNkg2eU4p1nftHfRPsPhwHKcvMekDQAHiabn4s9Z9yx
AklavL6MKIHT9ToOyW/jqaj+qPXPBAxv4//cIHH7dI0bfjfKEScSC/pRC3Yktt58TP9hD7G9H6Wr
7X5t2pbQy5pB5TiJW2/B2Y8o/Guki3dSDRh5/2hRoXmwWhYrKxpj01Or26RFD24Z0ECbkM1Vhs1f
AclqMzNk2L/J0TBaMnVrZ1pvKb9OaAnADrSg7H4If6xnPS71C522lsEF98EO7zXGaK1bWybLXaZK
6wchsGYBg59iXmKoBQYF66QvDm3T4WfO3mvJSZ3gEXEFWm8p3MvvbDRDvHsnO7/wfJPGNOrYgTxG
H5BQEeiVacaVhcXnyFdonnmJKmn5Q9lY/87iHHgDpTqD6Zcx+A1RnbHl7foyS2PJmSTxx19OJPig
v86nnidaPV2aSwHxJ6BZ3YqG9qQx+mdyPaQo/XF7q+CfqNG0jTdyoeEsmBtjbOl4spIK1zsdGUIX
6g61PISU0bjSifYnql51NGT8Tk1a0BocL/ojOpIkOIBmPWJYF/Q+IujpZpapKMjM5T2XA/Xo/Rzl
hvb/tp28fmyiRSmSt+NZDKnkw2st9QpjNg10g93/q2LHJsl7gZ+MdivpI92B4kAGPZLDcJmA1w+t
Ie5gHzBHqNqJ47i9dv0V5TGNtsFNJx5URNbCFDsKm3fBU92Z25+0+0Bf2DUOhDNDKkwVZO0ItsS9
C4E2bCPko+iWDhapz9svEOp8aDv7FTwtBUJX9NQKafRqlEpLlUTJ62fyW/w4IxfoHIcfyuNhhr9z
sx+ux7SJkRFlRic6u/Q6l5Wv2c+HOHzXxPmjFwv3eTvjfVqOoZvsrrwMe/rBMQ23RdbWXzndW1+S
PixFQI9bijoZ17gU0zHAFyVIxDoBBiQ6EXtuF4RhaqskcTIl4QqrPXfoUQpbOdlr2IqVswkfJSw3
DNXCw8mWbEVeGfHq97mcQQitPB5O8ssIAQuwK1xzYbRw3WHDJzsKuj06xc6k+Z82cMuH/1s0Ip0Z
sVaZsjvZ+ensofcsnTgQ51AhMmMWcK/XO3p6vrObzM+1V0piFZ3hpchTTW1kGo1NXtYWSIYBBx8X
58pYhNDrcj4laSUoFBf0peARmSLSCoVUeOHX2dbbLp5L/HKrua9EbXhHE0q9qcNY6GsgMTL58H8S
zDnggYlqp6arY06fLePvSvYInoOz/sO35Fd6py4x3TYwb3DH7cvB/kYsHgukz6gf/rQpjbMBUdcm
QAEc9EJRUWJHXOT59OAZD9pNO1SP0V4EDdxnwfx/J+lsMtJuZjlD6LwOUbo8YKSC0uSdLfByHGUl
McO24xUFu/7eiqNN2YcOnI3y2Jqq9wRmJoihkaOsZSlKVn+o2IzlNXxJWCp3bMKis/f+HVpfnqH7
RuLu0LqkQZzcGq9LvM3EQcnv9cxrlHvKdtfcfzrNeu4TMLv3mpFXf8yvARn6RIQWBcs+j0G7J8f5
y71bEAjRb26KvnePeZt3uFf1zw3Ku3z2Wl17FGrDjYE7sfU3w7LqvdzpIp+q69N9DpxfpiB+Iv94
NX89yxVwErl2aJQqgUcIKlYWiw5x23gHTlRpsSox3QD6WLpgfuRRKNzflkJY3hRh3ROLevBvzUXx
6DpzHLrNGRk6glVMf+MnvdE2I292Hea/4erJVaBrJGkoooQjrLlz/wYs/zSgcXMsLIuB4SVqi9x4
0O4rGG9Z1y83NtcpDj9MU/kIf1MQaj+bSAEDDq29+izuQHXnlG2kf1KmOTXJ+H9hFGcDqYM/uB6U
v/CiRk9tCHNjn3VMtt1ruGFdYZ5q87R7TikwthTeGEY51F+u5o7IES9mHxSpUfeImjPZ8WTpNSgU
PkAIOHk2PcbK86l9nhWwUe21VTRZWVuoRmA4z8jLUrXgNs6iW5o0o2lpRfKZPdzXWimyiqbtJNO+
Ov4NeuS4s1lND0SajZdaJX0BubxwYDqRIexLmmi5CEJNDmn/MW8+poN8ffstTkxE8u2ZeYyzC679
eF5xPrvfWZTZr0G8vpXILRvrbyvmBMIf7+fHg4HWhB03A97AK+nFwVnVflho5ednibpihQowlvfp
fPhU+ceZNHO1wBPoX76IcF8jeUF6Ufwudhv8XffK2WQszzL+vhMQZf1XzS2LV2TPDupLRAJgGpwc
RlG275fn9cx5iCnu0M6OlWghcZPujwKfNpkpkWDEQhoMQcjVd9Suz1vdrhrFpZcsssP1z6VghyKC
jJ93fq9asFWvzWwPzaoNh7qIAqWQbD2ZemEu/N/PEcEc/6BWg3dkyfdDmsgfXaZH+PLvdb9w1AKf
DBj2NSKF6xstoUSDagl/k2bFA0HCSujNYmoDjMeQ6qMcx6cGMi8C+Wj1d0dkGKsnV23JPjNtYr6W
6Tl0Wcmp2XbEmP0CKeXW5J3CReA+MIqIck+9+uVvJhZuv/7LOsiMyQIVZ2OD12R6i8B7fP8iYtKp
e1La7bheVzQrkiLj3Unkcy7XvjPBkZL9Vj7ZeTGXr6LHhH34DCxfBjRAxzPej7HzJ/N4ehl3L2N4
wGRCMp/TZQfVFknUEn/SmYbDllm9HyDa/WXbbzfeTMvAJXYVfXytUpj26AzIgPk1fyaZGK0fLayt
Bx+wqRZvW30JD0kHTmd/xzqLj/pviJuQ6Gkze+kUM7s22bGSDdHcInF/YwXQrTYF1w3PMSupSzq7
X6/mXR9xiD5X6QeeqFP09Ugr0FihgrCzi0AwwlSaETw2Cl+jnGCwDD5hi29seXg5mKl8hP+uqlyQ
FE9BBF76VjBWqq82DtN7VSwmatdFRvMnRzvrPZ2fex9IB+dOjVlhnrArnHoKOc6lKIz4RAuuGMKl
GL0nCp1f3a3E0HsPKPRfrfTUOYKM/m8uAKC4lYb04PPd/y/ewJIr6OT+T88l3H2B9l4kvOFy2jib
2/9+l4p02kcm+vJxPL7WPt48butraYFRovG/9QdxkYfmJ4b2g4C51Vf+naSuWlFJ+AOwYQar1SHB
f2aowfVa1Tnsg+1eIEarIZwdWXtZQeYaznWiMk9uKd7kLYVu59cyLJRpZ2MbSab6P0CLbHayxV97
IESV08Wh/DGoUnSb/RAL3YeXVeBkz3I9LKcZ23lFOjzewaPL4jwgcXkJk9kpiFYL6t0F7dIbZZqJ
HoYKNoGQrftRKwthFuQqwUHZZfYlKqlPanfUf8AY0IFhrSkTMQHctxgCw0+ug7yrp7kMKqCeL4An
I/GiogSKv/tB3INQT/Wnk+LWvOnuKLSX5+Iwjqoo0PYQjlCRedvQivVR4jBh4DjIc0Ga2kXkiWkK
kle3uEVOJ88dhVsfXcTcEPmLz9Njf+jf+mJgBoATjJZB903fp0S98aqt3fbUsQ00eLPbqX8vjOVb
z1ANMcEbXUilW9LLcQ964XtH0B7pa/KKgnrKJE0ecFneMZa2x5iL9URolKKz8bLGM6fatrRNTEzl
w1ec0AExxx7VWMA/C18yeXhAPO5Ob1PiiOGZtJXj6CKiMN2YqItj5B79F7eki05FpP34VZ/xDVp9
m7smQoSz9eoCZ3HoW+s10/ZtU2v/c8VXaf3hJeSHblSf4IRQwxLc4h6nTLLwWbiJliftHAF3W/Pk
LdneeKysMMcb0NUg3Amls1HEvJinAmRs9WDhWpyzCAn4kB4mi+3vzE7yPvkwRt1Nmow7PUbLqpiF
BUALEjvCYMy4aGROO0KJDUyFHa6iSDG3AvOVeHjZXTeVnLAxt9NDVz3z5rbmU6nplMEVZDPA77DK
wz1dKh4qwxdmne0EyXNeCmBee973d0EHC0xg8B4ePKCcoFIHg5qv92XcwkK8Y1UkcSFPI0ARX96z
JgSjZSnVBKs71COAXq0WF6VC/xlYl7t8YkF1K6thogu7h0JGINxsO8rdlzEMjcRJx9rGVXS/SdX5
sF26Y2WjMFMgH5QHKCnaXRF0OnJECWvTlr5i4HQJN4dYLJvDG7mQZC3OGi5HdbbOu4gn5/1oVgZU
h0lP2gItnzBCjV6YbOqh8GDevA82wLE1/sjTVw/S/0w29uodMhiglZBTUPqYfrjteVc1vl8Dm0lb
8PrxxkoCU1Y5gg5HGffaWEZ9pPbqQB7rME4UJoFQsbHdO4b+t33NFPJbWn58oHPsErkCAgLJUHK6
RzNCj4ej+rD+0W68VOUXZArDC0hGttwl8V3+zVAMiworGKwypcYopyg3QeaY8GUuTEGV1lcQ+ybp
cbRE4t4CeYfPmEk6Z7vVj+JSaB9k9QatmM+RD50J2VhEaYr2WnpVMMuq5117u01WPyFHEzkhBgif
7mzX62OAfeKMDt/H4h6yf4/luiPRi7ClhA1upEIQ0uB+xnKspdNn3zcovSuX5fmTxBvdY0p/TnrF
G68PTEooVGlGzDsMYSI5bctcl/5baMN8/j/jWNkytducIzz0849rHuBElMq8KqUGWlZL7lYPAw5L
7Lbyl35liq31chdu7+hz/RI2iJmtgsHNvTgkGj9bQWk0xCfsPI895t9rfKcMcVxKJ7qgMLyEfeuW
xX4YJq6Va7JUni7vxRws0UHH6CAtBRbepHO4dpTo5jRIlsUQzb6imSncIeBl0ep1HXpSPP4yXjAB
vke0b0q8AI8Qy69/bN1z1oQNU5/E5ipgOJtAwglf4l37/xoX9i6skd0oCZg8bly+/5GHEY3/cSEd
Fub5+ZuGIRImvfsZKNu8QXUVyVyiByeWG5b4OH/jfHhozA9FnTE8Wc6e/3gapizQXxh1sD/F64yj
HPNI+/+wP2Q+LHvF331IYdMjO5hGVpThU3Ov4v08KLMfrBUehRVLNIDtdVBNJhd4HGHe+ynSjAef
HY+TaAytNGs+oqdHo8ExwQc/xJa75NsJHvhxD7vSSY7/Pg306vNFtPxl4v3K4yzOsGzE12bvGuLJ
xl/eitqnTeaolzZLc54NSjtg/jEjk9VBT0WSB0dJI6H5kei2S0JFz6PvCBWFGxhmSDNqbUpGIbkU
9z+JKn6oD2jnUx0u62quTzscyv1oshNC5Bl3Y7mX0oE1V77RJxf+txbRvKLsQYc+wH+XzluD11Bp
lMKCGGRd/4DgMGQG/+SrVF9oFv+8xZLnHG5FH67SJcOZEl7s6wl2vLXWRwroyyq6oWkXZn+rbCD5
3dNpNpzXzB/p4MSo6YhDgOrzPFvdTgWW2+ZQofDnv3gbdcax8wFIhR7zufHmA5Jw2isWvHjWfGkp
pXxt0hTl4yd9uBlGJ6kC/68gGKk1DB61b21p6a15gc9uZv7aDxKUKLJeWUfuRTSn2UMZNxX6xcTe
1dWXnRQSntX2gze/n6q/meQRqZP0eF6Jcc6CgSa/m5w4j22JFiv6ot8YB9NeXHUPzB9jLC/dRkJV
LE8EZXuOPSBuBp0BrXr5ZBqRsMQPepd550PMJxJMQIThfFmHv5ScqwxXvNXcHy7aRj5d9lBuoof3
up+qdurTc60e8sF3gqKBcSEPPizkh9ZsVmHptZ2t28g0Qq2BXNe3u+hGrBLHOWJ1wKtg5PQ55cTs
VKPn5HmKi0GI76NbiC7m4ILnryCUWT9g1UawHu6Q8g9jAWl6wV7AO6pI8g8czcAAKBdmWLeICxVe
hQFAf/w7D6wsADYbA4cRuD3ftdGRkDcUrwmvqyqCNy8LduOZNz4a/of1knGsao2AF2SSizv0cbLV
HCKdHmC9v06rWcejYSSj2FXhUvgBambZ/4ASpz2vrfizVUue1xestgfrJekbbA0WXThKopSUsjRP
nUOB3QbkEJdw4rDiPRNF4QTmAORLy6eDn0T8K0/gY/aElWl8FGit6GbW3Y29UmEO1u12NCEoI3Or
gHwXeS54Qy1i87WyBnxU+15kJqd1cHe3GcY4I2ZIO3cqQRZSmG3niQQVZEY/rzjqldaauKlwq41/
MN1LXVdzFksoH48M0B+NCTQP29S5/TMefRo0P50uU428QxczdCTYKrRDNb0FlMCU45otGZpmK+Jt
lyjFdim5IkHL6GWOo0LiXNYh/weUJkjX4jYnyDEOlZhuCh6PPfODVfnQTjcQTF4EDJSuJgy4h9li
kgMqFZCKokCI8zmSUNYeuZBXF1YhoZ9GvMZ8seZq+TjsTELtWWYj+LM18A5cFuDADnEP/l/BJvCO
/rmgpSPVfUL6f46aGVJEl7+mkACe7fx1LLTxEKIrCUfYezfMcnKlG/Vtgwm4zRjiAfEcb2v4rGLC
/W7kHch9Z87zAHm0QzFbDl/JWEv4hBy6a4D9EMFJHd5LpzZ6Lr5Wr9/yUnB+ILgReVHFYTAZfhm0
ZqrKPc9kTJOf7FGOjqqmARxdGdvOsv+p2fFdrDDEKP04RoXqOqseKZHGzLLnL8F12koQMHjWbNxh
LpG3wxzeeQ2K4nrAGZGR1UGQsBAQUD5E53ZjUOl8rrqVbjRBs424lD//H86H3JlZHi+lYhhEa12m
V86gW03d6J1c9HECqhACOC/ttuYlkLz0l98hZePEgBn33Hr7EsKQxPxJCTtzye2E9nlsFoBOlGIt
VA+sfk6C8XRKgDfxgAQiewmiiOBy8TpEMa1uYMoHLTQij1KTz5+bgYMpBox52TrdHKNUuO3VhvWt
Ff7DrmFEq1WalUpkSZ44eI8K/nP/RKp3vlkA1p5RT8qoqKkrPnWKowZ5oWdChKYT8VpFma/IVaRo
e3ka5dU2Bl4ErYMMLx+A34PbAbyGEu3Fo4N3vaQj9fqv2QJ/2QqCGV19bQ9gq8EsUBkfIZ2/gsIg
zoTmnJ/y7YQveWMnmCZccOthzeH4w3XDXXA/S97dQ/CDXj2bsUvbTDvUzCiLGfiaVvKeAz5FdSjZ
POHKRIEwSGBv9P14otmZ/rnepqxUzlhk5YlwJc/Ox3xIXFfn/8R1JBCqDBCvkOxJN+cIyNRwOvwE
e1tIDVupytGqER7nqx1YkLHpKQzP59W84Ant5lwP673hbxpg+dO2y2QNtlxP8+Eu3i1NUETTXE1V
5/sAlrOb+s9sHNXzzOmx43dNtixZo0L2U9qLvBWfTzbA5xV/dXO6MdCJsARpCiEPKZpvBczyGATQ
or2z7ji5R4X8PkyXWSpR7UvYnUd0woKhbbSHvFe+QpdIwwG03G0o99titbUoxSQ4jishCp7t1Pm7
0F+MX3C9WlbJgZMIfZvcS2zMerZ7hrlMJRzCSB62jZxwRqliU4wh1NwPbddHf8AtGjFXbWfyEWR/
kxN37NY14Qyf7JTqYGWXvPAwAkSs7ow1NH2Z4T2wXtyN7TgWmmGBwirbLFxwzp5O8nG0VYnHpP5F
MIEFZSW9arMgiWPd4ky5U/mVFh8pKOW/TN+8IXvPaKk9CC509607xBZFPzEuujW/0yfLB1HpYUp9
ojzqgr6stWT3EmQhRmQ83oEtTIrGEk5ziQBLrwWa3vCxXKVfSlwZkI7xG49FF5HmWH6NS+VlAeNO
BXv0dZ9iSLhJ2lxCchLSteTSIrj4TlIH9pSc6oHxb4r6kt9qPSixsKsm4c1ZlEcRwS5rb9jWSL+u
J72BeZED40FSRyHg0l5qEZoI/coWez56LHFR5RN2xocQefAIaeir5qkQWeMIu5Pl/6QS1M5VHGDt
69M3ZSV8IX+HxmE7I6ims3PuXYtE/qMrx9d7+sBExgmT0x8Cbkn/aKtiBqgMr2eBcUOwP9XFaox5
8ZF8OjlMwJRofJtQiCApSFroFErZHoPJNczYsppJO8UC4zYS4l6em3RPqG/JpZIkHJFzxrn4pWcd
PFkrUYyNVqLTecA5qqZAHDmJiX1Vz5PqwFQfSwattGdDP3x1E+hFATLSddCpPJk8UyC/L72hmFt4
w/CH3Wr/FQIhalJHV6Dj5gw7FJCgOGhxb3+nryQ7u6qaHMcFArjhLsMR83epAzoeUjmrU/HXsiFC
BshOq2hP738Towpm+xb66BMLmGLJDocTAsnI3XedTYcG49MtivoyeYADnFtQvsOEtH8RszrqqXyR
a9tKRB2pMSwfqj2NhcQb8y90F8beWIKubeN74NTfmyr6pywMaleqVx5MqDVverSKBXTud9VwbO7o
AehWoaKGrDx9y48mS+LUa1OfCp6vbm95gAqD6cVsXuKxXn65UgMVOwKLrsChcFWwtMyrhn6ArQ9h
03FAENhWThdiHfVVhnt6Cn7wGEv8rvTD99DvMjOpFvu8h9C6X8JXqMSp0mkX+BoOgsdxKJ74yGrk
sO5tpOUqeMZuMy0D/EkOiWQjvJXuXFEX530/p9Nc9Y4xIKnUUC3rWccBiuAnUA/6vKM+stEjpFrg
0LTW/dUOMBQ1d3rTXOcnw9IltxLzQ+liX7yX2m5OtEO7LdUWPOd7JJiLWnnxaZkn+rVtZ+zFKRAt
uDieZcT/lwU0MB8a+HHY3vGpnVntmTcbJ0xgOsE5bZ7fc2r6PEhZYibUK0zfUUyXHfRC9k3wP4ZX
vn+EhdcrXBo8a1EIWN5Cpki4zasgwIcMt0qwAknZRnwk5ArhOII7ZW18bwubIIoJUfiTzKgZSh7p
F6E0wLstKs0WM1yKbs7PErukqcsYDFQOhegsA+znHetQEvWYcjnZ7bYp1vl04ULKzNPQ6JBIM7DG
TjYEMzOgXmz5jBjrxGPSYyR3DEMeIwMsJN7aDwIUS5MqFBZtwqycZPVZiLz05Elc3nV7cuhK0LR+
DzslDrrIeGAmWImDBzyeas7xMuiyRDnSIS2gUA+lQMhJpHEXJ7ajHrs7MJxb8yKMSxJnb+De1LhG
W8RZig8A0iccnxRcYsbPvKXb09bchbzUjTVs0cZeRBa6khKeTOK5gkshBed0SgxengjQ7x+ghl8U
+Ff+YzIzV1oEp68yvkdra1MNRdooDQFMtmQ+mQ4pHbkarrXFujlAvJ5m8Jbr3PPuOFSGKFzisDud
g61S8Bwe7yIYSuJM8OVLcHkjYTqa+wbk4felyr1I/aE+tHdjXp2GKivtUgZKS/n7XqRyzbl9n++y
TrmKhkIvswu33fitJBRI4psOyWyZlbbfCxeJ7IK6YAyW60Z89BJoIg+sDgCjppfjLvVUY5AUmEoC
86iUBOJVTYEo/vxJ2CDgrRwQCV1BkNXetL0M9YWR55mbW+2omPOkk9M3HbLfmW2UJ7qYBoeAN+5e
+mKdE+Pm/py7iwO60L822BdTxDqUzbHSP8djrRj7SHfNgV79nzgWfduSXeaQaljE7PupSxRLnQiW
rPOQ0cTElw+LUiuS7KsGjM8IRw4GHqrJ/8s4oqajnhYFMe7DwnVsg7fQQQAGBsthb3pZcoV/yZLY
e9b1BgopGntDYIHLgUiuflwfM5qq30D/MJjAUvKFbe8kDCTxBGmk7043ldot60SEnbyMNH1HpyUI
m+KHZjilh6pKnRqfYAgnzUo18krZMPaLYNdnBtTrlW4mQ6xcXc25NSFGAGIJJhQH5LZcoxu0WT+i
uAdtw9P5vdPhO96OBH6jW1QBSFbJ2/L+Z7IJQIepVZi09r4lTGWw9Rou83Kpbs4KL6vqxE1QvnN5
1DHdQbFUQeKG0AH4t+XE0GPR+D8H+YxGS57S0wskNcPlb3C+dWCqSdgDhzlc8ildOdlMcWKClrOW
bqtWQ5qQIg7CzB0R8EA8eepZ4wnZAm7sQ3ZxeHpunm4sVXffXaXyTDM6MwSSofcXCk920/JXIUVT
VY+8Dbb/U9wt0jp5Caef3XE+53iA8LUGpFXhROEU3fQwq/RsMg0IdD6S7vsTU2DyPNo8XFK2jpwO
ewg76eUZhS9ZgEY4sEDhYMjtXHAnyFH6PZSdCbBnjfffKhU1pq5502p/sAG7kjT5wDkIwifAKmlV
rgXVnc0Km16IM16bp0MvT58o2o+WsqMgR4UJkZ6c4XZq8RrIA/T+B4G5e7qSQx3tWvEbHmjd7yBI
8oSuRzzmNd7XSqQvKt0RLO3KA9I9Tpd1UinwzSTrkxU0IZYpr15oVrtv9groRVXf30HA0Cm6kYhe
PhwAZS8KQlIyX+cQg+2REwYfCdz3q2U5mmgK+c0RsklMz/YJj4MGh78ZMhwGsch0PjfWDqKK4JDS
Y2n3CxiCMbIwEjdCLen2hwJbGczqH7zgXJ5drmXU8ZDK6nrkrAxkEuC7xUmqepDN2ZjyT39RTweo
LoRvc2lMW/v+315tbzesh+jdLSnmWUILJAYUtQtFk+KMelzpi3sL7j95GYFEab8GG4XCCOY5aWEx
WIS6cJdeSQGJkKJvG7QiMuS/D/57kW04KAOLlT367cqE+G4pl2Q30B0FDBL8u7Wwr2n/wExb5rS+
utrifZGrFHNNQbUmW3bXO0HPDZY2dxmrGguyTwcUorxOEc5LZUQACI9zOkHlXEea0/pmLa5d8b4p
RNeRksztUJ70SY9rkYV7JLqGpOFB7s8Zs2PAprqldbzst54oUzCyJOuaiAqTP1oE+HduzaC6kFZz
7CiQF6e0krB0RIaJG1RMD2/Fdr3Yn8wL9kjcVd/H9iEuCu9KT46TmmczDqhWWAJzdhrmUbNKjP1M
k90uUeag7Z6E6WUdfl+Gjg9CmwOM0DGYdeeOrAk/lzsS4Dc6X6btdktn6Hugm/NU5/vfD5sOYy0T
colIcVkXw8sDiCgV86qwIM/95AW7cbdUjA1WxkKYytf3nScPzBhbNQmFIwtNNlRMQKA9zHh/N6bP
36KA2HCFJrzqBecFrM2Upb38Wnqq2lzAlNT3iyF+0lYs+blS5YihtUpnrmC9Cw747NLjtLSMP20m
exRdnoFSS1vWgIgKTZ9eOTAsp9EZYTn4Fv29Jnt1q1TRRRbE5mVOM32LsYYQS5NsjYzuiPTbv23b
zoIqiy1OczVPvxsIgBlV3iDe81Fz6QzyPc4GQkJWo0D5aW5rYh5f/Sy6P8cPw1TA7yjLcF2L5Sv6
j8iAFu7Ze2u1nnpLO7E20xUqKq1nP7gTuTLDNbETVERmNaM89mhqlJQ77K4L2QpWQH7HZ6bGKtxe
n4/h19vwlMBWhRP4xSMrytttIhX5S0zvTFNwvtQtKRgfQXqfalbKm+kiMt9UMqpGCvYzIHBZWrkW
BPKMMkBMzFFgDdnk54grGN3jZCnoaj5Xy8zUl7y3pg9FkpzctegrNStMcVWPJiUaeF/fZLM1G/yV
geMSZeBLWcqFfKgK8J7Xj3XLdzsGWMqz3oq+iGNjawpL3bwGn1p0WTye5mfCt8irQG8EHvq+qd6i
GX7hqSA+hTU/hDqYK9J1IFNyjbV25+VjuA48IwoFgrK0GNoxeQfm/1/OHuvxzRgjaVJXh7N4z7dD
3TcpEoVGot4gk6Pb8oCAPWXtUY1wK3UhmBYA2TV0HsS7CkJkP/m2ub8ddX1tNNOMUoFnK6suHeZo
CHkAxdMYgNFQCl95Mowv0ifYteUXdt9PvkNbmVQA8FkcD5TRZXLAi3iCJbiSG7+cRSBrL4QMgPAZ
iR5bMczS9/CjoqWiws3CddzfBZbjJP9AN9/sk9io/j2+YVb0asHARm1UcIvZ4N6vmttjshbjGUKm
WvBhgpTobJh1/y3If3QWPJb1oIzrXIWYNq4wOHP6fjoNY2jic2pSgysJP65GPTcKvZ5DlmCIThZ0
KeeVwWjfbSu+R8wGdhSI6kY8x4RkBIwXMbuf6bdKWq0LVlP2iykxpTNqm+X7cbZhb8Ep1/pg+hGT
J/CjyjFX7Yf3CiClHzZYVY68Q+Qgx9hZJ4knE0HE48weQs0d40IiFEJDwWmncfWE1hArasl0ABD9
yoNBjZZ7FWNRIngwJm5oJ/9VIkxgcuhi8t8hEdDmSiFJglQJ4ROxlLgIBKeweT25pkkO28h6WuDf
YAX03oNzu7s7ep1LqH1kYLKEuEdsvUMhpmxo1/0qs52SPBTHjmkW6Xf5REbtdwMNXqFhL3D5O55D
pqks04psEBwwf5qA8Ic3XrRKncOMWYfv3H2mwhxXGlkzafs2bAEj72HVrGnGQNFpOu8D4vMCI5D5
jMGT4OPguVSvD9UO5NhrH8o6AltUQ4WGb0UR8MJbrEsYavcmrWGPb+dljtdPxH3T/CozO8JlQeMd
Bd0GbunfFn/OOZgc4JhJc8pqLppcsDgiwd8GUvkJdWyzPGeEf/ffOorGeTaQ3rMvAJhq88++3AaI
a4XyRw8OU4yfxaQzASUD4mmJTMgAkPNslA41qf2hPRzg09pRQH5c8ek5MoYDaQeqghUbo+RN5A6p
7gZlyvlu5mTSXWKV+KbqYgCKkUZqIqJ78rrrDx6OBRvZkDiNjMGH3gvKvD4WvXBfULqrj1jkIguY
fmrewuZM5mvtEtgNi6M9F13gewNVNTvT779aq2NWwMuvervKieJWjeUnXKiSLMjp4SRc2RzdRCKS
+1zY+JjIJ7mQKa0DoXQZA71qvp6o1jYxG+n9zImNl5H6hdbTTtVAjIbEYufupQ9FE0OxETJI+GoF
aVRFx2L0sZiLUNWvZKg9Nk9IUNEmzXiDi9Hlz1AVSW6KKu/80Qn1zWLFRN5sfipA+GFQZmkjZOG7
D+SJou4yijXIez78tKNMBcZjhLiyh7fQ8MVE0HOCHqQoM5EgLH0r25N8p8WQWsAm2wAj2l+k0Emj
PbwuBqzmdMN2qgC6BXFGXHAoIVi7vAxhRmZFTXB0gMsZIFTpCHnUvpNTH3ACeIdmJhR+r6NzoNT7
d5NEYf2MqT4+WW4iWZe24DMkc0BAO4wP7I6/GX15HZX3fFUiv67e8tsavZhahGgRPP0F4BhvbbX0
xjICJBfxueWaWL67vBHHNFrhnVrlr8L3mLEaNo2YVhvm3B2nCISzvIeG4PmFiDV+VdcmLmixCIxd
L/HmK0zZ0y34cuhaNUkLsQVcIW7Yeqm7cHTBSn+LTfr6nFbVHqYVtfP0D7/uf5F93iMW9KUTeL59
Kn3edNUgo5wq6YmaG7qNkesHgROEFoo8zhi9H0nYmszByeE9VmvVOVWGcHkSLpvTeumCnzGtuqdB
bDS/LYgkgdu8fUxIo/u8LFN6WdLCKrMozIIs3g00XQYTyT3VsRvuKLvJzM1xQJq4HqOIAEJUNjUn
nM6tEVJ1evN/iuVHNehObjq2B1a8zO632ieGWATSIK9RsE2AW53BcgzAQx4uz4XdZgIMw5foByvQ
Ce8GkFAgfUBmtKOzPFpriTvFfu+wrNjTclmQ2wlA0eCldQPu4Afy4FaTfxGYWqgMRWM1+ejrDU9O
XjWtjQ8x79KcBpastXgqIvgttTyUEOJgI5Y93xOrHF7SMF5O3wNfrSEQtjmil04LxycsKeoajfZe
dE1n7krX6SMHMB79DPfSNTGkKZequIic40qL0cU+CyIvvA2YupKNM4IBMS6/h8b/cGLDNd68QfAL
YOoybcjroVt7pW7BV/fcpW5S8QeDusyh77PSRYTV6+F5rc94Zx2QyDOnOUXokOL510Nak680NCBW
rhH428SbqHyvY3Z/M7ERckNPhHudkq9i5wwILqu//WpQPC4pjWmDp4kNGnYvQZmhPf4dO3G3VSSm
k1EtyqOG/Yf7S+bwWHfm0TsfCAVzQcFAmm3aJifpvZgb2Q2xwMCjmQNHhAlhZ1eiJTsf9hqSbsx8
Qrl4ZV00qQ9oOZjzPwz37QzhqEjdfyxu+d1Yhb5Q6dAIv6LvDkOJX26CPqEG3PaxJGmQU5iMnAjc
Fs6PbQ+MeS/GagA1WDd4Jbt+pl+XLzHTZbDqPksiwlyZMpfISgfYdvrCS6xm0jjeQhtHV1UdpFoe
3QMPzfT5RycJBVmSiARj40jQdqNaJ7+YTKE5zdKBJ4AhJmdAv0biBRrJOLKbuG/iW/rtELx6z+GG
TKrQS776gNmw/s7tKQdCPlSfvOv6ozJJpRk00v+XiQpqSEU4BxhRbLOaIea9JEIwP/z4F6/pwBPD
BxxDc/4quwzLi13AO1UWEXludMMH3VleXPNbXQ+IV8MzRclIu0MgxksqBlaw0ifh3+GCqLKQdEDL
ZjBt4mH+H3M+W1knzOSuy0+Wwl0FB2Syk+SLBEnryGMwGwhFIh7z97IQ2+fHNMQMPy/EPZcHxQ57
Pr1scWBFtpxSvNmUx3oLKH4mjT8DD6U5JIoibrJh9w5qQuVw5I8YdTkhVhfNL4T4Oki8Lo1+9340
LbAhTkw0vSbA/VwwKq3n7ab/DgnJ47nmsTFxS0ov049SJ4PnmA0vmgmCLuiagBPFxy2Sv0om+dw7
Jw6y+fV3wf23X81g5oDqTrK2YxqNxhTln7sEnu3BrPUODI7SLcxWYSubHP9xrwJHCfsFkworGUc0
QrNL0X6kdoOiu8vOPQUAsO5Tg9EAoXuNjqnztT4pEpAcAUNr49BZbAjDZ5QU3FsF1pQul2ka6AVf
MtsfCX0OHcUH+0ZSatAY2NCA5aFJmkRKmMG+6AuzB7W2Ovxku1f/aYUwGnMVpikorvqufRDGbaBn
4wV2GixJUjrFWuXrBqd1K5Gs8F/bU0/yBD7gHHbyj9AJr8MTuohK/leZ2brkQecUxT0J0r4DyQmP
EWBAts6P1nSffBrKaj5gBjF4CQARqL1ovLeerF6BuZERtfxfyAi249T5oOnbl0QU0h7ZIwqjTs1a
oOXWxxpxtbxjEpl5rLQaWYTjsPgnTQOEBS++HIglzAYTAoDKHqDIrUBM8ntycg4YazpXXXtIffxr
CChuurJqCJXqD0nzVP+MILZSXUW4bI9bbNPOSfXQOa76avTU5oa+Bhyix6U0hMFYprQc+Yg5yand
31yAoCKybN3X1Am31PFnrHutXsLNPBqeSyQXexJENE/AcBr468cAan40Pl8qUvAjxQuGK5VavQG7
3lY/QEPx4yKJLdrBdi3UeRUaTOt5QmvL882IQ96YKl/SM4j/sac/Bvcb/xRBqwyW2Gp1btY0Fedy
nFudXgf9nOw6GNkd3ejxpL7OuUugV2xpO+NFzf3LO6ihk+xdfTgMfymPCzEAjCFS+eTt7gqoVvlr
8ELGZ2JTIfHMBP6L/dNWsvjQc70dc9OCyBiLMw9CFs46boswfTT98e2Fdl2eKnkGpGCUoUI3vzU4
zLC4Lm83MM/+oAfh3X6shYO+YW7f9mpa8Ot7xCybXUnnE37s/ft3gGLU8f812uVaUdFx01y4ftd0
Q+VjfpBvzFDt2vKxOP06jAgLlQeu6avTVg1MlY+cqELjpD/Cwrc4XREGA6PnEVvyCk72zId6YJOv
l1zJ8QEqKBdAu2Qt8ggGHSJ0LG8K4HAz1gs3GU9WWj2TH93CR+hPbPLn46E+S13gWUSyxJ59Hy5E
apaavJsAWUdbsiV/AeaXQYesMonvtIrRnF17uzcNdZsCXPRqXa4BajUNaqyQdveo/YpPXEWuvnds
BJv8D3YOUiH65+YeySzaI79jg+ESzForG7uOPY+kDynfWAbiGXMS02BLWOFSrW3F1p2lyso+FzGg
btFl8/Sr1g/vh2x5A3Sh9rf2ZvMyzmmtnq6nSQ1KkWv0o13wZR5GlPM8qLEbvmfM6HsYxK7QmyZS
vEFNQAbAPrSIehi6rCciVPmDduNeaol7Bz4K4KWpuATRNApfa7O5yqiFBirfJIF+zqFp1YM+TPCC
Y+s3wRRvgfl3UWnmH6AB47s1scGrngq0/K9X0qBoxwc2hYT5pRBmcz6v1/W/RyltEw7BIue+z4Vw
TT/DldDfpfhDoEky3OYi+4mXwZ6jqvoUcE0dMz56EsRldagP2Vx239NHDWepYwzEFkUoidgjp3cg
76l5FPI4wVZcPnBS1yvtb0PoM1u7Ov2nuZnEmOtJfeYmGyqymBoxA3XrfAYSXPlexW29RFdw+D2N
nWhjIvGuPRaCEgsbgUzdIi/iMr0qgNUO5c8FSUZ1J2AeDx3EI6cB7t8zpwDDgsYLqdN1Bp4x0cG9
+7zkRDsGR+QBvfi0r7UztQoFaT3JAoULqTVbhTeGnChazFt8k3QszQuCZ9/E8XrrXYIqOayJzZcH
/AAvhscjYIQvSFulWn8FGX1tq9gihKSFd7L3bb+RMYHf1YZrJN3UCODQWhhM8+QC3fhRJUt/DHZg
3vBTAuc/XtAM36kLtUzUel9EPm41rZtu0MMyrwrgcTldz8pvoUPC4MSe8qesceYBqDv4vF1f6V33
mzGkSDHKsT/wMPEs5a6Qa32kEIgHPa5dJYiLUTaua5cgtLOBdwZlQEhy8Va6UP2xh2ZDxorULSuU
ENPm13GymON5BAaYrnZoJfkrls5MYpRq+FXGyfBPKcLSO6FuLTo/w/j4Agi14b7x49Kh++VU8y6J
PiamgxBQPAL+5n1ztSV+AkTwGnnntlANbObLaiV0MKrDnEakD683yHEiiz8ROxrkVHn/joSw6f/P
2FDnBkouJb3AyNR9swz779XRgh/rZBwojPfWfAUiYF/6bPXHBMRUNxN/Ybd+QqW3iK7Gwh1KAjTE
baRpgrWyZa3oV5XrGOPu8TSq3iSAOkznlZFkOC8l1zY1nLzx086lg2XbWlTGGga5gmCJelXnf7H0
raRlQP8YTTCJ9Cz59ZjoU3iLuO07VXfz+LLu3yL68Ip8gTJmJU2kSCNKoJ3rNXSRaxb1I/cvkiL6
HKTFRXplGUKoIzCvQH4/8gIRoXlWB5bUdRQm6ZxtKFh7xmpjbjmVsaenUDpESX0Ry9VgI3mZ4iww
twkHfECYoi/1xMy5GhXTJbQnf/cpLGrW8Z1DFb0BolQJ0h6di/W+wpupgd59D9lUCNa0b1eGu5mS
t2YC2ixsO/oiqGyMGCOIfGUvZF3X1R5kkaiAw0bcYLhUTjwkxM1aRHoCcrrEatYahs56m7oIy/vH
8B/0sWkD7TG+Q4IZRQMaDnYSnZOk9wYgbnM8gCgOAPBU+GhBntAHNAafTpab4WnSnX1ehBwQNvm+
00/LKAflK0TSWk0N0Tu1ntHZQRS6sscSYVxYuX4dLtFbhqyXlTgaBWfxCtYd8MUcOuEIUsUYATvn
PINT9ZzucxbGhu04xztXKVS42/GFCC8soSAfJh01R/6qwJVh8tIH1yNzau8BAe0emwTCwN74U7Qx
oCcaPXm1UA9AM6l2+XRgIHP2BIMEBcBGxsb7QzZfReZR3G7nPRXhVOWQgrU/U3Le2mud6VIwD4kB
CYkUgLo62jmm3Fpo/ZxbDtWcMr/p2MxCkxBa77BQzzgr7wA7SnqQQ+W0c8kafsQos8mH0GVXz+7f
HlYBssv5n9Chp85Ol+F+8PFnEyapEm6/AoW7kknXGcvW38KQcfPSRi+v0H3/t/Z5Z1YXT+LOwvGr
tW7TzeMZA6XX1SKeeztjw18upfD2sjYjAbQG4HhQPQVYuNhZCQ676P+fFtJgxqrew8Jq63I9XXYO
Xx3q5ML1DW0z2cyVAOA371wzCIjKfGsShGmIQU0ip2TEdiPdjG91ZO4WPvpnAAONTDOAw2DziCJ2
/8NWB+RXgJX/Ukk84E8hj+folSRxE963uI10VMX8zK+taFExfb8No36x8L74fKfqAtfvu/6YCTOm
hqvc230KxbW4jYJwPU+Uq90K3n7Ud9lphyYAxg0Z8JoS95Sn+QI+bFl47CsxDR77BwHy6Big0Ipf
6f6v9XHhJVGI/Q9lW0wx3qU5UjxQalwPbhxTCZt5N7ITBmyL5pWDi9LsvWrmcoeqeJcJiKH5t/TC
vj8ql2jizdTskQzBaxvEkyWCBPgMbvk+zzbA0wqgBhEdLdm3OgwuSA7oHBFenPnwG8hMz+vkpTWW
8tNOwFJHGJUGfOv6u3W9dGYI5Hx2KBH5UYOo9raldEgQQu9iRu5SiHO4OmKauB+Q9fd11xXAinyF
4UjO8wgnEgudlsfYYDgScL5O0zhAqMdnDTFnd9IasM6HinRPO8MNiytdMChcKur1nl7nMSHDsaoG
X1OAQ3k1tqLGuhQsp4qZIYJ1bQKMKezJmB3tly0qjwKMpS0ZT8BVNKAmKfUaF2epLU6queJI4ahe
MOEl1cdJyg3caBvfI+/suUPSM+6FgcA9m2L76yvby0DR8XXdyXC0SDnE89PN43zQjAlx+B2uZ9kO
+UE1QUIwusORYJ6SKEbXrNTKliPznUID4/S3DO1bglKPG7wp6gmzw8tM+pM4/jmj5UgGAQsD5vqq
bhCEuWhYNgHBjkk95e3z6o+5C0VTqqvA7inNql8xPhmqrzo6jDaNeJp3KCHoKjOqCSUkpgFnaTCr
TrAGpI/6viz4afGpSoLnSj6HiRC7G6BkgzhQuoaBqIx96hnMI9AFlkRVtEMzc99y3zfxBE7f00Mm
wvEl1H+AZcgeAEiJxRFxxiSdrLsxh0pj8K/iBb0JluGLQcdMdvWC4U94aZyKZMYNwwKY4hyXdCEs
ax8UQ+J6efexQLdfk4xGLm2AZ+3znViXcRifzmsW6lBxnq47zOB04mb6VNWcHx/sDGbgsxrRn3rp
cNTPyRPYsfNaVQXoy6NII5yDf7+D2kiUiqYZd9rR6VgyD1dVoOJ2w+fVjDXtit+gcnhW/Wts0MQk
Z45PYBtpM4+fnZU8EvIZqc2B62Fl6bfjgdx6kFkkf4x+T0StBcYUM9UKEEA/YlgOdl3G9PxEESKi
LoK5++VSxNjeSu9NyhN5c6NElXlzDJA9d1xhe0WSGPYwtwYdkdrTxhMaw6A7NaImHzkRptpJee0o
RQvx3hsDZMNlcFspbX0N9w8E43FLiUY//uFVpeSYlN+N/QzLgP6ThU4gNRPKEKcmcOH9wFITP3h1
obp4Dx7awnGVNidCJRwvqIWKvGJSbt5sCCnKLnIRTpav9jqYv1wq2DWmaQV0jnMBEij3Cbf6CrNP
QIelItDtoxOqfYYuUif1xlrewjeph6giLTA6xdxi9BlgRoQ9cx0JGjUhT/KSAJYkkFCwltSX2as7
lTzxs/2ojiRiHElMSK3cTEAuXIvFIG/RAC+IsO93eEGLuKDhiig0vTV/MuFtOKypNTVCf7A7nuUN
gTPPZcrNz5m2pGbwZXereKTBryZONOW98I/5neWcof/hRX1h2zjn5NuKfHjVMKM8o2tTXhiEFIUQ
IF9CK+2NS6NMGYdk8oxXu66wzpfr+rTAjbvpQuF+N9kpbLR2/Z7GWWDvwujt7wEUWLXwJdBsK/f9
wKsA42xEvgr9fULuagkZlOyrG7dMSeXV7u9IrVy1/FshQhA7c8ZirkBVcIyfgBJsaM2tL0tj0+I5
mG1uWcuEgZ2xypN5dqRxR5vjo5CBeKzUH2PSF+YRedNt9W8t8qNSwT06KEyn11eW8qmlHTSXahOL
FOTOO0MndbDTgeXppEOJyc7NNMQ7PlefDcZ7HkAjFMrmjGWknb6K2AnOL5SCuG3pr/IdMjrKWl4V
V3OVyTh4gPVyodnaQDpKYhUqGIjMojokz09912XRcRQXLbbC7IR8jWZUohfTLOXyYDTSCPL0jC7F
mkILlxL0k6pDbWyHvUz98rsKCLAm4dkeF+wgisXYD4aiSzkcz1mR7uCiG9qHIK0w5Q1Vfa/9IsNc
Ovv4l++/VZmLnAGVXFzU5/B5hUQEOzqoMzolMGmvUVxeG8KpXUa2fQrEwUHYp2yjwEmp/n0YFibd
3nmMy+znwWFa7UzIDnDm6p939AMOZMGjiFJGGom6DNMdpY85b3UEEyb5iD7Aq++3uYIAq90JzJF0
p/YUL1MhQgTFrYr+1WAILjM5KLvJZIFTkDNLjI/TILS2kaDdpgYkGX4Ot/SrCr0iLkybu4w2KuhI
i7+prRZ1PmStiHc9Cu1CaiyfP4Ha8ro9JUa3raqAFK7d8reT2c5eAQeW2gQsnIEol1LKGqQ5W7GF
ZAH0KSANHOLokGlz70qFBrBz2GjKhdjND3nNAMHORCcCPGy2c8xGTIOi0iMxrJuX688KAGt2XeBs
DCbuqXTE+e2YkMhEn6/xCD771PVcFbk+pbsheE4OU7sIg8WKdZ3qJvspu2mvAFqppSjjeeWhyPSi
XnoacGW4/u+KeUzutRw/sdOa89gbs6+AlkYhAGr37TgowriDRMdI7pchyFBEEzJi04grcjbdAcvT
fCSIqb8cCU5EjyC7vi4I9oGyA6aAWiJbAZ3RNojbOcTNJxodfZXfLYsT+N449MwrkBho+ADjd7a3
eThNMFdZWhxJ1kQkfDmf8ZIWS8+uiZYj6JsBAJict5iVoBMDKqgxxgp6g18n5S/DOsXSRol9aBVL
OtaIdvcvY44WFapMYZLf930Bjeq2xr+TN9f5GNhegFiMd5GhJJZlQZCRxsjzWJoNgatGL4ORsMtC
H1AHxZWTXfHjUSre2TNfgb4dnL7aZiiahH0HnTetZ7MAAG3PFwLru3SNAH5CbLyI4WxE5fkO64w+
frLnQeZAsIZb6y80yhujgqiI+t7oOSZkUZwLebACp+qkvXhdkzGFE5Ish/j+/hN215OosocCTmgZ
lX4/vaA8h7sx9ymeJE96wJtBVVI1QSLgdcm83eGhdwJqECyJG1GJ+3JlAu93ET1Sko5hao3G0q9t
CGas1w2UwVOIuYyAXQgNEFYe5Ow4ZHIemue53aoCZYp2Uy909MFfCNc/ze+BHtCv8j5I8utsRh/R
ti3jeRWptxUOzMhclGCUdzNCZYP5+ev19G72S2QeVh6+EHRTngtzPuIhIPgKVO6BU5lsHXjQMRL1
pfdze3Sv4yQORiCxKs39MjMpFLXdjcNbvfm6lotI4qSQUbbxqJKL0YwUk3KlX9ve04MQ14VOsqd6
wyYb3YWmp5kJeDL3MkXX0PSDyREfZ47STyq5Fnyx0JEYF+qLfPT7ptwWMtS9ZDd7Ec619CYRdLM7
J5T62vDQff2Ys9jKe2cs0yT2VdpkG12alps+xS7Y5B4UImLu4gPDXRBFvUFn/mttDO/3kXpdi5Zu
1nE8e+r4DBXabzTVx01N61rqZu9soPXMu9ylfopfRZgpg1wLma53nyXRC9n3bLAI+gBxRWVFX3rq
8Xn50z+m5qA3Q9PyKeNfwPtG1Y1jEK5dqLu8hKINTlGLLv1yRSLwAfPPncV0HIES6pNlGBQwDpJZ
chUOrYOjN3BZNXlNZBLrBnDH7ZXK/kMnRW+2Hvz2whT7ppdQwy38cxv4sJOoInUxgEq5EzJ2BAri
acKdAirGhxKObUO6XRg2eFH+MkfvSDF7l88Riw1y+lq/snogA1dguaPIbvF/DEC8eJjTJBLgiaHH
b+rT4cK3PaaiAyeMIZZ/rjm/gJJmz5WmvIupd2B7HVzs6ZwUaDsB4go7YVEAxaeFfJHXkaeeECOr
/ze6LAor1cVqSI2eqy/ifsS3pwvch8wDA0dqaM9tfSf2tWFWV8qL0C9RHmoFLedr/OMQ1AhiJ8CS
+7NIZ6XQE0omVJ0a42F20Bc8Q6kFSKzVPrp93c8lX69HW0Im3+n5bYSOJnE8B6yy+al7pY29i/z9
k0M3SdVxoSYJtXsHpKcD1kvoWQkmBfH7XN7fzX1qaaUer7iHWwsIFFJDag2DyUvKZZrSZ2MPWHqJ
w/tQ4/zpCZ9/pntYdyL1uqDmhs7OCpUdTeWg0Q1JD4kpz+/2mLLFcQrFuwkqoa0rWmIQB1zKWSwa
QSFsa/QdQguQU6wRGv18VUZiYT0ZvMaOdakUH5S2N6BiZWDHSlrIekGJBfsz4xmptgtRsMGA2Iqs
Uddpgplapw0Y0G4ZbChdHrr0UWoCfAhjB0FPm/vlixu/sE6Y7zBe02hOtIyWTPimNEWJWyF+SoUM
G6E5BSN9BJc9urTAq6fQ+0UdBfQX4PIbsLGi7bNZL+zifoXvg4Pfm7kGI+DcSyu3QSxqZTqdd8e2
JYYrNpXnphHWGSl+VZuYUoHDlr94zns2VDWKZddkm5BMPp/Y+nmvadVcmbmlOzzWFo9LsGA+f7rI
NZiTJxg7bJB71qLANqKEMQlWvE6RCicxT4Gmgks987H5b5rikl7TtL8iB+B6KWi3vff1QgvX3wYO
gukFzi8M57cFDgDFyCtS4MbkQ430gDj6S3miJ36XysP88G5+wCZHTTtVJjM7IWVrltiRVKdsyuGM
tstgL0+hj/UkzJWw7Emeeo5nhgH+4XtW4AmdIDU5LUx+G7x6WKx2OMhkODyfOWRRXZCJEsge1xM4
709vrtBdSEL1Xf3ZN9V3SN70JMI5fZ2cWrzXKUUKYnt2nOrpKohMTEMOe7NWPmhOTXxwSxHxMddB
mO5CfwBJ7XF9c5VTqBVzGOMwvo4lzO5JfrS+feB1XuPCwmuKwdp/4yX60qtmirEoh2PpQshILZ+F
8smyED69ItVE/RNVDphxgQK/XzlTDgloOm3mr5e52Vfqkxp7ThhZHMbhJa2zVHxJSTDNdrYaaUzI
TpqQG8Rl1KZYQoSjLHEvG+kJj9i13b1u+pWcNkdcH35a1bkumoN8DY4RuqVmzrnaLZ6KfWOkXTh1
qU74kM+P3od5VmSh6L4tgEyEyF1WUryEzt4xnj8sm6JXclWvdS9zxMlrd+zXbBfJ4Foh9F00URpz
vWwhr8lCt7MMgXOkc56zsNd2aYD7tAEj6kClLD1/rOHni7HkP3LwRehkJrd5lRt2/9llewTtPtA7
BWXS+Gk5cfYoql6CigGg8K2JFXKyFBenH9+7123NB0FhN10GyAuEjv5ZL/bSLdHHDPN8Op4qTT+H
vSxRL0aZsM6QvxHWnr0FTtGosK8u8NtiQhU/gktElQbSlKNsgX/ws3Jp90RTAG/r+t+GRy1QDJ97
tDTkc7vuni1fpA3GuzQPQ93Kl8MmWD8pgbTcEtIqhD9mfaw2FpojHjGI5X0211E+i7396oFGGatB
BbK/Ir36W2fiY2EeWkUzNBQjo60s8SOBZb32OroWsv1qBZsoYaLPtIcUv6Ov/OGJgu8f4DAu4qnW
9hGsDwpRQ88FJjNUgp3OtzuxYHithju+lhSHLcM1RRbNqLRYUFDwG9459krstBGBDLSbBZ6n1r34
jnERDONJmodbnUatVxNAvGvBcpFz7gQi5+3RysX7fBLTdDdoxZiY1RgL778LPeiFCoTecFhfaoJ/
o1NGJCjS8TXrLcQwmYwIsCr/1Ixn3cgUSRViGmhlpPE6fDIcn+VFxf/QY/8fYoElDP+geV1BBnSJ
EXaHUrLMkKrIed3a7lO8vSRDDZ0HjWUX8emk4WkGpi8zjkxu86ehvrOA6sNVs49uv2F/Pqs/ivg4
mANH+QT2kuA1B+nPkuZkteuKhfiZOdWfP1HB7i2dsx5y5jIJukwfhInU3R7Z7gpJMCPhZDwsXs8K
NZ44p8BpvFuro9P+DdRQoNWVBkKdiYsWSDli5SDsdJ5kUmpcJoKp5hBK/YaMIRLmvG0OYos7wkn2
/Pytw+o7GswUOraKzOdVHWY+87OuiyanCoWHO2UpmYYHwY+29F7Am4r/d4U/P8r5b0qEJmL0DIZB
9FdCfPY/vS20eT0C9WROkZ+pDJKa3/SOwGlkt6PFec29lK19YdXCUZFWPO3UznfTnlc/7bUarVW2
Fm0vObuPreufGS7AopJhIwVH10y0QZsJVfE4ajZaZNLLzERvGpEO5cLvrawoQucL/78VN6jscjTK
bD3j5fh8kFWGONGvdbd8fQObX2gq5ni+a1PJzrDbt0kkZXgkBYmezer1UWdXx+RNkglrgPc2PJit
YQppEf1P63FxCrmK6NwU/GeKg+Q/iAUcqlXtz98SoOlT/ZYEnusErhZeJ5tNN+RcpYhQMH/r3L24
vrN4X4BoQkVYjLaA36rSQawQ/ALM7nlH5uRqJnp43fnOcrmlIx6Rj4LPw/rczwQDdtPcR0ver76p
Dv3+s1mdMYcgtjOOoh/PZD8DEaOkDD6Q2Ut8O0KWtVEJ9CRUWN9MjOpuw7Mgp9qVo/+mFcLv5rfd
BAwWp9qcKWzmzOiSNjVApxlVVZyVs6HbhVghTVoHk9z36Vez3SreIu6kPiuEmR8/Y1+9P7hGWvUY
i6vbaJXFaO/uMi386J6mmZP+NNGj6mc/IaOjmpdRnR4U+G5G/fNcBITnMWH0DJ4cPhSixq/U+EFm
EwlJQez0Vyz2TbqJXPygtpQ+crjiG4DEjVQ0j7w5ikisOOcz0pD9NQQTcLHNMM7KkSRvaL0ktqc3
kUOej7wbXLE48LQIwqCVJ4jYaFpxajN2dIawU1o3Lo66Yi5vJoD4itxyPJ+azEUcsMsrk6hjVZ83
WOiHAe5AtGjfpbvea8cUqVTxRrjKQLnDY4sTZ+Suw8UB+d7pm+aKr97Sj9dSIYrX1VvdhqpP9YnH
+vx/R3mwFhAHI0k9Lcxvwjaz5tAPk/Ydv3q44vtgRBWlkI5MP4mev+onsPHf5Sjv9FNodZdo3f2v
lMjIeYlLUV0MRJRl3aWY9yk51Xzi0rSd5+7Z+1Fk6imnAZOp0fjfaxf1pJLguaFDilekNCG9Jn9j
O2LIpMqSHytFYu++3DB/VwzbLE4dl9wRYooFzoj5UGztV62tDLf1VeWREC33yjatlsWgUWTaJM9M
c8Gh8e9e6jOca2stshJfLq78ZvUz3mPoBlz7rHoSBvkjkwLOMBZX34Gqu7kz+dMOc46NocdXuzIr
GoN8jrKqnkSYqucjkBIhENzwKP/s1EbpXrfVZ20fBD3Hsr7ljDKVr8+bxCcZqJEqcM1rFYneSg0d
OAMMO63fybNAQeUREQYEimJY7I0DWMfFdeOGcm/vxLGLWPtGaeg0NCHYbdkvtdh12f4SUWdcVsDe
Dr+YF2NhtYWryJU/QCiR6WeFkxQkKbDpeb3wdrko+HzpWKiBrC76i6M4hUTgVJKxaAUZNXhONNSb
/qvnhIayiQ6+WU5kBRsFEaxnDTLX53FDz4WCr4sFvNpYAVA7UOiDwhKLDHzODGoEKVOcwRiAquyt
I+REZVPQ0QkGSR2LvrzWedLR9jT6RdKpjTcshuDKebG+tITHPz+3mbJCnjnqBgQjP4ZVDiL/9fNt
rxcI8I8UlFmFHx5EHK9TelL1FdiVE3aGIq3bewfkzFWrh70baXjeiV5hJhU/Xwxp5BvabJNDxcfM
m7hrwJZu9u7naMr/b3vfz0gtAcK6z+fF2R1rLpWiir/lJE5IOHr23LRcaRQ4nDjRF/2AZBEQYOSK
qzlA4xiCi8gXWauINmkmiXQKSRebOAIZ9v8jnLKypGhXxtHPXEJay7V0Xx/nXP5fbq4joN0d4YfG
qpZejLw2rIWrQhyxTeO3EJhR67Iq5kyeqM0hEKtVgeFnyEbzWFO6R43AkA/X8TWiMLNVltPOUmOf
1PRm+OSgjRdIE0h46ZIER6FpPhSVbhiXbAelH+2qNwUJfg+XpSmXjrsmbDbefqNmEzVbmAFDRu6F
bVoEvRqSH6LEAOS8QJrABCyr6HG/SJ7l2m5uvQOYSFJfZKcu5Kp7jrJMJD/7g1EjrfEI/OIfZdLV
6oaZbjw9Q0Rs5ntZqYEOw+IOGftM6qeNXnz8x3naalmozktiY/bbVrV2VVid9y853VHOdtBA64RT
Wpp7scSngCjlS41zTZDmoPnYDCa8gZXnT9Fawn0jS9gXNCfM7BxwkepB6/UsR0eMFPuvGdxSTB25
AYleGmh1AWCZJcPKtqB4wYxS9t7l7xtF6Qq30HC9Wj7WAXumVgJUhNSMw654zkPvN4FWMpzPT178
szc+S/8AEnXVqIZWCgF/CNpAr+/ZSMRFFEGBuC0qR6tjLDJzFv5PuPbVxJ7KlTTE3Jloo1LTEFQz
Z25rmS32B1gtSys+vyfA6P+dU+CXIniQblJ7OoQ2sQqyz54EB5NQcQP4xFjNV5u/ZrWQWIHLPqVv
IdvnWqDmPQFR7ztCsCg8xqzVDwixR5gyFu/lPzY9gjvBbjEKMjS9UsRjUnYdX0xDMTaFTsuswinM
uxKmUds1Gd8zCrnMSg9oJsQLHLiksjuCy1iCw2HK7kRUxGRXR5SB7tPB3iGjsrpfvmoktGRFNEPc
BIktumNhDPzU4y9EiBieXYiHoalt7CZxvyPjkoevC/YleeAC9HgO/UdwAPt5FzcOeavUrG2pQtSF
1KQLZdW/AjAE7hrUYapZllg7bPEVdppMNndUTGeL8uv+qnbT9lQlWAiPGdDTetetXPLzWbqEfzdS
Yyev8hg7zEHb8lmQR1Y1lVV7p0p0WgWeO7xvvpfrYFBwY0nqU/Uoi/wjI3z7DtQv6l3YlTtSwpSW
Rssmhvh9TJAFZMPEADqP8gXL1Vi98cVuH1uuqBgFzrPOaNT//+8gF30Qu6YK5vZo3YBwwAvekENJ
ixpoS/aLXgRCfz67fPmGcHDskfnrncFOOZwqcOvyO3BF7DyaR75clTDhCiII454NAAKnbO41XOtd
u7rLBTciH993nDcklz+HWhfHOG96gvQmT1WCy9YYnTChfho/snYT0rml552iosSiGRw5ANwJpD9U
3sLwaZGuifC6hnPXOZFXQrbhtivdz5sN4ejdyrgwlH4RbkFddV7IehFE8r0AHP4QD1Sj1rUipa9N
37wPH2/dZe1mYPA25/fndVmoQBN72x2OTuBJsst3FccPVOyEwnA6bmoxRuyzB/E9XY7hGEcW+6Lq
LhxwElOioYj68pGbLGGl8N8OFguVJXttvNED9YoAUXRblfENys/RF+F5nM+lBt23+cqsHfM0KXdK
17/9brmIzp7HY+90YOGQvHQiWAuoeRcw1eLAkwCkkjfUc+x0LEzsFVCQHMf6lXGCjL32WIv+sNHj
+67MEFbUOMuAW3yNUWHEaYabWLoW+TY/RLpQyv7GXg8ZGbw4xoi4Yxu0+uQOk9R1Yuy2Yn1KAihL
t9RAA8bbRCejQ1yveOYkOSzbctf4AwtUThGihZ1JTcxeLPNwi+260wsMW50n5flEp7WxrxtCwbNZ
T0faqRo3EywcBZyNDJD3heMbhAYeCwdpS6qO5m3b2ul3Qq7Vfx/ABufNwg04ExJL6Dzr0DBsz3OQ
AoOGcdwFDE012v2S5JyEMLPSzcUP4MylpU/0FZaQdHlrO0Nu//iCG51XC6wpT92YzW5a91nxpt8h
PNmD1kaXNPVKpthiwbonlpcAMOefcJw7JY8jaUiQDe+KWEyXp2DZL7xXnoj0wSSdprUZJ+0+cUId
+zhbEjUzdPevMf/ugk7xTUXh6dK+H+eWsQeh/n2PlKTSc7NrX/wFt/YbkQvMiTsQCXVkIaevlmfb
Jn/lGiKhR+DQVmAZRvzbrbVuXrEiSRS/VedJYFKmafg7Sbt9PKflaLThmcBGAVTCmN5Xs5vIAunM
3Z0pAHVuHV99VXqJCZyZ4uvwhcsoUzz4jlkXg14+hmO7EOz/SWpDL9r6apBGBsFn9+5WQu09ime5
QIxNICViX77E6HuznUbqLK1s7y8RXqLn9EswoO5gg3E2f0pOBBKPTN5YJBJxeJVdX+wfaLacfO3q
DkEb7Ids7IVwA6TtHshWF3kqpyloaQBAmlbPmqTeCQ6/Glvkhmm4VB58SBVs041iqatfu3Yk1k7I
XYt96un+MiFjYgaQ8NO1zd3WDQlKqP0IiuV2LZesmWRC23iPi9FTfN87Qpx4udf8FC/FszAR8Wgm
ZlT/5qGEu7aCJ/EPU46AtyQrVRygeMkfLRuupyDPEhN+4CTfTfsnEi2ja19zKLvbOVCuCtmmCZNr
PTOiPsgsQpxxQtSQJVbt0g6Vqq0xofa5BgrMJB8UulKTssG618DmI0JjVmmJQZINTNK984M6lUHD
PEursdZh6gI/2iTxJOxS0Pb6DQ0hkZ3UBM/SHdcnsqdn9jUSvbeJqE45KYFBcZUEl/PHRSetPjU5
mcC1eap6nEJv2OQnJAWGbDfazJb41j+mgxA9ZmtZhx3S5tigmkgSU1r6p/3PbHWeTeEtRy0Mdvq+
mMw/I21MkZr6bfuTqHBCUuYB6YJMf2Ji4JELuIXR5Kws+GlUKwkEhZ180AK99z/0yy5BcWllnzet
IXnENp68BADA7xkMR/4bV7zyCK4RVvMOpAE6aaTNMizhwo25ssTlrh9ttz4Mil7sC7Jpg6v2UBQq
6TagX3S0OcglNU+m0vsZ/i1U0E3BZf+1VLYHzfCayxBxhw/zzcws0d1DGdgl5+7BjrEHkzV/d12i
j1wdXulJArX5w3KFtJSW7pIVA7gXy8+tyqHKyt4byVknAlDjNODahnlUUx4gy48R8KBnmfLzBKHW
+288hdn3GrGlevaIyKz8NEE5ueeIaxmE+5vjOCByAuk7lQZj43L91O3x038ClQwiunk9JKKyC5FZ
yjpTflNR8XneuaK1bWgO3izTU4R3A+Bokx/HTab4OCPZwnn2QoInyHRcrW6zAqRHFxquCSVOMFOP
yesqKk4i/VtJ4BhCe2xF0yD7clrC7KnB3LTFYw7iJt4K9j9lVD/ebu4Etv/uweIblQWpcdMBX1e8
z/6pZaQlqUXmH5QfBUOHKhxg3u1HRU5GXWk+AAxDDI2qdmIyFqpwusNFfGDe/DU0VOiUjceZLLmM
KCO83qLCrhGTovXFj1K+Sb002/mYcUpXVeYjtz2+StWgjhJX2QaBxer3e2rNZ7y9i0a+GDyMAsd3
WcHpbXdUyhMXRKASgvJ9Hec67wPSt+p71dWw8+xRgETzJX1b/g/lSK0bO8Izo6ZCW5xI8fLhwLUx
tW2lqCjhn1NOiewMvBGikHw9mDj3R48Ldk32N0ZZVgI2onNs0Ggf+9MAwDLN8hn2niz2J1U0yOJo
a5etEcu1iPV7piU3F5yth8pkCuEenQBX0YF70NYJi550O0BI5pwwZoIaJFst49yfve3rJrQYMPmi
KsTLxYnWqcoZoAtlfXA6VwGcRVz3WREfWsL0ffuL3BxRCzwNP+tsc8j4qyOTdiqMDI/WGW74fXui
s5LCXfHLtA/fDbTi917uTLFggg8VGVlty4bknl+prVV+4u1bOCIfsLbM5KIw0ZBoHh1UDzplKrLh
O+x4ZID1DBP2fP+ldyqWBtxIV8gGvCPbph0ytGDNgUwQCCA4/ue6LCygUP3QcrcSYJ54au9D4NqK
2ih3Z35mC08AjdUKTxKlea3X/OIf9+g4rJIBeNPES8BnFYtr5SwQYFbwjlY9T6aGhuxrHIzMl68o
qF0dBSKVEM36sSVmhgNfILmNyaxVzMsnMTH7Ce+opYef15XcDm1zzm7wC5ROooXh0WyBAybnuplW
ZGr7Krn+S8uEJPoHyrWg89DtATD+cmkUWo1//ZPtHnZ/l8YAqFQ1QuBlh1iztZUNRX8gz4XV+bJm
8lD2Mejg+wo0PvlX119i9+mmBFUvDnaRU6Ugr8adRGz3qxUu9XM46An/b/CspBPb6ISUQKem5fwG
tL77QGI4NPVFlrGkxiJ1Xjq91FruFZEvRA19mFvW/cCP0qXj54zQA5KhgdqVm133dgHf5hb7yAyM
lcp56/XqRtqCaxWb+QYKWslf5FfX/x2/qwd5DEVc8TsQGHg7bRvR/RArz4QF90AsUv0KkZlzl7rD
+USk8hFgugxzhQLC2NNYi8F9mnzfXd31fc8Njr7NBQq6+33thEshHYPiz6lpiTXkVDXseXBjDyLM
FJjJskjHwcTMLvAALfbgwTnWejGl2ypjEJIj+J3lqkV4RI3Kh1K0+/raArnayqI9+bneA8sI8LcH
7wuO9fxlOD6SfXNO2JELax74t1EG3MdOUaQS4ca7CxIvMcTilR2+sHq8ENQGEuT4/1nMl3VuaYX7
fQVErdW3L3fLh4u0zzDaeSRa7pzaJjZYARXpK2KZRTt+cDDRenHeGawZOjP1bJol2Hvl59s6st8z
mQYx2Yf2kmru7g2TKjsp0GCuJr1fE+iMIuea2KLuBFYtZWvbMv+hnuNp1IeYi/LRDK5pZGdykzZO
H+Du8xL8fi2osXyf4wuqcxbadNiVcthRbJJgC2pep0gHavFja3boge+P/UlnxMt7GMCWOOWI9r4A
YahFC/Db8muFzTq3DduIFaY579JFOshM4uj4dyODHhMMKFtE9Y7J7tm++caiyBhBhendgEv6Cpg+
Hnmt5TM0A/6/0bnJGG+o7IeLwWX8XzTKR6SBbokYkfKsWvxQawx6uLptaRwRs2lT6E2ojPz8aWMP
06OP+oTiQ2ZJqxwyGOploaaStzQ6Tzky97hQG2x3raK5wW7OU19hP0zn3RXj64ePPmYxVDfPOc+1
H8qYlNw1WQ8kuy9yKl/xCRt7/NIuhvdnlpylK2WoZOMG0tudx+xuuqA78jduyRn3BkAQzkz210t5
3biZqCteXsWfWE43sDpe2bo0XHyTZI9HWh2NrLZRL4RWHrHrkiXHr3kdoW857rUrYX0MStUTtFoE
YILd+iuEECWeq70yNkyoKehnpuBsHOz+XtzuOaByVskn4vfWVGQu7eedSO9xtIYmosccvacEZnFC
rja4YpkwQDhCNkMY21dSfVd/6Cv6VTjHEfsp93G/Db5RmILQGeFu8EbXYO987uw7fOLcDFs4y6UY
FXzPIGynIJ3KqRo8snuk5X5m522dxoMA1qkHZQ/Ouajq3huxgYQAfLpBmNky6kIh2XK1V1/WWlLu
yt/vU8CAgpkOVq5JP/E1NLCRJwFpgDXmErkDtPNvAxMNnoZgEmFzIt0BnteYxtLvs1riS6bhwbOp
T45ea2jsHvFpDEAsPqMdfkGFEQNjWDHRc3nblaNskX352tWWfq1BpRBDyAFBa4O7JbaCVu7lattP
fSegOJ4S3b+FmjqEAb/e6RZuQHfQCshEChpa+ezy84T+E5GRz87I29n4GZt+G9J/fCzYvtzW0oJo
6Y9r+zGJwJudbcBWdPdd4ZneUQRDiD9lWTadsrxF9OleN3bR4xu6oobRG+4/6JwLfZQxmqgYrR0+
gix4LJfdHRjqnLolMbPv9IWHIdstNSZGfN5Ai3I4gG54pWzrT3Pfe21bB11HRTWwXDAbfLmvxcbk
wjJQsx1Hha4xc+E9lY1kTljLAXJObkfjq1xAPLlD13YlV8IzRvnwg1JRcuPKVdt5SzP6ig/wz7Iz
iiDqLhrX5kCLSJg4TDrMRpvOYbFGMI/zKCn9+EH23/KKGLpH6YBKf3FybkujUE328RQnup0eSfKz
cdA2uksoDTWPb72Fpi0tO1/qJa+iUkEWumX3YnRKYiY8huYt8s42/KpqZSSMyxJVpr97Ev1CntdX
Tpjaq/n4YvUGD/ENJH2gFFl3lLATQElUbE8JauBW5d7mqvrHcbvTuDVVC0lQ0UTtP+lZqUYhEUL+
LEyUGUCGoo9Rp8M5voPhGXQqgtNfu2O6ORmkRmKQEnalpU0mg95Fe807dLyDGtWe4jN+N0tEIuJS
SYFLaImtMxxvGMyxhE4ruKPD+liNjMXfxvdeHvtPx24JbbtoPITVScaEhWPzgU5I3Opp/Sj1kTgs
NiZfOBovpRIVS1lVfC9VkSDOhgKcZO4aH0HEcVrxt9Dw1scutnMr5i/QUXcHHu+EeC/T5Oohihn4
H7yjCYDkRUY+xjHYjD2q5u81SPKB9+zSflHBd4uRUXee2TVhgAHFr52n4jJZLFoUfR4x9rVJHzuK
mSvNbCt2yTIXF7gHV3vNSnG6kph4EXgG9Migyn2TPVR3czI+hP7WXhdC+ehY2esoB09IFFAtzZrr
YI/ts9Ap6RFq0MpbdS7A9tQ7wOZ2XnZ1Je6CkGNKm/WcM/oHjOR9KHgyR/lFUA0bjkc9wAVi8Gzn
xGMxWpUS5MEY8nDtBYEcU38nNNBKbOQA1m/VoWlCCvtz2xxaW9u4x7IuzW0NVjmZ4Fq6UDj6IHUG
ZFMuccGcvx1I+FFLEckkV5YSrVavJ3Xgvg7hsGUC1S4mX43asBV0oDo3ptg8U7sSX9U7m/FCideT
UoVwNg3zPu5ya0i4tjjVMD+mI+XM670BWtpL8naM/IA1r7bTgTH0NtuA1EcJX81f7HMuKxVvZ7Iz
sB10wq5ABeX8Cae+EnoMwRgYhCRRTJrgMO7mDL7IV0s8atTaZqze+9itkHhUS3gtzAss+hLg+9qc
leO6be8Y4H4kcqL+EKu8TOWzQSUIg3ExV4P03n8zx/02cJVkHSOcZ2WKPGwWLULhRjBCLN0JUl3+
54g9DHwyjg6RCTgChJ1OWTnsmR35YcoPZgMfEv9YOCgImPtQap9P5EHKlAncqk/u9RYxeFfK3Jw5
+wS0y6FRPMnZCWtfSHUsDAzN3z5xjp6R1HuiyojHtYbwT9r6m8pizPgk8KBsHhyaM9VFKHYOFvSL
IwDLtvVy6Q7nIkw2ai1vA4JzGwlUkUgRvVQoflif7notL8ljQs3z6KB4jIcMG5E7yVatItCD/91d
WMKzkYl67Zj/yMEcdi/AG8NxUlJeTOnhJBYCpmGgPriB3i0TzjOpIQL5RMHWCmXF5k0LZ5FsyKan
HPeQg2/K1OzQiQ6tk1n9DpZ//NBzb+ycI0IZ9K+ro2BC+2BtZNRTbEOpMocdGGpQitxBXKWq9596
HcRP55Rz4mU7+58Rhk0FFasXiv+2hXtUiZvquWCJ5qODA5RAzjYFb6J6dkORSyn8Trbe8n0eVkD8
vcoTFsxR/oQGu/qkz8kOZ4S27TF5g9ENYEaQshZrETeez3Bu/1WcRjxiQr1PSiMStcNbCDKSGthO
df1lD644dkxC68nhgZh63BL91tAGx2gYLWw1rUUSgW4SEZ5giDD5cHgFTb+H3Y3d5bjp68OaKEst
resyzPZJBdXku5ERhaeo8r3QqwRQjc54WpevBR4uPmYkvsNMgLHoEtHMLIpiwACWr5f7/FZGMgVQ
e6rZmbpRbOxF+4pTpvFMKRQoAONy7eMJ5Z8uWhsoZ9QUuh45l6B4CSpPpoIYV1NCnRaZbaWbygD9
g4GRoDYMsYQgsZPG2Jwk0nin5uvr3yv/VsgmRo11txHwOpRVdV4CWMszumYNiXcw3+HPC4wP/nqF
3LUGtpUBc7Eop8prri/gzp+6FqzOAUm0Vmy8dsPz+/FShjoSsGW84o6xhHkPCeWlAkjByslAkdB+
zYPLMeZsYlvK6zm3HKnE0C8Vx/o3YDC0OamOam159KZ4QYuwg6JyJ0DSrJtzxde8tZ4klbEwBma+
49BLXe5IyOATn7KHKhXddTATQcYFZtdW3N6idz08HipdfR+r1AdOkzhk4WbfKmVbtc0wNaZ5hGVu
xZPbZF6m1Y/19Puje1Lo7M2K/szfEN0sY14Z0m4mvktNDNCCpHe4xlEbxl0Um345G4xNYeP8M/qq
DK4dh//1hOBpeOMbt72KB6h53iplGboS9xit15pf+RORF7m59O/tPu7qZrqB0E8M/dSRA60RwM0i
A8iLQH6DBgdIcNq00FVA4AEI6/rJgxFlRq05o34kB7y0b2Bj4k39xx5tPJ2efd121A19aZOYKV5a
/YQm0jUSr2toDgZSFwvwDo4zj/STF5dxKZfL2XVJPOD7CmNDxEJdqNeuBe9bT5HALCWSh1OH2otA
+F/CDCPagV/cuNjkCU80e5xULVjaPw8iRADN0I5+NA+No/r6Sscglr/uRQS4x10xseKvKwkp20JY
JfJQtMXj7mlu80hpJVtQS6TQM0iaUY/GQFeI15wKykWN5TYj2PbPwk7od7KVGeejRbKgEIEXqlhH
DgtKMP9/6ErTU8T+i91EU9Go8S68tF4ck+EbyYDYuuyxpOM5bOkkbIpdBHC62Ijox8OaTaqKeboT
eK39KFH/vyafozDfXesiGINDFPtULGTSxRtYXFeo56WP4twKobDcZkkP5o6hH9REpguJ8l09y25N
J7Ap7WXbsHAq4apzzWE5yskYridgilN5dvVeK1z/q8zlS1Z2QgqXYNe5F7PYJuo9807HoMCZ5MOM
INGkHfVIJyrNYpWWui8wFSw3ubLXdjTqcfO61wU/nBbLc6QSYZHulF/+mj7H6Or39S61QYL+K3sE
Elq7+2Gf+B8H6Wj5NscWnC6kmKIvYVDzk2a3eyyL0EgRMvkr39fF/dkGimOKSEgvyleK2ru7vFXY
GNeQupQOn8JE2q8ziWwPfOSbrpsIb/mNgV474AjdUF+vx3tetVgvKXXV0aDzX/mi98NFBWD+94Pf
HKO71AxYXkX3Jid4J8fojYBxpwY3uN8CvcJZvwrSD7xfqA8GbgaScCfey3YICf9A1QoOkd6zPyQK
mwT52Oo816tyPChzdVhzuqGBQC+jfpMjW/80Yzjxw8N0+wLqBzA2APLqVh3veEBOjQHAzYVwbg4r
s60ncYOYDj1hbmimMuNE57GJtDgyYn5baxAootAWFwy8ppzomxXC7BXt2Tcpt1x+mI/uRPkH8n98
U5oov9vC4e8KvQAyHZxLgNLNJmjWiKEVbThkY6UFnNgOOIQ8pOIilP3QbwQ7bUkFa6w7NwsaxAnT
x3nIktWUCjbbqQ5Inuir5Pub4o6lk7bOlXxlEpmXOQv8FT/51Vht4ZgtmHNN/TFwWft4RRokHJ8W
yf/OQE2ydbH976/ohn9lyjXmY3JjbovQH6hAcXsi7FOvS8yFcSvoFFsAcFpdpSaSISkcQNKD61wr
TDGRornj5mm+8jUtatGiipQckhRG3zcEQuzfljsTtAK167ydBB2an1bAfkEcCOdEOMPdfC7OaMyG
1nV2aRvLE0mjXu7tyu+EQatT6p8ZCd/dr2WakuAechhLTs6RIWtNeQBJeKt+26nVM6d0R306Nmuz
aTyB3JgMPnoO9UhKsxMmtfIGjhM4NqbbcAgzY8skQAVK8jWpPdeok0kndfYEM7hx4fhFHB9zl3AG
3i+HidJ4OSxPqGb/PBMV/UmMZZPFXXY9cUkfFxJDx5NRvwWIh8A5YNFWMBCFqx05+QDil8J4dReH
o6sd5OoByJjOPtR3MORJJVSxx3DktUPHugkpTAok6Bme9ic90oHJi8gAg7gkZboWGvun67tiYmhN
WovqtVB/nWeErQ0gkNfkyM6pJagPfOkPH2clpgd/dEcBxP7bvuULiCvoiMaTsE743tiWVC0ZCvMG
unIv7sUFLCkLseWyOC3+5dSAc9z25T4nA7JttFNtnatAg2YThHsAR4WQxKseAuYH9R6lsMhjvITv
NOSA4ZI3LE/mAvZ9Fhx6Xykyad32WOvnPqDD8FN1qu4zsRXZQ5eqJ+64Z4ydK/CcIbwMHIPswCff
yQFo5gkf0rZfqfSlr4Deceq1IRGcH/JwQSQhr72sZrQtTopp22VJslTpjDlJ23FQKfP/6KiIeGCc
/WSrqdsqC7IVqAUn5417srwPq1XiSeZi/h6yBE/LNVeS8+3YSiscd/mH1r77aR/uvfKtz3qVKQKD
nCuUb+DNCApjnudao0Iqtk9CYfxDn6BcECoEq9gF7XmTB7lwyOHcln3s/HqovM/HUA0lVGQOIkWb
6DO3c7tcyVaprcT4PjPR9e1h8GEYS2tcxmtZwm4MZXreGZcKYvZR4Z91c7p60I5N9sreEPDuiu8h
FZ3c9eO3lyBsCJJBFHsNC4lIenABPYUVnjQ8FntUvDUajP1DOPNvfaprLokYUMfg9vajSPL0wWyC
lKT7WAiF8kH1F4JT6lb1GmtPFbNsCys3xqYCua7kthnf1xYq+ckimsXM7dFh/aODtCUly+bWnd7I
/lb6sGN+uvUduiSh4gmpjHPzsNqMAq79+hg2TKiO6cT9SaRSjWu0ZLkyoIe+tvcX6jQWrPigZl8r
Xi59tV/nL1v4IXmpYWSMk9QMhUyigFyXDcWf81kO8sdHILkmYrynlTbVvjVCLGoO8yLyDFai1CWk
qeT9CqbA/5AGEBWW70Louoye6C1BPa++N7VVF0HeCsZJa/0hzsnhfaHoHCWRRcXEqWMO7M5Xpo7m
UTl+md8dOUI9ytrHZBD/CajrSft2eCBwHaBh+NHmHV8S8I/KQuaJFD5ruZos0bTqYdybziiGow2d
0T01ZXKxpDGcNPaa9vDGxxpqgQlZlQT+r+64V1Nd/5bT1/3lc1pERXvOj5x68kT7RZ6Ki967Qq/3
ZvLyPysePI9ZR+Z+RZVhKYMU8psBWKLxHtmoi86L2Z8Qf5QuJP1Xye38j3nE11YBf0tyydIdSWuh
Cr+j10RXq7GmgyHJ1XUhBoYbRWAGT6mkjh9bQ8fVeBS8BPVAeicg8oF/vJ9pFOiuyDfzq6N6vEcI
DmXE18llCOQfIUotLNsC+1Y95WjY+sSRl5IJFz7DhFOr0ubod/FOjT5/U8nIAzbePm/lHL9Md3hF
4nLvFEGNkyxTpnHr0PW7Ivytj8Dwpo7oJIA2ie8O2f25Hb9d08Uqvo4a/HJa5Qw84ndkiRHp5CSn
qzJgi5WzEbAeZ5UmSfGSu4ASwhspk374PuzPB3Y6sxGAtdcwVLAcrT14L7tStopU0H0dT50xZG6x
GSxIMXpL//VtjsgaMuFijxblF1nsI4NX2SJ9alDdgbZ8PXD9l2ekm1rPmNznGYzxAKExOHZMhbHm
MACM356jwlOIDIkjU6pFd0FPqTqBEQHbslap5wO+nbo2i4x7bY9FDLGrrN1FB7wYQa0RrqXEiqNH
P/PeMHnp1xf4mekaDJCPetsK0l5lpYGJRu4+dskM92/3sIzbKyQO1pBlV4jSTT9XcQJT6MOGgVGj
7Cg4ltBsedt32wYC8KVM2wvgkbkeANWHBTMhtk9RA8nBqc4hGkKSExF6Mon0yBHQRqX2v4eIG8/5
2S1vADBtRpaRiwDkOeHk5RDNU7yyMsKDCPwdbkO91QHc51KL9NFcwhLqUROqrO6Pa6d0EOPotqyN
43GFKyyQmlzAgNSWbO7nkxiuFWuKo79wXLyBkDne5XBed3UIC+WIDNuXSdLpVBxrIXFm1/MtHND/
z7WkHpEZhwp+i9UTgMoCOfYINsNMHuh7kH964dBABgA9okD5fYjuD8qfW7VsYQ51YUZZphODJJWL
Nwj8KciqePYoaPQvacDxXWjS4cP/KpLPNNsMARDCuRqRRWKIdeYEZSEO7UfJ7GL9B2agv9u4GZyx
Yt6BsYW44378FFf/2gwXZd7qnNpAua/CZyznvjaLnVWrQpznRU0Gb/Z0VolxFmqufKI5QPRlCi+Z
4GDDfQ1+fDDXinpYK0i4ka4xLIcxogAWpm2xSEw7grMFJQ2X6q45MbNhPvVGpDpW7g9Z79RwYeFn
uKGqzdKYWnNFvm2hgT2Jn50iRtzJHlGfXclixT3P4TYgw7zp6ZMu4uvdUCpAg+r8JqCv/fBOX5nS
8c/1Z8JBU7O97Kb1NWLwf5jzJ5hyyZ07/ggfQSUNKwVBXVkvLogmG+8MFLnvELFBpzCK4wBPCJPZ
seVR5YGHB/2wsrW1yrV616HfwFSOyhzUhCAXF4Z2KJPi2rgJL6u8Ntxi36fjzUSwffOHLmYfdD9p
qDjfDdtHjgIpwN4fNrVMQphBOfBVC9geq4DSOvsiNqS5i/rULmAf2SvE6zsnpEyXlOoFQpBEHSlt
Z+rFgrOAuUexk3vmP1mV5pyFpCH/4PVVjPO06NT1v/+l3pfYRyNALdLR6B7vtyPTdL9Gq4nth0Vy
vrg17uqMLhHSgk99MEecxtelgRsHkEMr0xuqhwwTegS6wTe/mPDvPfAQ02YtRZEdIm5ZBa/f4JwO
2C21wvjdYIiShx3hifXMlowZnXO7qPOihvedC6jL3Zz3ewga3miOVYx7XaA0AltqH7Tq3GTaD3u7
/k3xU3UuLaz+0iJrG2/9iJNJDneJSc/lvESNDcEpglokctmIcE25ZW3mhoZgvFODcPXJyg5n/b1/
BiAKf3dv7OCE5uKWpDh32elxMLLIpAv2dNJVDq4MiPKwgDoC6uQEsn9E8avkAAmPV6m/sEV4h4oP
ycqJIq81WW+RhxJfQro09TNvhPdWcJDByLDSO1qvi8w28FVKSbgm1yxFDRSbc0z0GWPGVhNVXcgE
4d0+2Vf0uCEi4Hwfaex7qYYw9Q0BEEGenAEV6kO5iN8uE6VqhRO5KbCirE2myFNgcaPywUb+QvOl
lzKLPaT8xG2+ayrEzS6+KhNrqeaSFlxAtf+/dh6LRbwHnOJ9F9uoOfaWRz/XhaQqxmiS8hF95BVp
gIMuVTVXRQKRSEH+uVXMwEglMQ4pMV2LJWEMbF+CeGISxNWdvZAhQy+YU+6AC8JaeGNoKMQHOBeQ
T4jNyFjQeGTFAeU/kkjcMwEeHueF5iOWt3p5mO3QSQ/QL+bdgnW63lbrnrEhzpmEv3YyUj7SG++q
oucc01q0QELF/j4lV/iYUYTidl4s4wGW9tiTkycnGrCOPfd8lpBSoF4F8Z4hvIPslVRtAezn0SWp
mFbR0PJZrF+tx5ik6v70R8/Cc+v/KXnIhqtzSwgN2cXVuYiW0LMo+0LCNJH/71FKJ8UyBGjge8FG
aGBpNgVEOqdcrencTd6J8lgNBhX5Kg8CeJK0seL6blys0heDF4HGjgVoxxfcD1Ai3xQKdExgICYD
HmtqXhFpiMDHhlsVVfnywFVe+fsXD0DxqAlbR/venLs6lT/pz8YLMfu6NK0/bAtYJI4bzgMKqMnQ
AE0RJ7PY0rpKRTKimz1jmXe+qseRyzWBKetaQAIQyQYObMM64y8V+A7EFqDV5ZC4DuTC1vxfh7Bk
z8kMFDgxHdOu0zjNpNPCkMEBi3DczmUXctV3MOpzwBxpKyuMMEgjfW//sxi+pEVNUGxpHyWuDAky
/6fFmF9BZwWt8TpUv9Yfi4ZKoGUGONWFD2W/V55D8oJjXUPdkFfUwohcINl9LLOD0FtnGHE6QnlN
2/+M/TdKVPXoMO5/qTlFEZkHY6QCnnpHYVURM1dKrxnEfhRncTRQ5MwHG+fg34dVhAfeePSWOGV9
p83WH+f+DAU6Jds3D8zYRyX89TRRlxO4W6tmIV/G1dntd6KHsgqDO7Cu67m6i8kgceKmF2iMsEQP
K87Rg6Kmk3JTGdc2M1Vzj/t870AsqgLTDCelpi/7VPy3i/3TnL+rIUivrHpQaadWCcbUMj+iofRx
UI9ejEoixqsLXcR5YTyvIB/cmCeHe0NWIzwFX7mxokJ3xr22os9jjQbdwPFvyvaOm9J1V2HAZaAl
avIR5F/63LlUCgL03FXM0i2sUDR727Sp5BkXjksxX0sylTlt2zRSMHYpHSnI996Sv1hP9detE9Hd
rIiqzniMsDKAnrJfXYobgq2MgHbYr9QkQ1Gl3W3ps/YB9f6iaV6Dlu3BCbHVn1YzaVDEbumcmcdG
Z1vcU0hq5u7WkgWiZxr1Pe+l6E8p7ukgTzQH8OYD7K8iDxtdFipy/MCvlJClnVRaWQj+7C3tL/Fa
7o8ZcmvQ7OvHbbEcEQXbJwNfZnCXk4RPrKfznCaVSGmqsFtRwuWqMpxVFZ6rgcY+GUqGifmddqmr
KskoPilZxAysK0u8idcHEWuPhLHbppAQiMqRuZxCbyM3YGq+r+IpWavebujboLfSkrJAgvXmeltu
iivQgFlbiQcEoL5G2/blf9C0P8rotvklaq9X5VCJFqgmMQn6b6t20Z0ksHAVTmWWbQhE/KGQTEvM
LN9+cRJBdHQHkNdrqytTC9v54oVL22AEenboc3UswErYWVmDW0D2Pq5VS4LdgZvZy7ioaJ/ou0nX
iiIYKj3Fg9tXYrRnFoDCH4Xx2QhirkYq3BNZb9nGvMOv5VWOD1KG+Ra8VjZygeG7pqse8algVify
VPRe06s8HJ4j7cEffh71dtf5LbDnT/wAmfPNuxnJklR0TxHM0mpR+pXyNhJ5GqzQRSBQ4xZH0G/8
gacjyt7KqjIkQiNuXW2gTMF/0XPUkd5OTHxkzEBsiHh4yKm7/5Hvx4uayTtyv2gcLBnMBjkS5920
3jwlgsX51LtFwCjf51d5vpKV4exF17Ml6k0lly5FEgIBxhN/pPnL3eG3zXp7epIC7sjR7IBG/mUk
uGb1/wG0aq7IiObA93fNFIfHMpBl+rbyKEjQbEfXpDyLnoSKRTMrVpYjWYhGNfnbjBOkDLaf3fyp
9lPj3wxnMfkicS6WAmgdB0ufcK6YEVbm3ZF5x1zQfzY6QnTxeMoKfTDr+kqFpErq+1XWrACFJbUG
kbzB3A8XMu7vLKOYx1eatI3Ntd1LpY0E/8AeRueWJc0Y8rMWeePuXY8clDT7zbgJFAeTOODvsoaF
9oIEO6R3I0ymPTQgJz72Z2DE1o4BPhgLhXpnWqj2KRTjRcW5vr+b+k1EZ6nxCi5yulGZamyqUZcc
LuXTGjRQKzJSE6Y4I15pRFuupaH3aJVkHpCU5u1kivtshL0Ja5qzEk3HaZEOGbxjAK2qs0tFtffH
igBcNKkMx2bD3+z1YbO8KPUz2H8kMZqkEF1wnhfxNDVBC7vmXRkPSA7Sj/U1yDy4WZaauti/hBzK
FAR/cvo5dSFFRciPOywODoEzDqFGH+nW2IzsIIGkBDJIb3tq49iwCu35IK9KhR/XfU3GXri42a9o
+jcFQi+TSx1YfZOWmHm1nNIDHqJrXjGe2EPCCkrx10PNjxuD321/wgTlRoeX+LzZmAzBVyR/C7Qb
xsRnf46OCPWWoPbmkoQQfqo4VwhnL+c8TrUklZXroDttZT8i4hPPg7uCdoEdB376k1FNqjXtCTJs
v5i3Tn62ZpnJRve88XzOzl5h2RPyzuVx39Btjn/DLOlm6T8oiq5p8346nyd8nxjAYem3KfcwxXdZ
sSJej20ivpc26l6IGIsh+/HNBfZ1MVELCDAV4uH35L19R6YCM8wj36RZjVlGZstIf54WL0meNiT0
fumHWe/AEToNYGbZPgvcQjZjLMeaXed75CVPm7kkol9qJxHxQFVN4mBdPbCkHDuX9m49dJGTUXK+
rZopId25fGHEtIVH8YvZv8l6m/idz3mJsv9/jgsa1X5dS1TF7/6flB1bTEDPg3Ms0I+7fBkOHp2e
mnySsoftFfaAHWCfQplcirpJuB42zfHempIrKI04YKS9lKSxPFT2Tyf55JOlc+TEb5PjvUgS0FSm
c694b1beTNOJAAXx24kEiXmP9TwWrvecuhAlhU7bW+Fk7twRvTg8y9O55ZDKO+jmVmI2ddMqWkXn
Xw26eqjObku2Q0HIddWR8SI2SoBHPnS6aRE0d4Yn6/KBxnjbg1Ab1HK4AYXlhbct3+i2qQGpti8Z
zXcpHPRPK95Pyds8Qd4RurgEn1qVqhjBxp8eSZ5QBBLJGYGeIMxHX53cBt43LtManbX9hLMF3mCQ
dzibSW/HTS0ItdjP01I8n/+iLYofbllQAyhpKfsgpWmd7jmJk5FE8Nf3oJUaq1e4poDjnPH7CVGG
EVGq/G97LjznpgmPzY85mLmUXaXAKssQcS4JEhya0KGWFSujCkQcJAV4QwmUn8jtvjv4j2uVDqCO
xwwolPVraf8p46cGVU0lKhXOi3Nqx29pCau++U4RfkW1kA4fO/zhBAUQ6xCtangAHtqz0Ci2cNfK
uOXVLEGeABEDQToxt/zpHzHKFnSUz9mO6N4UcW/I1X8yk1jkBHDXcjEhnne5HxnjSPp5uva4Hdf0
K5ZeZrmo0GbwozXMxGIZ6+vvkUlQbRfNFkKUuXTSaAZtNQZyNcI8q3JRJDjK0R+YRgR3Zj4w89OY
6K3GT6TOX6R30QjUTjxXGZWguoIeMWwhKpJoJPPT++hEPpccEERNpexqoY4n7pnHTt1udMz4nAZm
tOCPbnIJWGdHRKmtYV15dnPyvHR30jUhiGN9nl2hZWs53jRy6KamOCDZP38SL05POma3b6loSpT+
IplzBiP846toNEaclJ0bNeSDiVUOXlsaRM949CPRR8ytk9hYbHQ1WI4n61D6ZQgLp0qABPIttQi+
Jc1vQyj/0OCLVTp+BksalFQxpCtflDKrA1N/Q3SItKXJpHOPgyPbVpOocKBzMnkQeAuc/2chMgvG
z7QqHTDjpAR4zUhavmLDNoK6OiHHuz+yFfPUQxgcIzKGVzWmimhZQVuM5Byq/7BkqVgKJ7UQ8m/N
Ou/e/+1N/6Fh6mULXfbUH9mpn4RFYdGW1lMvYrcOEFpeyLcPODNxyYsT6AMYWEVPQm73ZRM2nqQX
I7mcWusKPumMiHYebz0dmjgV0zmOlmMlYO9Tjy1W5QGbugNbYj3VRFvAmXg3P56+pO3+mGWJpAaI
wyNWt/hu57H+nGuV2OJANvF25x5kZd9bf/eyNs5BeEAlOiHqq6bduhA6SS5Xo0V97E4CrEN/+psL
4jiS6hTG5jcp5LbfFDqMlwB4+CazOvMuY1G3iBW2vXWPRPywaj8Z1QXVZBgI3rsGFvhkr6QX9zJj
EcUea0W3zZe2mnQSZkXamw7PfHIRuQylT+ycXauWCeY3YCi0DWnitX9FQ2Qjb6+4t0nQ8p0iW0DY
1wWF2eODo6U2OtOmfjdMB7c5Sht1yseN3fr0I58QGNa0QMYNHQxGDRIc7JknQqd4pgOC8xN3pzFf
5wmj7EFqzUV394bQ4ZT5n5yKDBHw4PUYW+qvxtyOvD/MmAzsalt33eHorkruZSKS9n5ZFcaiFLjR
FDYpVuqp2aM9wq4iP2eL7NAl2uiJ/XGeT7mgegdFzgEHOBz34v6lSL9CqCNrP4kToaAFmRtdGLqR
2vnCDv/ZzjBNuBUJsAU9v7+sjOeZw49nx4qkgGArB5oQNLihetyY/LtwbAqxPRGAmMMFcQmall4A
ZPSLY6rNV+IZ9yfrsSUdx8qPVZ8JgxKtAGedFiTkmljLCu1k8G9hmIPlKPkD4mq5e5PjW7PF87GI
IfUegm1p2GXMB2xct+wWYGDem3r7e97W6Z8/NqJJZjyATfAfVygXUem9gRdLyv9hs365Ad7IhLZa
xmeXm0hgAc5+Dl3eSxtaNb821oD8ChTME6Zqr9D2vlFuzS+2HycclRs/Qp5UM5OjJvdV2KnkA3Ma
xocc51v21ErQn8OkFmJw7pvkEMUxuWfzzFSZoFPx68bqo4BssX8XKDOGfnwyp3clXJ5KwWzQbKtm
jP0kCb3mtuzgMWuZgI/I1+o+NEQCYd50EdukC/QSV3VbCMV9GWolG+bjklQpMcQbPabEFuQ8kau/
walrxf/sZgAbKHrBgJFRDtkRS1lraqBDz7HF2JNi2rSC9oZnql+LUxMNiKW1czCaxFr8Xm4O1/Pn
vNuEHS1iA4AqZ2Y7zMGXbxM3YjkKPiaGtagq383d5jBVo6ZHMcbDc+IriPF33m1gNzviwDJZqPAL
mZxrd2KryFqO5lDpwU2yNzUb8XN5q8NOAtmiYwnZcPv6HOb56X7R4JaVZZ8PYHeuFVVEvHTEp40t
vlC8lA1KACTYWG0h2/ORBL3CuPS7ZyH1RyFlXi/Tuj6nQrF7SaGH4ZdjmyNFmBbFxqnKJNezYzvD
ak96T4nN8qJ1clUVck58XcMzX7aupH3PPFrwplQ5JMImR6ZCEwCHB0hibdHSCYYO901nGe6EiQBl
6tISeA30oIMC04f2ITUAwvpjb4nAIdttMfoUSnhs8zZuWmuqZcD/u6yZ7PXRYyXc/8OGcty5jikE
aEMAKB+SVUL5xjxs6GFtIh3lImteMCwQSo7st1AlJACHwuQDQN4dyBd4t2DBNB011zgzAcYloK/f
PvNT5v1DPziUhxpTjKxfSGQFvY60Tj8fFv9xplMogr21FCX8LBGoVsRq+Mh6SvDFdciDOWnAjHNI
GGgC9EHRAbSw9zKdZmcft5sfBMz/2VFESj3F+0WjSqzVxH9TkEGq6hnGlZX1Yyjy01pCqp46mtLL
C7Lq1JSsBifmlJjwqyGTWEluonGQeOIZFVVuhz8Gxwl0drxZuEBH1lciEGUDaUnFFt4PUGfFVW58
hIoFpPKnARhpvcr9PrD7BnDRFUeRLryCj1NsRzOqIa9hSR0V1qFvK6iF0MaqdacGEa2z3FEDY188
InyWtuDA5IuBL1AtQLs2oPzYV5/eVbomU+wZyrAwa7ZubxaZJQYWwCO1x5v2qktbn78CaVJhtnuP
YblYmJoh2XOrWihhJraJ7qEFngVT+ek7ENPpwcBt7b3nfWA65+IV2fNJWX9YjnVoSp4zttu85qiA
gFUVK3mvcix6dILPJYJM4pUlIHQCkaQUdVoF99X2CA/TK5ujALWmnIZKgBknPYu8Jvwy0U2CpzCp
JSZKLyLWGmUP8JX6uEprl5X7aIpwGrYp+sLGReo8vk4PnpBYhIoD4SquBFgA8gq2J9Vy4T/ADnSS
1P9fpAGFhPZsZ1qQ93lyGb9+uzpwO4vL3SysG1NLxse7AQoCe4drE7xkCiY9dpC+immY9FQ5v6rA
WNM945L56IVdipd0T/WzPOWjjM7s8vIhlPSR/neQnRdfLQ4VR04uKxd8HeVKKapCbeQ3ROpz6F8H
Z1t8iSXBUOIZhA+ol/5D0SsuEkc2I/o8eQpZ3FWp443EZNDCt2hZsx+MDPBwOvkdfcas7KioBjO3
K9dWwZnvzqJutxZR1azMbfcs+thxEdVMbR4Uy6upP4FaXsbaO/GRAQhivHLAR7MPyjU+BxOLN/fT
Nl9InKk9roqKekNJwmN/458zheEJiuV9g8Q60g5mejQN+4+CGGF1kHUm2x0N6O5akEmY+bcGuxra
Y/Nads0J+nC4MCONCw+rZKrTZUNo5/s/sb820+ArLOp3TiOJUu/KXd5l5okp7J8yYvrp9GiH92IU
l9TtEdtxZAMLDUuv4kG81M3YdpeZRxz/LigMx6zkyNgMMTdvlPIl7vcbFD7gjHP/kHNfH3Y3lepK
Oj9T2Dv8ZbIKA+nOAsnqZM2mRN1/tO511NKUCVqaBujA6Y/VKwHXQXwmxDgqDBAaEohVAr9Hyo+7
D0qSVq9b4kKBlhUNO3iVUZLehVn3RW4JrCfKZCt6HrVmeY2DCiQwkEli2/+rK/hbBBm+KXodq8fR
oeTl3qXHl3yFMlu2rZ4gaA3ZPUbzDu0PmG2R0MMx66XbDcXIX0H6074T9IGKpBfA5ZdahcxUgEZS
rLXuNS8RyKSuNEfP4dgfqEZzsL4XTu53La0u3wCfwG49+5MjEDkeDGMEqrc+dgzNw+q6QePs2XhW
82uEGX7biA4kMwpFEIusWg5fU5pFEGuBF4+RebwXuHEUGpfMx5Mjzfplt0t7u/zp4+U6UQo4iFVf
8/SBP3+vt/wSHESlpqXEK2yxBuEAicsdWR9CsTjfhqDV1JwmsTBlUebele028x1OPHqA6+jJMnuT
kV3xoyoj3CeY5GFxjbhsMcScwo51gKYI9kw75zvsZdryMwL5oZ/gUbCEC6dL/O6dFjP+1p1MXndL
KbEBzDRyAiP7PcHi2ePdlTWqT5LcvSCY7fM/Dr27jI2O4xoyFiZ5AFjtEFmDq/MTnSqIO/qOVwBD
pGg9/xpmD4L95nZacpLQG9XfxEA9XqDbiQA1ipQQz3Q60R+nelM4qnElvZalaShfB+w9StrLgvQQ
hcpjWVfB7dyTZSABVAXOHLVvA+gEmUCmdYSeWAK29E7keAWyzSRlq1nj1C/Ojkycd7xVgUQsF3BA
UEK8yJX/FkxZ5xOpUJnyxbxEghZ4sllwiPQAGqh2wihJ2kexYI35evxSDBlX8shIkoeLHd10Quv9
RAv1cB5N0uQdrzotCnGiWlfQ7mB/33boduiuxMlMw3aSxv7MGu/ky5NA5nrj11vyGEe7QGbhdnFJ
3yq9uYMTcEk89kng6OOLH/FouL2Ta6iJffIIwNsUiV9igkgif1wO9yxIjrExh8AXIi4HqPKq9fap
8dBN1DhDoRhFEVL1vFYFQZmw75e2AXqG9qNaXmpzCdVwXkImT0fTxOZ7qBP28CArQ2WWqZm+wQcB
YmxL7+Wi9FvVsv/ist0LpRh7fpdKn3loka8iMGYQuxxJltC9H8FxgQzoI4A9g8UFfnNtgNL1HVBX
H4WLOfL88HkeAyN3RmCLXi6ROUDsNo+a03LaEGSBbnuVyb/UjIyvR7Zwo39pAPL2NSWWLO6cwGSl
8Dt6m54xqXg+TuWHFvgYjOoGHKlqKV4v8obecZmlpalUMVII9z+HZuI9R7cebXpiYmvSaB5L6+Ev
2JsZ6FfaFdDlNCEo2LLeA8utOhmdXdHxxpJawCZ6oafa9K7TIiqunr6WrIQBXoW5DuRD0U2wdnTn
L/DvQS2OndWj6m3eDhntrrZDp3CgPvR3EiqZmNqimwovBqdUKW1nZZ6HS4kujQY37/B/l3r3CRIq
dydO+PY5ftoF/Cg/QRPUqig7M0fnZFr8xkg2RhJOx/Gam5xBvDaqApLHsPMAOYgSWPk65UPPNuQe
qJ0TdH9tLZgDqhyQrra3ih7wBjFXDfUPB+5lIy/68w1rCLZIAsRmBm3xDq8W2Fup0RmljFZys1T3
LAoaNHJYYIzcn7eesVFaVOrKDPYNiBd62o+eMqWBkGiocG3i2dQDryGXomOr/LTnh380WLIggFoC
AYro3XKlGDgYb+N8MC7ZFxNDfHYNX81M33P0Vo1xDcIeJk0JWOqUst09wxp78zvrcejDc4/TXVul
9W1pWGze/kveWbtwrPc86Wc7AHdqCi4/CsP/sJo9d9wSTWthCaYwilN0LOuvBg39cSOn9FuQsDTQ
iXgdi5if259o9LdUpm1Hj1bVmtQi1TdbD6Q5t7bWqIB6SuCCJMJYqiZIs5cpqgR1vAu+7yH3/ojP
CurXECb/SGpM9ciYIq+/UALYKEXel4x/jnxjZcV/vu2x9LQO45+MbZNQpvufOgWTurzYsiuH7t1U
4A6hhGWqnRCT2zMeSywyA+kWizl3odwdYhVCkW87YzeYG552g0BbptjijMlxNNqHLOW1FW9v62xh
w1ajdZI0YwfchvY2BnGgxmoxObkp4p+ZjWeY56sjJ1L/Vy47FT2pA4yiB62QpaCFQ21mF/5Md+XE
aexorxQHsMpRo0rZqiFN1yZAwRIruI2tsOx8TshujZQ6MqQL1uE5/gEHBn9dP755CD/sXgdtovCN
Mdvsig4QpdMDes041oUjp1qj0id90s7XqqUEzaKvRM1cHoz3CLydAm6yksmzC/k37xU4onar3CWz
7Dzim3rt/FqVcqE4wSozJY6CepP4PtDecl7/TYxoqUbxbalX9Uz3xr7spp4JeYK7sCDdFhX909g9
1oUwcphYyr/T40z7cRHy7Wd3tysyEqXFVCSMFue1Kkv/e1SL0xmu9OGdl3Ol/n5KefyrheoVXNwn
PxNK6VJHPaknBuWUhypcirNiG4ZigqJeLki5aGbKRN8IoD6VtU5InoMSE7rFLocwKa6sDK98AITz
FTq3jwE/35EeL40BX5r91pj5J8OWr+xUjNtPQTDyBY0zMCyk5L4v3ynv+X6FmRkM+FFiYvkiW82M
5lfJoAm7WIlwjCglXJ0AicWL1PM6z2qXkwiGJg7i5qNuWV6fXEL1XGjfI8oXbkV+fZpJd/szSmt5
MkEzDv06NHhdb84aP9jOguX3fcG+lVbWs7OcZtmdwGedxqWMC4hheIXeEmG9knlXwaEQHo09wzTw
6qScdCMXCyxBQjy97PblsPOOuduz78h1+jqk+sbQnSzsyYkNdCUJ7i1mg67/xNO5EhcaNJV4VM1b
DkGWM8J37/1KcqMtqd5ZOXLMCVO80GcqjtOhryJY3bgNwgg4PuCadwkz+jYuAZuu01p9xjDLb8YV
sxo3pvh5TGUUYc5Eqtbq9VKSM8evrQdrqrFyLwFTpNmcgVKhpg6Cfw4fQpr/FxFDMJLdWZEe/t4O
AG8wBIH0cUe/dF+BYHjM9akOItz54pMzgQc/UAKY1AmXHPGVLpmpouoq1iSs8xa929BYuveYu3wv
sQMdjSbidi4+Nuy2v43LnKV0RonC4rXXaf0BQIib9KcSqGEPzHw+yPOvCvUlG0TLp7q9WG7ujjrG
JJh9OdNMz0YjPKSBenUmgfBw1LvzSBkZolQu1f1vrCtW5BrzY+fheLyBY4VigrSzl/iTLl9dkqfR
zPQ2/BY3c/Ej8o6hlfmKMrwZO8794jpb0Aa4c6J0A7h/A4dgowW6PW5bnnXowT+YkZ7IE6lgHcF3
ytNXELp0YI1toxustd7Z+RdCLtRWNYkdv47PmjGxMJBXeX0Nigzzf0s5FgrmFsd7FMct+jyfbMIN
h5lUz356cj9gvAXI8Xd48qd3dv5Pq+OuDzkqeV/CBIbyWtOpz3RWHVSLmFBfSbbbjfzKAhfR9DaM
bokrgHR5p+ZYHowg1EK/D3SJHbUGJiBOADumHUbABe/XhPKF8OI2tWdgLqvFKq1piJMZr44UvhZw
xEgR2yRIYF63r96k0INOeT0p5TBgFHenBF28OY6TyLkdfYLEXRO7fV04zdG70mCGpvyLzLiYZJGE
Y3Gx9L5T3nlmOOW19hO5DIzKN6U+5hSMGK8QoXC7FZQkp2xvd5FU79fOQUajIK+5uala71bHvQNq
fMhBotWP6DOXUP11nwFlKM3/dpqQhacB1wz+KsQsCUUKkDGDjCd1GgR0zGBF1snc2mVFTiyHWdaT
5lQ3419E4SX2++NzdrJzrVKzaHOw/PWu9F3YUpZZrGAFPWIFc1eWvzUU7QCXebSGESk1hsIt2LWG
45fn5lnGFM42R14lI1PjHqdCmxJTjaItmgK5rEFco7lkjdgwviYEU7jNA1sU6stQYxkWoGEr3YIz
QKu/fbU4BX8x4QA9Kv31MCnxlsWoi14DzQYYGp8cP31AuG1//ncSWl5iMoIohymnGMtka+IBIUOp
6rkCJLL3CyRARoAbwXOiWANx+lJnlUQGYRXbwP9mSyJ2pQVJzRABjVemLWfVLVD9dhsOOBJHD3R6
GMhau485PEue6naXD+3fGtf9fD0Bq3xMayFUbyml6i0p8oa66YzHl3zZf88A4LeBvIjJOE9MGRLk
ul0DvAmiZcSjuBBQYWk3eQIgfo2vBDFKtJcF3uL4DqlkE/oWujiiEC8OOaf+eYZ6rPBUmm9gxuUk
r7ziGr0Zbpbtm97qLNqgxzYAu+Uke5qqG8Ersq2GB/c9zK7ShnJkz5s2d7C0oM3rJfut5fF/W3G0
v83d00PILTZ3/0v3kncaXOvciXcSTdLEf+u5tlHOtjicCB13TK8xb487a3RGckrsIWoitqkhvxwu
q8FhhgAbxg9YyyF4nJ5zkpm5JC5m+HgY43wLeKQmTrmF0XKprr038oyImI3wEoaTSQxsYQsNVPTO
SHnCv0IZNctTuWwea12/yL1fn+G1VbPaicln0N9KVeAsuhwYVcLxgizkYIuw+ssyTFJfOsooDo/D
U2zKCMV/puA+UxCYosxQB3xkLG6opwUv80OO/8OxjTceFtnvb4asgiXWAVJHr0S/dznSXYDusclh
rbZuqGCrDpB3SgEH4pR0gLeVEZrCPVAgti+0C77GTP5/tMhg4oVkwO7QFg+b6DlqStZTFh44AzLm
TEsZZirtSMrlRwdGaWV7//thaQXN51Pj/OmCXr2T3ereuTfregBZk9v+P0fbe6vtFzyMG1KQrdAX
wdkBqqwCjEU8HTuaSm90kemmxgNljaLrRglWidCqKnn5bmfxIsaSSPtrWYjipGq3+8KPB+TuiRM6
fdiwMCwSChS3IyAUA9NATEDUt5zQlf6Vbg4B1zkUyWy6HpYJNMeP/NZragPux1qo54zOMpDVw9Bw
PznNEtAmWQJ7ZgHVJ92yMoBbVWM8XY+nduffLxccNkXst/IaCXC6Hs04+g9nXu9YxeBFbsz4kuos
lffrMbnZtCAxOf3HqC4Y9al3Dl9Rs85ZW1345At1uCRWnvnI4Yb2UecGjZSGJcAnryVkTFpd9nAg
thWo5Rr6yQEft4HzYxHyKLjxbabqKSHX1BP/iX9nXkiZXBPgjhAoX0l2mLWJQnm1BND+ZWWh28ED
upd+htnIpOsX42Yu9pe31L5twVhDMYI50bsxf7jJw+S5Fpd48iqNK6QnOZAqC5TuvJPFEfYn86LR
6EVZLLPgFFiSL8WuGKpfxk+52qHWw7dHWf2zoxSV+vDO5pGrooQvcNmwAHl6iXydNGvxUlqpt0cs
4+C/VidT0+aSIZqbrELzY0dzHFmy47pKwV1fJ0jXptj/4GmXwLKdd/qyByWBAtk6S+sILtciqaX4
lFvE96p2wbIqzcnSFK970/y11YgyDhSMrfCWxKldiZjQgO3GtqTx6cVHl1ryPJfVbK3BPZI67Q06
iiGFS3f0tezP9897PI5upC/HlyE+aLN/DC/qAqVOE6OUpbwI6xuTcc7+dsAa4TzPINMO65hzU57f
vozwCrkqYo5hz62AQOjLby08Z/7Izkv5XiZiulAnhTWmwiQlER93jkfxp4R1rQpVrGt/MjCUohyU
a/fOCilLQh3DVZ8K/54JmAWJleEfmWTndYzuiDfbHEvhobuoUGRNALM2r/X5hckuTUG+ada/HjMX
XPBPMffIsUkTlCW3ZKGacwEcN+ovDrfbteUYZozIHoKP+/WuXLkFaawBAd61IWrCQZsSNh9hL1+Q
ViyWCIrxpzrsDHoBaGUxrCqDkLdpCvrjs+aZnRoCuzgUqpTfZ43WnBVENG69W7K0a4xVuAE6FC6V
Ycx7sqxRi0ByuBkwcVBr2XtKyRABIMjxWycgqsR/kqV/56BVLxAwnp8I7Mnqz+2sUhxygvS6sCCn
BCTFy0E9TsXtLTCbOzZfq6m7PYTTV2OF2h4YO5h4/2YThLwIE4Pq6xbwtaa7Nd1PFeIXQ61WvFhV
4VrGljFSX9RQ5jwbsBR4yv5/SrcGSfbEe20nn1PMz+JPXuxCGJZPxhsmM7jTwNGKkDTYlodyIaJG
hFzIl8fTKrKFE6FJI6mCEjoy6hoQEunOZczbmJHW1PPuWAj5Z7JQnN551Qi9Q26wPIJ7rDY9hOmF
IN+qn7JquUmEzYeoM1oJs47n4BSSNSMGVZuB+Bt+s7V/pUvHq3NJugHpZzwFkkOf+Oelt4WSuvez
mRc+zEuNx1BCrhnEOrLp6Zb3zRjDigZQdWscjgi+Ex5d/a/LuI/48nTZmSjijWGLb1xpj8rxEMoX
kTrZYVM+cG3CzXXZX+lIu4IS0JT51vpKtjmQ5cue8AOr0txK4Eo0n1IPHmqf1l4dqMH+2UUAAY9n
S9U3hwT5BpSnjEE1GuBlRnaOgwAiYjwkt68jY1zwUxAXlQZHLgmG6VhKNoTar8uoW2Yk3QyIdmvb
GuFE2+grezT0dZO1ftU4a7i/7Qvuzpw6YfF6afhL4gAph0SEXIA4mSzChnzlh21fKtbtclAZiQfL
PBxY+PlNpZA659J5+He2KVUnY9+bN1O1XMWB7V4PesD0deJ3SDm2XRO+A7i1Fjzv1QOa53V/t2jv
8hUxuK8Upt2oEiDFD+AYClQkDM49mgcDDiCM34Z0G7N+bWjPHy5Ft4Z8+6i3mQ+ISPMs5lRHMLZC
PDbsrswylokBHAeZ0k0gXNAVFC3VlPjcDIjSnp15Ku1NymlRIH6tj9OGmPw5M99kG6V5qdVI3aWR
Gkehq32c91OXPHL8GINpV7PNblKZoFrALa85gskUgaciO7QHUq4Fb+rsuf746KzwbGFc7LOcrO5L
nTQ+YPaTyGE4K/4ydFXhoBVa/954BAvRbmZkZnGa70V2BMArx1m7idb/PZ7azEj9CoN35KUXVdsf
dO3ZxcQPmx8mx/4MCq10SZnvNCkIUC72+nTTrWvTV6x5DJRbh9DivYCKU63h949HScFAMbwNIgcG
fP2mkrNHnKjgDYxS9CJhWEmv7IYqCQ50aYsOUT2pyqYniSBkQT3gn4QQLa99LPlXP6/6Js6txUQz
3PeG2wUj43uI9NW3QlQTjXgLVq6Mv8SfWZF8GQdY+Fp9WfgMfdPF9cDCdY9kY4mORZBUopu6zqXW
1dD6S0FH4YqDrmolKns8xW65VpomfDZkTdtTs2HhUtPNM+9LtqdK9BFPMhuuiWfq2U0RSezeTnF6
K6UtXULTUH7leEZpw2VdswCIb2KMnsM0vWk5VkGTn/zmonnUe6sCZ9jvffbTgrjjiOyNKAKWc2nK
u4990tRKnDEDhPe18XKQCvnF87TLnxxQ4kIf1koV/k7FCvBtxcnZ2Qmhoja0KsDZ+OOKCm7OXCIx
HOOvuaj2FB0O7rqrBH6kYiUkDE84pXvePkjNFGYEnhUI+j2WlQRNQXTme6OcXwzhfCtkYzb0BC+t
UFRJ4CQIpK2UshDYE7Yi6Ew9JefnzvJrCI+8qaamhZWoojO8gbuWfdlYbL2UlC/ptEy2z8YJLPG3
0v4NqNZZNH0Aag6E8u0zdmW2AzHXgtrlD+qatAO5Z6M7cYnMQt1eFL2pJMPNGkZAhNxQDcLWX619
0Ud0m4hiJexL0fUY7q4y0Ins2bTF7/N7oDLeatmiK9LTpHfM1QgAIqWmToVlrzdgwP3c29Udiw6d
t3Gorf+BLxlEYMc056V1cU+4b2GtxqtNMOsEZdaMJawSMQaQbKgZpaxd6PQRyPAke97fHVtxuw40
enHzIzw8OdlFV6PAktdBoeClBC+Op1p0csQpcOj7+8vxDhsI5X+PI+bEaVMxLWRqpzEP0ENdRyEU
NHo+5bJVVS1tvQeNY/B6xNORQmYnC1Z7PwdteBYe1hzAy856PG82BwEXluuiKc03ApNdgZc/PmzK
us+gVrhctwulLq72jCrEzxuXcUDKVz4jCm/W9Tcq3AJvxcovSq3GZzCo7lDqX/NKSd70DudfBwSB
oH3p0GR5uSmvCmlgUFm83x/dv8u9vjkw1We/V2pjlFuAqyafnNRcCsdEkG03cM6i3N+4LIVSsk7o
R0rnvNtvd0fWuGIRhOHUexxefaB6u5UZlrf9ydDpWuh1gD4UYvST5V/u+bQayNFDjphgbLlAsesJ
KWYt6tAg+MfgAhs9fmz2WYUc07cF1SIG3suk28uKENfLyuAQvL6R533xrMQ6UCfb5TaCkanF7uYx
oqJk4ewqxF0nT42woJ7VHt8TtAwn3IZUMTUe1uVa4zo3Z6txHwQQwhGc0L9ev3XxMiwDvdstlj1o
14UwR2MCRspu2gRLz6YzfmLrQsNUBR+cHT3EGJG1PpivfrrEV991BH04RTIXuKmGfoT3Gwa9719j
rJRqWnFrc1X7dEb57elgac5Fl9D7BEkFwRNVxN8s459DzHsg/UgD9jHnTThFczc9wGrBgFz/ddNv
wLhWaNrpgPRN9OajiBQvHvgPg4SLyUWUoojD0qC1DuvktEOznI6VU+wGdCji4oNiYeqRWCPPq9ey
du9mdo1gsAxwdcOPGsx+lIfnZD7z4Z+kDmc7VG9uEAzcq5eeZkLetiF0zMt9X4duJ6yayavVVLZ3
1J8QDR4MJ4UDjgJI0SkuOOntskNU/yWGA1O2HMaeLY6qlRQjc95NFZYw1UafCFK7MC2nc+KqeZOo
OAz9nHF3VZ5NgD6S91nj4efivvSsCopvmNHxOH6GcgKeAZEJIZx258riO7iA1K98myoINUUYTdof
9Hu5B6UsWMKWzt15cZCTQqoJEC+Vv6i8DA5NQzqD/UYltJ5FP6kTcx9Q9t/2X+w/iGQXrPlLJy+D
QwuumQ77ULJHnG9saT3KVOVgj/GJLsp3ueXkG0B8fgxrZ2yawUx0ZyNSfKh3/X+ZDa+Pd1pEekpj
hG99rFTYYYIeYlRQlTSpwIVyXsxRlguMIA8YBXPAXRXd5d1oCjSTFK6sRpeabjoD1eIFZUqvH+SK
JL612DN7MeTHIzae/EnhYuy2FRMJzuBLNc+9NU7viOb8YY+hHuIG3ooOSKta8+839Ry9v/gLJEd/
f02LVmC7oO282GbMJYCUULwppo3AJsj9lQcHo5R7U0MbG2mgpd9qLlEDZbvGpVUQSe5gOjuXH7oT
NPdTZfEMsd3CU41mu3fXU7dEwzkKwNb4x05SHpLZoq+8vpprnJa0kXZnsHE3EfjlEf1imVNkFaST
EixXgVRTpL3eOemrIsfIx/ln6bGCmptcHU/DcLLmNl8CGNI7WbXTGaFAxNOgJOAPySCgF1Xp83Sp
WVXd1Vmue0YOsBljwBEQq29B+rGU9emIJvQNThYEPV1rfjF4n0GhbXjckRIt6FKERgx8IVWRcfOz
bs0xu1pdrJwb/nlU+RtcsBZSyBhdJ3KpD2gJbSwrqj/4tLWtlT2LgmnRV7wUbCI/U3rexwgE3F8D
HPRfZqA3MveFKFtMaK5VnKSJqYrlW8II/Lvz5lixjmdMUp2nkyf1FhWXL/Tffflozqtp3vEJiuO0
f48OXr0CJnCeNlXcUk2dyB2mT6WlLQThtsNimpY11a1Y1YvnwNH2VG2cSXBBAVmq1J14dOu1EygU
uwseNpL4qE+t2P51fv7Q6l0pHR0t0+X9f1ehaCQsye5J1Upf6WfW48QhTEYyLEL9I6KZplibgbVy
cWIoQyFwiFJLeGGdZazzgJXfExTWEx5mFV7D5uWakZP2euNrib3B26aZtk8EaMcalw/LnHuo9rwm
xE06gTsOsr1W7Ja8EILPnb675kXifNmVHwrRD/g2oJ+0pOElESsxpopuya4UsHbVdaGYwXwaXtKR
1Rvp78D9jIOub8/a4fDStC5EmIcxmqLW4oBx5QPRekuvVh6p3cdz+G+ZLMRugzrTFxPy6W6BDA6d
86k0EJ9i0hviGdoWvu2kUeqAzpv7TP2Zufoi0Q5EjyP6JF6W9hBNfFQyvLBTTNMrlFbzghHVZaRe
VRnug9hg2s3OdYPJhQrWug/RblGG6SPXQpvDjfXbRL4sC3szqJCf81ZR/hnYCi+LUyLd7I/no28k
6oKzlCa9TF6S+GbAMu4Ho6AU5h5VjEz6BJbwc3teRbHpmXkeX4Nd8m30tKhuj3Ca6BFggcyJnaQJ
4U5QRCV8/jygVW1IWvh3TjXBTCYsj9XYaWRGF1nJFt9woOZiF8DlZSv0JYct6U7urrSW6MG5wfuy
h28CrBkghtKnOyVPnbYslc913YtBUdoXFSvNbpMSkUk7Lq4/ErsIlu8Hmt26G8YUl0TYeMb67+C3
+3tPmyZSZhrtNvc3Jmk2lMCBKKSeca8f+PE54Isc2Oh2BKDYy2/HybjpJjF0p8jR9gvfWHBcLnWr
WCkKbtflI6UTjgn2fuFy9QYAhs1f2hNyk+Ob6+HLGucj6Y7JaoBlHOvtZZjZLRXrK228/iNZlPUB
X3rGvzQXNvWjLHwMIxvlUR3Wo3PZZU5oXV/LzKMHxx2DqBJlPHPdp2Pw+1QtFTSreoNMHSR55343
MppmUKnzS1Z62C4Q1eIUs7i4lR9jTEvU5UnH85ABIkDbYydw2Gr3/1V+xiZw6+6nxD22gVRHtYeC
mRv6Df+9/utg07lNdt3t60FM6BVzWTvptw6Saex7U2o0FhZAIDqezKIODXgznlUmRMe5Qgh7QqS1
tnhp6tCDEhYuYksQA3KrJfUw6iurnvDZ+BB5gzEWtHpXsuFYhB2j1NCokPQvLGQURTftIFOlIZoR
OTUqQ3asvTy5iYm9+shsPeCM3bVIhRAsP4nFRMwulG/4eLxXwGcjB9xxMd5eRMt21fhiDIwIGwSI
7WQoozHUM7eM1uz2+3QXMrBYUW79lFx4bfe4uoIwxyJ/XhiYG711KnTxUW0OcaeBQcN6Bv+AyZ0r
xbnmepzEwLdwOg2yatD8ArH2hQSxfYkF0ep1rl0IhsSjELrOdITSnCZY8TWmq5zYE94kjrb20zYi
Nl/G2SYONWBQX/31NIwyi4IEABLCDGWBrZFF78E7YICr2v3bIzilN4Wxeun4+hvUaJ6HGpki2kvz
QtbA+whi5bkzLHNE6qvenyULJhrcUDVATAiIGJmX+t8w1E6PrgyZSkDnQZFwawKJPu8qQa38nwyR
oqQ9Ea+YuejJ7DA3tVQWedkJzh4ZdGzKg1IvaRGjl1vwNgxsHF/nw97N9yd9v5eQx/+Mdb/ILphQ
HC8jX7gg6SNgxgMLnCohnA7QzyRdqyTMVyMyHIY5O2cIrDpany4Xxzk41AFTWLvY6XuF3/lxh8aO
XAhjvdxhggN2lVZmGH9/3EfB7QBUQe89fvkIyP53gRPXjBVj40NtI7fxlD2zIVR2t0gZbQHtvOUM
F9c5QAeWMddaj3n48V/gCJPaNe3yaYbnu9rgacBYn98O8cMQLcz4fdGvYfE1l0MzcqWzD1VPD5tZ
gxz1Ped44TQgG+t0VmmoMUrPNBpDX670HLjPl9ED8TP73D7nKixHMNvgoOFUu4sSHDQyECxQHfsN
v0Mfz2sBPCQt7m8/bb3terPs3VTmLSqhj7/h/SgmlvGlU8oWliS9DwDDMl+Ob70Dqa8eVmq8x4e4
K7JhRsPrHJoWIJhY7LumZhH2m8+aui6aWUWHidhaCYB869V9aPap4LUb1iW4WedUT+RpeDahZ+zw
iUWsYDM2An9StQZ0PiqC27miFxsQJk90PtJs/W+VIfHiIjNtAhBEi7wGwUgH0u5xsfmpfpiAUxQT
Ir1F14zo+6k5qeVc5w+ukJu5ZOAzqfsEmcNp6ErbaZkYaedFimaTorc4pYvNP3wjnB4QCPQAIlMy
paIdrgU3w6n4PqnY63Mh6GuR/ljjnBMhjVkHiHiykVYNL1NC3+VErPkdtR3phZKOHAS+XLfwCBCN
6WfW8I2bIIANsM8K+Nvpz3PDhCDGgJYxc7pCCBWfn6B8MvEQ33ExYrymC9iVZ9ph/eE55xIu3usU
WPdYX1Eou/lSsszPkBm+hSnaaVSAI5ozlJKO5dUAwQ/bGIwiWGUbiTZNqPRvDk9CirqwmARiSTX7
BIXf6IwRj2rhsiG5ZHjp8phDz1jE0UC3wL9xBk9hg48ixA8Sou2Hw1XCXgxQ8YCp+aBo7IFFr0Pv
dkluuD5pwTtgvVuoJpFYe7fST8co87w51s6Q3WXlJKier7p8sqwgmfreqv1186QNJjm71Q98pw9S
/uRzbmaXyBjN8/RGiYajfv9s4kSXxBmBKnU74q1wvLc2u3obYo0/g6g9bxVVVbq8ccw79+IAaHbt
6VMav8lVoLcFSfOgrYNZChwWsol6l3RScf2AdRSM+DTmaRtZX0SdHUpvVlaJHcE5W6nz1vSlf8dr
lozdCwaBRz3FQl5nfq4nIGQUrnpyEVjJ3+8Q2oR3unOOwoCYRXiYAzRhO32KY4E1ZWsZxLZCa5qr
BF5vFkXVZOIBpFvDW3vZVoXoa2bTJAYTaPXYS6SNM7YVF2nb8+RjV7/zv+5SppWFyy+eWwgtNew+
YQT12xN6i4scSPYflRJLHZI4hv5dm2F5+uNuhfRNirQ6Nns0MxO9X49Ty2C3SS7ha4UcqXoIswC0
D22g8wSDxgszPYcAaW7DiAHYTb+i5hvvm5BXn1f+C3SzVsLVl8eQdk4G1mawpxHNTIcU1jnpu84e
uxmcqRcACi6HemBIVBOUwNXu8VzFB1VzBRIi0T4ME1C4akXj9DQQWt2oQl7NNLbULEM7JQjvgLlW
9jyuDThFW+K8uXslHvuirViRrY9PLJrJrq3bTfDZaI9kGLn201mRfXvYLsD1kWWHJzmJLY3cs3y2
UKqY8p8C0BPKsnFVAicP9gdjf/e1vMEuNKAMlYYJLQn9DRN8NlV77xF38e20i0OaJ9i5r5Vq3Q12
Uyqy7dm/Uy7ksVsYimVozmv2s/TMY/gJsZCR7xWUJt4/dRCvn8+CkjDyUfv0J4i3/upoGyvGlg78
gpmktgxvtw3ifSAU8996IxGBVQER4hvMGmVlQlJrNTBsIO2vGDVIVgN0A2FsOuuBHT+T0XazE6Qt
rZUWVvlYvzTvvVkr937GD4oo+E3gwkUu1CgzLLLIVv0NqvclGeikbhEyxsoh1f6TPPrGQEgq0Xwg
BrbJ/JAB3RhFZpdjoarHZFeea2w9ItOUr/rleQM2ujkAnxUxh+XxqTQOz8ORq48MsEaaTRDbropF
AGMxXZ674040hkkMyOBpOQTajkthd7HPy/HKuPqyCR+Za44IwjaTbRNFCkK4Xg+H3NP9WoV1inl2
lh1yy7hLSqYKzoYV2j9E9frzIs3XhTdUTqTT3WqAwEIaqKFh1PT6sN/zgkrev0UtEocnPQEvr9nM
tSfBjVSTYAEn8xhDfJpnFEpD8FVx4qeKZ4PBACvZiD4sbBp7Efp4AQQ8UujUiC0L9G1FIkXQIGry
M5EdviZfcZGnaAmy6YyPKzvQON1ZjGzVjwqCto5eJ6CdYZ3V+zple/vgCy7gmEBbF9B/gvahvJGM
TgCSh+D9AAnaNOV4Ofm68jM5M+4iCp6txWLWkWCm1vGiQfzU88fItmaoEwa3R5tLUluSLZKmwJRf
d3oDcCL+dFYGcDPotF3+TEyf+eGa47SDdcUw6iIfHZ/aIVDZeymzFBNPBV8PtXLDj8+axnH8tIYc
eiOg8mb9w5wQ7o/eDdDwBqSjhnOmP+f1TO8Zu1NNWCLYEjRZs57nXlDAZdeQj0Ueqq8Rn84Je44S
lNeaZzFi3LEcIVglTbQhFav3uESC8t1+lXnlkyMj75bUHY9H6W5wrUlRe6jIQhofHGV+cN1RDBPG
3X27K69l503/+qXSGXEJCQEOjMD7KtEOigX3LS2/bFg2+ahUFleujX0zqfp8mjU1H20BjR6c2Nb6
I8/fNRm0t3/DHju4u/FqYwNAqsGYELxQw9Hdx+5X65eycW2LPBiy1lph8bvu2qA9ALqNHPSJzNX1
Y6OJVbKdFcb78BsV8HKaR7V3Dgl+6c77/rouJgmk68RYfDU7HNfzPjqrQApoCZbL/hU0QHhQg4ON
F1LTAtkoHpEcERS/s7V/ZclUuDZSWhaxF/jMaePJJ+qMBfNogTIJuDcSbDTgucYZcVTAccjFTtN/
a4JGds+k6A9GY+9CBB41WnWlV8xrO/Uwi0RbIwcI7h9sPCwEcdA+rmkQI9bF8b3g2JgczFzHTJ5H
wcXAcPW9B4GKTqHH0mZevuB1e0bhUX3lLoU4NRiNvrbO9pJHQEHkCpEP1/c5yUJwb/DfV8AshbVl
iCTIesBvgrtIFuXDY04Ejtrp/v1FtN9rNGpbKM/PAq9IkdDZRzdKpQUOlrGmyxG/hFQypTnozH2E
1+MH5OYDyxckncmIDNL28oGz6zy844eCH/4s6hMblf/J7yrBiFXlUoi7TsxBRUyiBn+ovstfKFDG
I5iwLOui/KCmKezMS8/NNn8RnbaeE4bRIoEVu9FssJYHdQrFwf6lc9Pm3kwCoOsSObH0gBAJemPI
1d3ygBEOYTbd8uPvX0XzKoFGygquWbZiiK8ICJImv7cazeNbpDTTDKIj2fcCt8GqUvqbrmg1gyj6
RUsji/+3oDzwSpt7mCKUYFysnlyIXidFWYJp7w4x0G5uMrYyLr5kGq57lsD7D1p9tH1DRe7zHZf3
7AtYtXf1XsmhzmhUn1aWJZxm668lXWuPHcmDq+KOrmx2SGh0exYWuXVJqrBXCjwTRkH8pBPUOfMJ
2mAJ2ADoWJogmLEO4l9obK7rNfmwRjvMB232xIev7iGm+RcyzckFm7NNKSd2b/1U0+DfOBBceCXI
GH7K//crciAuewzdJrkD162CGdRZihgh+etS+W5CxAkrihaNqoLxGBZ5thBkquVoDfWE8TW4p5K4
wysplJiscp9ULJSvQZ0+tx5OH7CC4oM6oibMcL4Dnr0VLH6TIJzIFQRzjpFBZBAoQKrpIgZbz5PH
DUVBt4puSUfGNKOlzSpNVNyqUhy1FH977G5JqqjZQoncoMpZoKMM5eOo4pwlnakiCxk595Z3O49/
tnRX+adcG0yvTcMcGyHkMcibIKQ8I/sGqGfR7JkRZkmdYImlRBDo3o5189BZP0AT2BZn83G7Tqk3
lGs/GT44xqcN9ODBf3JgNJu8qK2sUCIlIciOCMsof8gR5q9YTiwihEfVLBCXZyGxs4Cpxx4tBTDH
gmtmiygCAvrY0ze5r3B5RE1Hz5XPbcwQUUBQ1Zkb6fC0G2davp33bpIvrlNzynoci/a0aE1J4GU/
RM9d5V2QBZP60vc3hR0VY7q10ZgZRVLmKbwhRQf+WCnAQWe2tTI4hMxLn4A4hlS+TZL5/ceNBJdq
x7OrqLI//WIkNX/b6aIeFe/JT/7dbNIQBOPqOzP5epIbeZzuST1+x4fmLxlstCI2bRYWR7oLQFP2
ggHhim882IoUBB3goneg8HjLixX0rfYhlujVqG1MiKGIWAgtZHr5UyFP6cb87w4W+JOtVpWoFWOF
pB7OUfEDyveHP+5gT0rdFBbUeKqZEM0W5BVDBPTVB6NxTlhN0CDB9F8Ha4rRg+dK2mzVoStrVJ1s
4Cr/xxfD1/wKVsrRNtABxyybE8eqBQ34HfirVxxaALbO/zTzX0xdd4X5Dzd9rx5PKZ0SippFi9bD
X7Q3hOSofiS5pCIsXl+f7k91H8hhcdXLWLfTex4VIWLpoKpjNWINBBF8KB+wUorGQQVbpkunf03f
0TzlwAqGpjAEfqfLbzi8wC5Bjdrfvl7k0oFyw8WxNer46UfkGtwR1jUDyyk0LppWAcW2Xvu9x2hN
lgMflvRHmxvkeESBVx365F6fdSLuCisesszyS8UnDoR4z70TWM3GP4aDJCLEeVw4z8FTROVrfnLp
nDPcA4mEAwIPOF417oHiQnUVG9BuIoZ59Z2OttgygRio7/rB8XOck3xV2E/YOi9vVYN6GA4cx8o4
KV+C/uYkA/fXhT386Z2wQKU7lU8PFsiKnvQGO/5EHVT1qCdDwZcjTqGsTkYXPQKdPLfaDOmwJs+e
MDa3QZm7otnj8cG1JnzuaCTn6b01p9tQskhI+wfG6+ezgD7qh+7EEBpeRgVsSR9KXpchJS3PLGVN
FJPyQBXt1buwZRNTCG5fdYgL2RCgtIOEpq3ZNTY9ea7VBACvvR648GJdalTZlIItmMWwnMsV8RwL
qtwEbBZbkoHa+UURV2nFT0CAnrntdffyEaeqvWQqq3SpqcSYHC+73eu9tpj4uMXlSqRny0Y2NHj/
1eZmcsr+45u9g6Alzed3BCH+GnsiR9hS8kNynho3zGF592DMXNQBPWEfmBYNcGDNjX2s4Ci+3/r8
SkcmQigra10LLMqrCgjOHw4Z8xKD9CRzueq81qPXA6A2DXqz1Z4yBGdoM88dNdhzpmoK1N5yCe7w
/axCjtAGo75RiLKdq3MXL6qVfcadddNi7tLORxdTMYRtVC5E5b/g1mLi3J5CjFbrT7+IQ7es6XUR
63fX9m3u3UB80LGn8U3I5PhAQi0LXm+C0FLHFH1/OoJrSzNPhc2YHwgbNoOsnS6GwbJtmkhgD8bZ
0xylFT6Sm3/mhz6ESNEx+faxSg4yF+SWOGDVnM63DLuRTgNeTdPJQgQEXcshZZzw5Ip5CRFjbuFz
wijQuIlmBbGwsB/gO3C6aBc7oJUeQWVoRmzU3XFvGR3X3xJTZJ2RCwTTINOgL7GGnLrtUQPTffoq
tjbeg0piLvktZexRX6Cl3Fh5vo8AjNKeizpYNdCOCGfuMxaUhRajvP8aMjvY8RGXRJ2zTuXAL1JT
IO/9JxUbhEG+thrJITwCT97UIsH9rnH2oRth8FVq6xfYxOAdgHWzYnoM5AaNJI/VIoRKJvc8E+vC
dlgMJCTEuokogFyogkpC0aX6YiuomZIVt+nEAhhzeu9rD9YT7KNw5l6IMOu3hXZyyVTVm0UB9ktO
0mHYZWt0Ma1wkNskNwYZZ825OU+sxSD4WKU5iu7Gor4AAoqHRcr/nwY+pctMY82qPuE7wGUbtuEM
zoeRN7z3rYLml4Slp2yf35tp0b55fcyqXBr46CgqKwV8cQ366exxymUEtCYdsb2c4NELD2axrwtG
FY2kokg/t5NE5zArw4eF2o2emqiliPdvzn2bYDOzwECdaO+2mPPOkwuP2NFpZkv/NX+R7n5/q9f5
NSO0L49GWOZ5zIkd99qtke63WSpImTrh4Tl2hlqP5dVd2C8Opjct4b1vSE80FEm4Yz3a/TM2b6x5
jg4kc+cVjb2+VVt7prrdlbF+7sVV8P3ow6rXda5WYRoQ1UpshWs6CfGiMErTH5rLlM21FLKwLUcY
VwoeXU6NKEw9hnE1UQ+wSznaXypkyGf6EgqwoTJHU3sKRRK3tvtKqPGVn4LBgAz+DsgRq0s0Skqx
fzASBHzdBzEzXiA4C68MNLjMB08sgVTEbJ5dNGItghHjLLtWyCobHZCGNEsOEY+UqdW86tMSsFki
W9m41+oNfawBgvl7IwvgC8lKi0YUMCrBfhc5dMuT6FZXi54RBJUj3HmbncztLp4mP74enzeBlcnE
v0XS5vtGIXGNpA9bMTW2gUXjY1lMOOPNokliMNhfUgua8qKVqR2otU+xdY190oXy2b6/I5UrcuSE
SdvRRS5kiN3/sNHb3362nVI2ihp8YhEo3V8zVLaCoLFNxWz6pqNhK+kbY9m2vXooxg6lKMO5lXt5
wakuVB35N8sAsTqgKyrE7KsWvXXNTE9rsFhe5/KHuanAyLrdvODzE/W5bzUgRjzmJffxkkAPwEx6
iH8PX5XnivU8Airl7PH0Havum2TcA6X0N65jYTxjtVxnRuDZxaxPr60iPAqgu76UPchEvCREDBip
Fnbt9wv9V3f8tDSTv4e0rvn8uXtZQ6eUAr2/khzj5DRByVuJc9jXD6PUCbg18gMYf1SJZtBknTKP
tXqad9ubRhlXjVb69eoNPpcdQEERINWs/2i5cNfFC7kqlo8fn5NMV7zR9oN9K52w0mwbBPELlfhE
Bi8H1jYAVBEERLYFR4P92ZEukI2Wlwbs6XAvs/S5ajZ44TciKO8hL2PWVtJdCocZidBd9Cysa3Q0
DKXyFI0TuRy0ol7/1r60CLFHLxVSkMoYhm6HAP3fwk55FrSXeI/bQJCYfniTM32hjBRjFCvseMsQ
tVrJGmaJJz2kfY25kuce5AS42w3KrUK8Yi5o3dgqTfvYwgDs1IOrARZVr1y1MXU3AWzt8S/9GsT5
C05GAAnW5zYpohTNMDaPJE5BHFTMNB5UJdSHi0Ic1ITXe0es6ZpFRk7LVdX1kHdqidq89yGewUWz
9wZYhB0gP5VNLDceRcbR9+lJGop62JAKp+3Zdqe38SoaQ8wIXTrqzk/OYCHw3tkbqQxlwFaVTjGZ
ZmaAe/btBJfjaDlxznSKKIHKyU4QBae2iVONuxLbILpfz/sA2woNcT7dWD3I8XJmkr2+DP3Ncgsk
3+cP4zRZKI1rI/ciBJK0C5P/irATYbwbJ0ZmWHWHLqXXQsRyuPa6pEs+6ob4Pg7lyOy+vAXFZAxu
MeCYM65JBHusVWnntBzLDI+9SagiEt7FshuviW+qj5I1nr19M3P9ZEmQlpLYFVfkg2WP/LBDtxTc
ifcfEXdfxrtg5RX5o01QmJRLJfNV0H2riU0+oVKJib/4Pdu47SpigAp7JLcRKaMX74baHBWU6xw9
qTHKydpzgLrYKmnMKecpVVzoUwXkXn7UY45xlOllI28pUPcB9bhnr6Xgew5UWMUfeu16lRpu509x
ljSM5EMuxaKvALf6Sg63JqzwWxNmtNvRZb2vk8EEc4hy4FLtsonQbmFNeWCVcGPoNYWkhaarDI5d
Af/SPSInYukNuwjygJGsT45sxHuFr62FI+3TnNr8I0chHZUhjktGhGU+pEXTSnYsMPsDiVXaL0Wy
z/eBXfyNqdMB/vls/OgtUm+b0Fa+RdA9V7kEynQDS00oVMR2lsHMwWYJcVWnIsqxuFdZKljNKsAH
FOHhkXxuwRuZ5oYgp3e8UFQe+S9Z2xFTm447/xw7r+VBdwt4Fqog/0LH9Uq/YXVCJHNslAScdXSR
06OBR0ZjR04gyiylGzwnWqYUUEuPeQqr2SEhoVF2t8RFlDRsYM75FCSkkPiZ7NGTbAMxnq4q000Y
FD/cYGD77TFyvzHyheytqCaon55Hw2jIZ5p+aV4Sg89KGOu/yaVPjjKdUhNKETUhCXTjHugq0Oxg
UMQyZSX5B/2phaO3HHnBUTpayjTVY7naCdCnvheIZ0t1YN8scoIo5S1lcB4p4G7RFy/MmUPd7SLb
wnyfLxajY/0jAoR8wyXNdZsLciiQYpG2xiSbiRV0qUMuSv2ggR8hj0OiVx9bC1zcUffYMDuBugoH
+q1sVu1hsijIDmVedR1f1tVZbKZVF+k9xVTD4HSK7WadNDspUzElVDXTqmszruQoG1rkxXJhQbZt
H/S8ERGq7lTvDPD87DZ9ljQAzz/4xlRe9VJHSdUlG3iAYu6Pnu5yxD0tJ4ubCieQWvx/KuJFH+A3
VCgB6jRH2K1JxAmmV8bSiBWVmho+3LLD4IhzSzXlLdhmFnmfsgbtrZKq1fadB+qKRcF+/H+MZhS5
JmqvDqdacWV09lnEQXPYKWYt6CzfYcd1aYNmfDm5IkoK3jfFSwMJe26FZZxrRezOY+IjjRkVXrws
dPeplFbgZzB0/k6yVddcXNrtYHvbRqBGMujjOmFWbrU425whqrVhDqLHu5tUGAFNV9+F8rd8+yqU
7qI3n/FxZLlZ53IftkdesEPqr+G1V7+yJdCfCUYTgIJP3VRBzECdQR3RWgQZSctrijiSITxiQZsS
0Hst0cvRUuNDP5Vhy+hAo+lOQQlQOuzIKeyp3S4QvMZ/sI+Axav3Sr8kgvUZEsLEmEDvEmNKGwqA
7GskvHzax6ACLBE9Uh8HwGKZb+VB9M21D5Gz3a/o4myF8oGg8bC4wJf4Eh4rSHovfFRfVd5BuUbD
lTp2g1O3PDKvRtA/cbpEKBO7m8XtFpIMv7NfdHO1XezTMyt5r775bSurGdafqgrqZurIMVwKtcKM
hGli4h6EYj6/SeMV0Dpwjpwh3tuIm5pcmKg64QmwZ1odgUlRb2WLQy5n8Cp9Lc5kj+l1sxu8HBwM
z7NHRfVxAwimSmcqFxlccIUJw0endvHJqcSY/cQ7nM34YhojuPn58UN+Oho4EjSoC12JiYuUOnqE
hce7PpgG3NxELSubRoXES887+wenJhOLx9rIQ12BUFccwEDkVA8J/RCkYmOyG4yzr2PuGZh+b2JY
8UEzJ4arZlhh3tnm3sPMjkmRltKWRj+J50/qa1pVounjiW8pQvXBj9rOKuACVKOF0TGmSO7SRnl+
w7fkl71hLe+GUYem5Wni5NCWSCOfqNA+P5EdxsG2R13Zmgvsb/Olf7WA42DKYEXoo7afpv0p6wzb
UgDkGGA478XGg9pXmn/27E45DZjvqfvxQ0d7apIBAyEuAEQlEuXQgIEtesbHxGN/wV8WUwInpU4e
3xWj29VfH7eTwoj9/BbUruN+ITuRwZH903ADkUrE2I8k/jDn1Oja2rpCZYMWg18v6FQt4v+QjAHn
Q8Os97bfnajFcqeVpoj+3mNv9TXk9r9Q1mljZ8Io4mKKzylCi7IBV6ftqJgi9NrdCwbxWoy0XxG4
RP6VM3KY6UY5e2zBHjS2ZDA+JmAgsA0iYOeQ/z2D5eePMAJrGB5X8T8mVDWBhWguNn0ZeLPN8WBx
Uxfb635kyRDqh8BzK/RzRjIwzz6YXW0Jx0kUipx8DcvPgMOOJxJEYzqwuBTISRU+0s1Y5Ts51rkx
Smg/BWAhpkXtQnKVin1hv7DpQjh79Fze7I0NnpZcZeAhuHuKUkrPbE/KlImR9ogOtRMkEZ/peI2E
/yp8uT02THbLWw8W3adBuMrPX/C0qpQfdSlDT8aZC/4R2wabq1GgaAneZAb1+TpWvSs99qCe3qQW
9mA0oe0iPqR/UvU6j9R8+W9iA8IzNPXR+QTaE8SlHGkk/i+0Q/v/RzLDBAkxBR3Wwac0MKrDcBAy
JoQTMSHUhf8sAJuNjDSKlCyzZrRTf2O20vX4gJl13Ewox3TwSA1WIhc1ZlLg++Tkqd5DyHbMhYgs
lpYw0Hp7uOB6sWa12ay+4VxS/UgdGgSgtyLmqWGW8TCK/LZ7JNQIYFZ2l1tSwKlia3Zry2hyeHcc
nKShlQNghS+DSqgjU086nuS6JLT+tUj/yOVh/9Akkuqwe0qmk1rhRCQqVad9bn8X/zO+mU8msIgV
d6IvG4ZYO+et8s5bTucRiThdWvEP8J3dcfUhd1g1b8It++i2HFX9q2FgHbovbEQCgxCyQu4/tcu0
rkTNLKu6UwtJHDA09RxQwBv2sGs6VAIl1tDx5Hp7A+S0J7iBo72flBvJddY6P7LVmU17lvlyBhNz
1IwmjzpjrDmXeVaJ9qfhhRCuhr+RRVqZknrRZSJv5OFeexT1PiCJjLmrPyiGxW3tWdpKqARTkvT+
xatpewTWVoox9vbMoKrxLO9Su7qSdToGZw9GrR7gdg6PgPzBV9BZD9pfp2QbTbWO4usfdYkz2EDJ
quAsDtZth39nKJo9/N0t+xDMctbqxPu5WlEJ9Lyjc9iHH0NGzjNfs0sqFMCEr4TNtA2LC8VZDMHV
iNxzpPBPwY5imxfy4xGQ1IZneY7EuWuKe3MicSl9gxd3TNCVZAUJaGm/EY1XokY5kZqXd4E5AM3x
stmKKo+JE2uWRIH2RHN76EE/cCq4hjR9k2F4LR+P7rnO6rHW5wFCTfGcvy9H14EZaCZQCqwApLEa
JjIXJNWj0n31k/2/ayZoe+q9H/bAgFz666YgTi305EgV84xZNMONH2yc1ENYFMrYlFZ+JtC1n2yY
Bzfp6Oha+64+WEgo+iPWRpcSc2KFtJNu05lH1j1K86ciBXVc+rOR+9kcr3tLANxgsri292PrYABq
tZ/gJgpHiRkDr7BRfwVJtqskwTZshfObyAFbb0wkZdmdlMHnPq3JYuOOUSCdf/mGqbi9zsFHoHsS
aYXKdrstNY1YN2br6xVZdgnY+FaGoHbCKN/MjkJ8wdl3AHrvry5yCtQQ3dpixmSx84QEcuewpRLL
WgmqIKMP+i1SXXo7qFn84C6H+u2wq72WsocT7z+fy+MptpCPBgK0Zvr8Xw7vUDfZ/MYoFD2yWZFX
Z7Nw0jTLrI3dg23GSmh3inogb1EyV4mBCpkNdDKV7uMSejmgiTPsFFP028YFjUahj9bBPXds0hvx
fd84jh6spTXbHfRCRGNN2u9T/jYSjDS9VEHMIQaE38sdMidQWMEICOnkmTQlFM38ak8tcUe46sLI
gKrKRd5OXOjm3liWSiQNh55lJ2ObZLzRTyMz6HHlJFOgL/IvOh50QP/K2wg1NGfaRCqXqgN96oh8
xBJcTK1Qz3K4OIVwunNoQOTRRA1X9P4HAzzSbzaVHpotMH+P21EuPvbx/sdCKaQYXSknGkYCDokg
siJoJAjwKXSfZRBEtQPimS9E+peytpu0BpwLBMGnioZAmWT6Z3xLnGBnC3ihM1BtcOfjXX74unub
ueojWj1DltmVBP/SQSoWhrsXIVsJf6s6MYANZMVjTaszpoSWrpEHZ67DR/8dlqLhJ3pPijaNx/EV
qWeQF1rj1h6nLAzT5094m1iEvA3eWUPPVpnn2HIhIygTO6f/OiKRjcXL9LNZ9RVXaxKO9gYOz3+r
yuYnxCPro9Ljv2S3uk4elGDFpEQu8wdfpr4mM6I7dIM5BautpRmEeyufmnRk0wLwJrHcZS9Ak+wP
2jwgL1Ts48Mtrb1jlMkUGdy+ATItrKXCgO+fwmI0nJPyOzpg90wfqY87pyzwQ4gbfMFb4enQGOR0
DSYRZP85O7Ic3dEk/16+0lFfFWfs7S+Jqxm+gwvC9NYnjIre8tgI84kAlKCXEE3sJJuxkdmwYIsb
k/1PSNdzBx0ytZmmNttqf3b4AzgjGJ3HACX5PY1nk+MeF9JaGGYHq9rG2lABVKCUhgKSR+T3aA5+
c9MptAomdFiHMgrjRwXXf1SJ3zZ4y1dfUHMWRE8WmRUis6f2uTCfBTNZcgRdKLBJwsN7s9xU+/Ub
N1hlQJzZ53/bOzQFP7c4QTa0cUDUbvyGVHlFzPTlCSsK+IMR3t3D/NURUBuiIT3V5TjdzGjUjdsX
WJBAZ8U191XK/NHd7ugjvBHN3ESwCQxUE2wVE95+xbu8vpW13K1z1Ib/l/tJLrp8v92Zyd5PFh7J
s41hR+H7vEcYX87b6lprc+g7JrKJKIrOOmOK0xGZUi2MJ0vJ6GEeRuJIJN/v0mHOZeQd74TS2h8R
CopjZE8G4Vx8NtF1Xggh/RwMlXxka2G41geBC74DWPlVxnxtzGb+pEEKfjWezGNKi/b8psgOHM4K
Kc0Hp3lJzkvlWs0OGkH6HoqY8cP0MxVhYVZE9BfozCTsxbYdjTkIegYfZDHad9RFu0XU/O2QV+oX
DDdfi/XFmJMHffoUqWBcfGZRwA+eyvZsrgOE2xAaphQ0KT7PRyZYv//gs35GbWYqM+2Jj855jUCF
FRdHfKRXgZRPPifH/BfzX1+GyPMB94+9qyWwPRIyl+ba7s4PHN6Gn7qMdCrvrR7hPyB9H2B9eXt/
HgxnGpgsTRjt5AB/I4CQtMs7hdcNf5T6VhIPlNsTUWzE3Semwi02cN3RRylAOYQ6g4Ggd5spzUPd
Yj4ND8sycqC6qnfdzbI6WNTs+zvb3EdfpkRg3J96HvHah4sv6zRZo7aR4Tosht3lpA2Els013iYe
KaLkx4c/54JGVX8DIEaZSPR8SJlpm5tvQbQKlct14QxfocaRoQcajimv+3y8ED8SxwK4/2hWuaKB
ji53MWS1iW20BqR9ezh3LyEh2NlUPkEubZs2cJSEFqXav8ECzNFcKMy1b4GyrQHxLUHo7qq+HhLV
aWU181tDba7A8IqX6y1T2ou91LWuFgrvo8s62ejUjPXW642WAOmXdN3+shCYLnYvaP6mPlsK+ANM
PAWzdGEvTgUTx1DJZKZJvpVk+xlpggevhfFpClDCB/3vjzzBmjPlYPBjOji/MTygQsIJoMQyhvlY
PHYOL2Lie8fQIkwW/b1/abKwIx6ZNgNXQ3fCmR7PLg4IewBBR0uwuaAu6mT3r4KbBzn+bcBqJ2gN
X+UTr1yPvGc4kwzVPOllpCWN4c8X/kyKArXYuFgJfkQepPNk9wmK5ZuYgwOQjm1gLZ6PoU7Wu/2Z
h1fCgVQ+RulkdN682TzeO1Aq/vUtKEXKGvo+K3Ox1i7X70TwJVgj/fOoxlSlixknLgq9+aXYq46s
e0xvVpSAyWvm2AwEZXKLJCpPCpZ52SLODj+J2aetKmr3/in0i2143myT7bAE7WsJ875D7eT1mxQo
FJ0IutXz/JAiWvv8Zm9CmbgYEoWgkIQwlr9b6qduNDDGH5dAYZ2MzTYc6gImSIxl12FDzB8EMUNA
pWTDYFFUU8GTKrXt3qaxX9JQhdHWF9ToR70CKdxb6Cdph8yPsrdjrXK86/XflwnI6RMI8tzue4o+
/XrWQfJ9SZ0zEQZbJph6ROUIg8pmwAAaPAWknn3a+l1lF40XEdahGbZKpXkLyxINH9AcI78k4X9G
TbevPhQg65/cDMwKVk3/cpbfg9Dx5j9xWFA8VOap5RBR43A42AlYAHZz+28hk6rnoeq/U+W0WlIx
yqVZlH9XpNbSxKUMVUv9rCAJBXJqSbKk6DCBVVvYT/z1lR9SFY+hNII6Wi/JyvHp0yrpXVq9IPav
Y9oXElHkKG5aR8Es7yV/wfVNqslbfAC6+XmWOee/eio/alu6QxehA4A8dwViqTMMY1PDMLTDqdKA
YrbJfegoAwG5xop+UpK/5PK1KfHHag82SNStAl+a+emILqle4m2pjfJrcvbQe+LETy9s30jgzvy6
uhADJKW7K48VNi2VvDrEDrKrIxYRwQ9nyZKmJVnTSL0At+cXcb7bh+zVten0J4JKqsbfIv/GptDH
784wg9imGhSIkwE5phRRCzJLD1DZ/Z2/zIs9wcv4RbvaY6miXQMwhNqhdVOJMlshLdJICpEoaIqe
k62ocABHjKo+yp+OwO2Hxjx//q6NEO+1/yA0nAkA8ypeQSJLzszi6kEumCGlx4noypzdhO+C+MyW
fL8nA9jxSIzXV6taHHMQ5badgCMwGX48ZQ6jE/Nz5DHnXIkvKkcVMdENmfcjxFA+bngHyX2MbHTj
c0QJX3xQqr4kzwDfBQOrBPETdKAwnsErvvB8v4/oRsmyPxnTujab6i9RxBezdHYTJY15R9hlYflv
oKVoZj7pRFnSwW1YFEePo640iWskHgriIk5uA4JmHgu+wS9mxzCz37VBhLLJ6hmdcjgiNt1OF628
gxPXIzmW8kT4xNthh0PVQKyD/EzH5M37d+AdHu829sgi+jz/1k5/jmOxXGacWIaKZiiyy20s7sSB
kZEFJf/zKqvIfTJcMC6PEcpxaWJabfrNR7g5ikoMvX+5ZLbgYVal4RN+MBqsBFb2k6CTVwspeTTN
3dNQvSsxD7v5fwhy0k+DLhUsDfGi+rK1FF0TbgtRuvAx22jGjwtcjL+NdWC7lYJ70G8GiHgWe8Nx
y7DvKHxf4bLs73E7B3r2RB4KdbVRjLdM+kXWvGk9qlGp/5BUoviMWm7wX76P+2Ggxdm1w7MAH5kV
WftRHclo5po9X1kiLIQGdnOfhJcx+jz/tW6d2s24WEvNziTkMpr0IWjAwLsjuwM4P+P5kuUGB2EW
guNRy9wJO4SCjFHhgwQU7jDVBFAYM6Nu6AngYqSQEyewxT8YlDu0FaCgiE55GtTA6C6b1+0TDpnN
4VXtWy7W08PLVEwlRkcWNcQ8QA6NEiviKBsOLubsswMkwef0l/p0VFF0lLfsy7SGowXbT2WY+oWc
jkrRT/JZ9ekXAF8vHKDar44LYrz8y1QeDitUSVGTDzT5+Mlj2OsHupbCMgZbc09TO6FAyEjKXXEU
S8gUwBOM8Msq/MApVpdJnUjkHxbHLrHjWUnrn+PGQP+9FNJezzdLaJabaKHglVk+s244al0Bs2Tg
aJieEfnAIZhgt9QoVgDFw4mXjfFADX84T60+KG8fNdqXNKrIq1kT5xiUD9IA3kBuIO27FeA/9iIv
Z+dVQciQk2obp2wOLVcXlTFWIusoRZaLsYfYLAuPv2u7IAW9sMFgrSSJPddL92HjZJ3w8iZgaq9D
CXAIHssj/JgQAZ3dKx2VjjHbf4TZbf4f/rdkz1yviuc51V7uqm5ykYwhRzZZTVUGEAwDX8F+QI3a
CscywdTXPMKXAdaEBtC5LSkKCWJuLs4aOI6e8uz8KhuHbkqMM5fqESG9e6En33Byw0x7J4xxU74z
hFt6cW9Gb+3BRxM1+HdYqFgdvb/hBQEwwq5hO1humzeQvSnh3qKcHtJQ1JB6lQtW0HDnb5XLcnCu
NPk8DZ6QwdJ7/g9zzBTD4ZThnWrkI5fk7tSd/aFKiiRHfiqbvk2A0M70YjeHbG4PxEW6zdFGZP4w
U3TZNiBmaz/Y121sQ2x15kvHfD/k8Fs4dX/7x+qq3VG4iXft/OKkk35QehyBszz9D7bCggP8Ekc5
w1FQFPbLbqtuXfDh6SZuyY/kPRczvfKkV7MsJdtcJhIsPaUnK9KI2lDwhwpXm4OpExXfipLKicco
ck5g4DuAZPq1jsnhPRpGCXsOBdGWpfDbBYeB4YK5xFPg8QgTud9EyUuPE6ePM3RUiS4QCuNGRkIT
V0iL+c7Ml0NhMwt4o9aOiJYA3jOqKOvWkwECirjVUHn5mQXzwRxTJZrdEgLhP+938Q/ToyEmlUnt
3H9XzuxuinjLTsUL2y8Frq79L50G3TW+BgoBnnocFlOrrGEsEWB8oRYvFe3N5r9xDsqbIZPJgsSK
rtgDTDAk8cVPr/TFOQupOgAAjHE9ol1Soy7Eec+WzXWCFZjvgsrPNjVDv9uGQu6hIF9jX5Zm98++
sXvhS8yqHLUXQL8xTxuZPY2XTA/af/ivLFI2OKQ8ROS/a3fujUWxMfC+s8HbgGn79bvETsqBoZa5
B/ZZZU0KJOVgXQ8GMJNw4l5YwTIwyOqxWDG9A4C1OIj3e476hw5mMqUKN93XKW5GxyenZjexIeRF
v7FSusUUJ1NY5G9o4brpqweKG9i3vd/k8YB/2WD/+hlM/b0LZ9CyhbHvtFeihQFE/IB3zO99eNBw
qmW0v6CsqD8KKoJnKkx2hFJyGhAonNEVzdqhSo+ILx0YdiWQKvgC5wtyRdCXGKerqeQt/9Fw2Z+J
gNsPIy6rY61b1Xu3QI/HT4N5cUOhobdtlziV1u+dJoTkIWOod5gUFTDQiq1GA5J2JjMEoT9jwVco
2eF/qrNoTPJt0Vm8EyV63+9LoQY+v4ZWQxAQ/BhXo5An8+fKr13Vsa/wuyxOdEX2gV1a0Cn5GsGh
zsY1oxkxZ+vxaYyKftWFkGzRHdVIlOWosFJ4qX/VSE5bAMZJuIbc2sgaEQNd7fBeRf5PKLiJpteT
lrDYBprUvT4ReNdiSHtKkS7yyPTkt94UUize6ukikfMQfiROjNo3MGPF1geAyykkrz7Kqbqp8xKN
wb40FPNyG1P9uJps2rBJT03oA8KAEBH3U0KfPvdsRxCY35CbUVwGYANjIZfxGrRGOvygt2qdLxGw
VlwE3wQMRwgITiJIDdDJmQLwwGebcthG8YB+cW8X0RfzPhc1hcRCzK14m/VhfshZpCtfw8+D3l/x
rB3GryIG1F6XywxW38TDuPEDCmhTMR0+iXPGmkT6+0TriwsLP1kb7veDI6bPjojaTskxzxY+a72o
KLbWUVRnB/09YIwlOBTNFcHujwnIQ4q1p8l5c3wSsp2KK0FQdg3rzbbG+5vA/I3Qnf1CUh8R/Twv
gCD5lHwNQlPyLlC/3nAFyaqO7GyAwFIruP3HcmnlWwol8nqmcM3HLV1eLf9ZDMjCrkBo93PteQxx
ELzQQvbbo9uhcsxS07hvrT7Tj5BISlChR6bO/l3gCIT69cGitFmYio64GWwssb3tZGiud739m6hA
a3HzGVh/zuV4JGxvcmMGUerNnHwkWvkhTSzxDEpNOfrXv8ZTrUUg+49RND39Frcg1SXtG+aaSMJC
H9CXog3r1Ub3ayThrvjOLnOprdsXCB916Sn+RwKp0xG/cJ9NG8sKFSIdaqEhyeruLOrRYnkezjLC
c4m4z8ouOp3mGSHT4UhAWTCLzatFRY8OBmbPeACSA7hDLkTfZQFIN0520aNEu2Mhd+DTIv1VDWTW
4nPuVhWI/oBu+REc5Vf1rJeqL1Razdtpr91XFLLmKdtBSpcekNB2p41cWa+vCJ8UmOcwqjebB5cX
9YfTxkN3Vwbjdd88wv8hG5TK8zXY7kFfu0sTL4iHhicCdzTuWrzJsTJgWcZojWXYCsV0QfM/E7Yx
jZntmdnsezGkSQF73U/6n4297jxyH4WPAeZAhhcaFr6DoBfI5E2aCEcFfvsXOMrrcumncw0NHAA0
iYblJJ6OiCzz1reLh4qAb6eQFh+NveSZKMv8W7av786FVUI+Z00iVNRKvxZSg7sLTRrUgLPA2Bf6
LQBJAaHE8bR82YuL7QANiEb8CvNXiLiDSO0/uvwNKvkAA/qgpAxLlqMuRSSnXM+rx+XYNt/NFUS+
FYruNNlwt8sXD0epcb3K6eqjSHkRooSxzBYYenZx7ouEcpU75KZIaH6DuK4RaiMHXWeVXnc7pE6Y
2yE2qmLDlUi75p1j3NGWalYOMR5+D3ietn8Acdnp8GkN0Z9f5rVlPLxiDC+RuId4qLi0Zv7UvqxS
+eMiltK1MIjJwlIfGLfscHqY719aPfRu1OaOfBJ0qnXm0t6jxJBP2B+LsLPzTDTE1Qh6XGaDfJX2
f2XGgQDXdquBUejuURWjLYo8gVRUF3n+lJOo2RZFwg+Q1eio6fm6+CArUDuLRUMpvTqZit+30baw
Naz0WHELYP5RTX2eD+GidEaMEPLsI20I+VyLRjjA3RNjhD1BO+3pdmyRlLJ0uVXGNjQUrJ8Y5Wpr
DsVK/gKsWUYzBzTKIIs1MvkjhgngkizGi29x/cwa/RD2SvAjRx6/McScuZqQjdFOdtvQESv6PPaI
c1XbCrS7gL8zblbqI0pEbOO9v+nHgokMEgk4TQk5YJx6bqgxUVGaWSx7AvK2u52dkF8cOiOojzOq
ccOYt4f/QXcC0xuyfMA9QP/7rLGzyh5iElALttbt3MDkspLbvnptrjifJSi9hKHBFt11Q2XW0wox
ii0Kh2DeubAtY51kDmdKFgBFmBHWKMvQNbfakcg9xBNMRVbKEAybU+gisvzjreS5hsug0k57dlJU
w7K/q40FYsO4NRjaCUtZMb0RI/muOAJMVcxBLvvhBGxlFNbNP5z0zhQGlOj2WeYEZxaQAvfBokyQ
jORcjGOJvNeX+uPUfV9cziqE8NM625gqzbXKHyxjaoZHE5kR/ZjjzHvN94WS2ADZANsBeRZLYobQ
Pp92AGJTdUFRP1x8MY66eaSwkrxdmTDAtdx4zzQkSIRL/iMKb4f7Sx0iWrcVMC7b+XUlAhgtaSRk
NJe4DLfJb6bqH1Dv6oHk5PAff3+cqHyAvPg4I1XWyHVZSlrk88zL4qcUbt74bLWL1rabErptLALN
pUMiT6mjEIfQ+7Q/pPycB2rOO8V3R2gpy4CrYly23rBzmk7WFD3kodQJSA7klV5fnpH8FPw2SJPT
M9oxG1qcc9DrjpoWp8IW0sM6ti2gcppoy6iMSZX/OjltpqPD3GItsfW8VVLQ3hSMJddlApZI6yO3
kek+wsh62C39zJ8czZ/nZkaB2lznf2QHHkIaTIEX5aUTc6AOsx/Ual2WwFCh972CNRQLS3HI/0M3
hkG9JeuPsryUVcR0dlf1C0Us4YhljatEA6uA+6KYycF9+cbh4CslhM/hFXzyzD/HZQeZfCAlXVD1
Ec6NUEJybOhcBxmOqB9NkXwZ6bsw6/XNHYKJwACb7lJS8p+OBYvUrqMwPHZGk+I48ETnRj4hLSex
z2OQRunqwyTAh/sXxnw9aKlqChr+G6TUAg3pd8LneQxTqvFjrP5/CcAJTW+QLUJdNO720jKgLGXg
kHYXywX/dr2peMrsC1r+IhOGYUrwpn+hIzv0yc7BuEa+68n0VB7T/CeSsgYn0kibRqz3zyPv6oIH
rAZxeUv2s0HsBFW0MharCTVKc+gCyIn4GZ9mAAVtTYe6Jf7g8dOdIkA2wavjHPADc2UVcHW+mHV1
q70SrcxSpLJxSvpC09o+snU7v53jejqVmiY398eV+9G0jIZtoDL9DF77rbeS4/rytM0pzMLOEVRp
YcwrRJ0VHi1nEJVOdyULypc/iIX4sOnakqgaivEMKMxkaUSrc32Zf32itvTE8wRR4VpM1EJnraPP
ECpKt1uTcq+xGorKHP75T1YSePrm4jZJo2tVccSM38vPJK/bEddC84sAboM8YBThgmm1xPjruMzq
v3/4lLixXeJAUGMbU9O54PwEHJPFSto7si5tBbkxlA9fEhk5iVMGuZ0H8WCrstJiQjnZoJvLI3SL
xzUmd3xXq7uWFOk8cfXaKoHYsE0cWo6ck4ahLWJ7RGggIkX789tro0/wYa2A70Zb0L1caeTB6DBU
DKNmzqlQtOI8D3ZOnrIhHajara0pJt7L+ot4ot5JInqBK1WW62BbRM7gauqdn6/k13JekgM4NbvV
qDqEqp0FTnsiq06HATKnTEV77rt1W7r/CRCeISs8yFe1WQ9H6iNe8l/bZiW2YfzwHZBKRTGVY7iG
ICVzFXlEekgADedkwSoY5B2djSZVnNxK3Ukivv7Hty+Atg4fhBdjkXsAgEUaQ0bdJ8CGSu4A46hd
yy8iE7rTosPjqcijhFW7aept9Bs7SNPeMPYmt6kSJRuKSrnSxBh65mXWb4Xdg+Qgn6jUJNY2GHED
5cI0Odmeroli+N9Ufl8egO7oRbEleaAXbf722x+u7eB5B+D0TNJtRIv+7Alf8gekpAIZIb68VPDU
UUorKpOQJ9PhqvHkI5RTFCNyvlKrv+pwujAQqn71db8Iswan5ltmNZAYRrGcQdcoFXog+OlJqoqH
aV93emo9PL/BrYNl/R+ApUWJWsWICym4hKEYEyFWziFr8fzGH0+I+iKYBvETejPekkvEFgaav9WZ
UhpW+XCJkTIDGhWVkTMuQ1FxtN6m0wvS92hLyT4NoCTj9WrQVK1LwL2A7PVHg4puiOj7c74lD3jA
LlKngbVc9cp9u42ru1jBluDYGIYTG4v5oEPK1sZiYbeQHMCMaru8TQZEdiNjbLkHdS7b9KQaj27a
TX6M8p6JjIfk6Ya4F1Im/Le83SkC4HreakT4DZUQxQsQBgRpCrZfnDEHXJjdY+C3191IuR4epDyq
/hlb0CPhZBOKHF0WuwCT8g9ZQMNOwgCvYAUGkthR818HsiWJzZxEA+W9xNmxFmfI+nk6If4D04JG
0sqy0jZStwTPkUSjZskxRAXW2OVebezUlI9XnJviBx4cyJlm87a2Fh2POon9ux2LjZ2eGvx/LRnz
pwzMashXHmkpmjAGrXuegHYaH+NDw4BMZS3maa6g7hsOMF4XX2s53wyQRyMXGPoNbIwonhAnfA5a
ixa4D/g8jnCmkXJT8nIPPWlpYm9vq/O9MI/7wAusPPIwaiZRlJiDGOhJAVJwPmps0hUE1IkPzU/R
TgHf4lv3yxhYTpr9ntf2sDhuBTOGRRMZJyp3FCLLQT/1owZCfl9O7njgtTWUUSWkDbAfHbxNR1sF
eFqn/m1npZyESqtXY3tMYSasTu4gcubL/CpF18DC59EGG7uBm+4hnNbyDSr+dPiTRDHynHLfqiCt
5gMOL0KdsVOcJ6VZnt5gLroUldl5F0vOUgNksIVKHwZrOn1xEOi7Yjo/3dAe9ZbcXWdhN7WYxSbq
Jd/FIJZLdXnYYuLHGL8ZD5i0wE8YAsnFb7hIk/kjSei7DJLSmxd0vpMFE29Q6N0MGxN6Fgsi491b
URda3K7iP/WaJBRLAfraN2WIIvJzCmEM/GbtkSiTmYscEIN95dDwFg5DcOGA1sf6Tclg7d6qo1zH
nepg9zsVK2Tkf8WJv3vHbfdIOQMoSGCleBcIjrsxzCjesGp6HAvc9YxwzJK/URdjzR777kZA9e60
noXoAhwNjZxEaYHxLE1VrPaUSFnDEla3NZE3OfD/COGCgdx26czF7My3SjslOEZFNocwahIMEhlk
mpbJAXdMGOdqbuz1GabQDia0wQ17hUuokvwJzDyzViL5WCx1Qp6RjkbpOTdHwPO4RPwMJ6sHgVp5
8f3isLmF1h1JdupUoBay0GPCoiG7PGgGPnBObNPXyAD/4UUBXcO7mHjjchYq3xV+RhR/EnGG1NAZ
LZzzjbnRWmtYeocjNj9HiRFGipqWGv9nND6KN+rVNUevQbeHVr60CCYZglRtI4PuxnFeznazPnTp
iEg/o4sSq6SxColDfR5GSJlJ2Uso8pYR1qMHBGvzv9hHobqqaziVPVSaL4OpZFuWpHeAm6ej0UwP
9vKdho60KMZI1ZaxBPi/krsHyQqqFIqpicko5pTfkOnHLgKlPaL/9tCaErmDp1JmliPQqNsWXk8k
JNA6DYdismAB9c7juM6z9NXKASLqmc2ITMd1kFopQLq3XHDVSJzlnNmlGzNRRNFQFshQ4AG+IBuB
Suu3pRuCH23SfWIp2ZanDLwz4sNy07T6e//7lOi0cMMqE/+wGPJr7+Woq4tXCl2poGRtycFuDSxB
fjs6t26hCcfVk1SGh8EHdrvwKsSSL00PgAUvl3ypRulNeWrg8TgOFnf80bnWIdeoZXxwTKD+W//r
MYqyZWn9fzoLyFrlFAe4eaKoDGJU6C1E/iEiKzTIMPX3dZDXDuguBQ+ORU88908ZOkqCM2wP50Sn
qKYWjVVUNqz+YOz7zrBF+KIjKS1dVrcdQpTR0I98/W6lZ5usjJSrUtpMlwNHrKsym81OURZeL9kX
+zSUhmfAqjSyVdK4WhdZKmNwFnvEPlxfYxhJQXBtn2bJHuKjGKnLTCEkCgKsKg2vkaq4Cp6f5+qj
OYakgkUqSUs28W0rG7nHTrZrs+I2t4mCidhEcqYEpS+EVDXBilvKcScbbjvu5o5z1XACKb4p5YrT
LdkxNRUo2kVEvlYkZDeK6dswfzYEFvMSew9DPlVeRCBUkGlWkczeLNigWy33A5MMPQxEaepciuvR
ZQBXztV26HDmOSeDRkuyeszKYZBAZXzt/kvUMskCk+ryUtGP95i0dGMssoV5SuefZrc7NgRLdetf
QFeketW8P9od7D5cIkbUImgGjMd8/7kC6QFJ4Tu7Ce6m6yMmpTZfdMmJ/Du49c4/EG7GjiT0z9Lv
N56z/h4omf/VUYjhrYkyi3PkpSxE0Fbk9tjyV48+H43NzQofBgwL9yK5mSBoGYBgAVn7VmA+BOyC
9Fq6+i3yvZ1OwToqNxqdlzVO7G3FgkwlwzKmMTueIuML1wtwT5P6v1bFIP2DnAGx+NUxYAKyXyQc
xWz+yw0Lpc5KksuSe+e/8h7mMMZuDghyhjGS+CPwh5xJXifjOtp3pwjaR9wm1/lMSncDLX23ACV5
TTbayE67Gz2SgYGz6I5lMVSwcoiGsdNZxkAk6LuYEF0h8u4Tog/CLJxuoANYXYP+mZwPaP9WNGQb
7kP7+tnaG0bF0oVCeyQ+5MWkhjclzUn+qaLXUFc1LWT47hoFSAudzeatNJ0DNWVniT+28OMcJg90
KuzreZ0YcU51fznjRQ6xnvgBY8/LFK06Xh78XNvIhwBvlNuOoJ4E3MudR9O7Ba8h7IcRmFUeUxTQ
12XpmtCgP0zzO7y4Ll1dKhb21lgNptC4k/JzJgmpaZo/zNl3M9Ils5ppGX1TIOFYX5F+cB81TZJ0
h/QdVAQmM49Aqvr8x5sHOgoo+wA68U5VLRI5hGLB1grxROENGiQkw77evVUACylBBdLgirL64MJv
B9j/DTooeYl3eBZxv8gE7Wfl8CpazsEs2/FhPSYwJvi1KjRWFTED7pLwtUXd54AtBNXgME2rOgnP
0EuH4/UOsPQAkzGe9YVLbAEUfb4b1bD14fSE2cm/13rHw0pNNJpiVdn9vEw9Sr6dS5+r6J22r55c
y5mtrmaysU4tcfQCqz+FhbWx8qYyj1xMdUZVmAbGkAbvu0XceY66BgnBna4ZU26UIfJqo0EVh5bq
UJOGg9fSVSRnEZnBP7/W3EoFKVBo9mhn1ns/BW6jt3Nzhp2Wi05F5I2mpciLJQ1EWvbic2Ntm7wQ
R/VmqgwgxD8liS6Dovedo4XXorncZvr3vSoxgdShFvVzXAes572ToGbaV3c1od8a89UipKtNFKLB
ZucQSeZr3MiMY5c/g10GglfVpaPDEKFwg5wkDJheN4Q4MOa2pcVhUHcF1ri8SkrZ8o4ZDkU+hgSO
0gUE1u/TDk445jHMzNCzSM1LHA3m+moRyF8jMcylJDcY+ca17pvHt5BgZ6GcOAtDzp3WQfDSAhD2
tx1Ao1Gw5NSch5Vlb5wXHRGId5MYbPd2rSURTnLrjQekVAVIsEDNMkQv20VEiJiuO1p2Y7CUw56J
GOBJS/VkDBTp4SWLTLMuQWFQ4tvcoIABQFJ3lLar2PiFkjP3j8DtNhSsm4DDdhlBttw7hnmMkRMo
Jf1fxpMqMHextGC2O327tjTgY6TR9m2GATqwxZfJCVLeVCDBbvRCAdU09FljaM+umJhRX7ydf7Yz
Vikx3skfVxisX8pgQpabwY6qZt7Li+hepwrnxtPJ7kL1RouF4FjfIlRFsYt1rg8DDrKWKKCzo5vN
23YRVWw0igBp3gK8VCkfI15nSbWwFjhFMiQqR7leEyEa+TiNNcJCWjk56NZ2SbxhGmMmXn3TyAIj
lAieLivxF8BIzWsrya/ZR10JAV0agU6MKg7NvfAlj3CslKwMAktcO3DVbxxDlP+K7sYDyLqiHufn
DjJsUKbTtUorXnulaJnL29Sw9n+C7sYAVLPA3se5eRfYXiHumHlycgrYwsVRwtqWYxgcAUAZa9ew
pYwpWeabvhZBhhhsqFiHvSZLXox9LDASDksNMq3ybRpUqOj14EJ8JlHAtXWkp6iCUVNpHuLc10JK
K/fXl1+eov9Nj+Y2lFI2ryzRh2sqfCr5EPC1JXznzg4yS/wcVfm1FXU+LC7qiLI0JGnTQY9kUQhl
7iP8PNNbk1YAFYtA4P+hZp+ZPFXMc0q/lKfJSCGQzcIcvMflfLUd0HqFZn+Ln/SRAKbrgAGJVYwG
9WGG4VCIuahpLM6lyGgq2kFK7ADpSdQl8WhQVBWr4h18pyaCSXTDCCKk/Xv9JTeiOPLHBwhZ/TNc
SLiHfJMWb+UfMxko/M/TeJGscgoZWq+BMNZKSlVLD+XJ4SNP3osqHanSUNwzl2Cw37i3u1catDGq
lYKu5ZMcXp4Fpu63o2DYZZSTBRVv7zC5muDS5W+JGJLGjMfPqgO8akeqrgr5Yg+nUGqKiWYbKvSI
IIzoY6KkuqOJuQ7yj/K7LIRLw1WQBg70IDsufI1KbwiPDxoVzGOOpgWM2+Z8jQ1Rqh5xPiywnPf+
2ZLYpPRVegzpuGVTVWIekwPCqsUgLDt9g/jFYsN19mr5h1N6hoRxk2ctCISjQTVaQIvPnDqUoBaV
u0LaZdyrbsbr7o4kjIfO6b8OIzmofDl8LhT4/VWRNBFRHPFKfYrH+CnZQFwjEdNaxca70tDPdSEn
dbPvD0Bsb9crOKxA40RfVccG5KXc6wpZ79iFpGhYBUlYSZ4294T5KspFEw5dpNteAdKtmsg5ML/M
B6bWRgtjIyRluX9BeKZM8XFCTINfreQqZIsb5SJ+3pb3e/eqrx2703yiNQcAgU9hpVCaQqHACOhB
vP2womIWLNH44dXERJHmdn0xcSeqlO/9KP7RchNUqU2ikk4mp4RQJ8wW1PWtZ/fGV5sg+T6utxne
H3i0eOYdQrCsdC6mg61BFtDkEvf0tPtpH2lt91mXBrD2w0FUaYk/upf//UOFttySrSMujiDOoDuS
WztsSMX2XPQESSXtFL60KZCQtKpO1NBmDVsOETjF8hayXNoB3Msze81gvmnmeTDmmXxRLvWvrXmq
1Q15PmzUAviYsCRjhGQbAm/tUIRp7lLjw4X5L68q6UZbNXovMRM3tKCnr14hzd+wQDXakL7yFklY
L3vVNifZrh1UZ4X0livOWo6Gde/rPFWbNlTnxriIvyS7hZ3jIpOGHvYMMFtShiJ0tm+O+0ZqnkCo
dUgnoUiYC6Sm3lzyzE0jfX7y+jIFvyco3ZECqq0mvV0dto68EIs/APLGuMonod9CxFE7yThbvxl8
32IL0fNfKfKwx6uqeaU68mP/vr4RU2EmHqmzktGgNIJm9OgD+xUnsP4LdYKyAVaO+kkNIZhL/+9d
Mesr9tjxO/+kIvEcWxsb8DjaBwhw9jHOvp7CfhoiaHWwDdZnPILETxdqdioUbhRuSoO19Y/jgEFE
6Be3faM6LcLj3xLxQB2/OSuW+KBQ5J6N/aFMORVaLJ2B+gW6uLemujxbsI6MKXTJJ4HXhOTzZaC0
n9ZQH1lvOv+fyAb/YpAHnJ9xp9X7wB3CpP2jVajlfzSJnaSCjLIeH+XEW83s3sMF4ILvAIwAhuyo
ZrcSvijWUMRUUEMzOL8gt6oyUyKQTmjBsGdLNPBdwKyzF+TcKTslFkb95c4QYXPQDjra8vaa7pOy
Z8JqeHWvTgtQCVFoxpIQpF48Ij8UQJGlFg1yA+YwhiZMPR0jJdMsptjqc8eNeWNMOd/KMQgMUPLG
F57C3KpWoDY7nuNzpnFgTPrpu0+wFp1IRGAHQ7kDp4q5doHfwtHyb0Y+Jqt9Ip/AXcR6jTXMFUv4
bu5Mi2HcHrQXpbNCHLTYF78z7MGmUwU0hhI6xiAP7s74mJabT5tfywiloHwEaeaPCeN8dbU2IQa4
cV8GBQ82Bb01ISPfeQxW55aT1Kf4ltRebiREYpw/25Q8+gVNr1RNQIBdgz51/XM9CX6QJyUhBeOy
kJ2ppv34q34YMpzEWu++Y0k/nuhfsvr+vrYov4ffyqZl88dlNKPyOHt6H053hioHsSuE+5oxFNjA
e2CmNLXq6cHcE1SFdh7d4bvWPD28rEg+mv23pEECvVvGfFx+gcIXvP7QHZfAtcqtLavGS5ocagqO
MBozWwLsA0IMa4Qer7fjY/jxWR4D1f5r327OrOOrp5QKEXpsQ5/rCon84ApeyivGuqz8M438eelc
9TOJJcDLXfum7LCStwIZsDTP39ntvmJOZiBKX8xN7K1g8FOmIcagBRIk+xoqb4NXRqUCCU2lUIEU
GaC5Nn9dRAuTGhTbqwujAknWGo6A3LfRetVXsHuGkifYT3bkKehGkm7bcB+26/iga6GNvbH3ZA/L
cEzEq+D7UzNUxPHnrxvH11VpDH93JJN4I8Lf8Z6sLHqfAGmXRhRFW3oL7cVRM4iSbqVChcIglOzf
9cNOCW+ERV9nYNLjpiguUe+ufccqcjOiln9DzvH0kCVildjq2VDzO5uoq06ao0aleLeEvw4CfA7R
GSwK5BaNJXEzXbmVxw7wy5dCUt8aacMO6TIPT4MY72muAAcAI6BLuxZqnKGlN5eqtZRnXyAWxgdd
RbeR/Zjx/sNmgMhbF3psHX0eV+PdTiHsOaoXD8a950VkDes/gZp18L856OjGyIFxmwr+YPxGfbC1
mP0f5ZlQMUvzocfShsYVLmIb2kq8jiziBIipQZ45sYU7jXMMs/m3zQkjhbl8s8TkDMt/2mWkApY8
s99qAP47tOy9a3wWOF7lX2hYul8mIappuWQlP/cN1yRDmhHwObK/ROPju3emjpZr2qHZR1YP6BoA
h13X/twtcFxHFQQpK3PtWsiRE56yYnfUv7DWTPvWE+ZkFYPQz7RVtdKKW6XB/2ZwlZsJLkfIGeSb
BrxtrbxYem0NjqRtF+aJYfYh4lzicNV1Ri1OVwABePsMnzAGCSWR3/cJGe+j4vfeZUKnqL8Pd3OL
K9wDGri+BVmeHSw8cGefPi0cB5Y1JtEwBfprBQVKwePvPZk8DYANIAbGdyPMoinci+4TKyR/w3TT
MPp+ZCScONetve/wZhWwP6vzqrIkRtbVyr+zxIq899CMuwA2ZlEyHM3QKDnXgC76Ul6j9lNBl1pK
YEl1pCFyN9hO1XeXWqUm6EdVCO0lnMGkp+V/nDobTDwQzBdR9bvBgN+MpZTkcgZ/ZTSGDeKLb/Iz
LCKHxD8tMuyHjfoug1Z7+b3O7Wbq+F7Fus7irT/jpHnjdeubFv0b2SSC4REsBET0QFMNgdFJ0RUI
yGcY90EA0JM/+7w8i3emIgOi/nZo+s+hMrvAMQzmdza0hg0cU3MxkMKNX31TW77SaStvS8uc6z9t
zZLRFxlTRhwVH2S4lYsmUhK0/CzrnTqyJoaEsi5ta4bI9jXFMQM2QndV8yhOY92o7O7/riAC57GF
/TvGjW0kf9wiCo56YQV831UamV6VApyPIFFknCxafw10fFDQw6tv/rOU+8VmuPuYGU5QSa3Ao/IO
Mi2oMKu6+fGTDXl2OMyyTFVmBdUezhp4OFrGYztnatDdiVWnJXDA+R9qCjHJ0LZETfFBrtVMhxvt
NIZ4ARDAXEr63aU0Wjxwyuo2XbTcRVrgLqU1yHnJPYPavXW5gyyzuap3UjdAieCrJqDHRyQf9JoO
b6cr6fdQFodFP+pAB9eJEfVduIkxwROG/5B2gXuxTnnXJs0OHI+67E6ZBFjUTEplOyKLqKO/mgId
/DH2vvvEoTcyNFRYJh9bNxLVS5q+bxw6cGOkEPzwd7dN5LbhgBrXG1StMn2LnSpW9a5fIrlgOBQM
2FxyVAOe8faYjNUVxsRnNyS26weNwv3An0+L+l5jbdylG31vxp+Ljp4aWR0JF5IhP92PY/7o60Tc
wZljgDifs7/4TQApT67Hl8ZO/hlv3zx/8sYmSh7FiMJkLzgH8Oq0B/UdB0Gm6xVNEOzuf33iNmMl
fGxHAXvDHRHTDKWD7t1++gi64E1G4knPcsTliVnZ6qaRbfK8Fir8lGy1NrYjdALHCMwF2GF9XsEd
g3Plqf9xfL22ofp2Oe6dj187R6xaOESTjYioQP7Tg72C3CxVEyO/mi5Wn02LBDvTaSVnIt/cxMHT
+V30MKMDPoh/+PtaBGP6kFSWvLKQRPPuxxJzFcEuSRwsbEzimExcyfB0r+1/Mw2PSsTqimYuqWkr
6V7XspFBkzrsHGU9c6p328TuojzX1UCBG5Ct4Q1gJF6KPzOGftSUXchAx4YpFia/PLiLOpGu4g1k
TEltdv9vcnYax94FmlbwEPo2c95crfPZJnniw/dqBwPiWhRG8eRerY17pn8Bih/I9AaxOZOD8xZm
t1a3q+TXxzcxKbzBP+Qy2iM8pBkH5qEz1sDD2gtelfpx2TiKcozwEoSCw5JAL6Buw3eAc+S6hEWB
aDChPB3XFBhugdgFhk21jndU6MFtpEnDG9XbI2kVi1zqDoj9u7ZwDuTjL7IORpAwESxMkMdej0tt
YVxmy2wsNORoYT1G6cgcfnvd8eFXV9i/YNFECtraozphEtdZZPjyYEhtxsIvcjJtEFW+hrLPY2B3
Z8TGlWfwsGEkb0O1naut+KXivcDrYfktafDK8a3BDYnXG91nyn+P7EyXvWBn8wpAWE9FDkw3FQ1n
nLCBUEeZqFtR1zvdyh/9waaOZHRhw9e+TsCv97cuvCmL0W5q+VUqg5VpTArKZfCI51r37hRqzn/F
ehzTjWMQXDSKv36FD3z0NEOcK1I/5tyCfi9qEgOdjH/eUmW7hmtS6iWiXL/+M1L33lkdKVhSiGNJ
dPkHDaQclN/AGsh/951kFcu2PwO+l/xXEPJ2hdMDtfWMc+XWXzDWBlJI2OaeUCOgFD5aHgOFdR+0
tsOcJlt8tY3lqHKzBKkdY88eEGlgWcvbF92dTN0z+Js/QvNrLkGquwbiBGmmgzCZYSnNo6htP9/6
aMFFBE/Ae63Ob/8krJ/8YNlu9Ydp4uxZGQYia2VCEp3F5G0wLg2KJjj6ArFQM0dWzutXQprltANU
2GGNCWoIOVnESjjjl62V+iRybFH+XFFzvgadM6nhjY1i0jYHvVgCJfNuGgIBv1QbIbV54sTRZBNm
a+iJqM37dQ9Ed3S+HiMRTHsO0b6dAB8PJPlUkO7nN23fiUSmJPDYTKGPdyVcayOjdc9uX99gb58J
TMl2MxI86K6URn1KpQagrw9xFQxyMlizWcmW56juGwYjvuWhXcY1rPetbUYbMxoeXxQetwGu/mIH
rJziQ2OpUSNLsDuh0HIUCNv6XgVtuKJqLeV0mXDKw4EtGj4cdw1d1iGYDBVfX7wYMdATtLBAbyEd
uw0ibMDzd5J+bOCgG1yb4/v8hdLgAtMehALMzNdjJgJnaLMri1ApJ67MXUQgWv8+O3HjCeYDI6Ye
pfsahbUsRu4tIQhzezETHwQogvQcjiE/ySEjzuJX5ZhyRjegLku8ATxhQrQs7ktqMR9sbSod65cp
qs+hNk0LITWL7X7E73PynMwJhecTiViI4llRFB2IibJ/VwFkjQE5KHzy2HGK86kvHmaWIoh0JF1z
u2W3j+JqJ+Jys3lkYOwatP2FGPLwuFq2Lp2HDPEMTHDdx5kBvbtO8wP1w7CyRg4Rw/G7rnfsl+YN
yglAMpVodHsTNg9Q7nRWUN7Y986vO0A3RlZyrYrXhToqEdHcSM16WbG8pYmXHTK/WfSgKmSY6VXU
jfTEmI/9/AJKrgqPHCbkXnNgdlEgcv0eTIlgs6OSRg7axquoF74uzeAZq3fRSKdefbs5xVC2KV4n
FAFNT9N6SfzZGwChb7YlZ6LFmXBD+xhKqIVMf27JU0P+lGE47u5GxMzl3mjUox6y90jdBgT8KLRm
Hw49m6s26ZnorxxDcpuLCK1vA8lPg3u+apKfYO1ToyFvAragWXYgzAeO6Qbk10XWiY92dezwZjiq
kq+ousbsAPdculU0psvx3YGH7L4xB02HxqBNvp2xaYuR3QZpwSsn5SfXJHWQfS+iYuWjlpkZd6sd
+MkCcpLvNY+25AyPrRzlhCh4kZfLen/GankBM3YeFzI3wPYPB31Cb5lN1sVs8G17zFp3Ld320Gsi
gV1JeFTTr6G4qnelFateBTw629Gj8Su2YhJXsG7cGp/tX+C3TI9Ya2+I8cloQNy/yPEY8DkQXPgV
n/hqfViATywjy3M0TbXNY5LLHDBaGZly4po0ThfX4fb6euwlhMqvj5+hAa4guFRDPlOAAElzHGmC
9sX3oSbMFP8FnWRBQr4WR/sklcQ+uqWsG7eu66kqLDtGqZSTvn+IG9+3rO/Bcq5fTud8ZqUYqyzh
triQYffo+NyeXiIHD8/cJPwIiRpUxyz/ix9w+T5h2ozW8v2NaY3VXlagxjWUS2zUkFg+Ezks/Phw
cpQnYHJ8MEO8GxEeEk6RsgxpVnSNO49+oZK0c2wvMby8yJmf1WOqubDRUW5/isBDXSKIsLxJ99Iz
hHhXotL8TxOtEW23xy2IuT6YRLs+F6QkIBbSwyJVWnyfdgquSBmZW1jTUDUN525eYM3S9mOejwkv
9KYvf7uQ7PQF4o1d6Uvc4ct8g/Jj37SewpHPPCJ+PZouhIabQ1qy65BR8JFp8z79/y65/J2nbYBG
gxqOoTr576KVzB/DKAcZsDQMsHREFIcDmilCn4t9/4kl5S7MuYN5EmQKs84I+55HDE8MV2i70naP
t/kJBWuGxImESASDBtiwQKCRIH2D1A1XUlyYp9B3hCtvTcRkBAAP0xoJcillfxTDxjJIaiyS2LkV
ZnIpfUVQS4ltiMKi6EPHvkFkx7hlToPq5RooXYUZq9NqEnswU3H1ORpw/wxl3FlzstzRPKVSW5Yu
T2y9Gi8UPDHagLmEdbE7113CLgQ3LnLsw10AwdvPcv0m3fcQlegwkGYDXroCOUCAC2vf5MYNioz3
JaDcpsnwjQtQ8t3x1g499+l8EjY3MY3B0twY26RMxLfSlWj0jFmJ+7xTi92Q4gl1VlMez7kxZUNz
dknbEL5ibpA+SvUqLUcfp9FSrqk5CgW7ptj+wWbrvD16HOqmq5jfMJCQZfQgCFlTGCgIM8Y0rCk+
3tc6IT8aaHBJpGZ7im0l41eEsF+QqiEXlo0//Jg4v4syNo9bLOHhpb2D+NTiWEA2amQLFh5GTRMN
xws3Lrmgvmr0+T7hjuwSAnJhxaxnFEMbjsvFnJ7Qu6ibdAnOyHeFOwjZsfEj9sM2bzn6fCly3PUF
pywEUp31oZRvVkXNHk46L1VNptD+ztQ0eqhzax/vVClp6ef375HuJskULS02JAdlE0m8RlwHO6fL
fLC4r1J1msVueZLN0ZieVawsEFbvgx2EBRrrL+7C1TMk1CLQUZjbUKLlpHZcAXcJvZh5ZnxOP7rh
fRMbDXiVTulNLKHC2W0gOVryQXFa0OqgRBu3LXFoIFzF9WqWIF83vL9UKvarjgc1g+/dPFLvjkKe
E+xUKT7vTzlII6bGQIbCxWJTqw4jPm+Gj0rSQ0rDNTYv+W2C00voVlSdINmhUZVOk5hn7GQaD59i
TCXDaOk2qNLx1Z3MlOEdaqd8LSUCGCNUJW8nSrrbFQwvvYo20QQ7+6w6FB6n6Al7VzUUR7ujcqaz
nmJ/bAX7lWaU/R/19HQBXaUOv0k8mPNFalE+7mtZQaXzrCyNtqDdg0EwREr6mxoBlKf9SOa6RF+m
cCE4fpX9G/97baz5n4MEYuLFJ6eeM+vVHJly88zqc1TDNRmJ6QgonKYaTnArs/KHd/BaIv2PG9CI
s3dp+cZMbuhlf5O05xJ5NI0ZdFKCaUa7rRMtvwyerVmLy/YvjVJp+02HOLuFJpfTECic+cfCwnt7
8tV81wIWkd9Mhzf58pbNsrgfCXs6xhmf08EUvwVvHoTDOTJBi9l/fmuSPpSgBnPWpGNT7tZETMFJ
vbKDktUAd9hMQau9HDPWuaoS9Fv/xmxKgHhS2rg4r7+TTWgVdGuXIJpwdx/Hdd9tla+ZFJCn1W8/
Cwox7SF8XdHiiQsSL1gFCEy4byL2o1AVrVI0B0uIaLTEYsXohO6HIFK/lRCZiNLmNit/hjG9D6Em
Mg6C9NGEJvYLJBGLRHhdEWNA8sJYI70il/lOuMAEcuOimExpm7ZdKNKD1/8t2Tnu3iQTUi3Wd3Xh
u6q7mT6C2KXn93v8ZOTRxuUE2weiPuWJqfcTubUBZb1w/0S9sOdpkgubGztyxG2LX8C3EitfA+sz
DiobjltNytLJPhnFlDEZt8xAJ/vUpXbHGKFWxOB+cKIaUQXFsl33qh9BgIHg1CpFdAEPp/2m/7gj
DQ9tQtRF1lhmkWe1pw/bkH44XRMMRwIuzeRkFYWB0LG62jIiP98NED/G4uFEt4kBzPFLoYQ3p6Fc
gmkUskBSb0LTAmN0Xg5Y7q5j2lEHhRLEBpwNewbm3S7ZcWsaBe4QX9VombbIr5bmJLQmEOzWX7DD
vQFa468Gz0hKUT917fUVg0V7poVy6MuYzER2v3K8eo5PRMRtqnwQvW6XxyHPa0d8zEye2tjQHQuU
9ZQU7vH3FXjMDBUvvH7WsB7SJxbFeLXYrwJAOcmNWKUyA926tiNeyrqH42i1mU85CIibvkSnUI4x
GdI151xp3wTdy6N95/sJMXmtx0LqZSyRPMzGo1MLrAj0Hla6L8lPQ5IWbqmcq+7Fn/X33WJ9u1et
mcWCPA/Y8PCz5iyV92mezqwmnDhioxvcTxl7B8OLpLcqgB5lTzu0lsWvn0Q55Wasc/1t4pcT1kgS
PStuPNHg7Val5BR4CRxH0rXKZYCWog2so5wFK1Y9yUEpQt0IRwV85NZAjmSkPCWnLXa4lFC7I4Yp
sqNYr6MX2HqW3VHRswHucCjp/cwblxRCe13K0TmwLPfIzuRvRW2gywVuR9w+U8fMieHmz5NM2hrZ
WXyrbXj0xZQBbHTPBWN3ozwdPWhHt5i7x0rG+zqF1nD5OMNAOrMQe7PtAUJjAGUKFqQ3ANs3xsn1
diCIwk4/ntcd/WrpPFZ1dqdfqAiyx81Bk6hqP790+O2N3E9arWsUzsOcJDlWQnyrwcgr0W0QFqwe
/yQVZV8Llzc95mbYYYEFnJSkRfAsXUrLuvnMl6jxhcB3ECzNgFgYdCnxalK9B1GN45WZAwsLB7ke
MMluSQySYrvkfAm63/NBa6h7Rs0mJwihEm9c2H1uH93QWmZvtWLp/hhsjZtTr6WOIr87RL2StgZl
E+lXs1xFvJde1DiWm7dWTUgKxL9D2vP0DYggZ9SuxVj5oD2JqbBKVt5Ug0P7M9nPIzR7lTHvzX+9
dh1FetRVmHf16a/kLW4oOTjpcCV8EZWsjB7027st9rn0ycb8zlOigIuRquiM3WnRGFIIaY5aRBVi
upjAjuudEWeSqwfQXo4DqnlTpd6p0UCZRpB2BFB5vmynZA5QtwxRDNkxRTt0nf4G/cugD9/MKO/7
2ibVPOhNuqQkXUSEaidM+xIOyOEO8m6NIqMSg1Pj2wg27zeA1GM3Lgu+pThgAV19slUt3ntPIR4p
w1OYRHXTkcDJ6BQdLF6InwHFL6BUUtJvXLjzJBrZhIIA1w4llkNiX1MHUeQ3rNwyeOIVGeiQVeAZ
W87DFdxyZu2CSk2gtPGe6IGDl8HJPLcDduH0Li6pfRgsTsfmHN2IolMJHCRLhVhP4+rR0nHtASrT
/KVRDdWQc8L0yUYhLGOF9V48zShalcdy8Qdv0utra9k42AwZx7xhKtGVlrgElZwXAWZNeZApHeT/
lyHAw2jTkfpFqAadNgXXdZkfnkx/UsoY53BzC4YzlUbVerx4tsQ+Ywu3kX7tpMGVDvUrClURyxvN
LRd5YX9ePjq9us+TiT9zDl+MNrTiVaxVlwjzCQ4DezxgIh/lk0vsHHGggqteEKNGEJYPQa+EoC1X
dXr20nWZ15ZnHyo2uDS3tbl7s6pOM826pLI+2185eQIVbTJdU3Myg0IUv0nCS4ycJ7WxDtg1gzjL
B5wfCBlacQrkSDnmM4KQjOhs26oohu2bXDzWx8hP8JpKV9qSnXD0LpmQEMV+JpaIpRoAd34iH590
iqPTVt90q9v42kumkMYXVO1fHibe55JCG8GhzQxvCMlCKIQtzUKhMdG/ih+Wjf7bYptJJqxqur/P
vFw7TSVoMF8DUKaB+uc8ISTPxdH9yVIjiOy7byBAWB+Ys2T6EZ+QwzUWBCyCyPKY9emzvhET5mXO
e5IVPC5bXBwQHkuzdafONoJa6ktgBMr4LWf2jx+4XwXmk4Yh42nqtHxy6E+do4cLhGEzvxoRN6hC
dgfmuLdp+jtjbjhGSYPa60aH1ImmUq9s+3EpBlh4wEFR0ZnX9xg1ZXLr2Dd9LLu7PCGWK/1qc8vF
JtUsRdbYWoLa9t15ps83Psu2aL1fxZfPdQoHgAQKg4akyhO1jcWd8+lsmzy9H0BR9osDgWKPJb5f
DKAhDvuYdNJ73ORqkxTArS2RWul6Lh4aaVs9mK3DSJZijeEhIqaPH2pMRuIiNZDQhTcxm3ynVTht
RQ6aiPrU11mPsrWUkSjy0Jc55g4sa95u3TV5zePX7KDrJCor7NLpYrMejoOe3gTXeer+Qjg4icgZ
ti8pzQyegh6WTDpBnHgvUzLOEPZfYuc96HjJXSaR8goQFKjglbwYeoCiOQfbA5aqWq7Tr8O0KOFG
VdH0ij4eFkfUy30zKCJLS58mIoAsLLffxEZ4SR7y9yBVQFMe/LF38rVO0MHvGta/Hwks/VEQwKNo
eTa8xnlsOQ+WLURAKiP13xqvEFdjs2N3XXAhVsROM4ZLnvWBbXHrImW89WfXmwyuG7/yZydsaYWH
THOc3b7EOJdqb1UZ5mdSCN5drtgMosM6PMNjsk2J1K1hwRu8col4Hovbtxu2U2ztEUNhaVHF0tEs
1YF9yxzKW9evChtA0wdf5nC2iWFSg+IjgTOfZgJ2a9UJ8TGWbLN3ac8sAC9IZj1tOojX2q9dveG5
MwGJnWV3EFk+xu0rSPC6tiMzyZuStv6XYm0asI1QS0Q8eCX3KjyGF4Al95s4ISi5F1L9WOweM0WF
ilQKPIq1ZZvohkA+Qzl1panr4h1TZKUYOj+HiUwg4yYGv+TxfsaQyLw5h8lcl5G7sfg3zUoC+nrK
V+ZEWiKxshRWPv8A+JnxDgITH8pnCdZQgigngZEW6dpBNi+Fkkd0KC5lrOHby0BQ6N6wsiI0WHUJ
JRJwWtsgk3e61Gziicp5pxfava50K70CUoXmKJjXwy3pmlCC/PbLqqQmFmxN+yXm8FJoqEbsRrwm
T0tuKS7Z2N54ten92CO9O5kfvBIgn0Z0aVlXBdFfoXqhxCa+FnJ24uIeWyksZYAR/zdehm5c57TA
ZntjiNSczXhqI4yd5RBlt+BG36BNNxudJ8zhU05Dpnnd7wh+CNNxY777Xzp9ELHZLD7Hw4TUwFVX
4puZxCTLROQbHZDcq5Bjp5r1VrsQCBj6aRoTClwGR/X20nDrYJrmVThdapyhTLq8eDPcKfnsS/n6
q+v1YGA2/x7OGeFKb2BoLC/DWXvISxRAjiCa65Bln6SxQNCrWlza7lo17K+FNne6PTtIsCWy6l9O
uX4/dalSEI/ayFxQlncEhDwkRM3ndKcfskrH+tJNV8l5RNyIbBqXPLyuB8B5Jm99ds8J60k152hU
Xt94DTAS9s17ibE/41umbTMU/cMt+q+VXi695LoAvXhFH6p8QucPBaWx5I0FopDRTUjycrjvcXGT
b0ODCCIV9m34+0BQRaW3C5Ha9DELFNzZ/D+QkhMDCuw0OQxtWavbuPsYJVspeKyvpbujN0/BfYi4
CxPGAY0HjjRhIzB3DTjzwa4i33mzKZcZJWjb4hupyK2xbImpxHy80GeG6ZOv2aWLp8v3iGYFMYZt
lBdt6/TTQ/orRH+o3wnpOnx1OPQOzbDJMeDZFfLrCFVjhPQCmJVtdUSa89GbENmwjJ8a3V0VPcD5
Rszc+GjAmIBTUmL+0JzkKVOoVFzpkdQiYXGk/0LuwcZc2btR1VHxVFE7U2kvLaxYN/fiGAgpMx1q
GFKXgnZn6ppvwR+nIb8EJM0Dy9+QCPDUdViWqOSJke2Rwt84QGBGWzds1tQ8k0Z7/icey34obgre
xkw9QnnZBQBHXy7w0Bz2mesZ/dduyBliGsK2zgwMUC4fgSLPsRtHDAtRgBTqpQEIDJzncxvDxoNA
KQrrOGA6jw03/aLgErWCw7zYmdN6flyTIsHAJ/vcviYRsXnHFKfpBIgEO08ICoIpVW0ESvYxXKzE
T37Sy92B77M5s5d7UA6YYvwvQTZn1cyC7LCpuV9K6BNtAE1k8CYeZ1h5qn3gnfqtVJAinh/I4QDI
I2K+AUn9wFmsP2C6OQRDlZKxsV1d2caBjQpdccTbuAfTbuWA9hu/wKIH7+zDM0hK19IhYqgjM0M2
6gD96B+dpYxBr4BnyV3rRlIJnwWWgZcuDAItUwKaAkeg60LNcS2ofsGNVSX5cYL1bs60/qZQio8H
x83Zv9nxtRLq63IdIIFKpw9Kvgr8Uq7tmAFxBuDpAZRa1ZyX+6xA8fN9e82ejaVdcL/rV5tnAIyY
0UHJJsIcf7ulf114s1ZHAxT7nOSXs4GxWb+VNa2xlLkfXlW5IA+kGHJerkbSQ3+jHE8nJ3CjUzyX
JlSzcA4MvA5Xj/hVUe9dNIKWj45atCGZ4aFjZQXsmtd5EbHUgXVYzhNlCw+NeXc+CJ3JjhXkYX7w
IQG7jD9oQOtgi2zEo1Ssb39k3GnZYkjcZFr8qY3UbwsyQIvRajtKeeqZlzH7kjINFji7uJWiYEYr
AhchKx+mQcazUDDsFzVVoieCCHv9lqukPlGB8KarZA4GwlP6NUUw8pWA+zzu7FwAbxMldmuiggPO
wr8l3LBPCFqlL+D7xErBbH+EAg06rAs00NsHmife2HnJtnp//+T7GTv0qH2o/4q6Xf5GOQJsdHHU
fJxts5lfaJ4ZMllRCBGN7gC0eBYNjpAgny9zrIlmW5CLawxkAilLgkxF4QAWLLo3L2DaAtbuzsf5
rGtyVtbJ8MKrG9uTYq8HYQdNKgCv7JrubmVd6KeUl3YJYf6zU3/wxo0ribA+sS1b1zdtb/6eskEk
+xKiKAH+qt03H+Zx+rzi9XegCTosRMJpGY14Xtm7HHxdgPZL91w8PTggQJ68TctlK1ie+gqBL1LL
oGIErMIOXPqKufrM36QrOJXLeqOYbKe2CzS4eekDecSDEjRRsyowY54Se2WRicYAWzimh48qo6EZ
iDeSP068swHpG+uLSw7Juvl4XXfBewUOhBSH6TnrH4ilsumYJm0iMKAsM7y0he8REgtTo4FOYFIN
g1BfRjoGnE7sTlSdvRZVndUrXoBMWHTlXbSsSdmojfmVg8xogwbT81s8gOob69uryHSlY6CyBayE
t4QV0FOFmhH6oNcQdlt2Gpihcxp1iGX+y07xwr3xNDg+i8/3Xq+9grcO/cwo0QWoZa5E6Hv81bqp
vE//DCmYLBZiSKs0wO1FOrbTpX21k6ZlHjdW0T4i/iSivyndGHHXbqFYIKEkRJAEDKqVBGrtXXcp
706/mVfZan9WFu3twn6Gw5Sp/uBkDXYj0z7blnRN9lfL5KN4Qz1RXqp00r37LBogVNMuPgONxXC8
xyzFyJ0G3hp0aToR4QRG4wSh+gswIYRpdCweohfTctMOe3OsKqjvpXMe8GG/eNcUr9RF+dAPAbY/
Rx5Mg63/oWaOquI6qg9HLyTZ+AA66yeGFjkjPR8XAJhYwxxfCLtk7RdEtq/w3BAvyNKhKC+nhAty
rqlJiYv+goh3ZVRXKMUpK35ykUju+kNlWbIzd3NaK3H2UV45/C8fqyUOWpcj9zexQpewrPH+MUJS
EsvUHEalJvJ71wAPzxCKdatWNxUDe/T2rLPCi6KrRJbEA8/txmNGmNeIbn72HuSz1wvRUDSCDYZf
jGchEGTyqoLIyjQiUBYuL5i8tuBeIaptYI9fgnqLOHWwAGbO/3xUtzUiCr/YvnZMnMmwYPL4yjRo
ZR791aDXZJUQpyOo+GSRy9GiJTl+ISgpkoHf2r8qlmlst8/DacSStdczQGcBZG/hbkoefKB3QW/x
Un2iQtwjaMcQXhD4HO9AWwkmWv+X9HpTdCSGgmA6tm1LDCpHaY4d68YlH7lEwppEQL/6Udqyl3g6
52uZ33xU/AcJA7FlEFqxIvyQeqb1VgE/aJZ2LoLcM8OybCm+SJq0Wl7StiDdOvIUdwqmLHvg9rBj
3lAWPDfO3Gl7i3vArrvEPoFzBUGW/YSC9uBpjEyhdXaxtf0E9W6sLK0FtGklTD+JGyyAsuu3zqgj
+yVq81/UNQsJRxlvWwPDkwafWEou9707HLGGaBUONZm9mGzXcsnJyPuJcQQCMmOO425USfh/Bt6r
o8nJbeuwcs2KVQHbYOSNYxwShvw+pvs7cfCdDOHwVBTOhJQFEuyUPSlqX3uBdv8XqjmFSPN3e8VU
YyMxJwzAgbqGwF2O09U/4AxqzV5UBYMCdRqUxfpGT14e24oAfYkoMxb8qBCRg9OkLRftjwVgYH0w
B2FP3TgKBWS+7ZsdKrgczINyyHwo21ssk3287W8+hId6T0rxWKeMq5MziKOTQDUThs/M2hot7je8
UCoFSmK2oLVGwcoI6QUVGuCAgLIOpBw/HYHbO0CEWgpNABec0wL4YnG6iiLFFKcTQ/wkmCMIBe2U
sG0ugKxxSrqGgLZhljxF0XKgkgu6gbKvTM2KJqnTkl76jD7MIGK2iuIU+3hFBQCmTVhT61VdTzy7
+Yo4F+mNuwwxBTjD2pC5ce3/wuZzM1hg2HRX3NfsaPFAHL9kDc6f+K+sWm0RbaN4ZHKKraQRPWMQ
LZ2r0ExOaJHRREpXFL7x/Ozs4bLf3D9tBOt6JKWvSFXROtwGafT2eUAcR3TaQ5b3xqR9l9C89j3D
WIWHgIRdpy/bQtBknw8D+691XJjN3lB/kLKACXRs0wrpUlD4pHo+wuSVM8N/Ag+qPNmmgZk7+Kdm
kgX+a5T8Z2g8nFaqsxx4aM6rqMr4h1e7Lu1gQxRJwOni2JthOWoV0FjlJQ2M2KryvkgblD1qKNQc
kWAbMd+9wR6sa5B+8lWJ3xGogRBjdwoAISdb7+ggGnL898A8ODq7ihzSXeJNEVcBwpR7JseMiAWC
I/D6qJPhChdN7tXifZ5tYgAo3UwH+icNAqzcnYyFCpTqh/n44NjnrwqsMz1OKiKBwpToduG8UKTx
4aI3vY5kU++GhkN0eR27pb2f78+Bg5f/RNIYNYsBE6Hdif8J0qR80QZaejEI9Shf4yZHwPU/8Flq
IZyuvkEmaHa7XEVJgZLqxWPe9EYU0fXb/Hm/ai7eRHoJ4h8Y7Kh1gG6w+6j2vBUMIvrxU+h90ciD
CDR0kSsRkIOfQoNb7mDzb+0U3LGM4y+6yXubbK+KewxbnNRlBo9ypYO/XltyDJH8KcBIW7KM7No6
h5e4riQBwDyIngpTt8oYWCFnppaks2RTH+mjB2sT5h/+LIYs+mi62jGEjV43Myw5bohxnJniV+/V
BmpnQzBnSOcsmKTQI3on0bK72ds4ip2sjbhJCp+LF3MhQeLnQbzkSnoCZHCLDbYv02fQdLrgcWPw
lC4BsxprGU8xVf6vUX6NZx8MELeJnx0iNJiMWWYanJo83T+baMhmjFM639l0YsA/hMm5cPLjF531
9fl1jHlMcZZHfS1nSrBQQMSs3/JknINvHFBxS7IVveiBcjbVs2XnB47gsjNpwYjgLOK85x9fOzLf
j8ASujUbE0HSH3rHFEe2AYm6tUdLrDevN5PpRJbm/uswjWSVpjQtKjx3VjJmouqOUWr+XYQ8Tprw
Rc3fga6NgiddQmrfga7i9S6SGM9/24M3w5Q/8C084YMImPltYyoj3BmlDVqddhufe9MekeFe/S1V
5VlI9o2xzIyQhl6jqcTcRwq4sF8i+80FwTDdTcBFdpdR2RdAHB74t4obmBlp29hYEluNpUw4Icxn
JzWh6BJI5O4YGTnITIU01a0PJ7Avr6G9vfomtPyDKiF9TBEsd1RFhoBgh4uQg8RILXn0Aki/HWbC
RsV4JbYK7TACZxJYlAfBl+t3SsgJ5VMdZC90NYUXmk2/JjnV4zRSVE74/3RljW8Ih9nmn3Xorl/i
C2wY54NErRO5ff9UYezDkO4D2EoD0Uw3MgpH2s65f4h/UUf6NPbo3LsuPDinxgwIQNKm0lV7f3bl
KTvCPuOiyayo48tvUzSlmwsUnkYBtfiPJlFJ6P6+Ui5e+9GBIzZQPVv6p4qN5KWX7NXZ/Zgg9PxS
CtaMKkf1ld/ttA0cBHleEVadLlPWgYxp1xlHBDpk/MSU2bsxoAT9nUH7OQmBsuw0rHqlj9H+BSBf
6cPJLs6Ii1sRnO49yCqgm7217f8KDFVJXi2qR1fZTjgNl51+ZeaQq4mzb0p1hcJ25O2qNXs2jBSm
12BwU0TSRldFcgA8nrMWNIna0XHNBRcnQ/m8Xru/09hhbfpdRfGQpfVJCofZxp/qgNALtrDwp1ih
PEop5k2ciP2UlQraKadK1RaBXU72igIaZrs9TE1tt35pf8VR51mCBB92jAL8xDLQYj6ArlCvHYgr
Ch+2dx984XGn5it/ZKPCoKEDGwbuX0XF2mM2B7lR0uXnYYXD2ZvRExOu0nsQ3ENW523wYh5DpIva
nGw4XbX6KYgWl6Q3F+b7y1A432/5QPRKgR0cjPo2OXvCgOPIzyyVckUI7zG65zGgT5VbIhWxfJAl
Qe8qWGs041r5i66FZsG/eCUVkLQIXYwr5btJmwWNGRFu3OaYUE5+FSjlCKUIrQMWEXSrX2MZOl19
F7AGI8jym0caw1ss4pReUmIF9Wdf07WFCkG3av8TgKhraCBRD3jEtfLNkffd2xJmUdh6IFOQzx2+
6Uw9yq5fMFh2nVMKBxdCeNZWzAPuM1GUtx1o3RlquWB9W0QVzerJ283KEOYtJEO7keh7HselwlZu
PE1URtbt3VV1quAsuxpxMkShK3YW6w8Nhde48loMqCaTRVbV4OFnqnYy2NxSsLtrKCiXphsRPLx3
BAqrcZwNZFqfCrEgRKYBRQonO9j3dJleLuLZNhlhWgTk9FsVsxWneNRSNo8yZ0Q5fv9VIvgxACzY
BubU4GoBJm/E2Qts8jR4mGog5ynB8897z1gBambZVBkep2auSqecp3+ug4gvpr7SNB4NGANqeOT7
t1QCpRoJ5eg6YIaOdq0G388wEosloB6cAVudzFHLwuUwbRHRAswFGh9drWgorDB47TtoPqkWQNK9
/v5M3urir8JZjTq19xtGH3OM0DNhP1EBhgXwM+S9WxD91GJabiVXA2swAqoKp0kS6bujH9gtUHYy
TJR34GgAruaQMnq0+eCiAnuawtLnHoBkV1kO99LpkPH7sEF4MI1phYEDZ+0oq5SbAtaLJjd58v40
TOn/ltvkJW2WR7+HabPubZiAa/SU2v8mxM8nTqAaXFsoZqCjwzIuUJJUJ6N/yAtPS8bVbf0HJyAD
aZi79A7SdFEQbx1uCTfJ1ex83h2QgKGeoIDKKA8Jr9NYwiyJhzQwMzBvHqKNwsRethDKIsdVP7mU
b+dJ4IrD4+85kwaH4GKS7gjaF5UBKyxITnGdQDhfxrfzuLalktXbaBC3WcLY3aEH8Qogy49XRjCA
7nmIVnZ2+p5U6GC07x547M5Mri+fsDb7cvU6dM+gzRMxLUfKjMlUxcfN3Q/IpSDpBlEI65ZyUzkr
fJBIZadbn93xtrM2Bv5zIHeiaM6Y2oiDH6kAkkYsG0/6n9ECk5euxSLS1HH6/frLPNf5ssPHLXQk
eL5XaZpznLEA2HTdqZjTV2lbm/x7+KYueMLiWZY2540/+hXjEqq2/o3+HsXor7hQwf0Sq78mNSBX
3x8HO17Hn5iHLv5POWJ1CZhTwkXPpZJ9CY9UL4Es5AAOwp9RezoL4VxDUIQgypVWFnX7WOam6xHI
aUeiQz2W4+cAWV55tvQnWnvzDTLaKrUXkN1SzJwtD3fg338EIe2ct/3Shj63zpK4EzJzzC2/Pzyw
tTQTe/j03sGt27cSLFCCGUq0fvIeWot5Ze16mDG9CFsyLNNFiqwzfzHcs7Jv84hOmhbv3WrcQlo7
vfOrTdTrvw0sqA9IhrBeSUu2R7F9b5WmFHnaHhpWzsBpx5qSsu1ldn2OFCgT19zanNUUCVR/A2iz
zuuU5f/N9xAsPVxS8IkNntYwlTyLZSYTvhymt71elZT/JxC2mi3+Wn8B/oqezdWm6KjXi07QzI6x
o/dhreWXuhxecLno6oM+UVH8mbdMQTeh1nevQTI6dvGdK+ykJnHkuvwLIs3JrMdYg8hPgEsY6lmd
FOBtYwkZc74J2FmQWVS536Ax3Uh6sSADUTYVKKA+gYQ9o9wCoapvROhiKQeabuBxkhykxUsCKW0Y
i2g0EbsZe9Q/rE5ryLlvCJcy7DvGXS7FElDMXQUYlnNDgkGzk5h+rtn+8Yu8/cE04qYM82RtUI2p
RGghij61xIjVf8JvzZ9T/i4sVgvKXGH30vTKsfJcrKepE0PzjBTyJNmVFcgShcw1v7OiZMGwfYyK
LfiIZXkAhTB4Ci7j7nBl4YbHZWxVayIrrsx7LBwmTT6Q6DqWUu9PjJ/zVt6WQwG/AI17lB+ntrfZ
vNOKoZAY4wviPpwgpXISbyK71oOvQpF9skziNgyvYdEtYYh1naNtXZ8Lbz96o3XxRoneBnnXo0Qb
5WZ30HIXrQfS0OAwZ7fg33n1GV5yd0Nm43ZVkNnrwh/DqAwBjbkxkY2OEcSlSIgxXHcYSl5B5YXD
K+0VvXC/BhCUzFew6uS9tVd1QMGvTx4cI7HKtcNaeHNOFCgirTlKAvR34rHpo1SlHDDU+GRMTkpG
dPFAqUZshJ+F4eYO2Crd/rZWEwd7y52EOqp7focjKxkTd5Xh+zB49jMjjyKiwBIBNOtBuQ/h5JAw
TuD2ppWVuymUCZ2bDC97gwVk2uQD+qH6Rbub8lU8fcEZ8DqQs7LqCBnnyskt3ihbPQiiLeEneNki
h1RB2GXFR+sdCLM/JiMRlKjlvMFJdkt0J5fLy44CUGFpiSwZqLfhCDbH8SXyzcF/Je2mwKQSvRXg
LNGQzMa53HCe/HpsnmRQfYyAHr2G94mS0CbEG2osmo2HoQRFLOctAZ5UsmwVCpwiqefSAj5JGsTK
NV2kyOzZUsQ5ir24N2sVM/umh0eYMgWmXOIo6GEQJUcGwpUzA2SA8zWDbMzXIoiexC2M5BbYZ2lH
bHbTKQn7Dhufv335hvcBz/rpSwSioYV9k1naFKEP3UTuTCWMrwgUDPOVut68KADFUxp2qLCw0Upu
46+Peb9suGcF+8UL7BoLRSnjVlT6WtPtn/MUnOYAJWwbM3daBRAq9kqYbGX+zy8QVNs/EpFkYX7p
LShntZun3H862VPy1LV0IRJBuhPmto8/BC6WHaSiiv0Jb+eBOsRk4shtXM+OZnbhL41WevTj9vo2
ScqHO+EKibG60un6D59UpONRB3cd7TwhCeWhS5mZCbsQ2/JtfyIy6508kat85z4hfqsjlrAt5rGr
sQH/klFS+r4/uw1s8Ce2uNksBMaSxvZfRmGDdbTUy9e7FwyC2TgYD0Byl7dhKMSlIMHn4vTU3cML
j+J8qwmNwd3gPiM8SAz3RLZpVpr4fbrvzNPCwB6+vbsuJNPmudxhJwkIQc5OAGeH0EJwSLr4Ffc4
YDCCIiLCFniVRl1ibv5Vqn+Q1ZTkfUA9A0Fys94xImHcYPzey65pEytgfV3E5LCi8JC6Li+htVpZ
GqRaLWJ4NkSrBSEeiNB76WN2SVShKG3qd4xhJT5MruiCm4mUkA7Xmg88KiLQ1zEVQtWIb1bgD9Ay
aKTd9GsepV0jRSgtHC5NR381UejR3q9OJhoKeIvcmxDR1BEtvklP7dhoJ2miti0SjaH77roOl0+3
YyC3MfvN4pGxbB/BYHns4op/1SARr4G8U2tciqOGcVyRd0Yi2BR2UahAHd/r3HtBwbMU7S3xFdO4
SfaxN4UFLw3RenmfA4KFiku+UoUaamtaFEC6pX4x8p6hwXT2MoD77xZpiWIYDPOeYEFZO4rJvsJR
z9S9EMOhwyU1HHr4JsdX7WIz9ZE7xIJOYZIn01WAf4FF6F1A9xLYiSrWFHwXhHxBUD3Vymzz2G0o
8ccb4tctEUCXJJ49ZNFJXoUbK0IrqQGQ772unR29drxcIRVcpM2YcBasyOubMs0mrtVGxR5oQGXo
vRTVERSbgd+XXAQr8HCKm5u339wOrYUzxoT/EN+W4Exph8Li8sGSrtsFWkRo3jsVSuKW/7mc6uKj
qSx/UuQXSdnaLfujfpghsAC49+/HUSkgVkR3/yVSbi6xoHOciIkS5y0y2JFXKjSEYhWJrJxs2l4G
eX5njE+H4Gk+g+oB9LQoZkhb9K9K0MARRaZ4k90iSspSVBWqk+aXUkFjsLGDSXD1bZja/15lqS+x
jCg2MZZ9ya6JwchyvaCCnfLBfr5Nyk+C6wdKbIbk3a1RIb33BMddUwig5N4jNfkPqhoWSf+tBrgg
W/JoENqdAHlYxJtiR5uctoz6s+5UalK2C2HBN6X/bJj3mILeTrnDV3yYY5Z0uWDhWFogJOzx+Gzw
ggpRyyZmxFvwdELtVzRym9ns6jXOWcY53laV7z4d7bIPu9TQT1vPhqCiQT6KNVKb9psc8U/CFbO4
4MdzpbGz6vI11xdIVqxx/vW6OOk4k8V3FVIchXJT2KOpRNsP9PPwjKTHb3HtTH6r8gjXDSUSGwsw
emSvlWgd6kDqsZ6mqVBUG2tRQjctGgyn1nbZe0Eh4ur3QsDpvwYtjUbfwTuSThR4d2svfpEq9Q1K
5D9FURSzpat/ihp/9ah+k3JYQQc56tPVkpkOwplq/i6Oy5eYr9ZWTj2WcthbQeceBoH00+8MmODB
MweVhUj7Ux8er13Nj84vsqTgZj9hIh+8dXEHjhQXMorYLbS/1oTlGOkHgHHisuumuQOdBYjHtBkm
/sRb9+jLkvSGM/8E8mgZK88GyLNrXVcvqwVVBdrvyYOUGH6j41TNfLsFMFjo3BJf1yYKgKYyQHx5
yptSRQ7q2K7u8NJc2TE780KN+mC6YVbvyOMVa8UjupYD9s85mRuJjzSZ+BQBgIyyo6rg4KG9i1RA
ogcU3cUIJXwmIxYEfQbDceK9iH314EF17B3TmBrmhx6aTr5YZ0mVJbk4h5XXNTOEKJhkYZq8bZXR
7eGrMZFWCHenULUlEg442f2jb8rsVancc8W3WNbYfWVhgjfTBC0Wy2Zs59gExmu4YB+ItB41XVUU
1Ww8A26ZNHULqVMaUay/UFHQCBTIl/hft5r19i7YPGkbRXAWHsXH9CCxPcMZHovHUflmt5hBcqPG
ak9RV/zg2HNNZbVLZmY/8Qg1q0I8Z3xgF0jwj0zQzCQQK2OLS2Kp8/8fstVfN1fMoZtjkqFcqp1w
R4suNIk66iNGJooVlYmJW27D8fNc4CsqfPnQDVEA8NbM0rJS/fiWA/G7/Inbe6hL/gCj8Er7QeRc
OauyVfnTIhmCEPg9WLT4KTaPk0CBMPsnIa9fRjjxRsRCr+0vLEljCRa2Rj+3LdVsV5LFChDbocTF
b5AhlfdSQxElFDkZ5lnND/UKPHjyrrA3cDPC1B6XQm9dggyNiPa8TS0VTfX11ylcYEi+uKkpr+vx
ukpJ/LRleb51ud5g9n0c6DgXKXjyoSb7fzvbYll6DcdK3dVpueyyx/qVCJeSM+vtRpkzY5ASKCCZ
+AN8RWq7qIo6GvNtnb9Kimq/5XkcOKo6DbfnC6N/TXUG/idcfaD0k0qZ2wx1ypflvT9UdZY942uL
fK5yUmVAZU3sypmeQqUh7Br+Gbbs2++9hYVKkhYvF97/MYuI9nEibjk/BcvGo6FufdcDhrtnSxPZ
Sj+BdpWx4hrT+7adZbAr4+7gJBX7wN4n15t7T6R6Kz8iMklHFgWiXDMegz1FgFaaFkOHwnaNRyPt
5Do7Y2pf2xYq9N6+7r5ggPROmz9S/4lnqNspchRNKqt04T0dy5XP8ys8aWxfzrtFp7+7Gwv/GUGE
rXW0ZpJtAfj7cV/DguylhkNhNeSet9lGNrIsHbBO/Ifjjnu9+3BDGaBxScAeOdE9hj0cGyLKXmFx
ePYVCo+zM50fnSJOx5JpT1l/4c5gG/J5WupPT7pUXXCanCRF4cviMmLmzXg22YwkEVVjvk8QDOH0
nB1mlpFQ7iSiRsd1Zj3O34n4VRUKjpQQBbNnKKJerdt+rW9Au6jSVD3jCImLBr8cso4s4ICbPMDu
4LgenU2WlPGN+jFsC2j1/1HYENngBgKk4iZ4PkVI5/hPFxWmDXtIR2SBT1epIA+PosfYFMHowEUp
ovu73qnMgw4FK3AsXgRmshusR+MR/mEqDAu9wqabZPgVyeF5iMVuyD17YrUFwWCswu5Fyg1TOMHs
xBNQ2hADe5aBbsGyyDo7yfEXLMYLGXIXhugMy/aVXnNIBmE7k859ZCfDtadW+yycSmiDpTje9zJl
3XaCIsYk1XrOqcQcX/GFsTgdA+npT6zcP+HYqlU1mw645yJCPpmE3CTBRcEI823ck2hoEXIDYLG2
6nuACdCHw/88mX+gDuUVDud42gIhYMop8wBnT4KdIiv3NcsNcrR0b2GFgGbOo555PYEGpU0gKz18
HzT+JaLGMF7naviOF02Ffe9BxBwjBveZZSYdWwdIJ/P0LJZ9cf89ku6P+2ezN5s2qD2POEaNaE4r
AdntXxLX0Y/XWxEhaqDI058gaYfXbfeSGlX7Y2oKHWQgEpW6eezoH4r4sO6Lu2lWyLAdu/IobY1E
ewrA4eLQhPLyrrp3K/ngg74CNqT+M+HogodVkV5CvGbvljaoTDFaPpatGcdRIoTnYG3Xb9fDhj1c
NNf/Ei2HeriYyzX2pCen26ESiJFpLB7OdQXFaJF4Q71om8LqjoYZFxWNEm6xA0rCpTUn8tBCq6q0
+7K20TFHIzRPnNXFA5g3uYSY5MfIr2bEoMxVnXCPzLwranlu9abh3wEKsy5M9Exz3D/o+Qp8hcuV
Dvw9g5sEaeM7urKA54q3sNWPKIpvFLULzT6DEvyfmfW43b59yaDNt+zT/1hVtRTnfaH0CXVw884y
JqEl9wTiw5VH9zt7B7UIVIhfKDSWzlsKfassmzT9iMF4ipqXZBSjaJTtv0NOe1IbrCRhcvounAHM
7xQgidauJ69aizijNrTY1dbXCKA/HdCOhxJZzvrBFvehBCL0vd1JgT6EtApnTSweWj+Gh0bbFk3u
Vj6OaJqvKqfGAF1Ue9gCjPOI7eGU6W/kxrZavM3YhQ5pBNIZitfu+YPNQlI6fzA1V/fKCneTGrRy
qj4kXG9rbUgvEfYTJdau1YB1ncOosHH2gJXl+fEst1Odbwqx80NE+Q4sUdrxza12QryjXTJ5568j
NevGuIOfXnTfF/QLneaJmnoFgLQByMda6dmdvQSqPKv/ZEofK2LszPobXs4phYGtAThRcUFZYA2l
cyQ3E8MqjR5ZP4GPkMsGhG7/+RmJ6Qcp9FRqgQ9gG+P7UpMZoRiLRLcA1cDJBhjb9DaB8/ImGglP
+4paxFl4VUPNSequrlnqYGfd+T4c/jZQApULGJCK2LHINvB0byTcYY+hAp5IIMjC125b22e5DXcL
lB8ECJHC43Rk/prmIfPOETYvtENiH0VBlX1B3N1tSiysb4jR+m8sx6Gm8/+MkkZsA+9VkvVr9H/j
wSGMWljjARtQCMCIO6tNQxbwmQ7lVgGRyDks7Oa0Pn5z4aIy36A5VstYIg71/88ZkioVWjXAzE6z
bw7OyU486/ZMbyCPYAfWJaa+aoyic9HLj2etm491Uq2w8MD3Dox8mODnIjttHPEsHKoiYscePEPi
K46dp0QWQv+wpvkQzibQjvjK36fg/Ke+K1fq9OxmxRkNVbFSVzS0PWK9qH46C/62Odo5naskuK1R
J1OKUO9rFmDsIMPFbhDk2bKnosJjjXnFOP/pai5e1lilHP2vhA+CAsWPpVqVUSETIRsqIteNa2GO
oEooSapkY4MXanOiQ8GZtiuuOWvGQoPuMA6zPtPwY2xh1EofjInv1CRALeLZEqlH/b3lNuiSXCWW
J+67ooMvsV/rUIzsj/onpLjMy59OOvDm3c9/4VhCmZ7f5wE1Ev9XA13mnszdjN70sR6xfDzeJ0BI
ktzb9ll8HpGZhr072itLDolBGszZyJAR9P+8I/nE48mbypKnkVNoS3CHTPQ+S4r7FmsvVUFMzu1x
e/iYvDcnhXp0qY2jIUQ3mTfHMpYkfxClg9KskE60LsCTqk3KTLv5BoeNKtam9rnD+pH76e1EFQHJ
d48j4PwZkH03DYmmrqW+Lpuy541gzvgZ+W/ereIN99GR4DDUP9EY0iV0NbIusTx0aFlOIM5VFuM+
R25SL4oWpiqjWYtqibVDUWcAIxVRlvEE0aObW2czyDEPWHkyvlc6XdcDQcAjinA6TR/QEApx2Ivc
mJ+OG7JsBKMqcGAaxCXFHK7/CqpWr9EWBui1K2aEu3wUGI24+k9JVmkeKyw1t798qhwWdjxy8k+D
vTrZb3GdU6RbGSDUojOk/KdzgyHyyBsfbZ1vRonuIhI6UUkhaavxtfks12q9gmk6y7SB1zQqFmLD
p/PaxhoI4+BQFWTp32d5ZiVnGMGzXaQI5M9/xjRkBVfWg9lLbcnXZ0s3KLqDYoFmsMWTjecExd9w
eoI0h2a8QakW30fbhVj26utNJwEJMSotfUnpPfYFnEs2gUSclIyKWP4f4tOWyXRAIDaSWn27ocZJ
Hfd73uX8vZK6ZsxG8H5PfF4eVWgqZ8XtC1Gms4ikJNqfYw3YIkOXaU7HbvFqYj9B3XgzsudesTVU
QlAfSRnhUbksyG7j42I6ZaVxq99EnY6heGpTJNHTbB1GqZhDV8tK1CJbFKl91S1yfFg7qDyMa+X7
a3x5vntCENu3zO55A0de6v8cAIo/qvwnuImVSzHgoU3ZapaDA3vzBi8GEq66lwmzJ44awnHZxcuZ
Bj/xnB4R1+dLUtHwM8lQlzxDoaKu42gJXrVtV90oDeQIYsskTaEn9CNjNwxfctfzBj7VcgBKMY7t
d45i/DNsOTgOVaJWLw/lV8H98hYhGWixsJgGDQzlj63Ih5pOh9+QPuADMptmGcpeR6QQjBgLDcCW
B6GMyafgycq1Qz/QAr1FBYj50d+F8nSyf/pwwyBlYHpDVhJy76JpxfeUyycWln4krMnMogyiNwPn
CisNH/fX4/uYQg6tr5R3DtxYK+rs8mymMBaR/Rl9UQjAbeGGdhjFkhqoh8jJ/pGVF5tYwWNEt6+s
UtJkyi9J+YLLbHOogDcdw9UEAGYHiZqurHDELtJ75qDU6cJIy/fQFnqY92llDBPkaOATruEJCFcB
woTiYBDL1NdoYUd8fH0ydyfaX4myb/rTV347ixatH9JEbyKTc4i2QDh+xIm5mW+QQwA4vZo15IkM
xJDePkFfAGthVI6SZbAZTh74yvMO6qteHCsbaRuHklK5zkhNY7uzvY0J3HWtBCGd4lnhUU1yJzZF
61sJ7yFg1hwr4jeimsfigofWb9bfGpvqf1Eg/rodxTl7qIgEN2uDoZxTCIWhkSsykg4pWEfdlOSi
wtrAhClZqSbSbDCa4TjKW9xLJaAV9NAfdsqV863vYnJCIkKXH6z+K+Jlsn/9eTfQ8JnZFYkz7+ez
mJ/QPqLcPVQij3pEYQ9nhPzJ8zlEPDn74fJLo92Qc7BhqRvb/aUZzJqrQpbHb/0EoLhRdijB37tE
WXbRDEKuBBFlvYVhe+nzA60SPkntid9IxhKSFAcSjlAgJB6xQVMvxQkKmR0/KqTaPmS0Hxzmeni1
RkTJruJSfZsMFYOSSOmBQLePBjGWqu1u7u4J4jCqEZsC4r+zy0/3lI2KaYxmBzaLiW25+zjCDgPC
kmEiHJ247hMWtudKzq2ttWUwJ619sxksrn4Sje6PeTQwYMRk+7DjdiYtpEeHeV6izQcnpr9dg/YH
P3S3tv3hAF8ybwh0tKf0K4Vz/42QGkVFZQuK09KzbHtNxopUuUdVfaEfSbfgqmxqiuy6pYNB1lWB
81YptUsNJEJfoSRkFtGH6GJxk/PevjkwISKxgp+LEjQusfnmjBaTKkA+WXbmLJU5ygDfIzgQf2cV
3uIwGTSMMbw8qZS0wdng00rtnzFs8ulrPL5ptujCBezD3XvRV/OCVO6nKXA1KfcoVJO0/IWFqJE6
3kW46waZRhm4fFKFTZbJkNgjZBVcG366znfW56p1lJYz0Z6l+yNt3YLNdxcQtX853sc2zlHxBF32
JvTLdmSYRhuQyL7qykZlezs9Ouj/6OjsusUUruTbO1m4B3UvWOoB69zb67wlGdpjldZPVxODM3ac
oqG4HSwNlKp8rB542euETNBpHzjBHcEdPhis3iEHgHpBgG8JG+GqrDVQWFWTIEQYpvSSU87c1J0c
MraKZEN0fRNh30uJZqLhUmBwYxM1ZRAcRZiwsLjzXe1kJ2PYteFQV7kjkuqc8exSaI/6fl2Abbpi
PRtusUAJ2/dIVedDm2P6bBcMHGeop/Qx6rFkNVOJdzWqAoticjFOojJqiC3GCOJXKdp79R+lw6dI
ekG/ubDuGkyMnsLXFdcyaZcXuYDofTGDsMQNQUr4th62QWhBmSjNj5Q5nINJYzqQGxmpBlY2Upfm
mQWb9HU2KCs5aa6CMfTExBDt7uFFGGJ/Y0FQOHF6jFjuK6R8VAzI1Rs5J7c36PlD42uPhTZiwO9l
3Khn0THBGODEBNFkOsUroZycKV+0P3ZYBJ9Ij+IkAmw6UyLOBHs9T9IPbtgYpIDUPLDJBpwjkSCI
sGxKaSGVZ7q+dod63/t2QBt08to1PX0wmpbbSEDD7ugxVxyc620DTvyEWEEfEhUG+LkHz4v8bBs4
0yMyvJ0pIKTowL1JF1WKJ61iTLDvn6mZG9nH0L4z9DLSZLgs7CbgKS/IiF3+KieHs3XLYwjldCqa
bSQL5hXUE+jilyFcIty0VsdEBjlLN6A0NLCb4RMKFsHWtjsS6LlHQz86KOZchsJk0l51OwYZ8cVQ
dI38IWVxMt4KTCOymQf+SGUaniTAvFAhAMC4yF5AE16oDV29xTdMAg4J0/hrG8v+fBD/pSiSFLSv
sNIfF4HF136kI2vH8y9Y6KRQho0Th9E8xHibxLjLkrzvL/oB59pASfLP+UpWceB+6bmS82dRSzsT
ju8mS1n0onwYAUFZpwVqYfwEoaN8Z6Z6AQOCMYLwURJRBfNzhHCOgK0CuMWrlgnFi/jMC0doXkgQ
ywVFwkROCUjHnfNPS3IRCzYSJtd/F8X/zSKIkRYaJWiw/pZgb4xOsxeVWge99k6nVQjUHVbtEv7h
3aNvsmpaXFWo/z40sU8kG9ZNbdmtgRiXIN8lqLUMXMOJgQnINjHYJyo3s9mtuQg2susZcbCXpQjp
mMeoY1zPNUlpoxo1yAzqiKlujl8hX1zRcM+yjdL9nheiNF2itVyKJQca5SYOR7ytLog8F5XFotzM
rT+HW6THJz7oh7slL9TqILvtj43+yVSI377McIk7dFi0VGZJsulZT9zNZFGx3BD5QlW7SJacY6ug
VP9OPzA2zHLskMmilfDyCelEaGxhFqYhPMC6bYisGQVXPykndcJSixvuIuN/VSvPto/U4Dylmaz0
b5dP4Hgxgh1YcB4PixPlx24LkUbseaStsfkRr5d8B+Ej8BVOWH8Uim5D5nQkwaj063H56KFv8yGP
pg2BZktp6y+GX4BgYrGlprD3QvHnxEr9Mw8uUxjkTR7+G6hWoEIWBurXtlVXIaquJJdNCQR2AIt0
1FZB6JSuc6o2d0FmrIa+WcmiAICFUR1MnBYWRRxnm4HkVAEDlRBB4uoLDgXZQGAyz/D2qXITa7sA
md8iFz5jaLrtxF0IBBx6d6jFErOWTwcbT421FKuFpF84F4UL4+2QTvKozo2ke5TgNt6HP32TY8T2
3X2rdZwitXoyzDSqQwBS3aFq6L0eTVZxxvUDeAm8bvOAv8Pj0iX+KuAVfja/770g4eiU3W3bhvh+
27bDnNFWRe/58lXyOextzfeDknQVTw76Zxwg/48JBm3kWeOBhbguGAPcWCwO0KMrAI8GF6IYR9Y9
avzKUE0Oj0XwbBPKGQBSgIlkHxqkOPi2YRa8mY0YzWJThyzzxb/0BPLGiiNNmu0hSnQc4Uetn5hu
tBGHnXPdZ0YaAK4SfUKEF417GdCZIKEDj9TYIVZdt/GLNFTrFfxM9+cnGDlipix1Wsfu47/00pCx
aE2Q+bE934XNVUnKa4uy2U4jVXzHUOkvawSxyqgPgRMTByu76ABqrgpxcwdAzdqvmIa00Wl1LDBv
YCaTsszfrmxJ8idLPVp3NzJA2zn87EuDPtGS1wNTIkI+u6YuReZr4+iKbdhxEKpHd+Ue996ZGX+V
R/nVAzjdcG/LmpxiqQ9YNU+uQ2YCsKYBmXFdCn4iQdUgHwXk26D9M8mqP89w7BRRWtW+Qn1bQ+Co
iQdmr5k1tVkyPsw1rtqFUOdKdHlSGL/4AreNN8FKS5AMZGTU1sVtjA4pIrkD5nkXbWzH720oJc9B
t5Qsc4eoJPASUgxUz+qkcvQnGEH8WzNxDUIhNCpNogJM6AcO1BIhf552Sn16f6AoFZOZmClsgQOW
/wXQIqEIzj9nq+jxw9wGz24mbidaFTnCLRZLuLG1rAet59m11YyQUUpk2Tfa4sRQm4ISa3qhDDsh
wUzC/dQuyop2rjV4KRYaeeRM1sGSx3nII6QWd+5BUZYNVCDdbvA/eIn9jvn6S/Z+D7FmxuoFTHD7
gOSzxquHm5CXdJIrEuvKYJ2Ra2uLE+h7fXbszweaoZ2sN5kD/sgAfmV96sYfZjKTJdYEGsvz3TQc
xXvwSVm9huCaEAnESVZplk54S8Vle8bN11h4Ptej0WUwE7twh91CmQgTV3hSMyytgSDAEdSFU4DP
IWQ/CYRFbAOmLMdMkDPmBJPPnM9wfxDyeiB+pOib3Ig82vLZw66Wjs8DYluDk+DcstrGelXBsavk
zSSMLLMnVDlOFtawe5vTeiTCu0vEYbyhYndgMIBGgWW74jvhju5ntmIR3vsQPxXVf7mTXWnPhwem
2N9LfE9TZ0qc5ho7TWJcX+b/KxXwf6Hu4Og6Os//T41xmJMOjbyRe73M7FWk0Kq//J+m7xUWTrr9
owvhgxdQwQe1eR8ATY6f9OpBCjtiL4Z2y/pRQU5YezRcGD9oDd2R964JF3XgSXd98h4Y8BRxg0l7
8sF8F0cpeJkFA1FbvAEWQaTBuEjo7896R0kzjLsT5JMkkSHUypgl09rPiV7cERB0pYJg8DE/7gZ3
5HhL9FuIbS4LYnU8SHETyaOh4zyblHkFvNgWCmdfKllXZucj5ksCGaywjSvxqRgiTp9Sa//Tx6/t
Q6jQkuzjPSo3CitHZ8TrGtzKM0BHAjczjzkubUBghOhIrWqEiqE/5XPGL7yEZuk8RyTV+aGQGeFT
bhid4Ga4FzFnNBRet8OQ0wFbh1BKZ3rQJt7XS4uKmt0Y406Mizi0P3uSRUwvb9DIdB5n+A64QYnN
OGZPYKeUoJjOdzYUt3X3bSc0tCYqrgDJkmGNl3k3+pEX9BCp3ki1fF/60cNe3VvAdoD2Rzq/k5ll
anihk+63Eom9TWEt8d7RXOHYaPreSOeXE8SL0wNqiQULSGi9gjxp+Cgfj0TH/s7pZ1fPSAcMwSW+
cgXMCiSeBBSR0lU+V/pTzwXisMLmL7GOPdS6o+CRdkD+CmUhezvKRMBPzz8i74NgFP2YwVm8NADh
Yk8WRUjV5qKKyUw+k223eCnwmDSO0kLfPwiK33RSynxezk8+anLBGVK1Al5aTKymRgziv1UN6LFR
Ygniz2ARjDKLl7xl3W1lBhOb/+JhVdTLWihikX06YQsteuAzBmPZ4bjuykOwS9vA+bySiMTCU+VM
gg2mSo2xDO8okyXYAemPzD0IAdy5fYS/Qac41PpFuWkSY3qLsPhJST8zVy/gIhGJmZEF4NffRBW3
6jfm9+f3hGMIK4iS5gSy99RPfltNaR6GRj8FLgFeCrHKFuX2Uqu2r8dPGou5DCj2Z9r4eZSYS+pv
ihB3jklwvDJiQQm8RKkBPztIcNjDF1ccjvfQA36QwJt+s6X9cLD0f7mEfQIPpcGMwceheeO8spwD
PWiBVeU5jWJyK/1Qyzv6nyq3ZUUZ80rDlx3eu/41ELsllvviJklH3x3XRXSym2v8byaonFcXiGHq
8CpbHnRuSExJAtej+NUnwmIlxrJ/NnGabCXhzlGEcXoWsqlXR0Bhb4GO3D8tL2hlNCxqDXskh7Ri
0I/z4XTRQ394B+KDUHAhFT7Du4QVo1tAO7TvTCcjhGwozHvnlwaN1QvrvVO3V0TXu8dpMnp8Pzn2
XFMTZV0RPSjFzuj4cOBI+g/rdtZy3DUg6T2Sqbt9lDVFQ7tMiV1Z2VjXXXiaTfD+tgAGl/pY1+I6
UKlvDLlNkQv5eMRXITq20/w4mhEK7Jqrnskw32m4ldoFeZ12YSHirKuAh8OEu43gUPxAnf1FN9y4
+JPm5XGxCWG8J7vFIwMlfK48nW/Q8myU9XCM4CrX+OiIBaS+b1GMr6xX1yFHm8/kmKvbUQg4TQ+0
rU9XqdgXQLiCsx2Kkbzdtjxs+1WtEISWk7UgD5obStDW8tEGYUGbY4S3El1zTs5EERtL2OP3tYAH
4hYWYCPo76QEzjWpCMO91p7xxaPGjhj7/17EopwQbIjNveVmnHF+4JqIXoz5oEmEJo7DDXoQl3LZ
xe7FfANKip0HkIh9Hy788Y6vpaCOPGKV3/TkOvusoL0fmrAib9Ofqa2bLLNVxFfXbBAtR1PIQ/Iw
ATC3Upci1R3fbzNOwPbEQD4uz4XXGYmyAfsjOWrudC+9q/nOVMBaF5RHkcx7x3XFpkO9CEjykJEp
bkgf23tjVRPBSEKnQpnsRdsCchYt9ko+wofFgHqK7BSw7uU+ZGOzMpSm3/lLUIRUrVh20lYhlPx0
7Py8ulkBUSqHMsS689RjTuruBvpEKlt5V0a5TUTQedwDCmKsYlCSWf42IdVSNVu5a7i4C/oev4yZ
1G8zdi9oYSWhFdpgxU3S9nkzEaDAK+T/txdWNVX0v9QO3GF90AvwZ3UHB3KY1oSZECid77yRxm8+
7eEWCDg+F9RO+E4hlcqi+lX0l3H6jvfJHopIXFVBsQkzCLotkA/sR3/wvx6UAo5ZOfat/Kyzsezz
LX/ypGIeTeyE1c/qv7zYmDvABoUUQ8r3MNBGAJ3wtALAahM3A6YM3Sxz0fLm95SSN36BJUnJMwut
Ao36T998fQLlfaqnRfNEcCPzNpDTHR2zcvj+kXh5JK5idyT375myLUQ2/s8nXZQanRKd0mZejL5q
kAu+/FbRrl+oavQ2SkOBWVtQ06JsJxmJw12QhkrgF6Fk6I7GCOAOHEloC4pByDcVeXkDUsMhhD7M
v6KDkpO1pQQH2jXLzJeS8T8lLgx9G3Dd98tdvwhU0oh0AxRqLsNm2ndlBQuGzOVq9C/l4TzbDAzD
rXdvzJ7BG2PtshW+czfzP5c9B4ndp15uIoeWmjuWWADvovrbpoKUEQdxzJ3uPnr/gSR+maD266go
nY3fFy7HDa91cTSVC52GaAqb2MNHCoNszbWsHEyTDpOo1r7VqHKK8sGnnyDy3Iw9C+NSgGGHLRhn
vt5n3aSxtcGahVoYsLj8XDbGgqs/sugXndtCRcnms5Gh9PX+fnn/zgCcEtnuUANobjbkAprznn0Q
nc5+2pPVuu70xXfoSkFXNRYXVakEM9TxZ8RHXL6FX8DZAYOSrgOAtCv1zOgA+JTU8jSuY4CSSc2Y
pafhBh2ZW7MJRBmWpUi9XAEeVB9PFN76wSZDszHd7r230EHFI7tcvD86QvsJr8Pf3jJpDqXDwQ49
rKXFwIXpRK1xkk8m7H2VuPoQ3s69Uhhb8MAP8k3Punbk1G2yvudoCjNRaVRDER3OEY/T/IlZL74t
eLZYoZZt9AaWhJVHZp7tiIZIGut3DR3GneRe7JUQWKNMK4IdBT4L5I0lQMbVKUkW6Z3571UTlaaB
koa80/kF/nbUVkzGuw40pqYbmoikBQoJQ/HQ1c7Bp3jfpnXNXZBBN1v4HbacP4dTkUgi1tDRiKDJ
Db4dfHea862KVphKnfD8HrftFYbvj1Ttgsguo8RmJtxFHxOb6bzy8wT8kP9+rBaUubqLFKs66JO7
KWWCrToBmeSMF2xpnCeuVDnk4aPIKmNxTkjvE3zNhlAWQJUPG/T/HBo9VJhZ4tinhov7ICmaT4rB
8zw70hA8P6BJ6M1ZGpwrTZMPA6ndeEbpxxM9gxwjTaQ8txwVk43pPZEyR0b7T+8nos2JtfusNi4P
/u7UgBwICI342v4MU+FjNcTPY9UI5toCzzBwlay1lSZzRFPbv+78vFdmGd3DBxzaPsBbA0+PPN0w
wbZpC+8K5zGw/VVwlT+d0UNIHojmatVqgon0zZGlLF6EK5ls8LXjkk4zHZ+73VlfZz6jGMI9r4hR
QdQP0z3e35+t15+OMI+6Uh2gM+lsCQ6q2/jHbyI/XyWpl71WxmPPaUTL2MZyV74nnez1lSyod1Yf
M8z2cGaDv31IcCe7CcpWAsMZMWWVvGWL99F6qR/WWeb+49QsTZ9RwqyXSzbRBiQ9oxV/Paa9rIK8
4M8vKYD3xU8XjTF73o996uA+eiOxD1T5EcvGbcLtsdxM1+ZygpcrQY9GbfChEcQ0flCNHD3ey/el
Z/06roZ8fm48cOUr3Amhewj2HOR6MGxJs/CqEdbnhkUH/C6u1pm8DxuR4YcVjRY25M9PZTnbnU6r
sv6B1PWmmksXzvpSIQNlKAQ718G13ogOmfB8fiFhHXg8DLbtALNk3M7POzVq4R67ocyVNnHF5SGD
Afbb/M6Efkw+2Xnp+t0t5W+++LH7mqbbvg7Q0582YjjZTRlWV4Og+uDaSfA7+3IpeQg6dynbUByG
y75pY6bEyf9GBMfCXkah0kOao6nOleg2chHaKrjGxyIgemc6UcO6GutmBn7zzkifUOIWh3v7ov2g
4Ok05fAlZ2ldUGuCTxICcT4jCT61frSt7yIAjdS11OAC9K1DB1FIySjuCD/JOJUPJe0/yasRB2KQ
ASoj13yMCP5Oj/nL3Fo4PL+rMfhdnJ1DTn71fuuGiQDtc9GEBEZ0Jaq4D+UL5JA2rPoqHirjfv2E
1avrZBqP1CMMOqxurdMcuwRxNGuq2vN0+k7IJZpz1J5+VR5jZ7ap0wXgHGBiqwYLSGBVCZLRrHk0
KhEF92JltSbKz3Y/+Gta4VHVymTMg0FagCGfbhBSm2VJEmHrPOasc3mx/0vY5+6fNE22FA8av394
GzFnLDpJVemxgHn3wZuHNsTDXN9J+xdHiE0z3fZ807lsr4/Icxm3Ccv5aSWKveyyW1Z2j6y4oYut
TE14G520pOOxr6pIicmg6kxur/D4bupnAfAxl0ETFWnTcLIMom2DZr4fvw+mk6vR3GuL/okCc5Tn
QvQsH1nOAlgNef3yUf1HuYysPYdz8kjlmvVywhjiRkOH02pzPFGuaKVNYSYY7c53bBHceR7b3nkO
sta1VFjSMOxAsUwmqH0GC1DB4qojQyCCm22L87gRKUCFvtERaeXCHOJJL5+3HSAhGf1ajzi2ue0s
RvB2L+uUzvVZD/CZpjTcJ/teYBsYVea7v/0tRcLawoWhXzI2zoHbtKJThW39XGIAcyY39+JibLso
k+sIyUi85L24Zo7xQwg/DnEBiaBifDCIBmOOBg/XuJgqM7sFgx95VZbL2T5As1KFpEhWdM2Ha09D
kkOvt9O0TK9McnGhbksivpF+CXBmABsMoHmvMPUIuD3u0IZWC/amIBu5yt5eCgLOzwphHnhVzs+k
kEEclDGy1harJzpjL8pIh3NFeVi+1UGccomJ8OA7L9rDkS2L1xucSMT+2XUU65g6OcNcSCR867Ps
+24S2+FVAkitnt/znk1yfRBjoXtu+eZz1FdhaH9+wTFGvXc0J1GbELduppgFvOYRILRjmiwJTI6W
QZ/NHjwm7w7YauyW0VYgRO05FC7vlTvGLdwJNsdmRRSRtLQQZZExPPNdalY3ijHTncJvq9TuEZjE
ZFdE4+Xs9ZNE5QNNR7da5sIfReci1k38nvpyIhvTBvXeTJ86fwMEqfO+Fsim4xcCuK/deaD3aGtk
jEs6zCV1T7uzmFj9llDDYH4Ucy1wzpoFlV2PKiJVP7W4ZCsLFYiYWPyv6hjSwJGTdVi6+cl/XkqK
dnu/u6V7lQGY1rF29ZnvT/vvz4d7bCp74JFKAEvqQc4Cz3mecFnshK1qYGQifkz4KN390mdd1JHO
hVm+Tklmgrj+SThP7oAk2hGqNtOhf+OjbSiQDGeR4opfE5k0GXxmHMMSgPfiEpOVualC0I3U8kpJ
/rH/QOZ9xCwg2TSUGATItZsSfRkKMZN2RE94HA8XdR1XRqyi+7xfSy7w+ZcY1VFycxEO6JBvf1Xh
M4MTJ/qINF/U1Te0nsQMFBBizVVpcBM50vba1rCNqKVyCft7qXAeuwUNCVOdjTpU4cUazW5OCkUX
rz1F1QMw3bTLffe3WAkUCRuzV5j+dZrmhzHZ+JEerHDX3JzjBkfCdujX0K+/PhLBJkpbROKHx6Lz
Ww7I8F+4y6DYEXP/p5q3n/8o+q2BQy8Vw/gFBXv9u8myYOENTFtMMoyEyFzNquXiRiVbkE6inqg2
/Sj7eyzn8fM11FeKPJNfywAqAxCloT9XxbdO3m6rf0QvZA0DGK0Vuv/fWVfTS0Yhgd0mmsqJp6R0
3EdGMb+BZoMWuWZRDUO7nmd2uodFAFy+jskptcFskobJhbe0wUZGitWeNpKelLT9xGNG5MJvJ44b
StXt1ECXGZkinNRVl7+178gI/VQKsp6mi+Ob8T/H+orx4fyOAQnTtWAL9XAFDuC6fB09W58HMsjK
TNWvAiPUIaEdfG2Pss4MFqqA+c73N2ZHWtADMCvMW0giQ5zn3nZDN1QZGb/prX6iE/Ps484/AIsl
iZdo2WJB76GTq1NgYfFh3HhLkuFUadavISxUUVqHrtBsuxmk75m8LmDATVFi6HNrOe5mzL2yF/j0
Br/spRsYRZ4e98IaOklBSNMjZa0TzAhRKMheChHV2BiuS0WPYPZjZGWWkwqrrsySI/1Lg2M75/d+
N6EK0J+buGCLaLaAUkro6HpQdG01lX/HY4L97keE4h7QA5NMv9WhkkyR3t+wKdiO5ds/zfbRB7l4
aF1G5kHPQg8RmWdBEZCvXQgWO98s2Ae3STTaIzW7BvWR1mbdY1Em63tXCf0U0Yq5Lyd369T8nTeX
Bsc35/6F3tmuA1bmiGa5y3lo7VJCDh+ExhBfDsxL5JBQ4AB1X6yIVEVlq1M7EO7TtUpgkwGLGjD1
wrvikTXWpa1I7Y1iHEey+HOX3HMK2eEXlqhvl9Oo+fHkSuo0THsQZzvqAgiAanaoeVmtDVDQMOLq
w3I33KnSzcHO3gVGynlrk0aCqtaOx05UWj/Qai606XohS/CvALta0aI9c2w62KmlCfu2iZ1R68SL
OGk3/F0NZzo02jH3sK3OAs0KPQ2oUV8+0sjPrzZtJkF6iZ/CPPaWJdi5dFZc9CGQwLqNnT9of8U1
g+CJiRjswCqVQaJlZh6/0EbzyX7WvQ8jLs2Emzu6eLGwq9PMQmtC9S3YtiJ29Yjz/SiFuq1tls+c
VyMZy8T5pLVo3E2IAmJQYk4L/TRiLBQPq1rKSKzIqP8nh52O0x4hTAo42ufpshJxjbRM+IL14aAX
l+dfgjW3fQ01+OLxozmUitj9HGhbJfZh259Nnoe5nVFnNq3yz2uVoZRUYgvSGSk2qqQ94zBCfRr9
TWo9+Zauq9AUaQadRj8kXknx2SLxqM5MMP2bUqVmj3raBOzODcv6JeH5qYap+CxmYEZD6F+38aqS
crhXCQuycN7D2o4g9x3leaW1JNp3nBE4hl8OgprTHpwKPuv48iqsVhd259yA0xtfBQgI1wVKXkmh
s/iU+0ntleVE0EHAnddwZDb8rDiwffP2QZr8v6SCiD4g4Rh0eJ+LScANeWbDmwPyV/ca5rnihCh9
/NPW4SLif8uJ/OjJwrBxLODwPhKkjt5646qJA2tF+p45wOhvK3HaMXgqIolPJMFoi+tEKK7NjvyM
u78cQ1OLXQ2E8IP5EMsdDoxfv0HNLkCt4B30Amgr3bv4CfL4zD5XIsnNFxUWbwnFqp+m/8ZUCM6B
alBxlloaneXXRLLc9F93ZEahxP7+1KEdRCAz6laCMo2WPxof3agXa31lxOYkqb3GCYC9QE3CiZD3
idV1Cdd60CL7zI9V4GaEys8KZ+F/w2QgxjDmBszs46xImoHvMZ65e5lgv30n4QxqV7b3U+/B18vi
cs7ibE4zQpaug+mjX762Bqzmg6aPN4HsNL+xh6iK+mRIPH/2AqgdJHUu4POC54J8qaQGXkmqqt2Y
SEPLG5yFo8aosUOOy9NR/sjKJFezKRhnZnWx/D1Zgb1vObVGbCTyjjVfAvo0U5E8foQ3cI+PUfu4
K2+gkFcHgffT+RRAKV9g75RVzr19NXdA99KPNC2ARdGzR+V/Fsrv5T+b9njZ/jQUxAlG1PhOnWXZ
VGB0KREEOFrpJK8eJGA5bareAetML3tJ2796CUruiUxCya2SZsMhzOompzikvV7qgWSaGJi9oaSk
yVY05IThudsG/yWiZou50EqnREBavMPVlkGNd9fRHJc9H25w0PuOKVUR2eiHPu2MqBKhXIPt64+X
9a2qRghKqo8eL3KiC1ETVtXk4V3uHeUkJDEO4mzFFiCPVl2eW2j81uGxKBjWtgbAgX8dO/H5K3wk
rzTzUa5pEHqks8Wi2RfkFouINuGQmMOdgxzWKMJr7DFdR1kK5A/W4+fUcNOWHK35k029j45JJxym
Pv6r3ZDHxt21O1bx5zy157RgwAarLfBzf2E/WltWUaJwcoQC2Tom19oT0zN+/t5b7fv2nvC351hD
lgB4pQO3RIlE5I9ZaFetWkW3xIjhsH/U7oG+nHTJT2+bM8WWsTbFPl0AUj9+YGsFp8Cd3olXzjm7
u2kzSHpQ4DVsq8GMx+hP9T1pRXRutOo9zYr/uvAxNjMG8N1pBftdihn61EEvcYZqV7FBn4Lc+5p/
YlmMrypfr36/YBanZ036yZoQjtRRj3dQWDSphn77unC+gt05qCswQKmUDkG7/8zsJQd2g0SJEufx
m57jlOkYDaIlo9RMQKJkPc0g7S/7uIm/Sj7KpoBrQjsjbFkCKXHIf2R0GMg25rgR9Gi0P3YXFYf7
QYUBNHgZ30edH+wRrMGJUZo0zg56TNGn6a6dgO5EadOXJqCXvShKZLB+X8oOJB55T2ybXPUpvdvZ
wpTlPvVyODvaeygQWiVRqw+67iL1mvDqc5Y4exow9zWUNxrrBJAYIhYrfVcFZlHah5vH6iC3Cuyn
3RGar4pozPvdeaCtqnJ5qvTUFI1Ozo8mhJ5n2LadQJp0SguhjuRfaEOIM3dyRTyJaUUOB/zVKSD0
FPlw/675C1hjjGEYX4lXYe4VYQPI+Lc1Dkm/L0mDBIQ71s0aOTMiMuRU1YKZw+5Ufhm1H2szIIqI
MCIFM2Ae8/GBVIRzYxWRfivkJizDHsTakYmvh3VarXDjcnET5so5Y/o3ZSoJ2NR3G+C6x7E53c7d
rUThiFngJZE5APbtxw9POib52qkAFxo9R0+H0We6TIkG/yCjlrEqvSJfFEzKYvgku9LX0gnpLV4c
WCdgTxDHNyDoBUlYinous2xmN0ln5nNt1ItglBGAXBSQvymExwzKv+vypPa8vcwRhO+O8CGJ4LLQ
82obp8BEikMH/aVMMzjV0j6ovJaWnDnG8ZYyytq0w+sCZja+yqzOHmPffcB/cRTOELXMt9BJgkOO
qcs4OWq6m4dWRJFzMbu92as/uuz0o7ZNn5UUxH0GFormeo0/2qcZjxtoveYM2O63fvmKXmk1UVB1
XWs6Thj8mKFI873xxPd+5ubbN9LIN3h8Pe+WCPQ2ORJB4et1Mtlpb/wVJp7ufDIzRrqbMiVOuIwg
501fRkShnHB5rtCABK2g/8D8KdxXEqDO7j/wE+kFQWro694JMJfzfKBwF1r4GAdjipEGk/gteMhj
1PLnBkDMD3JTVoyHUwj67rfzLXtJmCAeZblRVdC2GKrCxxJErgDjTYjg1Wov2SW8/vG7li2ZALHC
QmpCoGUjjTsRMIVyil83Y23r9951yjHmVKyrWt0jGhGF3ZAQodjw7c1F9bgVpYk88BdiGIi5wQOV
WRdMR+3S2sCF1Z0OtvzuM8KV2NigTvc3PO+y4PDyvRE9OegWTuznSTWSZ7BZtxXYGJH41FXl/N5q
gc/Q9LryF+b3pz8W+S9t8eUAwqXLNJz4vuSS2coXeAu5A5J0SNTUqJjvFOrXQmBCc8lf7Hzdjdgu
k1/IqyGApK/wljB3mzA1UX2ApN+TttdUYqKVIDtJ4LX9JxT7VFBaY/PrVOsy3rCsmiKGO61beJl1
zcNLgcKSUsDV4yg+bG0ptwzvnnjDvh2tKIk8t7XVkQSahMhuat3Z+hnz9IZSbyI2f1EKZEt2/UBV
0ZsOaWws6VAScLI32LzpE/7nJsc8ZRLwU/9SlZeEJl11Um7zrM3y13cnmYAM5a9xh6tK/1O5h3q5
7A4MQLWXzEjaxt5idPF3rtc4a6mNzvxDK/BhREiJXckCy7kq/wL7D5gRlrwZLLT1SrwrWpml2//x
iAnOqRsmclMRzPBQSeRYSOLeaXkXF3N9l4+Vx0zSgQPkGL7R4/V+oCE785U21dBs84xpA7tB16OI
imCk0ohw6w5pqbGGFGTPriPy4np7bm4cy2Fx4w55o4PxZv4wrD995SPMwnk5TIqr2jV8TqaQ+m1/
Xa3vdgvHObaBlEQOlPzFJs0h0aRLRFj5lm6NcEjS9JhUcePpCWEfbnuGg97BiW2QCxRZxoBs7/1j
ezG7cBM1/iqCv9f7FE5KndK5Eg1awGoBsy1Cu/ZdkUvpEzOkZISgW2CM4r26X4PXnnnlUWv2CIsP
aZApfci2gSKbbodurzOKRopoTgnHIBQ0Rl9Tmv1KuHhRkTF7SxuJggZfh890iPJA6qrSfZogZApQ
xD+vF38BBPpUb9oUfXhQH5SMG4sjzOP8kRMmNtJM6XgWYFm67YqqJ2C0+t0RMSyaCdUMHQVWg4Nr
2WlguGuhscf0NgKS6DR/x9NYWnWwnNFehjfwT0fc50ghU47BQQ6esZf/ZIQ12Z3ozGao/M+nJ3Iz
ME7WMzZDejK+aq4tyk4S06Qi2pE8jWQDagpylQYDBWywusdMyidSJwp67jF5NvVtpWWhR3SY2kXM
jH/V0Ez4SKdKWBkvLytuicANGo7NvxnznjXoGo6e+kKe2CMQ2JcUFh9rT54TkM0El+eMPIxx4SIj
yn9BkqJJ2BaXXu9r9OZi3rS3s0U+sAdx3557bL5uiF3bdC8SG3KW6cvxDpw7k5TBSstCxTDVrcBm
h4QxaQXBtTowEtKn7udukUdf0K78Gkv2DQfkpYk3v1Zso7vJE9+IE8zuBoo2glA+e2jLxBjdBmBA
fWLmvnYdOVFvVQxy5rOFFEZwdnTZioB4+AKO4fQevJx8De8Es+ZlN59ynRHR85yHmrhbiA8nT01j
sfzFwOUgTGB+rZFcwvn6gRyUhJGU1OPoSaMktR+3aD5DHmAQy8IxeZUatjnQmUjBkohBxEXAkCca
Vqd+LErKvw9Ng25XwwUh99rwCsxXwSus3QsdRkp2hX6UJXRbDRwFL3ZztinZt5/egI2REGI3crw8
0FizmWzW9sYxey6WBQpVg6ExelG25+6UA2i1VNVkAdNvmjAQqXhn921TkTaYXInoxRY4jz2aXTMg
uVHzw57D0QInz2r6+9UGRwWxxxSvwZCuYBl68FCC061VVhr+EUxDw2dPkBrat/EqSZk9hA49DazX
YB9gBDrLHN3QncZgIkm3HPFbZwMtm21uuCTQzeljjWCBYFf/GItzJSrSOkzUkliN+8Zhq8jQS+hb
y4cd/W68w3+jCLHZuHAzXnFA2BNJb+Io4NNMqSDr5D66sAQINzyk5BEI/38Rw6VYkOpNQL7Iar9A
WVWkEaD6L9SyEyTaxEWz3y81Xf5IgRkgA4Xn/GUAOYIQLdjIAR0OueLRUOxpsZalE/krIsvesamd
m4RGu08jrwj/JkTcsgxk/Vnu8utM1hb1E9ETfJSIuqugrX/NdGWMJC6TC12H53EarT+vEN17jJB3
C3S/oIYryCYWUxB8LxTDMFvHkkhK1RnSwBHcTrXEM8s1QV4PcUTqtVoGo0ypAm7n46/gHTt7cQMB
OfnjIZVLjV8Gf9lnfA8W0U8toz8k2pUVkAdMuFHZkDYB5TOJkSm75YxJcwdu6jSxmZwQJDt/P8Cm
JJU+rb/3YI5lV5BAIS22jpqYdijeV4KXk4ujjF+1ybUBI7gLohqICiem4j3hqt1yhSpWX32TpfmJ
dtzAzzyXSsYM3e/bW1Ys5sGUtu98pxGUb42b67TAqAuSY0CLyLVvJZwLm7hNK42eNG0iTOjDr6g7
U9hTKz4RsWfHaemYbR4Q9gvBVzVBZiVzEx0e2pHDTyvW+cvWXmKCbUy7Z4Z/FjN7sLl7hdJAWHsR
wc+36jUKE1JsuSkVz3BjS8IsaFgSCUlPx0QSqpy8XEz9JVpDPQNWK4RJ/wPs2s/0jM2HMlCE6OoW
+pyOSYCTyBjtYqQs1KBkeafIjFo8JtOfBRpCQ3qBWGYGShpDAAzODutC66XnOMPbD1iZxvTWPm0E
eQO8s1VLFcFwobGt7n7VW7S1TVZqDdOWIr9sEn9fi7BVTNAWA4lCstrTS7JiwVvAK5T04VXBUTIu
rb199bjvP9s6EIAFdJw90v0TCi52VkExRGUKC8QLb/tIUOx+VsQr8pXUXG4OZ7S+LBKsNadAnzwu
/+WGZd3kRIEcqLuCFXjEs9Nc3uX6t75IQv+7lAMsdw3zwNDQDgS7+AIROGRG+hpq1rHHYoIN/G9z
MXQwZOFiujyF0K4d5R4J/Way5ODoekkuk5SKsqh8hRvXXwe+pJL2d+ZpmaSsgKtcp2BMxYNeRkAt
fDu3//Au5lrhRMdfnzsyWLSkv9d3ujvNwkhhCISUnUaO/jfLQ1ng7hMn9F4qXrC9tnVCDlsoFq/4
RUpNW/PdBIipQtk6MKIu+E7XLBw6TO49hqjRrXsf2y2aZmlc8BpKisGwkWBDgfNqLFHtI1Ueg3gC
kgHZx1dT8UsOOThwyktFCn5e0jRztSopFhyWPkfXBohdVulcsg8EQxGTiXVoqmRVIU+2mU8n3rC7
9n34d7yATvwAweQGDUEqyGE7pY7GnmOeD00y0NdUUR/xi2rEIzWJ+EFv3EQ8vT5kjEhYJ9alTrI3
YQVs8L30SfJDw8slHFzc5u4jxsIYss7dH9jEZi9a1b0hQwMvc3SLaOajDxFMM6vnM/l4ygaikLzm
7hz65R3XSLu3YE0689vKdzEzXJ7kLmNXHMgazfMhI1b4bMdIi/eYsglHDYsKuxBbj/SmWzOoXIcP
98sk7McF5zk7fYOuK0PepaOEZ5OqwiRnQiqyRsKCTm6uj1NGYNYfqRxKYcZN9tJQ773p+O6hAFz3
9caGfnQv/1tFZcP/bS0ejd0LH2CP8VCGXw6Daw9VXHgOr76NALjkTscQ9Gjvozto84Wc/7hqhODa
fdHscmobk+71J0DOW88eQJEbfghy9SlYVvlPFLSzEszpHPGOKEJ3DmUXFS7Quh4UeoaioHMflEyy
lVOxH+nmEbJzsQHG12Csshz9gsqhIbNZltVQsHgN+lGiXBl5ulXdrHXitq59mYYmLe/FuVLsgOsc
3oJqMc+Cqh6JBVUELitVCAd0FbPoJHifjQ6S311eHWkI9PohV29DHyqADgCUhIbbEcqJyvDddEyK
36kpRC67BCIT4SjDC4iwpC+RC5DmLKpOyWfjIlD8+KOzZqWB5cmAFLg7ZY1aWmX+FujWfacbAJVO
Iv+4XuJEEBUgwBSKKxrrGUHsbRQMRm1TSw2/B06R3LTYE6phVS2SBh0v4k4Q8YqwOSLJa/49ViVx
rMrk5IX5v7BOOknBN7HmWbvVPFqf2ut+iCm86eVb4hTLTqLNDBrFJ3T5Pm6KPwctp826FqVHCDWk
y/+qE/4QEJQp7sIFSaW488u1KYefkFkMpS93/ZTcJDX9pjRFgJFtKmRpAA0hCURrm4MGYO79O7Uj
vBJQY0l3S43SYXjDmlzt3UPEX8XOfL0y1Fev27Qy6EN08sVPDpCJ883JZHPIIU/WUcUMDG4CzR9X
dCkkDgPoQOEC32IfRObI8cf4kmCeFubh7d3i8au8LIvAtjjYTxG7SHtv0m6xBCk5qw2JZs4THkM+
22gfU5tDjGj5Plq8eZQHXqHF2u8fZf1pcyk8JHmwDM5f/OP7Gmt/j2YXrrAUase1KwJYGfHf6jZV
sG4gTaBp7Z4ednu5yZMpGiwlKFsypUCyYSpyPiDlqfXn6gAJymap+FtKd3lUgVM4rUEBOxxNG+3J
fi+bJ7bnL4hGu7ntFfcO7+np4hNl0S2hLKuuMJ11rSDCk9hY1M2L2mssTWiMH1QLFA/lRZDqP9Fm
ESaOQ0FzGQzP0VC2S04I7Y90iD6quKmKgA38j20gRoeiAhjvtzBMdaccMY0hTsSYDfiGskwDp+U6
X040cP28t0+4JbUtVGiUJ2x+DXg83ExlBfCwx/BfkhIyBA5ho/bIgE3z9nn1Liy+mvu/qpqX97Zb
93SjTG5ekL+VCXTpJ4D7N9atQfFvD5HRhhw2/bnD72eN/5CfWQlFtyQaSypPC0q+7m4e3GIPq2R2
538Ax7jy0G/H76c1HHLUcxqTFRmzPIj/TbMFKu7/pxEqYJY89B4fL5BvGb8hgqsI4TwvUrHROkQL
TSSPfQ92M+ZHAAfRDXzcIDd/h3sNvfG1e1hD727bRwVPe76e9szAiIZWcCF31FdxjHnQKQ+lFXFf
zxBjRAr9j44GUmRdjd9zXcWsjlXGzUSve3vHkDue6oraIPbRtXhHUAE1nOZgBvsBTz2DhiLH0TrI
FUnDJDPiJOb3Og9Z5wyqjzfL2QXpA84GztiM9Zh0UrxCX5Ufe08nvfZqYHZ6m9qXUM6qwEs5IVnG
m4ndzjbzAqVtHIchEYKge35IH+0xcxL2AXMZ76OmSJTjeqZFpwGKW2dFTQ29PBAeM/I87pYVrCsK
9HR0JM1Jk2n0SoVag70fXX+DatMr58gR0uqZgCYLCoDqnO9f2jJ3CATGCO9oOck7fVBPAYnvRKxK
NSjV+AG4sZp2FwJ5qE3yiTW4XztFA93NS9JCukIEXcpGttKuN0Y27j3qrSiXlAK0RVPlORlkhQjo
Xo2h1IVKNTul84bJrV6+/7lJyGlE19R19WN3RZKtusgwaeMhjJeiw9QxISJ/2uP0LJtWvhu1Y6yT
MaAMVAPFHRtyGEtEj8u3EAcSziQrkEyGZgzpUubeJ22QzExmvMnlZv0q+oaohqJCIOzfmDV+r/Jb
78HZACx2g0OyXUcwK3yNcfaI/F93IXjoFUHxBFwB7bJ6qt3Nag1aVLlpVW/2N+yZy7EBwzhQZ1Z7
Vdse7dR24vNNe2aboQ1oK0SfmhpIrC3jWYNWZ8/6kPC96yHniL13IMVFLmcraF8FtiSSd7jKmXCh
Rmx9Vx7vxGZ32l2g5IZizznsLC++Wj+LBRnXSs+/qA4cW3VKp/aAJ74Vtz9ZZ8tZ971HgH3a1wv+
S9vNvoXG2e83EpQUcmU9wZGdMJwMuPTNKCfPZ4i1f1AmxFZetOs/RqvTRxAQGVqfWR/jI0wgBN0s
+HdDjfa46SuJcNX5i6hcIAwv8f1JiFaxumpYFVlpmjpGu0rfONb43O93D9yJsl/tC3hs+u0+dVnX
d4T12FJo+QuRtrumQHhohh2MIqqkURdlVwuJJndEXlRWlnASB9lGsxVN/Mcor3ijY7NfmjpuJ7ZH
2nfqmYepjRnrRCrZTDJV9AdxQcouj0yZg+um5BgMKXH7YlrzbNS9P6skhIbW/7+Ql4+KRWPhxDT7
bP5fqXQuCTUZjfQZRS8rh+Pfgrufys1lCoSDOWHWDEv6CPJRBmliBxakFjsv2apO5CX2hrNBSu+d
DH/w9V+4QQoKQ/LfGZxEw5CqipUcmTWoLsxZKEI6SnNwWEP/pBmRvDe1JaWOnSUW22WJJVJvRyR4
ivtV0S3EWthGQWynYwApOh4ZlJRKWBkH7lRLCycGQnWCBwErrceIJ5KIcoYRec/cC1rPsjIIqspA
7Yh1ej3wSIt06Z0yqboxm4pIzpG5eHZXpo+ya589iXElOaNHKmkXcJ0EjfVofAmULL7Z3fWn3G8u
V6WkQmFv4GiRvYMJBNVr6H49HY7hCOYx8bINMz99XJxZFCLX++YyZHJDMukb7ZJIrgMFuIylmLXU
qC9zUIUGbRyXAAPUOP7GFB201Xog8Knk0Uubri7roA2PXa9M1qP8VvkhoKfn21E+gaSwE+bKgmm4
QmGYmYeWdL3KCxc2rsPo6ImNAQfXrpNV9XkeJwvYtcyAxETWe/DTbjiWGI8zkuC2kx1udC2B+ysl
8KqEgUKrbv5B+Gk15c69pwbd4UU+36HB9prDhUCI1RBaWJTmiGF1SnbkBoP+Ue16+xo61Q9NmYmo
LeRz8cEmAXw3QKQaIp23ZSFgZGzLXmnDAFgMufEZCEaHi/Hcps2rhCfwasy4Einityx22f4nZF4V
88iuHxq4IdQslQ0MS4HKAwdi2PkoylsDfFtUXjK/mUcto7NICT73ib+Z7V2ucjzKt009FE8YoOrw
5H27pYQf42zRrxKpfBj9PLl/2nplhqlHxwxlTaXZNyd5aC4ubu/V2QZR7Bi6rv1VDFtVjAJnUvpL
yQZAVd5nQdA4kxV8oVhGHE2SW0qg9OM5XWb8gQmWpeB+O5Z0OSefPa1JNbFTibaUmFnzyahCdlWE
aHP7mA5LoustULJ8I/e2X/7qhv5fgJ9OOW1Wekp6G+ZGhy2wTQADDJcE44bjX7hqRp9uTyyvzfZu
fF7WMZdeDtPYcLZL098NWafHFBEvffmHvwN/pXIz44MPjxqgwz78rerVikCzPZmYig72v3R/YQIM
s1yV/9mLEs8cATFcQdeRNxCJ1LI6P1SejZ4OkpOKf6twsiov5NOUgtR9h6CgBP/ieYKZ/g6G2yV/
EE0RgMAYJ+ngKAtf83k6s+Xy9opF16dUfl09aWDESDM/oB8ZCJa/oq2gDUyN9tz5mtRdM+7KqHw4
MXWmK4zHDzvouRT0xh+fup7Cdih1ls5BIRGDOi0S5JpL7JAdGxieDApFfqX5sn1uMZYPb2ZgX7H2
U9lqFfI2h/aEZpl3tSLowkrtrhrtYdZpAgoMm7MThYPvHmF2G85l/hp2vwTdIb2B7zaYOaKNP0s8
mCgNhHA6gpc2DaZuxhg2pDzweSVTWeBbEgr0Zv4DQGBMaq99fQWdgGj4OqWxui4Uft+q3N5WxURB
pyejKbWeIy3WV8OcS9Xug0G9N/4Rkc4rGPwhbKpMRKV1J19PE6IovAuXKxE7LbowJ3K9L/rmJbZn
+gqFn8L9xUl8ERHC0SQwTPzPL3UpoqTiuOz9sHb6uOE97aPYkELW68p8p8lKJ2Kf+qaUXD/xJwWR
tqUN6ZUWx/D+4fizycSkcYyOz97GAAcjbXvWEHClmdarDzvVZ0TARFzVxQDwT4pmqXNDCj0f06A/
goTZuJARmFdFd4eJJdwu98da4mvrOV/yD7FSaBjqnf27Rno5JLg8z14de1dcweRPEMPktyp+JYFc
dRX9TIg8yAUyx3daseARdnUFpTqO6G69f/+wp4TjwYSp0OsGXYExBnNUa4gjMUpKxLexDYXoVEca
GWDVsGj3XQGWOrh69KURdkHHdUF3xbjI67d5vUGf92Gv4zPS9OlmwBHfgykKEe+6BFwbAMLyGLCn
35C3f+CNuBG9gwRopQl/qL1vWhQMm0E1sCCBFwF/6YQAl2o4VZyv79SCsVD/qD15IbUPJ2DTzocn
6EkV78Ptl7LmoNaOSEKDvLLjFWZcTprvKR5D+taoGpALOcdHOHz6CBUm30ScsvS0E1/EI0fIibsE
pp1xBy57xdWkjNscm9hOUylrnpcBG1Yqle3pxhqnRcYqMW0IiVgmN3x9Q/mYBWyGxD65iDtmWN+v
5X86EsiVXBHJOeWJY2HPAw2Q3zVvWKtF6/0lGSf9NqD1bWdOHI6zPaobzLnFqfim2vgAXr2eCnUq
LeSMuscNKGF/vA6Wmrm+LM49fMBfR9JWuyDzQrPcxp7yZcI/FawfuBEO+SCnCMLDqhdHch40X6en
+vr5B4yqyQlkGV0cxJe4I5RNHGI8+32rZYtUvjn2RgG/ohSpykK33phDAdI/ovKLN2lsZpHgZSGY
ogRJ7y4GMHN7Q9sMjIJbN47mYtk7pYxZqgSfc2XO4HgK59sJtvUukIvhz7uQMTexsZ5PhWaB0osk
qhazaMTIp3XL/zDrGggD/cXhw5C6kpsbSLciO93x0YqQHDrU+djJbXXtMcCy1uliHgY6l8eyOraT
zn4v/Nm6PEpW2klEDDPe3hdE3/3xUyWJzFpBXJ3JdVBiqk67Hltm24rKnZuQE+UUz42YkGn0jvgr
ft+cXy1qdXOtOadePNtiAVYkSnCp1zFTRNK+cMSxgT8vf6FpAKuQhbGJrfkKSaKdldgekmQ/5S9p
P0FbWWHnU3RBGNpeyPbzCzN6b9AMC1Xn/tDX1VDCTIwvA9RSSRXK3mkY82/ZrIXj4FPqWJ0SHYpo
7Wp2PF5kuaR01cQua+6UFGWpmhUpUzP/SIiuE1KXZUbBxp2fZEa8ncDgghaKBHKfU15rA1uai4E1
HD22+KUYRdb8uzvZLdgF6+hPjofGMRw5d41Rg46K0qHZTUXjQOA4LyZD70TleC08W5Qh7/4CRuDl
leIffVhZBQyFdEQPE2U1R2FnmCPOypIVy0bNjY2jnSubqL7Shd3uC5zraqd4fQW+Ef7OGZsOiaAb
8jGhx/E/ZIEWvirnXJBXQCmMs+h5WcuV9o/XneM5a+iNbZ5B8uFPZRLU2dCdbfPpWHrktXlV8/Sb
waj2LdCeDgSgOxYsu9cvkjBW75xt5sysk/tYD4M/nE6DHjW+EMMaSycfgIiouBA3KzEDyVJ1LwGK
lmdR0E3IpM6tUV07rEUWpJhliGtr7dS8u0I36m4HyXmyeXVZS4Z1IGAcpt9qYschmEhIWaD5FXaj
rJvw5HfevuNtIKsnGqx9pEzXLTdEF76kRaIyxu6f7uaVAmrpI4z40J/TtgbPpMtwtAGK57SvmOWZ
f51vb+R55/3OCXB79CdlHc9HcC+xJnrm/FxT+BMXbwjfrK5aQyy3a4X8bwNr2q2nuuh4RGMaIpZZ
wOMTOWYdvYxGLQ1VmOZMRaOfMaSlTsgEusI/HAI0Jl6p8BOnf24WpQW207ZPMS+jwyXR5/QZCjhb
Ya5T7RU4z74LwMhyJHDoAoaKDF9j6IYneCM6SRH2sEh70o4K0e45z2Qgz4mRw0A/CPH23BUcoC8w
IQGBBUxnco5KTTX6CPA/jXWjxIvef/ARjMeFdStgcIdhL87189k7Z/GUuVqY25fVaa39SZ7IToDs
guA19cKS7DMyUzugi4hwtfSHPfkiNFTlWQ2nNNstVwKJlcdR7GI8vBUhx6PGzLRVquupFK7cYcH0
ZaVu1mb3PQOfWX1Ggg6CcXKFcSvP0jSzxKb06PMlPLg7gfXxInNxIOZupO0qqvUgcpgKpXeJ263J
rz7oTN/mW8oKf14Ob2cmuNhUQRpZNtfR1CfHWgPUJoCp27opljc52sTEM6YPcFHBeDSnPRLK0/Q2
IAj+UQl6WAsfTjlOYlw5f9b193M5zHR+75K24rv44rJo1A6xBJMG1EwPh1aLL0UE574vMgXEad3B
bw3MvRhK7W5abYwGCVVg/yVsnRQ7ywtJyklcXea8+Ybo0vLUNJgeAX448uZEwolcKRoEYvLJ/cWT
5/zBHUY4QZ/Uy6yzzUJXjjtMIevWR3YoMzoa3A87V6RdB1f0EVx81w3Ljfx4oeePf1xvmhdGdm5m
ePYQ+7GabOBuMq+Gv4UJjahv/77xJC6dFnE3UWHQJcWbDmvGKP2/erB02g0ut4utZMcbdPxJyWOV
31hBr4snkWPi9KxYYbtTi6v9AfXuXv+dMed67XLfOHgZN+Sq8IOcSj607EYjMjL13rG4ttQF/RDG
Ook38xLx8uTVNY5vYoN+vLVCBO9DD++sfje/wozpzK5r51Rv+miI4sbnqn2V6NAOe0Kr0BCZcHBe
GEniR4dHjfiM33YiURoJeIwmmAHvgTub84i6QZb3c3+KDka4HCDNUgLAzcbnlYHR3+He6YEq3t1O
BQciKjpI10jQIo/sfcM+L/dU/Lt6KZorvpmBaz9fzKYtJT3s4d1tYgepbl6org+Z6qTCOqXcm45A
M2ihQ+8Girq4Le5appUSeXnTB499rHH5LZzD3/dsKdNcXt22E94l8gTNRkaxYi42OfgIlLeII05I
2myMUVKbMEeZQVYZq8/dAmL+4fKiFCsEI3QT+hiUXg3IAUh64eOozkKpfiEcT9zlpzMENoKJgDOZ
eYnRUPwOGnlI8Mrlzzkbucgsebao9KcEexY1P8NFU+dVnuyj5H+R0JeIggZTMIk82X3y0pZAkkix
iEi1r/02fVrh6lZLyvbxU2aRPIvk6gpxqPrdVfu+ZaYAWBFC1Ty6ge69w9v+gqPX+2hGWROBuCAZ
ujslL8jrQoT5Mw2PPfnM3xjiFdGrjhcaRwmXmOmkYp3o/QF7ugPaqM98mEkBZjLwDmqQRUVudF/f
Vqw0W+xJ9MVYuOecEl7HBuuaukvhs121yCSvRaqxfIP7IddhEV4DQvQNWlaKutEqdEiO9oeQYZ/k
+t4NcSKpoU0kLb9MslJ8Y+vq6Acne+XYWxvSgtVeux7DyyHfKadL2WSBHQ/8+5TdOqiYYQ2Flufu
3byrMhU1rNJoREHd7BjIbutuNwiNlmzCSWhvrglvkxObru6y3Iq2DEGrbuwy0ppGcFvJK4flExCI
9cNxX+ld76jVTO9AgtkKpskh/oDqCvTPGMUkfKZwULn3z8lpm1URB7T3o6TW84O4XyXCYneITBwV
fFJ9umLAiPEwyt1C9ScPs99QfxTzhb9UAZKMJ7Z01L+GIY7NhHm3LONCkSiqjG6MchdowhvuBilU
/L9LM3S5boa6vdnfjFKPVboOVqKKfB4ZUYWmieT0bjATB2DH8xtrChwSqWbgxd9O1wuW7TJowtBe
Td0cKTk8g+WcaaodZ1Q2S9X3qIpLgT7XVk59+k3LtX6KkgMeqCfAARnn8WfAIb9PFEapajdQ8m4Q
vnzqSoOBsllZO9y9JsbDPgzNv6B4P0PO2wEhr/vOa0wf30oYH1dVaaV7MjsUUGW3REjagg+lobyp
F5fTDT4SU+8oyJotgXjyT3377gnB0eMHtW7bWEWXdfJuKdg49jvlCoHb2Kaw9ks2r2IosvfDmUIb
jKwDSg6S0MdsuIVUKGyrEbqxjuwoZt2dQhi/tGn04rEqbnouRkx8fWgYUrWLBRFsZ6m787O8mGjT
GLl/9s4PHAsnTBfrYTC0nsLmpNElWdwnOVaWi8pXapvMV+Iacj0WxYuZjWRTxwZN94Bpp87sbtI7
StZwZptbhqp5iCWh4aDWrYFdPT1txtYJoG8PUHCf9DZCdUf8zVVd/jbvPoqgMkMQV2vIGKAjy6UR
PH7hexExcXmlUKNqKtijNJgrxSAq4uPQjfsAETISbZ3ZAhmPbGN6X3Lnonq/o6B0tpPLX5a8m06O
KeGbMn89Ghrlo+CI9mP1zZ6e5iBeSzEVsociFKcAbrE4UB5VzwifQrGqp1qbZb6u+sjO2lkPiCSc
jUVsFo27DHxfAdlri4gTghVUKLLHPvN5M7kZl6wqkuWo3XCp0cmiU7//SNalH4WVj9OJirAJc6Zg
kFo/pNMYUwY3DHzk4y3zZmNfBdsk8IAVTBSGZFrxBfp6hH7TRQ65jdmFseCkHdYJ8eNJPio+qlVj
IdDRZWC6hlt49BRov1LKqfZEdDMImfO7wcDptp6k9N8iWEg4mQh+U8SlMVhhmlxuNxFsnH0zN4Lb
U8xt+1slB6nR4Bu+SBKJdu0b6bQsUHKjx3mZjdMjOOmdkkUd9eHFeFDBRnCxeOOXSE7KzfLQnGX1
rtKf1fdj8dRgJtTuHgAbEW+vsLTKe7qvwXt9rHL0I9x3rS+50YK4gl5HsLhpGhPasQYRWKwwSMz6
sjtbvvzXX9UJ3t6DzxxmpbPE59UEiNcjSDhMowVRfFI2fAzy0SIAEgXADrzhAD4b7+N23pnf7FBO
9oxp+USNPNuUAxNXD6lcPy3YtZS0xqQTnErCyGGgnO15F8zMXKafQhSJ9ooE2UH/zWiwcpkG5b4S
k07WguhHM6+GHxSBl/k9baxJiQAApcnO+zZPnlwVWSgFPX61a9CdCwQAftr9HYGi/h2uyziSxjBO
//Raoxmi8SPpswmerzG94upjRG/z47IDlMfiT/hEdU6Rkxb5iVUfRwsKEGgOffas6oFvwIIfIS0N
b66fJ9A683WBy8aql+FVautzRrm/sPqXXXMIKP6rhYX2Tfv5b/r5iZpbsYcB/RQwejSWcko3JnSE
PRG2d8RoCDBG9PwDSn1UrvNgksV2HP/IbXr016yjsUpZt5BG7lfGbJyMNMlwS82e2Mm8kiKPidhS
lwPdH6WhQQBF2ccshG8S7miZukeq1R1mldfMPQ4/XkZE+Pbl9/5sJmY478rn0LCMpAgbDPRd0SA2
6bDayRod2xUdonMvRswtNpcWy54nsVnBlL4Ua8RH+/1EuvCAgI4BZhIu8JS3hChgRa0CN3EPS7yl
klA9q3KzBkuPWOiEsFCKmroC7bTzDA0/8QsjVORHvOP/TofydKlJOZlUGRC8uoWqp/L9EXbPZeVs
KjHpBuwd8GKva1Ao+pWf6gEGlP/nK6IM8IL8O11ZD5EIETQMpZpQn9Z/rhjFnWv2W+czuuuwcapu
d/actSS82CM728eB3wRqr2yMmnTYKi+AMKAWb5+rTALL1b1bb5LoqKR3o1IO+FSv62U5vAAlUXn+
KztSSSZ1fqejMV+fTGjM6hej5tLHD5fnrZ/uw0VH2ZVNKpR1T/A+zJyoZgPO0FM3wkqihBFkxjYK
oHGdNCmDK35ygVtbI4qPbCsCOq1U1wkWmTrpUM/94O6+X1kgVo2Rqeojvsj6l1s8dAo/nDQMMKPD
Bs7HP/b+nGPY4S1fqa3vBz7XU9fbonhVMfr+OAeiR0lcezIuAXwB4Mclv9RjWZV6dQajLV8Cq1ru
HOPgLYbGCiL57HtzUyBPz4+kAtM7LBYEpgNlWoyNRiZq/wXloXnzZxYIQtrlsUZricjiWnlx/Iud
QbXlBBWLQgqkncNc4hkQBVp3EmjnOFcVSk6pR6BbmE17PtG7j5Z2RFfU5bS9+Hp5vZ5GXjj0Rc4v
eUaFQd/0ofAewdKx/LStHDWNIkL0UzaEoGFroJc6xfO1eJHMk2G6wGGv1OBA6vVvrSIFHkKi02xt
qGPNqQpJob+7Hh4EIf6DwPtmZDQ4F79yPSoAdOzzWj90Boj+wlNLu6+MqI9d4QBbD6HQ6LD+y/F9
vfBpa4mnE7lnMTvuVQ20v/NBGaoSTflCfkRxY4BTXGhs2JyCDtQxJhJtNzqIfvHdP16jl4QU/gc/
58796nakUKzoESEWJBJcKK+SH10oPy6Trhevya1rJOcH9hoy2x8Yr1X4qSg6DUEuTMjxto5uzK5f
NGAcpkTo0F199a8Ui600KNKGkaHYZ9F/S+EGLf6VfpllgeeEuUwgoT71YNCwgyazhdP4CAFIZbx1
KsrMQS+921+Gu2FZFYOjKrt20n3VehehRRe6WutfJlrx+u5HKz14BbWfOwE20KVziClNsLJ3yi+X
gvnDCYkOKT/1KfOJvdN3KLg6LyC5QWh/R7D4o+D19Gqt/NC+K7bYvKF/qOW0IcKIqRn35Ci/tI56
4uzM+HYrLN4uDHbpJqoDv1SQ27e29URvLvnGtnHzmzAT1biJYLygtkNo1xuNwrBHdDF2EGafu0jj
XM8OO1rh5LX1pftDXI+HZLo7THHh59mij9H50Mbh1totQCGinydCu7xoeh4vbKdYHMbe3sF2QN1D
20V0O3HFPjnVhUuOHGwrcdipHfsN1MJ7eUY86xfzRl5oFefZt36nIUM9bTwP5cbE/Q3TmTYEaFKZ
QJeUmUv5fYvIDEGidPCMSPwAcDqyh9/iwjmBfaS7J8Z3UzkYav8pFdN8nUzCXcWjuc1KBUDofNqy
rk4sqdZndFOTqO0z+X9txvkavcvdCzGE3lEKioyG/bjE28S6YkakE5BA5NaoCAE+mWZYk0Y/v9Xy
A4/R8MMMqOq/LBDkPMWTKNuMQUFJlzakeKhoa+uY22A2cl714XZLLwjfinJKBS7pw5r5IBu/uXB2
QunyjBOOke3b3u35D5R56yFQJe1uqrWUCNdsI6unl2nHPZ4Qf35BhkYjf/M4Q0hqH0E+n/zTLsn6
Etgusv7uXQU8aANnls0AgwS+eFFLzD1YSTiCoqnTX6IEgIttWvSQr3mJnb3pzVCTenaRr+F9QrJQ
NLX6vPQX+4VVL1eB3g9a3zVOhKdkpBdoNqXK2+eRj/nOXxZDZvg2qZaFui2W9MCw9YS90VvsYk+V
VBUoy4f+8AL7DXh7L+32ltK6mDctQKnMKDfzwbfUG+TfqdDTiXsJ1db/U3l/MBxe6EgUh2bvR4PQ
p7zVPtgAYSR8mtJN8QgfDlVsdBLPLra7HfigXqdmg9qK0pKNUOmcO5EcaQ82SN6KV4/zhC818b5z
Nvn7wZDqdHZU6tIlfvoh/ShJNTL7owhg38+H1ia6Mu//GDI7kzQ2jG35QupjABSYYsax5b4E3+Sc
6k/u2utorXhOePit5V+3mduRY3BCrw5b+KSriNFOmEQwOPLxj9PhlKthPlrJUJEyEFLwB51eDa9e
nGC1cp9Gmb31PWr2HD5l2cLdyU3i71ex1VNqWqhkJqiboHGATt7C59ZmW2UMPHT89dmdDxYdDp+8
xnSLyJ/kxkybaILtjDfvxDrxZtoQnWDsPPut/g8v7cj80R4owoDJHaE223Q7PKNtbuqtaOYhAe2H
FtOjbFCJKm2SupEzrH8FP9ehcnhcFmkRRqXo/dkvZHjk7vaucQrINDNgRA4Yq4WNshDNeyrQVnu/
dE42yPBOkOHwVJAxIBuIvIQUxJFh+Whyp1mhZHN8b58AS4NkB6Y+pOTxgnYXkZq4KjG/Lk/bJqyO
KWnCveStS/sXcPbM+uvOf8US+yVtiDTuDpMns9lKOqOE6PR0nnS5sBePcIvV+fy1Bj+KTjIb2OKL
nFuRiVTdWXYF9yu5cByFsgKwtQPwzF5rB8uvDah0E2gszJQSE0Hm5ody9KmaEBQBtwuyPechtkRS
66TmG3jgFCZumCere6JXNM6zrQnjH+4q7jADqJwMfM0MBHzJHHYeKnSZLJa6bk5XHpfKghaYbkjB
ZYUfsEQ4Up1NuWJT7kMFvIdLkykM/Et2rt4y/6imsUzSe99opC5J78YRvKvkQ97p1F6Edal/brXV
DZEuMZPA8ujbYPnr4pkR2H8n3mAkN/QP7AFvxMZRUinaBFtKHo2KPpDNFJlhZv/6cDCz1g/GU1Ua
QFYPQpHd/DDR/0r4Tnt8TE1onIoaY50CsmQTNlGWZsMcu0CjF/VKLXfAlFyp+NEMKLkgepJ2+7dJ
xIDvC8D57RuyI+5QMQUM+31HTp5HrPqkFZDbNxYYSvEAXAhM+Yd1GVKCt3iFuJwPsblnfGhwPMBc
CqlfcNvVXpF45TGhX64dATM/1MbtRtEH4TaKOamMKmNFyMK63IV9G8Q0YadZ8clsz6oCjJOIame0
rbY31ytjpXteKddc5uG6VGWX6dFgIeSmpo9/OUxSDcqNanv5vOKsTesRCsWF0UBONF2+kkHPMgFD
VvdrjtPFRVooLVphqxvGqqpUAnfl7XbxV37ijXCNUxEZOuQkWK4KzYQBa7ZH7aLEg1sBf684GK8U
Sw2yqciNbJDykAPmGRJL3NEC/3XF9oBSb9ONpjwIwcamhJT4csfKb7sfmsC5kF+gOcdkStAPqTlq
JpazaTjB+6gV73yzX9auYuTmaaL9Iza0hmom0f1IEpKk0Vd4oPfIGwNNGGAlqMTyya10v5WJKUk5
HViE4TfsoZy0B2LVkDkogicFWK2xEewzL8nGmCHpCCFDbUGnUDMSzEQjNoU1Z3UIZKp8/e/Z8oUC
SVaJJyNIv9RqxyfCoN9DBhMBuldLya+Bt418xjJ87Lb7PjiihTEgJNDvI7Zy5KNl3BDhJqXXJkok
PnDN3LaBdHesUM3xLn7gnplVl/ZVY/BBAll49Qbgyg9vnDD+Z0h5WIm4/oKbYki78yj5LN842pX3
6C+ZgiMesFavQxzTjA2IdwaKtZME7Zth5lWEgPMjvjIJ4MTPgMy1b6Njh00umwyP2fzpKzdGTPc1
GDCgXlkjQYkze5WBDtorNS3oWGRbdnVMaOTUs0+HAfhTkAqiGnx/vhqdGVxCijEmyDSp9uEpR5s6
a2i8hR6KPWM9l2+xOt8pyVu/qp3KsMnE+Xd0vGzVyt+S6PrSjlCsMgOqBRqMfAIxXVpgAh7qLrSK
4sJrHrd4kv7ZUR21RFaV56afvIzDCMtsOuZ+NGGVwKNSvC16W/VSl143v2Ol5fg30UoS3kSeOzVd
ALOrQx1HtbP6lvHit/D57+/2zwUHt/P5eQMdoTVBq/F0wiN4NjZljLOgN5MlCqkdQnXcmcnFzXIF
FPX3oqIQ11ZtrUgvnFpVYmcBRmIxVoU4cQuE/8DpegT0tTJUNejG6jKUXlE5Nb4D6p/QRMEkcbG9
xnmy5ZKqD9fr7TXM80jAm/gO64pNQYS8HHzDla/prCT6wiKZ7WlWcoU/qCkjiFL82oFNfWurG16T
grLcbV9Eb/VmYScU9P/By0u2cC/tl2kM6WTA1NcxYxKP8WNCP9TMrzB0xjRzaYxFQs/7VYvE4Klr
nRYcIakLqJMzPKjfbJWWsznK+/8E3qCsAVp148vk0D0qTCKjutF+eyoTMAuL8OyLbMA/abb96l29
mFKNEVgnLlZehyWm5ZZzpT0A2eNdWcsUozsJYJRy38HHZz0FZgv6wJ5JvpoauuLKAL4Uut5Dh8PL
V+J4Pt3NpzUEdS8rRrcqUFGED8o9v86Fgp14/e+4d6HUme4FP8qOAYMeTP/79Hb5rL1a1fRQ9khN
pxqrvywujv1/nxb2zE6rLByuU806O3gt54WG2QYnwEtMwmRykxkWKU9AwUWgyOvPsGIAYA1tjnWl
+0xb4xdWnGbSheu3QyPk/+FMM/XLzc3wDRIzLu+Ixe7w+GpNHQm67o1//3AXvdUsSpIuhbp+2l7i
7w796alxmwlb5hWlHdf6+iZRgKuDZQjellFzDehPoqwkNrxz2xsMAuqLN+Dpq3+2W+pFwG8UZjTg
7RUfWDicUUZqnTXL/TEAtBR0nU2UiSiRRI3Ofu6VBvdw41Me9ai8xSY+9NuSJjS6eXq5UcPI9qrt
BTlhJiT0CS/IGyi2tO+QIvIgOiWCsp4HPNXoRhb+KCydkVQPBbLSzo+LupYntWIeYyqopdaS1Tok
Pd9qFJ1sLPGHvX7kJX8pCU0BCDWn+VrF/nDTpdGswMzJ9opqCXtioeuPhaleej48Ztil81A/CHre
64OMKWI/iW88z/ZuoxIK/Cfs+RxK40hENsUHG4FXGkLXODILKNzsFhUncOfwOO7TQSis8IW+D0ve
7pXf9yCaW1LA/aY4qmWNCrnJrH6XJp6nQBXWHZqr7UvCna/tOLO8UuBJqK4L7FPP0rF5o2Oi8Hx9
BrxuvvDrWLxgs6axwH9xKIAxZVcsaiINBU6cFnh6qSLRogxRA5j1MqC2WLj4v0Ku79Mqj7tuW6cq
T5KuuiYPY0lIMkh+SzGH3NPhBwVAOzWAz+mnTirwGrj4X07InlmHR8th5WNxgbPzakuP55fwdq33
aHAe802ecX+5LtMKHrAZI0QsZzR65YTZ6vQfx2nVHZdvUKVye5lhvzn5YqgXiGheQzrPPMTz4wt9
51trvSTu6IPO+H23ig+uWhaGFBYYK5BZ7safvF5O+xRkWzMlinBhq7W51AC7KHcwMrO+1um0RV9H
xq5A7VrDaUUf1wB0cUl/rmqiWPB39RXv5zn40Euxa920vJ8rV5VByTxDCPR4GBwq/67dDWXxfPzJ
WSt0tDQGN6ssD8BZUTOBCED8Mq3VEaljA8HFGm85Hjz/UU3Rjoan4uLvDbgfdnuz2hMTc4u97xss
R1u/v+3BJc/eefnqH2AdcK+QTQAaNGH4kaOq0+1U+HgqY+TX+5UfDLh7T9oYyXEUOPmWrauEakp8
OVAImFDL+XSJSWrSxlYNKHWoRpJC4bSbzGY5xzHdEmitgUHd1q/SxgGT/+OOMlbvEfpzdlgIjmEU
WGtKfQ0Pc5/FZkGoKnoxntRLqmgPzJzhYco32RdcG/niNg5bkVRZQuUXEf9hMX8fgKpDkUs1x4fJ
mbzJYumqERZnuBIC8cwxigIwzjaxBEafEm+OMZ0EZsiP+lqfDyPKbhlvPsb13MWQvMWi9DMU+mNS
qYZrrKmT31uy+gr70tb2QF/ZmpZIej8zmwqPSjMcKceCKvLNE/gWJ31Gl2DoDfg/N0xK0tufF8A1
2+SOvSfCgjdENFhFuvmm4IXe/t0V7en3AwW8cSHtIROyWuuOabVHRqlmi4YmDym1GGcXSgv5jPMY
madGnGYwfVkNX6CyxL56CmYYoks2SCnv49iKWrJfEYeT132KV43CqyNne3qQWcIOJuK9hl/aq1iR
9L8XG3w7gB4irRRBXCav8lDU1naJx70jDmauVP1RzlGRq88Y6CUfoactJ9lKSaEBpjGMsIH2UmXt
Pou6Mz5t//pSH4uTWcfKkyFTfOknDBvMrb1a0lsUlWboF6vVCenKer1kuKD2XDO9BiOL8zz7ynl6
KB80PApjn0r7V7DdaUzY9eCV8LUJ1b8hUwvnH+yk/n4rqhRIpM4x1Pz7akcjK3LWrRnJjoGXBMVm
cugBUiTAmBOWyefg16mitmpTUrmdCZ3BwZy2AZF4ArcykZUwTwuseFJ1it+Sw5w2gs0TI2SUSVVf
0uTsmjoheAgXQyCmvfnYT+E+5gMLCzYxAzIGHbgHqQeYv3PZ9T4EUH9Ssnhn4/6Be7oWMBnnazlp
BiyK7F3oZMl8R5pvy+r2gj2zFue+0+v8rpMliY5lGg/arjCFc9SmnAYaZk5xssfFHD/RSCdOglOB
acXsNRbkCwhX0/D78xWx5rThXlE5N7TB8yAJoKmsjrMMnLzSP8hTos8XBS5OGMfDUC/t8hnEhdF+
RaBwcHQl/lEwdGzBwQAAZkOS31Cy4Xu3jdJFVPogTt2zihmb0c2dfWKf4Tqpz4Cqzgi+H2ff57a9
+jEiwsDSxeA5DyMdtVEdI9BXY/3ROjknSXcWMajbJePCxtiw6YfJQwn5SCz8C0iGN6JshXbe4OWS
d46KMHuHLBsXuTRPKVZ1SBWt1ylU4x/yfiBSA7RwuS0zhWzI53wWlybhA06W9v6ZKqHmtjYpopOx
kjXYugreE3Lhj1AYgXcCMJMvpUr9d2MOFJbsbXYgphGBMmp4eAAPT8NXjx7wIM8I/BSY+YUqLDTA
umqAjRG7QNLprKrMgjnp/ThDVa9WDmzRhjFtAm2MdeH6KoCUdEA7kighTOKdF2M0F9o6t505RDwF
eJv8wheIlzUcmxp7TwMrXpMec2Jf1GBjv329gxlKeCJZ/5/j8KY2rpZpkiDEzjwpV7iiLVvaYYhw
Pol/l2jECHA7+3DgHToGjgpGTYL0h1nWD3kAJAjZmf6AcjHFr5bZU7JAYR/GgWD5eRy+glcf9Tij
86oQX1ZqDLlLnkM+oIho5NbxYufJBY7E/evIjyDyqez7uhNL3xmH8oYe9neyrv8y9H71ZKp6W2qK
gEY6eMxPXbGpeKDOw4F4TEJpB983LcZ74KxsMaRr5ksZ4HiUWxQ7/MEq1pgLzBIrkW4JccSrC9ef
HIbqu3UHxBt8rwG8HOMco+I0mBJGoYiXmV9v/d+X6oGS4UROGoxJ0mluSRyT8AYR72QIv8k9WVLD
eCXHKOZHA//V037piRP1Pc0BUlO6TN2E9TPEw6x6jXXy6bKgjItmNhbuN0ZTK2k44bzK2Yh8f3ij
EJg6F7pXvEYQ3CN2pLdodP1rRl2kyx9yRO1MqPZ5ayzyFLA2V07p/58q9n+MpocUHuHLGK88vd/z
3igEajAd1oGHSKsjkXKMgK4a7O9Fuyjsk1lQWkBf+zMSobCKaLjsiUqtdazXQtHLbg863sI9u+/0
aquMLEqLiP1QgKUD7DxeOaXxnOSzQPmaSTn2Y/iIAzzywk5wFxXN+mRCo+Q/8AkjS8gPr2nFrQut
fJqzkEaVhBC3c/Y2AKsTGD8+HBrw/G4QEplFJaBB0ybxzFZPs/VB0l2hAd2+u6QTejX0iHiSDRDy
ux3IMeBlIVb48GmycQhHPuESP3S3idLUL0usEflc6+d8A0jbQiuo9b5Yqtj+J08Qw9xdGNUTCe/z
R2kXTqv1KMkPaajSw4v2f97vuDAzDAo8+6RNO0yKOZcgpQrrl3PJXemE0ROlhhIscRFi+xdbUUEY
XMKy/2BP2s7wkN5iUF6vXprPveWwGF+kDZuClcxAKv0m4jWaCYbG6HCDhWrbvxntvuKL5McoJylQ
TEJ0Lvc0LWhdBzsDaDwg+r++rmegUvMu0dHTLELNq7NNztu9iy4U46mahIk0p/kP3UWduhUg9lvY
Ekt/yaj1u6M1YXS7jDvZr4Uztgn82KRWNDDNUX+E9qlFKP9N7YaZPLfhTFHzaZFhlDVQdpYxtLzm
8tNmTGM280JNwRKov4h6Kebppx+LLLLRpkLyIIVDHgLSB48w5i+RRI/q6vzs6S1DBwGxCeYdKMEW
6fDTxQtBtidOtU380bo2ZnnWe8PKJWpl6VaAZortsTbYb9nO6Jyk00xx4falBIrBDscL8lKV5nkw
w0IIxLsdz+MBACQeoIPL1VPao8m3ZhVxFX7IuijsVT4zVJAcs5wVVpmg/JHKpQa8yMJFSEvRPITj
JB7XmJTLQDPuT4h7V6QezFBwwJ38LfHaky2g5E/YdFGJgMq2+c4jh+OhQa9Xz/YnOapik/QOjlIC
YqGRkLIRn5zjvHkV88uxX1q1KvfsA+tAxtt0GFcr94gdPpXnpKiDd5raKHJ39BvwZ0DlsW5fWGc+
sK/DUVzbN56xuyC2sQIlypn6qjga5XgJ1HCoet+WiBmNYK5WwJXtJ4xFj5Psmk4CSBNe6nqqCi2K
MRlt9SZQnzrA7xu7+r1Flnah5Dsz6QPYG8xszdNBwcYokiuhncy9udnebTMWNFB00Vcrvecbah32
hCQU+bRYWDHFn71jKAkTcPNOAbXemmtYwPqKmtOiwWPesZA0ziWEdMEVsmKU1gUrzb3vBq/SzWhb
fB5g6x2iV7nzL5xXZMwVEIYXRbyVZ570XNuKMxH5LHqkKotybrMg+hqC+d/fTs+48BncoUuNl+sl
wbB9d2Lj06yOyNuVz7bd4/c/GbNkL/ziRDIaikoctkITcXvmGAdy9lUSzzCoRZepCkQsh1GZpvwi
wY0m1ZmPztm5okPMnm7mmhIXxrZ2+H4V01nt+DoFTXBIN5Y5JZwBXbdq3/Tt+F4LM/NfOsNB9gTt
/MBExa72zZhTfaczboX57U9P6Anza7S67sfQTKR42cScJ3ejVRJMg3kRS53g+UwZqzcRLzEcEZ2M
DUW5oZ640wt+NG5M+tqBmWNrTqFTO9sarqdkeEpQOt8CkXcb95dyT6kr4y1/MxqxmZRTidVMBJ0m
dZGNXikVto0FULKLyxtbRPlSQw8ee9VslF8cjRhjy/JCoGuVy8T5djlXayT++z0dFTvNDDdP6cAp
cMJ2eugEtRRBqRfuNl4vjjFSZKjg67PB35pAfiD/Fz6+Qy4vYI8UHGHGJ0ShVThmiYjehttjPYHo
MD8Xg2ypob6g+2eASPN9ureUX9QmDdCl3woc+3EHSp5AzfIQnHp/WKKZNhEHaZSdZxpVMjhlbKat
9soleJd78EpwZC8R+K8+jkx9Qb0Q/YjGicYpS4Bt4DztYhGDOdLqvnimAWTkrCRD6r0zp+/06nDr
42P82vLZZsJ8fpI7mllj1Bmso0TzjVBiCvyqreRNsOXLzKLr1mC31QvqdB2bGI/aZc8cVGKKz3Pe
hzYI9hyMC0zE+S7WBDY+B0YhlY3wja9GBvrGu4m8gL00ez+XP7HQCP58kMckMUoO839XL8h6P7vG
+/vKYjy/TjK4JNFl93gqdGv1qLXvK0LX6eQwb/FxT3tiB6qQcPWaAZ4LOj7dJtFA8UXYGSljtpyB
RFFcoqMbzIjK9eXj5AWXpD16xHBFtjVHpt6LQOjt+j9G1anW+4y9qRZFWbGAUChLda+4AHBWcA97
A2sPpLcxKeHRyhzN2xdL/5HyHYekuYT+MHxGObTTHvEH3Yoky3N+2vSwAdnU3D7kZYHI9SjmajRQ
5R7jPedQVguHy80jLpMkX4Z7ggtGPw+Mo8NNFCgVZedHqcVW+eEex0Gxe46Gi2GxIIBJdeMVAjAX
Pa6gD1hrNw5QTdNBbTMlFtBdu/m5vHG4owxyEhO20bJNJ1B27MxPOtsWTIw0x8ggvZpdF0M1yKE0
GvGmdpYjAjf2jNbT2snKpt1cBjlFeXphlgnt61jtzk2YW053qtQTwgS2l1zgidEJ8L/8RWFaHvVu
23dpC391bC93LZ9D5z9HHZgGN0IwH3WPncZouaXBV0lNUSgj+JV09QhydjqxHymVxv1/GNPJgrB4
dvZwA1mbz3WV00bFSdg+G3KleIDeopj0EbERXYPdLvge2wWLUiMAn/cNXZLx5rpIpWIjIlz3Tp1h
zAV5/kdhkG93r7j11/1SMqVztdbXtUvD2E+T7EWpXuktps5Dgrkfla8qgN+6404XyD9mqLS4127u
zuYDkXiDNR591VZxPYMolLMjN9dgPAqJGqv+m3gNXOAjt/RYFp0FnVkABnXP3/xhCo5kWlS9IX87
8JzDvRZ0cMxBh40ydVth5vDWqjNDBsilMaOQW/N2A177MzMkhrGXjeOnoTJ8aKD71dGwDUzqTAiF
tcbJzc8IkGqM1XnLrdAJCrHpYHLeTx1Mc3i8ow7SZS1rJwitD4TjEcszE4BvEBH1ILaj8rlrfpgZ
D2EAJqJq9AosMBC5E05XnT0Bk+4NyUVbrdL2rPtNTC17AU172MXtZJR/gRn533vyWTuZbI/JWc0a
twmHMU0gW3sbTaHNCI518c4Cb4cGEZ5A6fhAs3et15exvID1+jadsKBQirUKgIeuslrJjtSYXDxu
6M8dvQYwZgHpev4K/2VWctQNbekqfiwdVPXt8J9lbizGzkTjWdWuqszyBwUGr9Wow6LHv49/wzEw
jG+vAHSjAif/e9xTjj979aB2FS1+24GvAXUueuNOLOFyd6d+5VCRmFZd50tBplsa3FFdWg1NVJes
tsMX+ZFrs2XxZM1mIYRqLiFwcZ8Xrr+MdfMCKuZnzaFSr9hUx+4srs9cA34J1UR1Cz1waTOChpEb
l1D3SwV9cV2g4ie9UOS7S1KgL4v3i2rDYzpk85isr4ts00GCM51u62JEjEVpgFWvz5/1YndK0tcj
wv2EJbYSvP974PLnhTZzfhAhvH0iQ3IBbwEqtlw27a/1uTOYl0owPdOxzZzh8zmNEBYrqP2kfpDi
NVYLNEheCpJRnMzBYXWQdLqll/8hUb/uZG9VNPab34gU/s3M2MqaxNEiNxx80MrDYu/rCHemWkTq
H6vafYsshWYGU6j8WyiiYzBmvdFe0AIlbOwaIbaaBxQC+a6IGstb4tybJRSNU+lidgnbbpOof6Jw
rCOxgB+Mii4gzrNUxVYKLr/fqEZF+W8LnQcXaVDekkzMGBRUbPhjAkVRSuF1bvvMGp1o/G0F2nlU
O9ImNHyPh5QWk2H0mNVZJQ0UVw1ALS54S1EplQf/+13GUVPpBk5s5+daPZhbPXjgYhhjO3lY+pJ0
ayVKrDhMGV84zLjG+FN/ggST6AmHUX34IUJJOuZiOkd9MK+ryHjo+cbO7TzQSD2yjNE9rP0E2ZcS
6K69SmR/ASmCNcOrfd4JGAaOe4Dzl9WfpiOOWBqo45UDsiCao0tM/Mq61AzPvQY2M1Ny7G3/qCuw
VTFnrEMLLWzCIHPAoZ8Qznoy0xOUyXqYX3FHT44ses94jNCI9z2fYxT3wDVg3uw6W4Gr+Gin57hf
8ecwypnZ9bzcAs3GS2Tt9XjnZvFhmpcNfDUFjIG2zw3bPOIUvv2HQLuBL6qKZeqN5DFGTMIs7cry
RJ4Pp5P3M1Kp6EbNWzFdP4+MyKxzVeiQX2Rp10R13rj37DSXfZtqfggidbWcHotYRWH37wSxUTyQ
WRkM5Uyty/KuqcsWR4tuJ8JGZxVoIWXFtkvf/Nir2GgWeDxnHAH4PpTnYLnkOhMLZqd00+QH/2fG
NSI0NBFGButD7Adae634MaaxcqV+42oZxKyBKgl/6vUtR3rWnBefO3ft7jlmnWbRjiXi18jube0c
qQ9WBEzH5uKiidyWnujS8dUPLF+zICxn93UmzM+mqrNKZVW8unvBlsQihzgCDhfG5cBRHSaNBPLh
u3vS4nZuBZz+Gsnlqjhof/sBw5Qqew+9FVBqyxQivWnZdSN97CfzAp5VuBYJsuQyX+doYBTX4qhy
4IZc7cktEdkB/Uy/CKEivPFx09mroTQ2NXw4GrsDMF1L23+j9Mmn02b8VU297BLAAgdV/k+SlU66
kQjJOikqo0fi6s7dnsqp0PjG/bPa+aXE+guIlVGFPVhCnkj9FE0dweXPkhoyaM8jzydMleDfd5pL
uAdp/bNEP3d3+aNcE1SBftYhBF9X2gG7BOQpoUi0aKWorMLRy7nDQPhDuwWvCZCmw3YhoqA8hPxR
loXA4dRPAxzfcBT57cV6zJCkwzxbldFPYpOOssEW3IPWuoCLZM5HU6InOZs+Gc36JliT7Wu31b+Q
TQo7jhPWX17jqnLoDjxA3SLxEHuG5bd4L4hDlGAe9heb0mPKasqlLvdk4hhf49o7c1n+4Q/BB/Uk
7plrH/fpwqwodLu67ruVbiotASeikruXGDHdL7sG5VLn0kqN0sza5ZkhGMPI+bCoH9/ysiApo0T+
RO0JPSDJRmLJN2jU0NhR8wi/2uG+EPv5XX65Jv+nmQeNG1d/mVbS5JnIhhkca7ACO4wBlsiZ8dP0
3Mxu2aoITVuG3wutLdCyI6yqx0faS9z/buQb38wejaIlVyaPdnFcOAUW3cvoi+NPKmonavaIHL3c
uZLcCSqc5uvmvZB6epQPCWd4UgLRhuIIgWDMBmrrtlTlbJ/hGsQwecCQcTwW/7Igneje8pNlYIiE
jmCQ2TJdCZpVBhdBkO4lHzEjDmMEafxFYapJqLxjH1Hmiy2kLZfeBC/m64pQnV0wgODqAqxvqNmy
FV/WadVLjLCj+vOJwfJjRC2NLGTpjPfaKxrVQcTnF+nyAknMmqTKlUqL75iduXFy+Baud0o8ol9Y
PIduv384Zza9oJXVgbrziLAxcd/4QtZWQDK5VxYXiuRPvMJgIUP96ihPavCF++8fr+CVN2ZLuSCU
rSWNARrkaHlySjIxWY2KaxLqb+LW6uBXsTnseX1AwpQz6pqzSVE8XXAt2BSdev3qPtnFDMqg5UAt
3/lKcIeUkQAzygvJgK/6qSMSxlelvkALdKUo+EfCt51h8Txl8sd6/EaX0HzUMtJYKshj4adOyPSg
+z0n5YxaLUF/RAfCGoYT5s3APYP1qU4jN9wEYvgkGV2ZSSNO0r1YD6VK8u48GxNQmM/PTV7Yfl9N
V+NMvnf79vzO/blKfhsZFATjf/gwo0VKAnVlevQjMzdDnRZJEJc5mlRGfVA5RgC8Jbz793IOiAAT
yiY5ppAFMQ85UhsVZB0nk9qQDQ/Scf9VH7cZB869z8D0st1t5jOmM1T79Lqla7nzvHCGfhI0o4Sd
jBtJw22NFIU+XHL+0yySU1EM+hTVA+pVg2Tgp6OycX+GoJrd480+c2AsdBjxT7ty1WjfmuEX26yU
UIwSadUgKAU6t3mXIFWLmuTcDlDuKrI/+9z+d+x04ndY7ud5Yqmmz6TDOfvFrjausMKUdtOvyOS+
rnrCjnoI+d9fvQd14gZEZ7Ii8g/CVugmwFB79cJjUw9g8vqJOrPdGHj+k+QGOKsHm22CUaNg5VyN
G6ONpJX4Q49/EuBe4Tu45hx2l64sVyVAQ9ypqq/NI+yLp5a1OrSseHPXvq3t8UYpDvJajNZxFBhV
ERGeVU3ZvchggZWtmcS/QaB1K4oEg6g8v1nsg2xrplQQeRu6oAaOWeZpuVd9ThZ+FlsuxamZSqeu
KedApykCiKnhDUabxbcyi/7gI1datdwcyMAnlRwffyuBco8T6IMwt5QL3Sxf6IZEkHXdW3kpNz2X
FnL+ssc/oam2kt5LHOxAIjD1a5+yfoCya/j5WnFBMq8NvJHOLcmEgXHlMLz90VctdYuHf+E1tbBg
92fqA5ofDP2HdNETonNDD4RvDViGd41jRwWt7sceE5cRDAglHelxdNo8pB0FCBw4jrywEO96A2uI
WFqRqIMfTiFPiseq4UGcStcq/7uamrg7vtcKuVi74Hh+WSugsZuoXUNKqdaC5L1uykmWeuXStLcu
DAvSNgcjmLguOnFTFT1UDCzzLnu5jg6GoX+qcRfxbM28mcSBC5AQBAKqpyc+4WiPXgV7tQ2ATY2M
wRgQ8LQ5Og1dJUDXNtk8xJSiyDxjG2XqbdvrxSzrfRcqA85kROnqKejHxCwm4M0qy8zgkbVYFysO
l5AdFCYnsiMGIYlI1KzWqSauMTG2Yorwn7o2T+csuneQdRVK1P21llqszoWeLIVTZvkc0V+nxS5B
mharV0dN3m/lDyAgQzBT1UBb1ZH5jxEt2GdfjLR0IWOTw3NI0idxtl6rVTDjesn1Hr2hTlKEgEmQ
mZ2uy8cAFM9WKZUFE3Ft2nwccjTeQvKuXqrPX2PalhamK3g9rLLhJVd9C6Jc/ikplgoohbgTZQob
O+DQ49aflgSdP96eCS+ij/4fr8JPMQtu01AnvxC0WFM1ruwgPfAv2oCWXz6e7/TscoV2YVlFAKDM
Jxnt9srn4BPfl1qIOtyY1lGtbifUCZmLErH+YLscD6+p65itSkbD4KJYoJmQ+m1Z08lEbOgrlJeC
bSoqwtE1vUpb1JAheL08SbzqLhjbXu3bzt3mmgZjqVHzeBjyKr43XR4W9azlcqVESK3ILHCkaQWE
mzj+T4ongAi54nwK2pz7bNy8JuM3u9UxYP4WBNtJmVCzA12JijtqUOizv+MvSJeSiz2aXtw/ybi8
xE2P1P65N3sjvEFgwxjnYd6E43ZT5FuP2hB3a2Z6bCWGNzhogxIMb4O1tFlhyEt2fcts/qOX1Cgw
+WQ4HwppZ2LlRPLNC0lnZ5iGJTdApjP2FsTY3Pe86KQrppQ6ubYYPt5TpGLz43kPFPk964L09j45
I+UtwxnSNTbomN/PJrKeT1dFNmj7QCdE+emelydSWoTeUcXomo4U5Q9z+Y1ti94iqM+FwN7bcV0W
+2aLtRRIn37yHoE9ZMA7WLztVnK5A9vniDeRKKJRtoRsE6V+R2m4AVANbLnGAuS/nt+TNMl4r6bD
8BG6JYCF/cZNpYPvOs4I1IK/u6joqDH+x4PMXU4s+nSZk1pEZSKmJDV81PyzNP0lC2IiMUTfiABK
uLnEmtKbzFELclyW0JV5i0+ZMGaqtFh4bI3ctGPMUD9c+rFFxLTcyPHRbj3BC756s1SCSAcWA20t
Fv6UVLoUTCy3Xe5OoY2LIP2FJ8lXo4JEat7zFh5q3tVFpuaMBh44tAV7LB6QQtAbPXoajs/2MKqY
iCUDEmn+akBYjUnShG606FHIj2vcgX1cGlsgYNdBLB0sFe9cnGJ/aTEb/jE9TZBrlWc3EM5sJhF9
B5Q8OHdXDqGR7NKbTGOagqVSgqPLF4owQRSQYVQf7ICuxPtlKn7teEa8VjqN54W1YhU8Rs5twkoq
tPXev0LTyuTD6nJFjsb9oa+aiuVgdHDCQRmfvHIHkK/d67inWPm1Tg8nqCe34im7orsxZ912lwNr
cOh8UvoByUpe6CStE6oW8vHwZ22Ff9mUWXfu9guZovlXQ/03luOuGbJk1Hobutgwm2QTILfgBMp6
lYDDZdt0JuupUpkO7LjXA+MTt/4zzalOZWGsRX1A1wqDC0DQ9tHK5YEnEy09n808hxh/7dACsqGn
ybZY+nkaC74bQZ92oXPYmZvPnLqmD8Kda3RygMeZqpzR8DwZv2+GscbykWZEBtpYW08zfiYlY0gH
cd0PzA/3mSOTlvXZKnpgV05MO9WV7U+EqPDlsUE8/FGc+gctIxsMa3guBNhR0pfmyLUFbMysFZnS
nxum13fFsZl2Guy1o06fWPOEIu2Y3UKSGEEy6ooI8NI6zvQvO6xH0uaorE5nl5mFVvN92snuLmMa
9GAp94Fil/tBiguTx5QGKz0S46LnkhrJUIbEHfU+gHKsdc1eh8kFAFLRf0KzPuDDnTpFcWcZjlCF
1D+RhX/91stsm+HpH6NIaU3HkEX8iGww1SVNHzA+3iVh9fXaduGGn/Jrx2B0b06HrMuV4V+/o54V
7Ph0O1/um+clo03UyhV3xu3DFxTrXU9v2iV2Wjl1NVT79w/k3ltw6iq4C2HdOPbul5GBQw1MlsJA
zd1dErk/d5a5PTkS+x8JWP+KnqaKY2TidEnO0lQ+rfLeFMkvOvY9i6Ej4+Si3mYnwx8Qm5VdndDM
abFKRpPjysMQQilWVEptVjNpgadAXrxgkhDBcqjUbIgqco8+pF6agvCdHT6Ica9l+zn65NDXf0O2
3spWFZqqmt97D1/3oI5bSY1Atcd5pE4qaTvViaXtTs55TwjkNt0LwrXlKnIYEgXcAbHCQoyoHwzJ
S24bewocm7xWqC3NqdNHFkSIWJFU8sFDw+pDbq8IDX0J+6jfnBnYG/jyYMpbxmbaMHD6yI39K2mf
iVI/LwUGUx1IZuim8fDgFla1NqdfV16bNdwJOL60SDdp26QPcLypZLXBEHBMBh3MU6JlUZqYj2aE
D4rHqDdd7FYhS2uufEWz5s0oRFpzXHHZL+C+dqyzHmPERxG6xOq7d55cHck45N28TZnbovqK5nv/
JrmR6y/iO4iwJGsBqe93CVV/vFaruhVckmQ10tP9nsRhqUDu2xbY5M6LSszM+X7Sn6USIVEDkyki
jx1IaA9wr7/aYdqXctafxgwHEGA8e+fI/mMYtne7TAUMn7XOHQE+wB5kEyLykOgntcHY59Z7Slng
29+53xw4hHtA2bX80LSoVvPinM+UTdHsHnPscN9mkYsaTGucLfCBoMQoGfCD7V6neES/IDk934Ky
IGthdhij+Nsi1KOyrO/wxlJ/l9pLWemf9dDWpYz1O6i614LwaW+aYLUVFdjZZZmFGtujJW3LgH+W
v7gPn3vY3EMij903T3Ph2PPrAjdtIEoBJq5cZtCu6Rv1fIbN0ZbUnpjD3JINyBG41cFdR/pugXEN
N/oS1zURqGrXMXizV+PWtzTs2UVF8BIpDu/BSc+xfCE85QLj4zgDECuqmCd/IJK1KiPYqVFSqZ72
6+Jq7hFy4aqmQPi7RARrUhMT9MT4eL5lDTq54qtE6w8df3SY8mNnn+XPJ20y7P5AF9RV1q6rA5BG
YNvoXF/u/nGB5MWKmaamSJJ5F+7g2AT260/ATahTfBZvjyzUMkBMIB0EUVqUjIvRvaKfDkmylj1U
AZ6CwlrQYXn1ZVsdkw2wtzHQhaA3frWIuP85zQ+DTwZRVRKJxNFKSFY2ZnMLPT2NpoeKaNGnJbxa
rgWkeCn8alN58eu6OgDl7HbhgP3IfSBsVV2xz0Akx/etvFrenjFfzFpMKjRVk1RAv9tB2/n4mukH
uCR/faAgfevWkS9ES7sAU4EZxF1ORrJmg+9crvZe84odyY1q/QtvTOHga6ge1Rt5tE5dzDTCMhND
tc+9wvsXrlsqZIhdf+1ohLVmtZujjkgLP9TYS4m9b7Njo4lcKIznoUa0KoclVdMR8GjeJCzBPcW9
Qd65HU4wMeIgiT87eVb2cxayXsgHtU5W0k/c5ziQmF51PmIt7MBVC6Ts3nVt9w6/9Qk8mLjx1tP3
cirkbRBfwC1hBS1vnIvylbs3IMob/BPvprb+3i1jgZGdFDbvThAHADiVS8lSU5bT0xcOo7j4To0Z
U0Sz4BB/M81EXwSTwyqbnP4K6qA97JALhTOamdfNpRw+BoyxilaWxGdp5JS2fxnDIxPDJ7BMwhrv
SQFwmrrzldV+pr/tor3R8tPIz0iBwN0Ihy+92WbcPEmkCoVekGaV+7B2QPzheGp9GgG0oRdej2dD
7riLg5bO/I6tnN1MvauUzekRn+8fh0MFaVtrEJ73g81WhNXYd4+x/CbnuhynWyZLhYf7zLx//15a
pzzya4W101vSGC+mdQrHpkvCdVa30v+52Eo29VL6s8QCtKNmKcVFTWFWqGTPM8lWhTlkQC+3LBu9
BFRs9e+naTfaqNub8/arVW0EkFhHimwYdVsY1+IWWbcsj2sLBvAWRs4CcF9GMeeB2xs85KBYdLeJ
WzJiwX4st9DIjx/2MnlurFC55PDj1YE2sHXqCXPSWUAXFQWNLYJGuMmgsFX5phiwLC1RUEFu+s/g
MUlycY0WtnuqVjVK+cX1+9bUNYWBd15YQahGIy8QdGWRplfVXZ8bxGOi45y10gBaO5vBixkdfXSf
D7upMwB8Uol3u1oiTQmV421uKk/sUr0rJenJdegmbJX2iSGx6elDBdp6ClmSMXnuHnj3qJqcWrIS
20PUYCR3zviV+It2HhIyzexut1vR2rPG54t6+3C3c9YKbOxdGbuBJBNKDETz2yDiJpZc0t/HITfF
j82qjIW2OWFhCcFu1vBGxKFpO4dLDCLLW3/WDtrVB9dt3Z+4cRcJQWhWPLPW7krEPz2WkWbWyGRQ
eroww+yv14AvstAWjrPV82M0opitsdcQs6fGrHrruok0t/QoZofJEHInepiFBIcGLPDO1upn5l4j
lLnmjqz4m7cx5wArQuXsXWUEEXiTEIgU/4ulM+URFWg4vG1uCSrIz7BpA7LzjhdyowsepafKnH4E
eH9OhFo+yMLCol/ejLlYdBi1g46uki02VJ+QcU9V2I/lSuOxzNqEzwA0VtOb8mQXu+uUZ7T9ZBwt
AFTZqPAvM0+3KxhAUThawPtxUc4kcCkNlDgWp+sfU+96FYd0McH4wQfvtKsx7ObslLNCSWFr7Xn/
jOg/AUNfzGetorzdfU2/jCrvsg1VYZgvnsa001lYawQhWgZZ3d11O/YioMwLubGXglj6kD0Jord5
O6zFHO+Ml2LljKwNrl98D0rINXXoRIjhX7SbT8jmY/KYtG0UJELmEASVj7La4IJzDhxpqOj6imfO
uJE6VaPsRkmatroDOxedQD3pIAhhak3O4i8i5eB9wAXMWE3p825FfvA+v/40hIMxusw/l3Sxv2aD
RL5B/hSk6AfnkYRNKkt7IvVqbStLfx0Bxnqdv8f1Zg2D7gm/9tj+cf8X2lB8/yLswrIYvd27SdoO
F4ZTPfjdNwlEWvyAGZtktp/o3S+rK8UuVc4AzuH4/AS0gKHQ4tBhMnADs5j4Zto8ruv/smbJ8q7B
1MmLjioYSYcWZAmgO19VaiAEkaukPidBG7cgFr7d7JConqysZbSh/hKeDHJ8pqL+A+BK+65Z7PY0
+93+Jt3dwkEjmUixQlTRizcR0030e3X70wBbmMcoztsPZllW+cO18qOnia3OrYOqKWE/VjjtCnZb
/0Iz4ANbSVw2RgeFFUpiRnv0r/38Lh6dPNejeg7V+r5mLvy0WMChU3o2l3fI9KJthE+n0EtSptTb
hA+N57MK8E5ogCngWcEo6LVGvEDjafTthFXjpRvUyfw5V8jVT9bW7E90WwxuprDAN5R4BjgK1mo1
wPm1XaYFavhNDoj1axBFo0nI3dknDA2crS9kfcx3t8pLLbhgWHMmTV1fhWeOg62HL45msitQ2wot
eY1akFXq3WgbA+12ZOhXu6u2W1eTFY7KzFMdv0ZrgGBIm4pVPrzxYWbrWzcP5/T0iU1PhZw4nS9K
OElKptVzY75xzgNeoL5knrsdaCt+YqbsH97FxmGT3TGrOe5415KSS2MXZgMN61J3L5BjMNBe05b8
JZnyM0gz2mtPAYNYQjebX0n24ATgFbGnQbCDuSqmmF+TZqmb7+HH/YE0+kf9XEOZ/4Bf8oGAeWTH
xbr5GuB7iaw7e1pCXT0F0hJ31DEN8B7Jkk1QdfN9Lui4BMI+ooqB6etZPqbVe+Uuana+/9iPp4v/
nZss2HNtRD+RT9kkIMsmVl29UYlo7CAuhQRhOrzSyxr0I7Ymr4groavdF074nwWiw0ZcTNn1bME4
jwaQHXGPaSEuDhp7URr8zMaonarkl05ocuBPK7TC9XecNVVtUF3Us8xYCIwUJSU+cYW3pwvST2AF
uqfa3UwHWSqybFBzQD3M3jU9kqHpGfIX6TbyGYoK74lS9eIWCCMAVi9xPL7VWVTdp5qBMVLCW/uA
kQA//Sut2nRv5acdm0rKsKrdHrV6MutArvVzxGSGsMov23IMigWUkBv68iOGBi4KUmZUk9sjzJRG
YYnwhPbdjokAgUNLLW4mbOOl+lbD7yjNI6ymy1Kl61lXCqsxkBL4Lh8hgpE+vZxQFhRzkFJjmOt7
5q4dxxGjmweimXCm2bdOlgxnsAKnPSdxXUWfPd4sIMXK0c2VrljitSkuov2UOIXIKfGuOCuI4JpH
hUmznrPpa8afBCmZr7SXrT9j2bsjF3AMRGLU1vHBDo3nov0GgrxWQ8EQQYoM0hp3vU1eFBqjIwIL
jmcLzVumfg8bq+5UVB7cervb15iytnYWXo7T/Wa/RjG6EY5M4iewANMczlOgUahd7ikD5P1m6epI
b+X6mjd9A7T91iN3pUxoOxHNXXG+d9Ge2gJc9FjPN5G7cNv4kDqhoEPer/ngOm0qCgiZlPlOvf6E
NRwD2e2EKQeHaLMdo4QmBoTEXXYSyIcYHqzng5n97Rg9Dt0yDYKp28RQB3h86czYNYS7Nfy/H6YJ
KcbF6dPhL8mAuZQpS4PV2xTy8zB/F5He8F9G4Kew+eqVts/ez+KXI02LlrrHOOKGAra8wVDw2c+z
lKQlWEu8z0VXgn3VtHvLHL0RNLhK64g+IrShMbAZ6u3aPFLEsrRHNy/xCovucINi76e1PlbcVd87
6YY0VsqgkYpnG+hB8cn0aBd7Q9zNs7+PlGCN7ksJdEeaEVXQPDKx5Qexxr8IAfb7yg07dBufF4jl
NLJLw5payY2+TOvOJvgZHtjfAA4akn4IiS1Fv/4WIjNQp1GrTzT4NY/Or1kp+f/CqGT+D7l8ERKZ
SaTumFf+2jCNr1w8cLo2tyMtQTX0+lwAAZ5VIdPnfW3FfDzI9elzIQT64Wal1kZihlXWzO1+9WBx
bjZfUqOG/cAWxKw+Bw1SmMA4DZI8BCPn8Etn3B3WkSccRYRegDMRPPrOdzB8Cu1O+8ZqowGUVkGJ
INOfoEtTFM/RK7ylyn+pJNJVfHXDQ0Lj/CN+BfNWxb0zsitHFf3YH/wJ+Cf72kXVqhirrD1Z0hWf
Z7yaLTHwKshpBnlHZIckkmQ3rFJNx/bXocWo8tBmBYWuXzd1Os8gDZOTyqE4GVQNTy3/F2Ve2laY
dyeRKPrdp9tt+8Fy/tbWRktVsL9XDhvVzje5qQY1THgE4Z8WOTfhSWsh9qQtJBeKcKXxfC2NYzlh
XjQerRNf3BAaEnHvCkkLf2ICjjDnEs1NNCl2R7KwFR5Gwcj2JaYq5q0Ty47TBY3aCbrD+BRpBaaT
Js6m1ylmuWpUlhpLmFKH4Qz3tr163mVMi/kIkffgQb49BFTHHgFVipcUrBtAWJF9frmgB2Rl/WMz
IM15aoScdHEQNihe3aMnWvLfA6M6rLwhO/9QDCxl+GzwoKgNSFPatft7SSAiM57PDGA2tKH+1r8U
SYmSVNtNV9lDevc7EOvLgoevK/KhKZ+JeKml3vxDvkn+pE8pF/Fj58FWEAN7NflGGZdi5goW1XZT
iZIASMHuPEsJfTPKVDO9IbBgIJjmF4bWFg//gckHN496I+pYnn+2kuwYoHySeKod3L1maTHb8h4a
ou4jHzDRhnSIkLZO/MUFaAAKg6cM8hRa3pzpIAcGWu9qe0m2sAvxip/Kpx2Gz9hDESKpOiPdRD0j
5zswu1wYY28Di0XvNyDbCl78nZQiLGpvBhd924Jhy6WUPK8cEKiXlj0PIGCfHR8etdq3rIRBTPhg
J4PyyZvnDIwuZq2SHxSlCiTj8VEdqU7aU0IeOXIOaGrvoCle9XOWx4hWG4sAAvsydOBYqBp5zMQs
KUgLdYqTkjdnUb+NMRUd8Cm/uDjkInjDplW1Q+Qxpz83js5QBOodNpGoDKBO+GAfFzkATNRKHEYP
6SimsnYIfUwd03miSDm0KiA5M2WIrVhWtC2EphhI/AXI3ObzEfxoMNdyZurhlRHHQkWPUxy95F86
sVm4X3iWm36lLNPRSAMo+ZJ+M8HU15005T4YHMfEYcfOqHUhQmPy2qGrG60eFUxd4J/LENcKq0N/
+EdwsQQq0KPMG3kRQYw7AGYk7odUY5j4WKnxH0E5pdacV6tkXzhtf07FESp2+CPu9nH1VpU5pWYR
253mTclZ4/PWnR44ibMF9CmLHcgv8jveGFqZbSmCyiug0ZDr5pEymhDQXFZrZAOWdCVmQfQqH+Gf
uyAV0JXzf10GQFJzSaMUxlKmVYqZ3VgWIddqg3scAZ70lnBz33MiP7qMZM2aW8StusgtiU6hfmMf
Q/KVfbrqMkvGaSvc6O77p852aj9XD+Ysg9QfTkmoyjJgzmsNtrv5YHNNXimFSI4iF2e6z0HG19g5
QTcsSjsijnfIVb5UV71ras2/Q2PycW+79xT4gyQSOMJDLDtLUAzxfeOr7uOKC4cn//G7Pfm+tMju
W7SY8mri+nXplRY0l51yFfW06sWe88FQy7sQx4eY13xQ3O9/sZakBpfJpKyC7EXPu1i92QzL/HdT
7AF3f1pOMZpFlCiM0/JO+xbrOzR54N//czeXAOtwSGq+EvS6Xd8LzpvusKe/dzUoxo7lt4YMeMSy
l3DGvSnP+FS4vRvzTflBvxV9vKuLp6ciRlV/nj5JM6Oi+oHEnUZGaNUNhOFR1iFGCMc7ZEDoPAYP
GUxrz8zChpmFYEDPYwgMhqK5wVbjGvOXMu/O3edr4oEHHzAJD97s+Sp9vuWMukdChaErzGtIXSVq
7jdxsJEouHUEd1YJ4qn3v6L28NntTeRArqMkhJKVLip/m60yQ4VcsdD1ug4DczpS1IRd6Sa57nV0
GPhRdQTzCTH62psvPOakB8Fnl0urWgaRDyWTRthmURTsKZ4SNFUkvXS2Fb2g6utrwhIW9pmkZvO3
rCfAKW44K8H22yyD9d+aemhGSwkc5PMdug3rt9NtvwU//CoFfex21XOBRLgcptxm1WAdnef5l7ES
JQVzB3IAid3hhOnhqaBsJ5p0Y8Psvj7yrLs2V/sjzfDuU1hDZ+6OWY1OQ3LPWa5izD3Nt5KR1LB/
v7Z46L9whr7lD5J3PbW36qr69x5K8BAiY5spCR28TZ9I8rfu5LuBT5bSTQq+dVCVBRZuwuGcEn4b
5mSHw1j4Ers8YRnr/KdeJJJDoBOSDnRdKINGIk4RbayFfM5sU/qMUVAKEvyWSjpAKTWWq71TRq56
7kHBLkNW30yZUDv8W5B5yZt64uf55/1MG3sS4sd/e0lUSZ8x/vZTOudGikgAQ72FIz9QQd2Vk1WS
uNM9AasyBjCofqgt5iBA7LubwgGF4KF/UoMcEnvVaTlOYzbq6OSX1p1CkhnyyePhqjbv4vHcf+vQ
+wlz6yf3UucZ0SUGYKsr9brFH7Xo5xSFwt88pPvjMiPjY6QXEIrXbJY0wZJtxLTrY3vwddATMzgZ
8Z0jqrhskQd64mnd7kPIhoVs1WAGTO+LhjX01YZmRXwQtIn+kywS4KXjac/YuMe33aF2dso+ZhrH
gxWlHYMcISXCNHO0UyRrNbRdMhjHtfLWYH4O6w5OQEOjD29YnL5DR3Ocy9weFxUfkGGI2WGRC6VI
/ymsYAE6zfxhmCz0jo/dGt9GWI066CjiamXrkF/8Y72X8g0zdf2gn+vL/F4HoOpghT7n4bdkbL1Q
nHYyDYPRhVARvTmukDOU3+HXKusghMiSirY9ijB4yRJte2VXaACdQxkMr/nKC3ctYdwfGTHPSdo9
GzTPH701SinEzi72B0kk5l5KzI80rm8vgaigic+DwNpGz8HRCJnKmD1B0fWLFwASPfRQaabKBGjR
mzvghnIpLwyBcP7kbinZz0ehlDEnZQIpeEKVxSEFpwre03RcpsQno01M0YvzRactROGxQvp0q1sz
UXP2/APhy6xT6HA78pAHTGmilofFXm0AyRkLO9I/J2OnkYr5xS/88QKoCW4m1OKOSMIEp0YiqSww
JYgHyivW6FhGueDWi5XXLeTERBiayad1eL1pf6XlsYEQ8kuEMoIwgCFgPH0P9tIjlneaEGjmFAJ/
M1/MtSl3qXciKb466CqZCjJsl70hTHmRTFmlXn+jviu+SQzNWaI1dJoZqcYRG15xSkhiX8t6OhIk
xvU7N7FzdpP1bw7sWW8uHKvce8+xrhjFLmUBKa8Bn6B0AN5F4ubLfuxPeWg/UqtKu48EDEATMJ3m
l7X68h3WghRu90+lVkitiYiGXyuTeppsitX5hzDNAMYFVqquGKz6D7XIkW1eKsH5UmXQXmPZWCDq
01j6qP1A8/WnNGQtQ+I9E2vSDPIkjtZfI+y9po6s71piSpNmIDqSaWPqgxO+Ky/orpnKtZXHPmI8
iLcz2Hnq57Veh2WLYDUQs3LWZGcvGcXnvO3mWA0x6RlvOzdn7upVpQeKnDtIOThF+FeBqqdpI7VZ
aRU9Vk9TeXGUdT5wprCnQ5F7aPBx5bp9/Y+re/l96y+bncvTXqIRNH0q3elEp0fwl8uRbrhP8PP0
zXHuULjt18SlbatUyOdhNFeky7FUQj1047uAGvhJUgr6r9hkTau0I4YQCwgsCnJXBB9gMYCpcm09
0A1l7lriRM//IfGEIKqk5Ev+dphAacjQf1yTzt4oPxa+U1cHVBNIfgeak62xXRH6p1gznNfYWcjw
DMQBD+RD+KVzR/iEpIhko3TZueLLgrrWqKnEA4HsPeJkfdc7naTmVdSfzcHLb4998e+r1+F2p32l
TlMeGEU1EKAf5U37Y3TUwQUmjf165zRQHDN7k6hBESAi/3cOvgBlg61bHhmosXbq10Mk21eSpjTh
92GtBNv3iDLEpyc/WeHFpnetg1ndbTxHIoaH7k23Ulp5MaP2oF5EnewH/EWqoNEau9w5mCa9rsUG
e8PPecucMFNva7iEwFUf0MrMvXXYgSrx1EPR1GKDtdlASqNJ96vK0HrtDy+0DL7rUypQuHH/y6zs
5QFzYJNdad57q3jC10drH9GMIpDyFCvZ8OeMU/Dhs309DStOi8b2CreJ5/sI+3ii/MLWjzbkYCBX
0F3OdGHzV/ui1OX+/pakAbHEr2683TFCqSGYSCfIeq6KsWrK/67BIog6mDKYU/d/80mwEDBDoxwj
jlA9Qp2L/ZaSBPe+mXkT9y0qr++IR/9vUnAGZd1p44FcOA6KMfj/ohUI+rSKYwn/j3N/m3g5i2CL
WIf/rSaZGMHB/Js7isEmlgwrphGtK4GS3KCiKTwMv4+HWU2ZGKq5EkOMqbaydmcSqJyDJtmYBV03
uJsZ3iezWM+jKtA4VdinqQRgZx8w9uNtNBWL6O6lfTNCtFgvHIxE5GIUjhKS72+rkxMieXGT1oxd
VkmE9UiOPcat4t1NGq+ffnO8afN6iegarbAtPWyqnVK1V7fjdACpEPu2TCAfadPXgWbmHkkVr1tn
hkoU/qnoTrNke3d8mCO1gJgOG69Ixoe3LH+qYrrwweEpx+dVrl05g4qjCjUYtuzxkfwWUeZerZmd
Bl8fM3mGSm+J0l/RH72XOxWJSWyxAP0lzSyskR8WZ01MB34tvxMQhLx/i8LVVAAY4VAx6ARb/sE3
+YDTyYhynx6eNiJM6EXgFz/4hxpAuyJuKWLwj55SQbgNDjUE2ASFAgW2e5IAWysvxg2ZsXwTVdIT
NPffhUTX1f0hilCdWmZHUEluc3uyEGJ2A+ZCCfEpsRGdnyW95IxdamplW5nFcmyZmdogeRH0bEj7
DiL+SCFlIPGJ+Eqs9a6fxvbU1TK+7BSkNyNWZZiTWG2MiHPFFAEAzDfscEsmZTaa+wWFtOpzXOLs
cSFNibcrQkALCydyI4qYKgV7WBYh6bH5FOzxGbIHkl6w2WfiyRIpIQgGPg/GHDglxC2wpeG61M8Q
gXCUfRMJ/amSsP//Dq3S1rhrljZkj1V5hDzlWwDYNgn6oqfAgNKbUGIMJzaD7NBZ/XuPOh/nuCoi
oTKPllfWqVHVNwtfXBM13JdrP9iN3AASd9kimVIC123lVOhiEJFVNX81Xl2o6LTSySdCxUPVZA5I
dVEXbSvHOPmXpee1WZZ1H8ElEF3T2kFEN7iphdAXvplQ9zZGa3bTAwT0V7epXtO1Jdwf/+cJ9gq+
WALByIC/onUID7bUzmV0HN1EcC3lx5aHL3ya4Kc3tgQ1u+1rupjKyMFIK9TYE3BsDCxN7gsOqbjg
cDrSpkztuyjPh7z71jndKNls29HKiBGYFSGnWdddu1g6gq6sBr5ElBbqf1N6x/NKt6Q31tfdfuV8
f/QkR89/7sgUPv3d0YznDJjiIQHhGu8oKKFYpgC4gSxzM/u7QRjGVaeyu4XvFI0IRx9LuwSdULK2
C5Qhunp9DjpMNZycWVyva52GEG8WkbUUDZFMNWidGPrc4hHaCQ0ZNRd7X7HWvn1JTa5jFUxosVFc
2oU4Nfeazz3s8vDHG/uR21exLwm9jCscA57qBCIwY6OC81XqpQn2hSl/dt6fvvowrWKgjXVTz/JJ
ogLgo4qI8hB9wA/FQjvjKe8wt4MmiyaMC6Ivj76TNpL2VnvwXG6ZVGg4ENpFV5ZM2+Bd0n3oEfv4
e07126vKp8h5N4668fA9K9NC7Q+Kh1t3wqQKxiSsheIr+OQ82AsPJCzoQBN0GbTD27fOY/gbg0vL
diwU4Kkrjk8Pr1yy1vobs0VJoGA+6rmTvMkK61CCiBHoam+FUgVZ13w4v34mwMIKDxR2Lj4Uh/yL
f3v0i1xrt5SDDFkNkLL2yBPiaGNSEVWf9gjDWYAyOdjTxrvO+BPz9Z4SeYYALOgBZLxj88ZTykgy
CtlOE/Y+rWKLmg2JhF/Q1l/5a2pcEUTjavUvnTHpPMU1GCda3w1H7EXPohBUPT6RP9G6kbmIYakC
UOoxzVt3pxiPqDVOKPJc5AYHoL7Qybsi6mLf/ahiPVtMf0nviiDqrbJBHo4vaF2v5YD8j/9a+ThT
82d3orUyxls9Mti3yM4GCpZfMcpDHkNNwkbPhxm3ggFQ99FDr5x/+a4dNK45Esk81gfe5xuQjRbL
FaqgrF2uLw8auV9MvdJOy+mnHlPBRxXFue650Bnl+KNBhPhZ+3GHYSaXo5opLBSJSXu2wS2/Urnx
aZnyG+QvM6bAPVAfoRL3yN5fbiOhEGPFYbTFDcfibFGy886+wb/V13aRxsFjSwaNVnXdaGed77+J
2zwdAchoF1/J4+A+gxRNEBYd20lFW5zJIXYmN3bOoe6tKscUPqRXccqCDijK0fabqEgtUDiaPRfq
GUJPWsPhpomtB2ro7jOPiq3PGZ70tab2xUBRgJ/JD4kMN+mg7y66h3NgcSIcMb6OY9nLZZNXyqzM
5Jb98nTti3j/khvSpa9i+6+xAyqdVxqzXItbecfSxv4o9eD63iC3gI7bAt6yeHLuCRM6k+6rc18R
rdowNef4NvBHpAifbPaIWRHYxtwb9jWCGfiPcQsuxfWOcTxwdhwZXUj+F8WbPPYLdreWUtQlKjN6
07ZlD6ziETsRCqjY4XyXu6IyZguVJ2x3vfaZv4PopOtkp3OII3sbDtVV+LGUBTj0Ac957AQlUumh
HMyEA+ZT/U3Ko43+9N0JkN8IZ9asX+l7TQBZtBfzaKYbnF3PRon2CECtJNzhsPFiKj/Ar+HU5oS0
DS/v2E9IsZeV8f1+QM9u8Qg1kpW3tojkw1BiGH5VkJ4oXxKY7sWz/Hfl5dbOTQu/ogkTFxuOKo+B
OhI2i5HuFtp63F8Ns/DVbb7FIDdCFwZlzOAE4jd8Nv/SeE+xiDBb6cqOnpERUVZ0LpB7kSTaWphZ
MJgIOqkdxHsehFjIN2xteT4jHhjH1p0CkFlBeFoCwDOcXT8B+O+K5jPTLVv7rSpWAlqDt6iR7LD9
FquD2QK+paVoIkS/7rXGRp6FOKxJWn260eRzaN6z24N7PvpE3rBGwNfGQEPhmiqIQo/Qzd5Wo3lW
k/S2eLz/odmEa8qc4trMZAomHxHtyV+crSqQ8a1ADderJ7QcaI1on7XNCDD/fCBl5r5SPo1okt/K
MFXj59aj0U2oSGGZyHkwDecuWy/Pv9j+BA9VgYo44ZplmuGTvWmnT5G2/2PdNShms6u5feBeGb20
+Sl+ytM80GomYlmKliLHrGaLz1rySVSB4Sbz3V6ZIAPAPrNuM7JMT1DyxKZQY+6e8+saOT5KTJAa
ehe3HiUJ3AeWSzT6DnAVEbABfybNk9EGKOB3gWq3AFKmiFKGKciB6EEc4b5S/xLtH88R39ErcWnS
4MEJfHerJWMyw9PQbSUCkKoGGYoRDhJLEQ4RQZFvE9M9vDwoqy6M/ysa0KDzAD7n5B+/kVG56hS2
0KDvM7kWEUnH0baM+MIXPnFJCEHzGOnl3LUB1BIFN8S7tN4bjUlO80ZaIk0DJGKPoBM95QEY4nui
a2K/rJn5ypSfEXmNfiFXqhOZq/C0Te+NzgBODp9qEDBpszaY7JYWFkWKe9Omted+v32IdfEOg/ua
7ytlTuKuNnkyyucufcWJgshJBTLBTwtC0Eer9MWvhGH7VeNIsG+yhK0qdXPYrOEL4IZTWaiX48hL
5TVyOc5FLFyriI5+UcxZ2ZuFi7SShazunE2rcuviGhYWcUlKs+zSZkgCJIng8Aut7kuxWCIQpGWt
O9edDQr+ZtGhKcfF4xQC3ThmgWVLMyPn27SWPMJ25I+XPtRobKcBrhiSifOTpEkNHBqNfhVYGc5T
5LP9LWgivapqDZC1ndba2EXq6w7xVTko6SaLALs5/j9e6Vjweq4V3z6gDnBFSKV2H22R199+nGFp
fA/IVFNN1GkVXM+b3mDUy+sj4y+29wMKb24OSsOw1vTY6GbVRygyxL7TnQGd7wj35G2zEOJ9Wwgi
/e94uWmGVRVoWdDWhlkX/BHyr/VZlnq0y33+/c2BcWuPaQS1kFcEctAAJdXTmGAQZAT2XKQwfukh
QH2zF2a2EOB5quQH/8dhxl30KIXYmefloqiqDPRW54NIBAn+VP6gfnkx9MwglO5qme8T59ZHNHzF
rI3T5Al8Yde+hSqvCUPbRtd48KAuRRzg9VRqYd/oAWVaepJnDueNE0dJaPMhnlH64KbRpiF9MJgo
cP9dDh5BdQY36Pp20lAQEUbCg3i94AOStzuVeZ5y7qCvEx+rYSJMuu+AOG1v9h555O+Rg5vaG2mO
dcw6YLgu4gG1z1wzxeKgdQQ/EIA7aRIjqqehYmsOzheMyeLXyvQB1IcmHGn2Tj4JLgTdSQma/7J8
an/+DQUT1Px1nI+xBh+4Fw+0O/0YT9KoXO6X+EP+uGw/+QhxmtR5ZYYkMrzk8orm8suN4IPt4F2p
BmNlQpxTlqRG98j+AXrie9w3Apby9Zo8IOja3aEPpuTJmW+eSdVphvbcQlsVha+LVac61ESvwP/a
wV+99qjjOrrDn8gR98auDCOv+Oz3dcNADfE/LI1YQTHWdS17ROB/b5ehyF/w4bs2FCcSRX8gAUVV
6CwaySelSyn0tsIjIOfX0GNQUg2VooD2OHA6rfNfPYSscFAgSHtPEH4NCiTe1U0r9kt7kqExQepJ
9YKhnRhmXQNVLw3J0ZV99hqNiTUMIH6enVQSu2lV7wFfurmFXZm68SAlV/jUM/Rj1HKNuj+Vt/tw
2VJ5gCAHoQNYT38LjPZ9xpINmmVwmIQYDKBsrlapQB6D1pZBlx6QyB31LVr/GSqQATzqCTeRxiHk
nHphN07Mu6YNJNoXY6iPVYBNwr8Mb91VO9iBpd6Nb1WB/QRKlsj6H6rzJs3urbnhRHMRDygiuQib
ShfxQxt0zJzPYLGoNVREEu2tIHWKLh6W+tBmD7hV3Pt6NKGQndDTscwBtBDJ33++/O4y0LsrZ26c
DHbrB9UZvX9CeGUtgsTfczsCx5yNe5PVqrclhHWk3mB8mK2VVWQBTuo8U/ex3Rq6QzfzkpD5wjcF
U+FDjvmJbx0opQp810BwQO59pVG63GN5CKlI3YZXIrE3RKRibmcNalw1jGfAzAJ5PGka3s2YqAVm
ph8AM5nTnKk3nQUYUzlxUjia3Ed7rD/4r/4VH+2rTwsI5CjTDsF141zVyzo6jvnUdJ0XMgtBxydG
L8XFi5qd/E482RgVNoX6t34PphQdpAHtxwBAcDhXVhamHHwbU/81nCUwwHzVgccYmY5CH6QpdIiF
qdkgWahTheoCebYrgpsVMjQ7Fx3yFQelPwzVOxDE5EwhXCZANc4tQZgdCb6RLXUC+8aiTOo7Ebqx
BntpwddYf1oVap03P9xp1uVDn9pMxKMieBBdTEKzFM0xeX+klMtpRHg1rT3F0Ao8nG2bEcwA1LO8
fXFL0Y503Qns1Op9Q4lciYVQu4DTTDSDrgtr2qGAeXBcKZy2TnU0GDWJmQX13uvRlkBhbtS7TVCc
C9RNDlBjEw9gjCAhAIx3Fbxtrgp/aHZiV24Hs0s4yT2Lyy8zicz2A5fVihMblOJLat17vrB39Ozd
agyTvgptyZoTojL/MuKWYc5q/pWYcuz95oZ8GCLDneBU1n5SM5KdlzYnXB+lRqSe34xR/W4HdozI
ho5GMi08v+qUN7htnt1GIZ/Lm4yBbdT+rhR8OQv/sVsqnKDyYqcEwD/ZAUeOmKwJjkOmJQkX95rT
LyXDkrKDBRxHYtD5f07lcedX48BqexoV2O5I6crSFzJAlO9me7vzLDDeSRnz6dsvuput8dP/amjl
/ymA39XiFAX6ewlnYMH+otdV8OHEfRdGdIQeZluLuFg5pb9mNDEsuHiX4BAUCOm64pvbsaMtqdgL
UyN8Tbt5l2CRLJUfeSktggVPjPoshPuaRRxuDHpk5J0VA1NNnS7QSZJguXlOJL74Q+hqVBugYyCY
knpgst5fEIaqx20YnCEHsnDm3AkI5qBeQJh0bqDr7qiM+zXxIiyitaekvkoGL/T89DbKwSEk+2lE
qr0Zzq3RFgKTg1OAaWtOSA0G1TspSERhQ8xMeWQeTjCJYG8hDSlB1Y4jmdgIypApLZbB3Dt99DKv
/Os2nm5jMDx/AqQkJ2uROe10ht8Ujr0S+Xri3deSRxrgkVVD94rZ6tv0OqAiPxoJ1OFS3ypYmtmy
8cr/3LHBibZoGpwteGTVeOL9c1crCb12rqBWJ/vSZW6Rloiq1fe26mpFJORRSJly7EKZVs4tb95t
i+NncJ0WwHPldyR+vft+uypgOeNNBp6CANBr1L1TJSfJ/EKuncllumh2VqzUCoBSwhM4VKgb9LAp
F30FIG3X1CO8z3rwCxV8Js5UAyehsDvCUQVzfng0edpCqccJRkr14CAX7nsWBEHl5uLI1HNXZWFS
ebbxVyPsQwH5BUyVzHmeKRepk7Lp1tIzUNwSGw9bR4ThDB8gKV2Wn37EZYjkqVoC3QVnlhiJO5u1
xJC/BEHXve6cPtZ7/oF63X/bmVewHLKB8A3463uqTC2dDbRSp/kFR8dE6wLxKRn1wKAf08bHGp9+
KuQA42OAvg6lfJvQdS05N0WGPp2PH5ZiaDIL9PNi8jjQkKKao3V4ltahtjUfa79akSgVoYBRs7Y3
69yFvgsenOKzArysweo9nDr44Fw8zXdgIHnCzf6FZglVuJH7WnZXZd+EsDHY4XaKx12gHAif4Pqn
ForLYBFJIwQV3dAETX18LYIVXzau44z/1mcI+0Zhp+z/sQHKcjAqB+qBk9CSqK1eyRkfo4X5MT9s
Fa8NhXeiWtRGT+TSeqdfchClkhbiGzDuLROsrdMdnXE79rwEt2gV3L376hW9+tJh3f64C2SMD3aZ
B9tPPe2dvw9rI6cVohMu7o9G4pOG6RXS1J/eYgzZUbhyaXLWnK7MwBfjZh9siqQ2+4R5J5UQfK8b
fH/BtaDOddxz1lUXh9kO3sCY6rGlsh6/FE50J95ew44Cy54uyCGUAWMBPwU+jdbNqvV8LxCjDMjV
CocPD1tlXJBTGEr/0T5/OvBQ/ojmLojmjkImDhhkUAKA4CDKcUIJF8M1M0J+XYLmASHHP28nn7II
d4d2nNwsx0EWudnoA5dAhCYvvJoHpjLsYxUJlB/tnSYpJ/LKGDKNLePZghuWHw8M+5V4tnf8sZ3b
9LG5nnD4k2dR3UeGzrmcp/jokfGGkM8uk+haidM/TrxCVTSsLCqhl14hoxk7d8Yz/mknzGS44Ma8
0JmmCxm+GFJ5xTL0SfidOWkXhO1x3Wfn49CJP5VTmuIOIOjRDptGpllXqu7F9m9H0QPELChUy61B
HC1zAHduW8QllGQme6XyD7jNYGLruMzgRDtB8rbV5znLzSze4tpuEzW8lLOWFv2UsAwhAKWGqeH7
1CNkSjzVzTFRWJp42QcHcWsZS6cTGh9cpd/zs2MChBLQpc2065SSVqc/YGCMmrMWmRuLwi3sjguZ
Jau9dxjHd67e6tWLEtQ4FFH59V+tyXq5zJv4odMKL/Mne82765+KS0QzbJxtYL9wS0qLOaiTaT5j
f3uVsyJJ8IOwvpBMUb0p2l1u9eoocpYqsmrQNNjQNMuOy3YAuB5n+Jn7ivkxxMopnfB8VR3V6jnh
Fl3B8LN0AI4105NG8SvmbibbYPoyFFZVwBATEvPMAKUKTomja7XFshjR7e/o7Ts3DptmGOuC3wOZ
e4D+zrONx5w52A4itNlcZydvgbbWbXn7OWBM6U3pFl2qetXRIm9XdFHn9wt/F73k7XY6y0qNp6yw
Kr19sDTMv11wNip+zm6zJ99fRWSx4oFXfb6eaA5wFT14bzolBBktp801LkOoHIFS3ITodEG0UVyn
hmrL274LfyhsKHE7QVl5GCjmKYQqdJxjP8eKbyjt/Lfmtya9qrzkLSGg9mytu+g4tS8c+w+czdaa
XBXB1av3Sv5d4UCnP7/gModTruTcPnu3rnsVaUZWN3FOcgvPwZbENOcXDmy+Oa+Y9h3qAlfkqvId
vYJIjw1Qlkh8oiawS7zW2qjSolFbXoASXEVMltZvcIENUH+dpOXNqkYeyTTy8LqRgGTgueJ54ZV6
BqukCZb8M6VUOtkR8jgqpAu6KN5f8c69tkNRbsyaV5kQeDlEtGFxiUC5g7UhCRJC/M6K0esgOrdt
q+SfA3rXYBUYBL0zaWdlOLM9Hcbp0ZxrmEeMdOdNZakkCWhM1jfhHjNgfp/Wljt0v/HzDj+gr+Wi
w7KzPtYJm+q9ghAx36VjmPLjBaH4G3V8vHKW8YFrEbZrnUbQ8vWSX5N2ZRwpk6oYNVTzw9bwpr9u
n+tCBoNW0VMjF0Ga/2oAUgq8mrFvbB3cNojtDOw7j4jP9ra9mVcYW06FQYw6bnqy2AY3PO5EdUt9
SkGxrDRLUDRsQjsx7wuIFgGVsuuHtYOnaHBGhAQ2TAf+wCs+tyNf74IaDAFVD9KKI8Tb6BsMSPjD
6ZazAXOpqsS9Q1J1yLLzA/zhOGgWt6Wpyy+705CynPk0KqV+9jv/lpPgRF0AoG62iFs4oBAY85eW
6qZh6ksogXbsDW2zIz/MFxOSlUJf/XMUArBbR8tb8asSytQ5iOYzgpqociVzOZE+C6zavulf08Sk
mjGYtLPWvpwzjXs688YJGN11K9QCP18qXl3e/NOrL9FyIMF5nK6rcPaf5GT02YAoe2TVA52WbQ/7
i9Sr/rmN410ln5Jca7Ze3dguTWVkAkOkRMpxL9X5LgcMTg95xH8bghjGnMcg09kxsYo7Leh37V/H
kc6M3WtP57in88WbzUC1uuNbR8MRJBfqUKLauhB+TH/uBzGQFZAbPktkE8Wp5JhzBnt2MMHr4AgN
7qPCwRaPme/yXzR+616jlzHf/EHhYY52kXccVivWr23f8cGIV5Tua7Jp8z5YugDwpsYbozqgetPJ
H9g04KVECPIqrIbAUE302u7c3FX2Uvx+v3hSSIdwtNZPlKi500+kHzr1/FaUlWM+tNPBeEnFQJdw
YxA/Ppx2ty88J/7ffJoqnzRDrOK8+OfX6iXiw+lji9Ut5cMevx7ezSuVmjmPGq/EUmkcPSENOywF
T4qINClsgLvr2S+lhoAvgrJ3eTCkAvTTmmyKLVShT8nKgUczUoC7gTwqvhpjy1aFoV+n0N/fQDH+
p1hy+qJGCrbRHG3cYC0R9zTYzvn8jLrUjuzqCqLVGQTXNe5jY/l0hRqBpu+YCl9J1ggz0pPvMi8w
dtpaYifiAxSE2WhznLLFuZ2cNkftU/W9kZ/saZyvdb6P5DA7HTnYwhc/Wer4M7Qbku/f5y9qT14b
XiNmkzaAl8gEd1fPTOfui1ITlK8WCm+3YjpA7RVpN3jW6Bont6Vzt37RpsweGvogo1MYLtY5Qf8v
3k8fXb7XCSfaD+25L9m3WCJ6JWDU5dqbAhKF0+4YWzq5GgzeUkUY5a9gQxo1UJiQgEkfXf8e7B9J
kLTlU28XnkItTxIgf3IzrLZ0ziv9eZLc49Lbn9ZYQOAtNNklJGa9P06rqJ/djgG3omRIFED/A3vp
+6GWxl0ZeE6gZI2Vcihxus52KfgaTAkaaJtlRc9B4rh3xQ8qI0c4I/mEn+PYrezHRQSp6MYuUXcv
YNn5S1KoFN2CZjevHG3XPxZ3UQ8VQPcmra5T9YJCnH2jlloxqGs9zf46RX85aoGV+r6kdX0Yp/pb
eRH+9Bux7jjrp4Eb8uhW5XdkC405FgqPyBiH1G82aj9xM+tMKnjcMNk7hcOBGVtiSN0jBgG6CGuX
Koe4X7Pi+HAv+9Jx3L4M17SpNOyBumDfVgXlKNPXBoP4ytByht22eYLHR9cpGE081x9kkH7Hx82F
RLncX5Zw/ZviajXmEL2IQv+2/BFa+QTw6R/DHfj5O6ThyfSeY9j9h6uaRDLd7N2ZZl7Q852Gkv+1
vT3I6I7OnXtyFevJHNRu06r0ymb0EDFh4KrB/kHlZct4566tAzdNOB0kQFB1NhgCUZP7AKZ2tnsu
+1YmgGskOLbF97O3Qs51P3YdjfmgIyFQAEFb+RRaOU1gGPOjSLQk2udAOJ72yM2sGIo9Z7mCPjOI
xRusJGpNqOAqhdwvkABD7JaYdforyvnDiPuM0hslu9G50hK+aWlGqXPqtv+itBPV8Ke+clPmhsXj
1+Wk92SBLSFvblsgmIfKWWmJhN3b3NIaF3ivEqRubUetivCDI+EwtyUHuF15mQ+owJBrqhpbnsjl
hRPPsHUzYAx5puFbpnM9efKR1930YJjt3OPUNxEsLYp7hj/CUpR0202iGXMdVW+ITrpdlzC98Crv
AI0u4FCf5pN5cxUacT98N/70dVexFYJSoRPrRNI8jysS04g5RzBMAL87v+Dv85hO0SM7UJ3q2wr0
wEA0aKrRbw/mJASdGviLe2jYD+MCGNvlJoZ33jFQqX1tQ+VkONOWfajl5P/EPtewIWSCGww6zIvs
lN5lNLjvN6H83yTeilJk94kBCcvcqlq+NptM0Pp6CqDtXM62H/5gsmfoRsu+mAbOPhI5j81fpn0E
Mh/fs4bLvMQ2HznFDEox2b7z8O6kwoF0YpQf5Drok/72zp+HxQTwF2mV/oTMdXoP6teWD7El7XWZ
hrT45BXnYPJ2IKDFwlqDeleprnlcUrmB+J2Es7/RXavh9HvllaZ/cjwZaqOTtgbmnawc90j5SF16
Loo6Vu3u/6A96ph+fFEJZlTqAIcXW4a8PVVtGkVgIIW4GOKkWdsWDIutVKIIv3bEmxNbf9qpt77N
SdUwdir2N0LsmCRlq3ISb8ETVi0atULuAbRZIpSDvUKgMtS/D/4zVvOGZJ2mDWiel//VXA9W4/Vu
52ZS2jQw2nANvETkb6IhxQsk3CN0axACZITlDeo3OKj5I70UIgtVAcNnucI5st/NDta5cDaNv3ec
sCTtKReenYk+wnmLUYF4qwgi23A5VY5FyDxHz5MPkNWgDhobcuaTxBSDdTcVZ2PHc6UBmb/UGO0Z
RzbCOYOyUds0sYu36RkatuhUFJXUF02ht8rPO+ChqMKfvVplGPttHpGl5YJYY+E7HXwrpObqgOis
vULW6ChHkI4tIXbTwppVa2Ud2MEjVjAnVLwVjDBlXMyn59Nswj+1SailUp3MA2Wl3iu0wnS87Z6s
nwycjAdgP8tguzwKcbGyq/QzzWBTGOfsycTuoAX+lW848tRNCAIF7/0JwhboxjrlIbOglAhdLjH/
8KJTMzuedeehhp7wcIrFTYO7YU07wmVC7MwGY5dmlyZ0j9vnqO/twKDtny0b+sAaiUKqzMBdJ6VL
ggNPIlo73hJ2kvUGlo9iAXVawcZHp+fp8T+m2GGsN5nqhvvn8+90bBVFWR5jM54SDA3mSk52fmdA
gHd/qzKQc2RMWqjv4cE95A/vsAMjGioqv91zGTxe2DAHbvKMH+Aj8AKogDgRrmnYry7AD8esGOIV
wY3RUVXAZTMY3J9fBqiLZrtXDRDJq0EPhDNvRZtBexZqE01g1QPI+slCGDwujkdeU16b/E5TOBhS
YHJhEkgEFuhVxdz+DIeqHIspLvjIEVDcoXzAOWGUAIc1ITus1clIm+TjvafBV7UHIUN10sDHMhKj
4uQJruHx+yne4tcWf9A4i3MTVuuXo/7fyRt/v0HLk8APL6kJCXv2ChTK86qBwUs7wervPn6gZD+x
aA6vsmGmnQrWUk1abSPXtc9ZlIyafcBsKvlTzEpKSb9mmFPaLlyPmyurRFAqky1mt3v1V1myXwIj
Uhc3GtS8frYDUpJU3ED6fdHzucs7CR9rELZc+4fxYjuSb2ZdNLVmQnJSBE4SkAq2CLsDlNYNERUD
shV+4uzqFio/FpXbtHhxqBA63j357LA9EyS88+NXSOIFKrZqMl72u0G5ULq9PuvpSBbkONOjo1gu
kM2UG8shgtkwTU2LtKnCIkn+I/gYtH3XMd55qDZyfuV9CbANtHJAK1o8bqNVxK9sRGDz6xd3zFXy
c31d1mZDjB7ZB5veDf9FBnTuBTnEY++9iA/T57A8OjgZqOUToAOhwlCotpojyl20+H2VTwmCuSex
pfFfQNpRQaEl5FW4QbffhKKRGlhP2vTKSk0OutN6uJee+YxQyYzCSftWo2bH4PFkN7of9JaeL9Az
sVd6rsal1hVVDRtk3QnkQTtip4aL9tsQE6StvjrzT7IF9kdYlRhIuNNfN8MRjxITtBuc6LPVB2/D
sYMhGc369pmY4Pd/51rmg6lpq+598a+pPO0sHSaP4atWL2xsx5sagG+pVYI1paHM7Y7y7G1IbUdf
d7b9EaCZnydQDrNj0fC6xnRnA1RrhyEexqUfkdeT+SCD/vsntvyqM3VrNGyQmZ7ntqUn51qAujoC
63zc6QptFu3v1kv+yYCG3Wzq+ZXQucDiAyKU9M3svNUeiYNFlrnVoXEHBbS64e6ZY/BYqwJwRSHb
659cziKFrTyAIRtJcHsO85DgAHmbFY6eJ1WMj+eP5YZoS3ECHfVQ8C4JZnj9t8U9EOwxV76B+8dJ
GiAnD/2JpdkN8dUNUDUJ5Lp9yz1BzND0cuRZ2NDGuqYBIwJNERuuQrE/BYUKeoA1CK+huQUMGjJD
dzXUtKC2o+tAuBXJCMo3F9G83CgAYgsoIlDEcZpwNwCdnpQK2tRbKFGp1dybMdb/jjFoA/s5VnR5
moSBqQAESxSknnQUz55T15rnksRyktHNJMQz7UR+pkH3i5v2dqFSTT2xCWXBvmNVh+RMCTVHyqob
FKBAci/5L3OPSgf6xwm4yAQ+BwvwSxeHSW/GUXyAlK35LBNJZEK4jrpwxSf1Uzi7OZaqG7hGss7c
kgI8KDdYn7TCsJ80lalnyGx1naD41DDgpcGeDCYWNUWIY+Bjj4ITUBFiMr8vziK9E3dLn3LLyLzb
0t7SW4yDkx5o+PZTiyC6cObftjiYJqYHy2d7PsT2ko+//lP1OwG0SbOL1zwNUE9SXQVzIMHRrI6b
leksWLzxzqrzDZdL4QU7noH3lK3lMOEN5obC7o5eX0O5Sr3LJ/a0QoaFUrFM/41CWxcb/tJhMGyW
1v1KZBGuJwuut+eykSKKht6HhC/kZVdMXL3TUzo/pmfEC84b3Jc8p0ESzweu1oWy2aIlt5zvmt+5
hnws2glHkLZOoVrw7eSBA3F4sfGAvdjcVGgOKx7Uc7Sdr2nDBtnTz8g++LGm9goNM67th05zU1D4
m6i3g+qjtbm1Ir3NGcTnivyPZ0Uzed2ewOp+lJMwE0ETYGZNQmSkkpst29LOcNZfLaPhL2I3jUG6
grlqVhjvO16sIxp4xFJfTwFktK9ZLnB7reFBW/ZzUHvCcRL1k62hA4cbAhfVs0hvbUzRFSjHyE8V
XzQg0XCvTzVjaG14KJQmRn8Aa2q95so3ENAFvmwupBm/uQ/FNpeLhYC7adcGEhCKGCEY6JB1O1XD
5RRKisq7NO4YQp+Oi9ZFy1C6Wa1rCd/JLsm9UaNqNEMhNFSBMijc9GrEZiapO8FpAsUKmI6D9evU
0xsaSE88zOYVaNlTHOTYRdMa8xvvtpEXv/TsxW529rJvdRoN+XD5fqWp9KU6bjy4t4jQw2iEycs0
H2UEYobUT+j04MBkxLwtP/rfHCJtvkHmrc8G57dguM0FTT2otvK3rWKmrXfo0sG5vVcxe9HYOgaB
6MNyhQQDNnxM+MoDDXQgDSLsavGRfUNZF5GhcUwqMQp0Zi8YvYVY3CtpOGb5iZHtLZtC9Pyr/1Q9
wE6iKy0cOKA29ttnbEM72a3zR0x/5ueeJeiv6md3HscW+KJHECLIn8VCsb3iiTDKu0QmViefEpL9
E5h1v/0Cqi6i1Bhk+JWJWuERtHpYnrakM4ueAu7NB7XpwdUgYTAtIfoFLtaW1//I6pUbw7v8/k+U
kXDzMW9IpFlFwYiI6NSDffU+ACgW04AAFPDl7NPer0eVMbnihMHV9D+XvfnTrjsZ7SbvPUrfHhzB
XHMrw28CsvETtZ946zTix0tRtmz4arRu843hzIaWTQuVo+NtaXfHlYqcdh8fKn3vxyskKzqRkut6
bQEaCmMeNEks3agOtGdgV1qocuI9wdEhi+FwczrX3v42PNnFzqvkpfBiQbJrI9DcxQ7mtJztlW2O
+pcphqAHixAltx4P9mITRi086+M3xn76ubtE8ytdkc9gU4bWVID6sQs6c0cSAA4MgYgEWXWQomY3
hSLTDSMtjnx9bjRD6kZ10OXKpqRv2djmB5RhH411AJPIOH+IlTxkpEnYOFI5hkbcB72jHrC7przT
GgOHNdDreq/Hi7EjXx8/lmV+DxHq0hu2Ou/F731wPFEnnHr+MAnfOWCUKvFLJJo0S4DhzcSEOeOA
FhAacMKl6UfPqc3bH1urUnZXmoATuGFpWcMIIN0Cek2HRlnx+nF0KUj4ovP68KPbyBTjmak+mN05
QFrgJAwvWYB97ztZdV0sVkn36guLoK50nxZqj15Cyu5ghU9HUBnBLKq6LffDopNT7Kyd0d6DEl2E
nXwaxILN9hCNKMa+4w5cDkn+6DdN0I/7GJqld3N4krS7TbCwyr6R39msI9arP4+K3NRdjgxBns1u
KghIv/vm1H/pmT/GuE1R8KzHqOZsBDABla4RlbDT4ZbgiK2hhE+95Uy8xczmSkzQnQzsXTjLkoC4
RqIlGW2cOIPpHpR+5aQVyI4gA5lFrPxWzdFry49GaIm6LRsvjh914RkrDwuGMyUIw6xLDckrz6nX
JSvImhX+a6OCL7dmLWSPRl8iezoS9RGC8/hOgi3FVO4JKgJ7C58YYIp4cW2mBjFYMf9agT37ZYF+
ohqwZ7hZMzbJybhmZLHHyymiOW2DscgTeiN1B5Io2OAOcDG6OiFE4IfvUeXG+1IXvs6MEADCNz7L
Ohvl0tZyNrUaWa1RuRMoDwf7tBfWafDyeZkU4bLdidAQ39Bi0gdA5wHyFQAZavjOOYA7Q8ukw2gT
X9NkF0l7LFiTDnsKzUojX9+9PWxg/IkPuOQDHfIsIXdqsZurfORw+s6UdfmOw896DNkJlho9FgiL
e0ZgEg6e6qgbUVeqFg/TAGrQa2vthH6DTaQ9yJGX5NovWKQnkLGk2blzj0qDajTuEhaZzi15sI4D
s0IrRr5n2STrFi+tvqSTA2mto9qiJKjdGZdWN9VLXMt90tJrpOVfTu/3ipnatiWY2agwyq1fSNit
3C95OX540uU9Cm0w1INWJueJTR1p6hyImdmtmzCJy6roIUF9OnlOgqneNSe4AVZiE+bfcz1tf0VK
qA4F4s4GnYcWYFeYaNDL/C3CMMRhDVwyFG+OQr9RgtpEROLvSN6lrrO5UrEywFfL6R0yEb0zEm6J
rYSG0FbP/3/Z5EZe43xtcvRtcUnpp6KE9pEtN7ZjSr4WSlNCfZYalmK9mYg9Qo23UhCw+XsaPnsD
UjQaFEdYtc/8gnlO5cgpUKt/xvIq1B5aAjfKp8SKy0EDwvlkPqXPrXyuXNaw0gayYhbWmPc+aUy6
CefiUoRYCM5ue0EA5KFoBUj2QHAPyV7S8GIY/XzxmwT+uNwHOvNvogbff3kFq/G4nu3n9YamySat
Xsv7/ngspAVp5ime3AaEacwzdj1vRgVrHR1siFciVKiBvNTmhgSTe41tubtQSq4e80dmJWCYwUUO
9ziiiYDdwvuoyHU33MRVapwxwHjmQGNMMRZctICEI+JA2rBRoVUFjE7zUlb4bEksg7EtsbUH5kAp
IfEHf9yV9qdrGj2F5MQaxQW7SViVAhGlC6W4btydworwDHi49e3uPnw5WPT+nFMuP1E5zP64t3ay
CJL5Cxvlg8rVF2QxswXuQp6Z5mEYNlldaMiUPqR7UE9WYnaOXt1QCxDH+alV+LGzWjJ6kC3FpbBj
QS53SKlxAbzeaDLZSBz70cJ3SKADezIQve1/m2DSEmVwE2cHIkCDoOiWlxNG1y7XEOurs9Uar9rB
8hWFZiHObKE7K1PP2vFVafAC+ECY32c80B5LL/p5FtKOYhkEz+OFwRC0Qejato26ds0Ta7tK+0VX
Tfkpu8m1XhyG4dUGmmk+AcNzhsWqdg8gnb/vJkZ8JC28rsL9uPHqVd/dG8cVNr/QsTrIOxhr+ECi
lCrQ9GDpgXPfmxX8XT3UxXSgbkOTDADmAOnEnliBJoIshxaFXIwP7NrXDSNfNNqksgtOrriA535W
/IBm+Y6vToF9LPdqrfElWMVgaUX7zRlfKAwlxh0FpIv1QD49wI+dSWQlRxTflMSBuO+zq/HaNQVw
LzcrUIRYRSCS/MzvjGkkV/wXb7Tb9/5x6aZB9wtlFRdxx2698h76fDx3buB5sIJpuZ0SFWIW62xB
hZdKjxn3Vel4RucnIylqz3xyqFdfK3ttUjGw/MxZy/sCltqFumPCV6UNHtcnNG3pZOg5FObT4O0x
/ysHMmYrIFkmRfJsCPCKMuoKeM0e4w4eive5H+O7a+ABCmIMmXJBjHF+xIwzj9PbwVXG20CisgHT
NgAgz+oRBNooyaBdbEuJkHcFzxtOmcyTeZLtVdRUlTHi0IpC3mOqdLEX9LEcDWkTMJ9umK+L85xL
5MXQWt5EydcL/M50dswdbxagrLKjLS/R6qIANjnqxKq2xdDxyVJx+e3E6F/vOVIKDCA+H22uWHNM
ht4mxx12GbEut9T33ijDc5iMQz7zp5gJGex+4Z1CR7daJ+61bUseIQYobglszIFagFPVW38Zoc5F
BAHxgbT0EHZZZOJ0lHXAmy054yd4kJngpW3dTqOeL5ls/qXi8jEqTcce94h2SCvqj7XPCG2f/392
yZZHWTp4wfBBRcFfgzlIrxCWUaRRw7ZcYsm/poF2Codj0IROML7Emdr7OEbGR1I3VLnd7imfWnhB
Xq6qphYDzRJb64L0t9YfVUlcFvhY+F3JI4xyfR/NDxVRA1biE7guSg47b8t7qLTIsl6AZ2zpOlf5
xskYxvkHJHe6+hIVmVKJOzafCui77OXxwzLEWv65hogmoo2z2VuWyE9xu08xcJoKmoBPuJJSjr10
QY8FJ6UYn5LbL2jVPgtLdW+9rdM4GSbnkgGqaxvE/rsgDA6PpX42v0tmNsUz/jOTVS/nIrolJ2sx
bTe3OysPwgVr1/4Cgshovn6OK5mPcgfPfrhonSU+MSdkfA8IYQPiSmxm3w7UKQTKmUwDOeIgyxKQ
579yUPsN2nrWs0Zb8tKpWgxuAYZyXr7UZzJ1yi/gJROOiMOa1PluXQhPbsqyx4nBKPo/FmerdZJM
v6+QkYrfK+dBAizolYLMx3xOKH2Id5yo+jX9+pi2aVngaUSTExsktWGdVfMp2/RSN0OkmQtpQssr
HcYBMwqYn2FmWP+P7Lm2CB8qQWCCAie5xV9t7oiSjKycaZw/CJuAVje7wJELN3TMaRroLcpOzCEm
SAu1f45jFlvqIhKt4Omj5L6DM9c+NBVJ7taW9LaVXRMxu3ueZtAMkaXy9yG73gGAvBJCK8kQmH9y
h5LWzRXAaEwLiBexV6p5XVo4MNua3m5aerYd7uijAwwmZKoW6zdxP44H7WiM3Hfc0pnq48nrMnhQ
VaO5684jn4U8UHnKg5zHCbsZ9v35ELGeslAsVUnaVSwJcYVq+noi1W2E7HIS8YggSM0fUECaxcZZ
VYGBEWmSZqlzwzIZ2/u4BpLaaRIYhVSyajancbKMEXDI25WPK3Oid9dGQGukwnvA0FC6rueYXla+
1IQ5sqdGEnJPtL3ILT0gEm6LVlD03lfBG5cqJEdOPs6c6dXri0IQfoywZRUwTR0EtgjqHqGAVsJ4
Rf/wXYcwtwwZZy7Nh5/jQ2Zb1pbp/Q1ET3r8pbFui6HjJmy/gNvwICjNJZX9PBXK312p/XsxmSgr
ltjkuxGImYXgTwuJBV3RF4rPYeQzaEKQmwMKsZTzP9GxEWvY7lj0MihD74sUiD2MHuuFs/Wyn1V4
aLA9JT4+3IlhuzZfb09rR16IWKpEt8F/hsdozuXgDMcTTMHH1/aUm0CMJftR1hy0z9WN0dtJT8cG
ljqfVIr+aCzRoCIr2UvOO73ATLWPJdXHCdmvVrOhGufCLbxTMDFvqmE0Ko2fSY0YJSa2yG3zXNfz
+61pX0W4/+gFIlplBFov91bXQjYiXhTBdf0YC6TR8MnIK7S1l7GUPbNvKs/FO8FCb2oLE6TlXM2n
1UG+7o0KKFfQ5nd4J6O+0DamFXqLShKMhPlZZfe17yl4rQbwvKRMyXoSqnCbSp7asoGgsoNmgLrI
XpiINwOiwdaUYJCFSYb21Y2d8WNo5CKGzLvm8p/YPCZgCYd2NrN5K9qamXaPHJnj6a6emIh0c6Nm
LvJvcuv2B94PoaGPTwR6gFOl0VUljU1iiLOArfHhniK7Jvd7rmxzHFQgRngkc5foqF5lENEWZX5t
YcmXS3Xu7iPrYJFwWk+qxRZGugxGmgAtpVINiecZW7zH7mJtKKk1CmKakz1AdhnoCQ+AJQ9vPtFw
21YVQ0UgjgY4yuw3w8Er+FIED9y4j8l1rgO6/RN/EvBpMW6jsGabrWAxQY3do/2+dE7a+HIQee7R
9pvRoPQ5Kd+t4MQ9SNPble78JwzJMKgzduSihPg/rv8AydNESsELnAWt3aKYKwRBK5OZAIBEH7MO
ry19m8YEYiHnZxGOdJbeTcTmLHRzspaMLmadF40QMstnvIbfOZBhSB93GDA14Hg7BEprx4IIdaDu
vaHSdTY0gFcJO2/zcOql9k9JDq4WuKNyieWy4w361/3d8LLc8XcMuGXRVetgB1r1nmINHqxGQe6s
jKIhXeXCuBJhR1ERxqEaK4/lvqpbYvj2+ET9eZmPo96dup7lbm9JxXMebzxf/+Hg4ktsecbYHnYf
W4gH900hkbaT1zfgBg4ZMEq1P30KUrOalWkrVNmsIbyAP5FeCMjCo9kkd/IIXH68mllvg75d5qSQ
ZxaxwZG9Xfnh6RpcdkWkmqppTkQP5HfSJlAw2BdqrwKRbzbxyJbj77P7KRCxc/XQ/8aXNJNgJINU
+kLDEgB+kkI9Yu8x+JynC1n9rxe7Iuvels+9wPz7f7xa85ywBhTS7leKH+/w4YIKM/c7mpcWhFmp
Tb7mqTgLZb6yBScWfwQGOVGwqVALbj4O9I/7qCzsce2jorfLfsHxZolyJ2UborDSU2kEz118ZnKd
2BoGOyZ3Ee6nRf4vpo7xEYXY38ExQCmcW8gu1kAxzV6w9QJxcVHE5hI/BearWJ3CKJM289FageEH
1VG1i/6/nwRAzouVRQUnvN0kDt50wJ6YGuVavGS135Z1R6dDv6NrxwMyi+5hG7BJpwKa6Fss+9QO
nw4rztzpYgjxLYbZNp0alcWSwszrZe4m6MQVHDjqeSJe+pQpE4zT1zBbEmHdw03AEE375iJXxzcr
nWt+86Mxqe6d5sjnOsX57RDuRNZSIijF9jzJQ6O60IDxS13jJ49q7AVYuo5JAJ92s8rSKCUK7Qxs
4pdtCHlfKscsLn9kavclP88hcKhPkc2z3gmnN0ySlgu9UgKERbmbQAzBPbYKbUTpW2jNf0XbRpR8
dFQ+4Dtygly3kz/YQ1vWharXSuWWC3PKkfr6On39/oXOoMWI+92LqUFQHv/NwlI7WkjBnJIgSS0D
bMafDjr1sdh5RFcdcJRBXlfgCwKUcpmaMPHEHkte4F9Q1AV+g3VnEMbjgwPBmA5aAnLqQdVKMHT5
nDTzbNdCg4tW6Owi7bsQWLHtGplmsUG4yixLmUcDEONyYqva4ZC2yQPeRmBfBY/V6JorM5eZBmze
KByYZFTdnr0KK9yEVh6DBL5x5a6re2N+TwCkQgwpKOMJgVUW0oNu7yO7EsA++h6Bt832qCgXovFL
BL2D2NmdyC5Q9LZtsPPgNHM2lds0UO8Hui6pJeq0s+CXhMqu6hdTogBSrLIihmLueTgoDu1qRVNT
EaDrXI0DETz02Y/yUMxFo3z0w18rgcaaiB2H1IGM/HA3ma3fprhHvQ5pK51hmUUoNjbxb8EM0ZQL
Ut5F/AKUT8kGeG8FRaoF31L+ACSd7iwNxSPzOeiKIT1YjOqSImLxRlws1rGeLkZ1Uw81ndaNqGAm
Vcn89gZf3o5gXxPEaee59QiH04hn9xqwSdBDF1Jyq13wLSdqR/EcfG4hzBSfC1utyv1Vn7sEy3nt
MP1OLzPHLKS4A4NvJoaK6nrvuBYbAq2JyCD0DzrgZWamDpAAJ15vvPdrDyhngJVnPSEvHGvU656n
26Zyq3B/CEJq/5cL9LGxbrfgcNOwPO2Mlok24Y4Ut+36Ytgi6iTv3W9eP7whDZ60EwA7+RGNWkQp
RehQV2nMPdzl6eDj46MSqyZQT0c5q/r2yBTNE5+r8kYowF6AUKhGBEXTmrgQe237bEAs0vFA/lNK
qOACGmv3+I8DMWwxdtxfcHujmIZwibU3Bz+twiBcFrSRoO855jGiFBz/CULYesZB4eNX2M5rRfYR
OQeNKuLvzIylqYeFXVGRF2UNXMK5/slEXDyboU3bTwFFCDagMg85nqk3CqjgSi3hWNLxnWhF9eNP
NdUjjSM70XnRfZ/J5eMRvPr1dq3vvcp5ItZbMtx/WovviSgZ4iD7+TEbbuK+2/Vc+QDJg7N1gX+L
GW5oHZditd/T6Vn/1tzzlR6wmt0TnqMfb8RUc7ARJf3+boWuZb+NhlopnyeH0XRoG+/lfQXutdmV
HoBK0eJLqmAOTwJRBBacUzWVFBqzsvElhWucE4iflimOU1BpNXheUg0T4vy3yl5d98XM1cLkm4fx
w+8e5jkbTBqiNv4/y70hDJbBWwKsezbQgu7cKxzznYxpZN9qidQ5uuWBKxxdHasIKEkwa8HDf1c3
AQV1YJciYMISkxLxKeAv99R3qqvgYi6Vt4rX6iPDwnqwlpNrNy7O9fj74rPa9w4LCGH76JDVIYJh
w5ujXFQeQ/VYCrSBIFb5LET4W7gUkhYaFGdleNZHEYkoouBhKsAL0kqDluHIbdvASGy7pM/qduPd
cr4Nozmg4z50MhT1JfcUN4jXzLzsNkv72vs4MFtkEocMbNA+zczBAemTmHkxAl/VCh8VImbaFMBL
dEUJQKuWVSvEEnTm9lv2jzgtTzpx9G+mbJP6xtpv087kTo44TUlkaNoKcyb1/KLfmv0TCb/w/kqv
zGJKeWEwWy7MLcSeEoy3y4+XSmkSG0pzyxM/5wcioW62ZN/HwYHoqf5Bss/OPQikNifAYi9gsvPE
8wgaDA2nSmb9PtRzWlj028W6taOAY8KBFXs//5tX4dFEv6DamAh9V4NKd1mp980fVcWLFrRBmFLX
knzfyTbT9j5kEWKUvmov0sQZJDilXNH1NcB5PlnB2mL9hZy6q/Z4iAlG8HHn00weJp5kZwSNSWb4
tb1uV8+xAtYEDccpwQ7AvyYSPUPpSHBdvqZR7nqtZt7h/rgOCfRqyeAqS70uiztTEZ7mqeR60xM5
VAvvLTE6EvGFiwmptZNlJ4eWARUej657oXy0hBmvIfZ3VfgPPlt1aldys92YNf2QJ4uJaDfe1Y3W
u8sbd/8FsJR+a0EI5pqxmVr5B0DzIShnfvvpZMN0UYGFOCSFQrR6WbX8J0sqv4XnL9RG2JUULqFQ
4Tti8+mQK7kbiZk7V/dtd8an80qhSJsOdRozOL246YLiw9UQo4iOvpmcOZo6IlWZ9ZYVydFkGKdZ
0Hs5YViiTVdhpvHTlFfMwJXsKTTqKD0vAL549RtbEBKH3f+/wtQaOwyztf51etwQ2MBSxJxGgqtI
Nkl4Z/DsfDbZ+hJIg61KyRFQ3JtzI8kKkPQjE0I2siC9i5jvZjhgKQb2ouK5VxCJN7ZT4zc5bRh5
ZRCirhou5h9/RBkFexaOU7Y+6cdmEA5k2e3qZz/G27rOxDiDH/w7uqeDaDWa04kPZNIfpiINAo/O
dTdvPAqXKtmuTm3Bze2tscf5Pi7xbzZ7rU2UJ+KZeO0lyNUrt35PfjdQdgH5Bha0fUwOFTIB0pQx
OmgbvWPgT3vlkvf4LqRncOP1Cx6cRa0bLKEcmkp5OW9uGNAPMoNN5fa5FwS8Q0fqDBds5OKfMGU9
nbvHc3hOspttDJ3ihOIF7cBOU2hYNVjA6/OqA/kuuxINWNk949rwtFZ/mi5kinOGgeS/cNf8EGOs
kzdwbrZbv0G48ANuu1TjG8dnWoYz4fUXJqiWMZwb60HfA4tscj9735EQGvlDc6UctMJYJnY/Iha+
kT2n4JNbEvGhq5rnRGl0ZjSATx6L5Am9ZC/1VTZxqg9DudX24/9asFmhl8ijZBPE33D6qhiqd8lg
oSAJU+jGRzPF88jEVD9DXRVGp3edmHddrvawYXieQy/T4gDnCyJ1Y9fea2icPvO1aJJsNxay2qOG
cPb8xH7EElPmI0q9EFJLCVg8bsZWDd8qX941wP4YjZpVbCcidW4b/UNdpnUc3CUd+/NfS/1XT3fk
en4XFS6Vbyt8PiYe+Y0BX9MXVOVXh7haP7qIePUO4Nh1B0aFzwfLMaF61cjwF3B5whmzxZFcs3EL
5H2VINeoZf51iTFaY5NPlBIjx+w4vECSvyFvN81Zuc/3wdFRnztM44ABneMqC+UYV1Q34SgTGHza
TOkd3pY3On48b5OGBYZc/OyUQhcsS7M+Fls9pQ+xLxLCy5xP3gr6f5AskIEPcCcEGLy41jQnM3RS
yG6lnloGqwwgvof7h58v0nloRMW4C5nLAQfElVsKrRBaFaL+VCOrAocaf6kFU3oZSGD2+QPmqNbQ
q7RC5VBmKy/lXHSuAmUwe5ysUaNqZOlH87CXStBZeUWIBuG9zWmxPxL+tebebmWz0KBAtlehmYOp
BJ43W+fKBUj/qsoVJYDXLS33ynNKwaMDdks9CqZbNB6HqKFUDOg67t+LD5gfBVJ90nA7ouW+LRTP
Ihz3sYOU8lpgSSMdyGYXm2Me3QooQ2RqELzJstIRycjr+THIxfQUGTkQl8LMLTkG9TNpDMHZqL/u
7wrUhq5AVvt0PUz2n8MaJQfOoeiOK2mgwhalxJyPBuGqAkRUn5O4DR9m+YstSPRJBrVywdEgUils
ALZTWnv5xJXCzJtlBt9YpJtObX/6JuKKm6PuwpFKt1sWBxrd111rX6DRSwHb79jPCjoKuIvvvoPY
ThM/wc1dcI6ZVmdYwkhCRQqjPm3Pi/yEuO3JzTJ9sLuUyd+eBdzs1jpwsee4zWQ3WdI1ULC8mVEQ
XCBF7ltlB8raO2lRaXgcWvYiAi8fKp4SMQhY7E4zh6EFxjbHhTqIR4Qk1ni+EBElGtrlrXM8hQtK
Jn24D/h1x+PnQyXLCYJijpk7XODb7QaHXJfBVAa1FZ9p0Us1u+g88X3+JZhk2lgAnoWozPpz8uxO
ZuQsG0IazdpM+OAZk/ptPVXkyIoJJAYkcTkIBPnONa0+XWATuqrgHSd3wol/6OguqC9LJw6p7i6s
tMcAjE5V4LKRD6Pr4aziI4SNVvLK+uE87PLVZxWqZM0G/XXT3qahlABLw7AHBa8kydIy9VDjsS8b
/pGPO8dj52RiQbEHXvOJorBnPCy7gMnrwzvXxR9peoMbFuSSdNZYkNx5EURb2X4y5QpYs0ClQtP4
WxMOQxBfx88x8ao+EmsqF2PqOG8iFAUACOLkurjKOUh2AeSg4z/t1fwGxDtzwAczQwtlGqx5DhWa
bGndYdO12hhEO4w4RKpelPD1GTyOy4js2b3oBzTCvag67fZJQCcXuJHcZTOt1oNzgLURZvfLRyqm
0K6SU3VHpqxOZxOSZ4YKkHJu9auOFyMmYTrbE9s+2FJeoeTWRX3RCZl2sSOOfZ3NvHc67NVCU2WR
ThIXdeIDCnWzqHV8IwH3r/cQt1ejWfor4vrR0xJ+MDROFUTCI3MvowfTFMl1Cwu6f0ptHmrx/WHS
mP58EzCnhW65CN4xeir/bI/O/wFZBUeG9AHL3p8Ys1eJvt9n9DkSNiuHKSV9EQ69AdPEHt5w/zwZ
1+87WD7aj0C9y90fEt0f1VjpLjfodn/AtdUfZs2nPBTr5/GaLm2VbuE4UNRpmZVGxerxC2fs2IwQ
sfgnlcK0s6WR/RAPlNDP112bIRT7ldyBH7+3mWJrg0P4isKp0WoRWs4jYIDtLRrqrdbNCxmf3xgT
sTgAMnt64It5vqDPyYRfbWUfvm+xneBL5e1RpWPnsoCFr9UuTPMQcD4eIQtUo/13D336KoJ0wgR3
W8ydufWC7XXUFRE2QSlqORBpWxWuNPR2tv57QuLiuJFdjN+RNZRuET3qTDVQojGxCZdO3mqjK0iY
fksDthRvPjFZ/F0xV23UPiaZpTlbk93SzlEdQfH6jDOIFLpFmBdOSkEIsz0t1JEzU+6cbU145PIB
JjEwR61JufGearDbbt4bdrJM1ndGPzy44HYn9qHEg1tJaYTbhjUimrh9zxzbfs4j8MpBrEKUx3R6
CmeeGymXlfJImjAh4mqSb56eQv8+XLD9/r1ea0PTY6ZxhI0jJ/zmxq4/oozdMSyUDaG7aBUyJhI7
Th6VCa/VLAeAg3Lf77SYrc1O/lPOu9OaHkYgwlHw+kiOa38cTXQnpNcZxthERdACdLQ6nUVvtmZz
8Q31GPuWZwEOGTN5W1XcTrYdbdXkBgCjSrmoJjgdf2gTbv7EvAcsWhy1POVmrrNt5mbsEteIGDrX
gSK2LjrHNBplp3WPmcefr2wzBd49SyAOrkO+I7EWwJUMelYb94o5WGStJB+Pr85+8zdqr40JP/5t
11zTDqwy3mC61kf5qCp7Xi1mcOEtKm4UhYRKp35DpBlnLFMxKrV8Jw65vUackwgoCuKyFpNOaLU0
3KKKKJpr2knrs16As9RBVEFmMo13WsoH50dhThKr5kF5NF1wuSOPCC9UGabpRBhHOWUCPnNjVilJ
ce9k3EMKerRvJwaN8sW+TzY2gXhCabLpLebKk5/VKNlOsJYUkw8rbzoX4kKJu3OIFEYkqpYeLqg4
Ldp2Yr1c8v7ZNevBUczHwt/ItssVeHIY1JL4f6huph3jMntSp/UkdRDjDnk77wc5hZkQbEy5PvOJ
nh/DQmQ80dCf+oIJq/XlMbvN4b4HxNbt2xOvnYEN2ZM2kS+VkEfJXx2omdFLVSxw21rj/D/My76K
a1tp/hdnWkVmhavRQQcsDLqFsgSVWND54eo9LoOwf9fyKgOHWxb1pOe+8geZZ1QCepSgEMw/thYu
50s8CTzpdqtCrfUtQ5lvcEbkZNtL8jZ5EHe56WbUHjH9Xnj5YjDQbS7eKGBuxeOPrF1LWR20EYnl
IdYHAao83sMF14rcbRW9fKH30SjGcTzZKTaeBDK2qo6FxNdvWqNQRHiPtTeNpMBys+N1DoB4h/0n
u3d8Gx986Y28uDh9lnr0nmMkTlJoAdBwEhR/soDKfeMt1hNrulcHe7i9cwBusDNbLUg4z8CUdClB
beC9JpdU+ofDgSuO1+EtYd4+YM8NpIRKAskHSR/TPEAe6l68YFZuNfuioQejc16R0iw6P4mNc6kO
lC+/RDV1IS3R3MT5bUbKfmXfwgGgiK4HrHRcR8671Gr48Wyf3qe0Zcjevig50Oni2mqyM0xuf9DH
i3Se+Ykim679VqrvCXRHG6Sw4sveGnKLzkyenVyCP1Nqp+3ko78forYvspm28VkWjaH0TFml1JB/
a2dRlXIWdvRKKzjUp0pUID2R+uKawJbBGGftCSDje8Jx5vv0RjBucuOcA52zdg2rXHSpSEp+KiOM
6+koI9RToLR8yAWEXLGqaoyMOYr3AqOGJPIba6+Q1Kixn2aOiRVhAHwrYsKWW42PMORX+Xw4/K6O
pmQerRD1B3tTD9H017F6x3eIAG9uUooAPyF3XsPKRzShP1H30V1xeFN85m8j6QRujrRF44P04kAP
Izf0IfEYCcKAXvWPl6jpJky0VKMKG2cNetapUrDPkl/sa/ljY3qN5N4bjdkbad09+Ou9e3uSFPci
nXzfOUqTZodgYXe9oa6WBiXZf/SR5IYL3uzOZoNxvfdVFvK0/7Haic7xDQwonztKo+BcQFPq6LC4
kFYEn96j8XU4imN7I7a5Iyj88RKdVzYdbTAYCK8GNMP70ruvWATilqWdpEOoKIUfJ3E1ArN4m1HM
lTxyHsiyrkb2IJ8ZRvR9J2f6DUF4oLxSrRxMkVTyp4yVrIEkaEJf5hO7NeFRyTUJLbVLUCQQxJoj
MB1WW8kgjSNMZHGSqbAbOGd7/bKoE/UrqyqdSPk50WWO89e8apM55Z+uBPrHvjrjm/1TOdQc8ueL
fumbYWMS0l6eU7+kVN6b3GwXMAXSddLQ7aE4aMNv/GIvEGwMxOd7p/b2vCSrMvTaayQCVDIM6xCy
avVsW1O98IupJ/QBofEeopFW/6EuYkOBQjnmzd6IAcx3Mt5k3pB7Lym2WolRoXiJz3dEkRRloiWu
2EfIvfewIxU9raw6D4bK+v/juKgDr9O0VGhQheAkexk+L9Ll1QzsXjDYUUCtCaBkA+W1iJaXJOtX
dr0N2EL0MiDO0biGh2eLabi/J4jnPH1onwakF13IqxsQvbOsd26s15dAWFPqztCryPNyMsWOLSIL
kme4jFm66EsHAFa4pck8ty1l2Gvr9RioNtE8RAeMtpIhbQ0sS/zesEHItTVM1kRuKte3oQMdlRM5
NlldjVpD/BC6JZZBPlwFhFhzIfScJTaYqabY96EAxP18seLxqAjU99Pf7KX9tYihgwO68Yxh7+b7
pPUH6jlbFd2yC0DYV8M+miX7vQOVNj32bAfBAD8cTuHiA+2e5kT8glTglbQbFTU74jm4lnePk4I1
zwD+fxxIJjmEZy47CL4DQTvfIcMdO0tI5uvqZJmv7jI7IBrYbTqDKQIXV6qh5LufwqWOEForJrhg
Quvz6qAHoj/2fx+6B23iqahz1GuelsV/DMZHx/nehvpTW3e/0oUFHDGC5GKHOm8PSuPrcOEdpXhS
iebEwINsnZW1mtdwJHeDZ3EWYlyeDmJVxU/xzHwx3prQBCdmiwz1YrUIJ67VIwuYyMS+ZOs1F4TT
/ndc2fSNzIMJIQmbj2vsSXWnooygW8HcpZOpXckjrLEp3E4wdThR/wZbk+dcy9fxTwT0zbwhltXY
cJnMrGXNBV3/KsDUjKlHGG32EuE8573GzdR0F5rM7MuYOVGgix2xlJ41SODs5UrObJ+M8nm0hml8
vsQDsf74rqN0BzV+71V51n5pXL0r987RxTK4YXdgiz1ODW0z7PQPk+ItAF3pXQiCBJ7/ekApv8MG
LSnUX/jyfVEd9zwl2Qt97vs5s9knd6oN1+PwkPv7714sXRdQ83ekhjKNHjiD5ngW5SJRMvM1zljY
JbRVFc0J+q0y2BXas8Nybu9K5hXrzfUupR23mrKSMDZ2ILX+8LaXhGXmbk0incx/fP9B2MH/i8M3
nCDz68gFhFOAWD1hLhK3dHUgtq5X9nHDijYkFlhPAuh20n2r1OZJo5BfU36s2xU8Ua5NErUA0c9e
jfig6e1TeneBaHKTVYoc4m5sQN23A8LF9O3v2AZvB+j3ufOB2HzOrhbURmFU1Y3zDBGTfWIiPVkm
BkpAqVpaKwocSX2e6Y9UAJIYRq4qwuL9f/FmCS1Z3g8/vVT6BBW0AitvVVYDO1t2xQWcengMuAT/
f83y0wkJVK7K1eYAkUSiie9nL9LQkSV9SenZOVfT/LDbkaypZyYpRYfaybIKtWV1mtMU25euEDo5
uBmi9qsKD2Bh6hRZQ0QHL2074n4lMa5UUKrZxvhLPQWA7D6PuV4gQN7wWWhIUW8Ym+B8V5za3Ezw
PuHlTANcfafDB8XJJgPzoVsiQBkgeatVbRSAngqpB7w9UuOwJlemx84R7IYpaENFNLbc6WS7L9bd
nh7Au/xHN8NEDnaAvsslG5Yz9MV5z6MFIQTgfMkNBSZ4rY7ISeM38sFN5GZiLzq2cSCfJwyQakQo
8Mofg3Kroy4102uFdfVi5YRdA0vP2IzVQNjcYDTPFvu80LxSkfXSLfAjZglbx477j6qTRZootF7w
72fJFI4jf2IXr6pOk7PNyNjz0g5EIvp2YRsSYiCd6Pv0RrR1buC/MhOyeBRl4NkuWKzyy/AOCHCi
7suy+yJuMxxD/VkRgf20Mx3RRxDNxo6+4N5CXv8maFhzbdKLdKwqIgWgCl+jYds6KiXTw14fR3vJ
LBxNCWO0Fdff4q0QlaDIxhI2/79pDWuSF8LECtsccv4w290Po5nfU0lKaTar0Qpd8mvaBoNScAku
efIXQ/MmiDv8vsitLjw+NRP4nabLZ3AQRR990zp44ASvCzgDWO0HhN28+p13D4xmtQxk63RCiVGY
3SU8bUCQ0ALFJg087lSTHU0dKFDzX2+5gDURRo1gqpDfmOp9fJChLwUJjp2WVBucqYjhhA/Alk4C
RroqNGLtCSstrgbldlSfjSjupi5zK78phmQL2Nm6ibHb1n72G7gUJgFQbYb45u1YGYVHLkoem1SB
IG6ZPIzSmOiTZ/I8H7kLmKawHpbxtRrt/Z1qSB34VGSUrX42kXf68lIpnPpj1h5XpLNBH56HDFUH
Jtr/Xkj8dUxxWMfO6Bhu/bvJiiHf0Bzyn+FtPBp7Lq+HTzfqcJoCZkE6YKR756yPXd0Q7kGqMzF8
uMSvprmqTH0c5LE+CigMdSB92i9ssw+bfc2F3pzMr9MgMqU51zPkdu3+byhfE7Ad62THEC7ttYk0
Llixj4eEFadHWAWPdBBgaqRiRAjM1FXVswlbZTa5cnzw1WvVAagkJC7SvOyw1CsD/9wpkjTP1sNx
0bBfI1g6sf9tpSXNwyNX9gju0XciM/yIf4Y6U6W60d5w5JAdE4S0lVZgja+S7c/cUlfDSIQ8AOgi
qydYex2APLn3gYIvw0CIN+jaDQArvT7Q1D6MOjMxGSeMomT7JxoeMHBtSG9nXF5EOVAIq9kTHCJL
E8Eie+QRtQE1TB1gh5ztRta6DuMtU6ytKidiq3BJksfFA30r5nTxoIADDTKD5uumCUsRdW0ejent
dwOMghhTtJxBvccbbQ7OK7toarjU7aaK+RZ+v0ir5Oln/WNEHR05poIN/bYzQz1driQ8w5Jujltp
L5+CsO7HMZWZsNmfs2tBM7bvZqg5SKMYlismZnIyaNq6zNgK3uf4Z9UiKcml8BbvMlq4nYX+YbC4
Fap8b9qIucbNagGhAOR5EnVBOFV5GLiRl2Ngh3EzFXBgf/HNxmjYxcXkZuR1Cjl6urOn6nSYpEB0
fbfdC/Jzeffi7ohf6L+TOXMqjhva/ohneTlCTPICyteJ9dcy+a6oLDJPElX8+Mo1rTlanZS6BFe0
ghZBcFKZbfnHdYOW27ov2ActbnJHJR5B4OWJ2Hmko8pQr/sN4vYOFiWXfKT5TFdVEtuRE6K630Y1
ecgXP+GanA5eV5ahOxkIkhYdUhrAwv4pyQiwXP9MGl9dw9Tam28bSs03acf4u44ERptgVIT/nYcC
pPJA8VsmzDjDsU5998/jW9gNRLzW1p+hsgnzHafVS0NQ8RRUMJRo3tVf1cSreUg9iK4c93Gqy/AV
VcjEAfSx/MEda8iQey6O6bI1xezSAZ1mu9wVrwdZA9mWeCmqYT7DdS1aZsxRcZ47GonQ+WIdo/uV
Rv6Afw4VFX1Hj73ooQ/aA1zrzU5cvzjmYcr2J8Z6zGOhFARiAk5OZgvMCkrfb49rVAX2UHyjtGlg
eTIwyZ28nsKKJVur8hhS57686ee28fwUbV0gIOaIpKf6XfGZ/L4OzJJblSUwjIaLS+6gP0xBeC2o
mdEDlx1sTsYWHH8BgZEh5R1lPMim8dkbyWmcJzHYe6wS/iW5KfejQsyM/Sxl6Pl77EB5c6a93/Bw
NuPeKverGDNeMQYmn2V4oWFznl4ksmM/rTK2vq6G461zSLhuDlV4rHLQAMZnN0pfoqLMmZUJvYbb
kli8Vr3/cXTw8jviqQEB4orChoLQ8slBhckW/XOSyviLR3LTsYojZHWyBpEjYVCYAATp5/tcvRt8
Z5GMtwdVlS6vFJEc+a1nHJg9G+bKJiC+X+tO2cQQyKKqgsrQ7789XvZEDxGOoDZ4yzUAgmXd1OZ1
pbdtSAhYrxXYh8d7ZUniL4N7nA0LQ4H71NHlZXKlPjQq0EYNtODUChu7LF/fEEUxOcvOxo4BD96G
EtDP38VSH0rEOuBlBQClti2jJv2yO/+YGRPY54ChOUB4J8iepao9JPHydp65YKI1aoTHaVTXHCVR
q2InY+XXiydWkZ8HhY5dWCxo7Jvw7wDtPCRtw20U2rAoN3X/RVrALI0oU/8ojvYCwTJ3cOcP7jUY
yT09OYEiztutnHJ4ZuV0APHieAVqWyo6bsPlTBzh/LyobY5LvZaokPCP7Dr0XI2TWKZaVZwk2/Y/
0s1uW/G0KkB1lCYOLbqMF+dMgrMC65KCeJc00OUrOtSrfhVli+Qmxhqu1As/SpmJksGRBtfpqWil
941+84U89A0YO1yFQUUIDAngvrCmIFHEIr+ZcsuvOdug29kz1pzdDx6SxtLj4uwoLuOFv/DTO2D3
VbL0mwB1xPsNLU+hK5ezO5GLJZ8dLgeIIw/IALtx3bOtRX6PknshkgYE+6AAdkbwoWrxvYw2mhp9
NA57jjZ48oGhxQtSFpnBNhEEgtE3599C2uNSKduk4kEJP/fDIf9vbhSjnP6wAIozU4y5JdrE40Ud
48MK/LuhKhBXlsCjMd/pyEC6sVkSyvKGXHtvjkq4Ky+qBnqhxr0OyX+VHLVRrblrSnQ6RegrCaaW
t7m+DfcZU2n1Oo2N1+D8aqu28y/9RVXInE7WxO/MIrxptJYiWD/ecgwo+bJpj3s/nk5vGJhMsXUc
ZKVS8xE9uZoiAHVzmWuJb73BhoIyGpe7rF9m6UUMbPv+nywk2UkfHVfU5hsYOLQaAt2tw1Ln139Y
L5w0ESZwvSy3YxhJyZE86mCGV0YH9LS47zpS/7lVPGi9TNEFtu0Tr/ppfTUl5RvtoG/+YmE3GFd2
4Y8dq+kwFL8CsLO0FJWDybu9Mv0u1FVtpfCtMxNROR+evgcEFDk7GkCTaJ1jRB/yeldGWe2nA6Lq
3mPIgKJlavwBpM6qnNeCzmMQ8pZO3nfWz31lccCRsozKD/f6zo2NrmeKjOQe1la/gDwBP/V2hf4m
RbnAwkJUG9paK7KdE7EiHH0K1wIjHkm/Pkigau/STFxrV9xkisIjRT/hbolWJo7FIkndkpfBtGEN
jm5Tj5n31FiSGLOMRqT08MlkC4tV3qQGVqWQC6iS+xuaW5mjMNt6zD3upaBaTzxNIjUW3EqLqqjE
rdtZwZL5bpYtEG0S5xZm3+nmhF3d2W7aasCv7BFasPRJp1zuZOnE5rxo/lhVpOmoOh1ou5fvgLPd
W0e04VHjH/GAWlhBvyT4kb3lsFlKAV0ELOd7eHcXJ+fbQ7954JRoyX68KvR43nJtC/AjpnHLwDno
WRA4QaEv1/F5SqcZfc9OJl8yv/ofiRqlEXPrF2lzRgtBRR5Lu+BMGpjfTm/hRDuQ5X0Mgw4/46Z1
59cSrJsSJ8MakPd8EsxKFKEaihDc5hwlzqzvydq9k/FsDGRq7xqt0DGmXns3lA19Es5CpbYLN8HC
iqYWMkXPdSdRNX54Kht773oLuC45D4PeoNCQIg4qp5C7nKbVEJa6B75Rdzv8OTaNB44QpX11uhI8
2a3XiMqd5cad8LpIffl3B5PBSSDbPhotClshXrLgSVdDuX4PfkSn6TTBIB2jPV6xeTMu6421guyN
5E3KNlVPiS96femV743edd5j0FHXo2NKj29D2P+ZFbNIceUAYzFCLtMNVeYS0fiGNV7eDc7cmbwX
qbibJe7BlG/1vj3KImioEYPnYAlqulPtjLulPVGGFriFAhew7D16FLlQCoZe05Ox9coYeeKpoD9R
eZcf5lOr5+KMpU96+2cbAY2hR7upkd/qRIZg59+VLKHgfvIHwULCaJJA1pg9avKVLXZmvlNIhNOW
8p22F1deIVIRrdv49HrtZ6NanPfAdELscEgf3r7+5Y8EDte1yTNR3Aa5fJdjpnhF+QHom9K46RMF
k3xLCDvAvIf4iawBqAlSPZOgvPb7s2mflXR+KrtS2ynMh4NxrPqeL+LpNCgs3lK/jVHt0AB5vEuz
pfWP8ogVwkm4yCqS+dgHhSPr6ZacKx8ZIe6uW789ykWc8DbjEObUsJGX5CA5EGTGTAHbM9x1T0Pu
qwlq7NrL56iYd2FSxCzeD8IfU8vj6ErkbKnR0Jg8oXkX6s2dk3Q9EfWdXWhUkvjYFJnxPGLj2m4E
LcYL2ofrwvSVxFYg3Js1ZUU+h4rhQ4T4ZOcJ9pb5Usx7qiCVdv1PONindIzWulCMQVlH3kPzmXRi
pTgAO0ffYwZyfcumMMPJjXUrnDWeFo4GdinvTa77Ro2bHoCp6/N1Q5QQ+12yPxSfX3cBKZQfxkJ4
DyspEZ1vC7um0Fj7vGJwV3i/mcou7hZdaqtMvPexeuYDa8R80dHcCHmwg5J1KICEjQQ4M2PJ6hde
vVmWkwGl7a7swopU6mF4UWbhMsRYl/4rg699IjMctJPhu6rYXUVESg9Rl9Hksc+iGW6Sby09f4pW
saExsyj63X2mHSVTbSF1CxST7eelP3YwUU2Jhba431LsQRjHpOCHotjWSjym47WL2tPZAz00BSyu
42R4rurpNQ1SVzr3k1w/LZ/tP2IzNJO1aoeVw63vpg5FLEWeW8QL0ygfte+IHLgB7+N70uPlM2oe
le0FEBPo0jR9sVOOWCvZnSW9SRcjLwieYZ/gC0WoCRfQuiXyeOWnVPqDRm/9WzRQ5UgqMHq6kgiD
35LXwU5cNc3T+AOgEQ5zeikH583+SbmrvyZVeObj9LaQlaj34EmxsyxWgFpoBBGL79a7w0YreqzU
atRqWR8/qADMcOeZwORqFa/1pn0Bx4OdQ5z+T6mO3g5BFXgQmCKkYIQ4XAmWKJErbs/Ef06KhQZ1
59GXBTIFOCs7QcDm/i+y+yQVGdvFDrXyFD/PZQBjKHK3//DoW+4qFtDWLbYyQ8r/dMwfCMusiwn7
Qz8H56CGUNM0LvKO4jW+s+G3cldyF7sajYVQkj3eZ3BW1RyQ5/wA0nYcEWgpkoeROn1xKxuAZUR1
JT4/ggaO6q+YAUaQdc92n/O0n7ciw2+ZWLTEWvEv25tyz3AFy+Xs/izMFfmgsxhJzau4fYD2eD+S
jHRppNAfWH6A/bfseo89NHKaqrwCPqZdh3Z/CUp60V1U9ydI9Ul/JK2lYscA2ZF0QA26PS8KVQqY
/Y5aYmKCoo8zKLTrwh7PHBTgb6cBZTUyAPJGv0AHgxtsArHLr+I/taFQgzgBfJ1ELOQ6u7wGJk2l
o/liAgvZDfiROl16DYq3Cyk+8T4s/H/sABYwznbCWW5ZuOptgd58mmk5XFi1CIwxw+ZryqaSsOGE
57iSUEk8cX9ybIHevkKaTdAXCW9oOpbDbaoo244V2Twou+SGwZYikAP2zdmNjiBUqL/T114kXgth
ELuLDiD0VtEEXES+eJBu65VZXTLs7wWylRViIJ0FrTNcsH3M/i/bHPmtTtOf2iY0QIc/f4ZZhEIA
77J31/QUNFeUYjgkvZnxkEPIcGLdjwHXyLLOaA9zWBbfAFLt/GRva0HJnWlPBZbjuwdyehG5TMz4
vPU775A86G0D27e/YYEzYy49cbunmziEemIXvTHsgC3owiVyvOZ6hD6XM0Z2Bw0ZLgzfBkutiaJQ
6gjGzcxhxgKl2UiIfJO9Ztzt9V9FuqFlNsnkY4fMOqyvC4qBwlwjaQMJgJgvhdo9r9dIDP0VFzai
ATod0nQp3WzkM5rN/djYqdnfYWHD5U2ZGRCCcoazWMHof6pNMskJj9SamCXbR4iqcI5tG2bQG2KM
gcVpRBtgei2c7Iurppkr61R1sy/s+6BkKROM8xFi7mucp7sCe5uMDWWjlompqjXaNYKwo2CPXqZs
/x/Iil6Buf0w8N4ylIgQPxhIK2bKRbRwAway822GHlFTLpCxzYFfZAqDDgPTKAz9S/X1upnH98nW
AcCU8BzGyvjVaboB5GRy+yuInN9o67jAStGMWkl69m7pMPbXfIbZvjwZi0ACZWYhJH7Uvm8sLxw8
x+yuPHSLiggWMq4nW4243yg/QRvIAQuE/vamObZevJmEXUpDLWgxKPlUNeo8vzfdMqDu7wSsCdsB
30NAXQ/5sXa4CtlndO0KK/1NBq0Li5+TNTfRPtg9abjeAkZsZxA8Jz2vmGZ2peqzO8OFXNOiwowW
5GgzkhTRzk0XF1XU3wKZXJxkdHwfLts7pRfp/CQdCjaXs7F13TLg/MTQreiCT5/aZWHUc42q/EXa
DyIfgSdogRc1rTh5Mf6EpJunRDSrLfbEW3nUwZf52e6BpWm2+Lcd1uajWEnRj9q+LFj3Mkwylzuu
LOtDxdgWu+BKLskrGWDKLW0/zltu9Mg8hWLTQFtH4faSTbXM4rh/gLDWpiKhB9rXL3Y5TyTQi/Tw
Uvk0CXqz4zwSFBuCCIVVVkn43bAQCG9vZWC0m16JvHZcDkTE1SqAKy34O7eVCxJOQNi/sAfj0sg/
PfSDisVEHJJIAstmtOocZC+TesAji3lcsH9ibTyH9+kzr1cw4LuzB9w13uFpR1GEZUJsfeArO0IU
7AX/N88fmocSt3ickWwXZdbpPBUeM/IkHoSHkSmlWVPu03CGYm7SSjrvvxINZ8uEiDGLzZfQlb6Q
PR1FssKufLD1dCX6NIwslz5uWlaPjvdm3XeHAd4qMM7SqLC8HUODgGwQLnP/XYPEk/XZDbAhCKlH
Mlq6l8iewW6sU3kO30U2JCQytR1VMgVeDag9LuEWPemaecVggvMhyiyDM8gO0QCF/JujaAIPhqaG
0G9O85cCZ+fjQgIbqAXG9eLE0q40Ko8rCl+hwA3LDu24coQDbmKNN1kZJ0/uJHT0mJAhPdpGh9He
XsRS6s4rNL8T9qH55vpVe+qoYE2YvObEp4hY2V2kyFWbYX0laQNRYIfUN3BYiMbjcu6VbZ9DV7jF
/Z/S/PGZB32EX7+dtwApo3uOpYcb2qTEh14s8XnNs/ovh6x6VqwepL9uQQ9KzWn3HuCAA/yCjcSF
YSoiAHaprRHSbzWe9slmTgkssnFJMpM7/tThm5cD8/I0GIjLYkPFtqUAkAs3laDMhB61PDJcecbY
wfFhe5J5ArlpWbsVayJzCfvhKCOkFCeMgEPZevuKIIkN4auwlKJK7ZEE64EHhr0N7nCa7DDHVvwz
02nNIGTNhTt3NopoFPIc21QaEzwFsIeoF8NRsRNpk+wiPt1ukkQRUhG8TD/zSv/71vTFx1hxlQVk
dLKEnPi7MyuETFy2Tc+RElmIV1tky91CtjTpq5k7rkDIKlKEcA+yZq1hroFLvmAL6rWD3AxKYCDq
rZ6FVmxJZpduxB/n+SO2t9hbSQKGVSFljz6cUHPNzWsVchCIHzLIUgUUkj3N40XwOmlwWAfT380Z
21K4qRHZsTMnbDwtn8Pna3seXrZAoGri0ZxBRBQK32ga1pd7to+rk7v08E5JKzUHNBnzLUcEZ8aX
WErCQf44Ka9zKUEU7aVEqd7wnxZuzV0JO8ExUNN+yufP2HxNgFj+uAh4oxE/WzLGxCyYiIpHm6zH
YByt+8ro4e07CbR1RKwVEZW/vqJXp6UOZKnCqvmLkZHrD9AH+r8pH64ffvSJ7Lu+ttyR3aXUR50L
Dl4JEVvJ2naKV4D2qLGKMbw/82pEFii05O1F0ohGuc0P7kROvkMnaUPjljdhhldU5EgNuGcIyJ2s
d3Cw3F6qYu9H11q5K1oCt/wA4BsnElns+jmZl2LmgTjtYTXbesP2bXjWesYucNW38/RtVKagEjSu
uclNgXn5km4SBikKJF8ZGASijs7xB/Zdt7TLI7R4a6lJ16AOx1+xZJ3+TCH+rRrM6FgAVPEyNzEo
ZtXestjMxic7cJOjpxMgjgAFXYtT6KnF5uonesr9Z4mRCxNLLUuOYksFqY9Q5EpH9hqb/2TsvODf
l1Hx+1gUL8R0unsuxBdd0C1VcIq7QSQvr3u2b0IryGEqzgnQim+xvUX7QVMCMEdoayigkOPnuu+u
EMOb+mzzn3wDBMl35iewhPpmQQX/pH+74+aEr0r690DoKWxQCZ8Krb4C8TjLrQkA6csOa3ST0fgl
tyqExufStGa5GY3ymLLrFxJN16HKd2e4MtH3gjQsyIq4PYsZp4cMMytdbfmA7FWXMFb3+9Lbmfu7
e0bzT6JcN3CwlxSYXdLX2b6YU663SKGwlL/gfwNl8mM2WRaRaeunJCaYE7GGWWr5TKx1X1uGs1kM
f2qSdJDPKSw2UrolTe+0DDdlTgxz91lI114KIKJ3vU6g2l1pRHSf7fK8bsGBB1CNDUghpdlTAhBq
gNTQEoTghSHTWdi4f8hYYsRD5v/hMkph505opZC4teHS7g7GYcFgmKiGmQzKWo9mHZOzuTvFfaTS
9N9yi1Ls0UJkYTF8dnZC35VQzIhj0O3hCpt/ZAYCzjk0RIrjoz0tcv1TRywCu2sFywNC7sKP6HBn
xJHoHiysK+YJjOukOrPgajfYQ27hdi2v1qWFE5ZMFRBjURW4v0krikWx495GxWLdYumFP9Psq395
lmE3Kk7o1PKqRPIPF/rGqlqCfud8EePt3wnBMq4LNXjtJ7eZKZesUaPL6T0wu23gcH7IP6sp9gnr
WcLicEDYtVMuO1sRybJ7n/tH9iL5GOQLGssoL1qZdRSl479Iy86uI8fCdLQPdqZ3HhO6mCsHwJ2p
YjtS/zfhdw5lc1ivcVLTQvm+dIfzQjB124p3uPz0YB9QyCFh2sX5dR8yjKswTEq5v6O3t7qYKbhq
eQ+WK6KM2DmFZNsypsIHEmUlOH2EZi/3Lh/0kB2AyGHWh4SDpV2b2rNQHtPzz+pQAh/OVJUu6WKy
zbIgczRreV5E5/42zhzD+UmUEv2s8Vyo6/iu1KP+1N7X9ElloA/d3PX8+fxqn5nLKXIZcWjn0dNl
0ybiYd3vRtjZikN8m6Kq6ZJ28PcSzxf/CTJVdNJUghxGLSLll6cVY9J8RKI77+WX5xyEeMTii1kN
EtNsXBnr3MLoU7asfjRiYvzJ+tVEpVtNZ6YZulfwKJunEYYlB78UatDktkc1ayNOQXgxwj8E5BKa
2mHR5/LnM5sBMC9OzmR64KavCuxuH9Pn0FICALIvmwi5Uij3mwfcuzNFQOQKfVeizdn82F65cEQq
6bOjbzYJgHXSeh1eNcwC7zHhTBcfy8Sph+D9uYCTqaBJwZwpYY+g/1tCEhad8DrIHmfBdbbBPX9s
KiQDqae/qS8ghX+NT7f0jJj69aw+VjB72ZFdc47jISkyq1FhHnjff2LH7KCWYuHasIf39IVhAyPM
4M1y/d4bgmq2UtD2O25XXdgY1FwdCIdHja9rH1z6TQrbF16O0J8SJ+gTkQEPMebB5A8vEyE9w5Ls
a8MD340lkH1WQknbdhe72Fk2QoP4ae03AGsk/uDu6bG5bg6epVq8Q3bDfvwNm7QoAN1StDN/TG3s
ejwGBNSCAONgfcgVub7bvhM6npf9VXUzBeubzOPcVjc3www8ZJ3BViN+hKe+n6WgBWjQCPobr36n
kdzzb2HHliuTuESXfTz4vtxFHRIe2y/i+TCaM+3XMefE05A+DwPaJuMDj5ZTZgF8AULj8bqGnG9Q
SdG9SDbvCm28gqpxB7fUOeN4LKk6fgG3kfb1VxkYyatb6053XwVnZBYw0QZ0yGPN3fvSHZQvCpvq
jq+C4zMoHqlxXOoKALsyVcHz3eOGBCk+A/58EHYte5zpCgulSqCh2QTAl3yHYNZVQ4j2+cwhhi1Y
e8X1sSFvK1dWq4oqhAWPrUfxoEZcU1Kd01upOr5sQUs4sp4+E4RnhW8SGbPcIIFskScWBKUGZNQn
bvUF5jbV/P0xtW2PAtwn5oac3jfqTH9Xj5QJ9B5SwPR1oDk7Fh/gxtlFcHrXJfX5eUVH8vjt+Eu2
4JtTlBCR4CUYxiFdOZiyW2FgM47TPm26BuFvdumTNA5wQhuJSI8q4oFJ5+yBJsajvzYlNgQDRaYV
g20dY5peyU1r8zwfSglYf25sDI8Z/om86vU4f52e8E39Olw23pRxTbztvlOA6xR/ODbMEXfe0ffy
UxqpcR+Kg5aiZ6gcafS4eedzl/TtNwRBl/9+Q9ERTfMvZ4yKQCOqXDHL8hSzFlgfpfL1fuwVv3Dy
ivH+UVMhHU4FrBowD1XJiMvIS32faN9/LNxNp+JXIGm64sJLGIcJCg2dqTJ1SVyvIvH+H8Ivbczp
R7Dr2YPULZwL4ZDB+Y1ePNuJBkGZAGTCo1Goh+lKfVOhQR2rkYPgdIW0SOkpncq2WYP3/6o03pll
vgWeQUzwUd2OMHWQ/jwXwogp5FKgsvscsYLxAep6UlDAOce7eJTQz6AIXPab4yT7XuIDK6XAsMwH
yHLo33aJmf21dd5Cuh4bt2kfAPRRlXZlxN11HFCcOZFzXDudZLBLB2yTT1X7R2kmQglksKVBC+HP
GeAf+GXB/DDxXRqGGBUvco9a0b8z0q778W89G90fsSTTGuJbI3snWQagX06rD7S0WQ0opYf+iZE6
71CQXcEFaiJdXFh6wD050i8luePJut8DcVathhlv7kZelVvKHpHwmIq1U89CpTQClqOD+tzj7xK0
dIcVanAlsVcpy7Z/wOGJzA4D23fnZvt6HdIn/KQD9iDu9fxCqVZnIV7AvtX1X00fygyLFbzj2ur1
7Qkl9iTsguUqp7cbBIvNbaAgs++3uTE5BQRndYZj0+Mz4C0W7E50g6phAOHSG2Q5UcA7Ta4IgEVh
HTqCLbUCoQ1SjUcHi+vv6lMVd/NooiZqji9ET4YPbVwYe2wjPDDtqso1fj2/pKG0VvfV+859tHCn
Nbc2Skj0vcMSbTjBRUi6hsHRVRmzaYPqPjbsJXVgbUXaUNRU3SF51qtkueDUWMzsv2JpZC1+bBzN
F7XGd+99UQ8pEWDGA7Uvw5tT3PLs5iYmb+LPZ6ETb5A5t0atcCitSU4ppu6pxgPQAidVviV+/Q9F
SEkmlAmMYO6relA5edXYRZRfjgHWcr749LJoDEpgQ2fBJNtfsjMUWsi2fRqFBmsGBfKGyhCg9Zn2
+uaDPzI4T717DwrH4EpSlEFvL5eiI1FBAjrQLUXSVsy2GjgzwrSr5jW6Pia99bTYZWtrhaxk/SFL
Wcnn9Nx8Gi04Ys+L8l76Dsn6FVGLtlGBJF159o4nMaUmDg4Ok3M4AIvXtT2WaLLFpCGcfdMrgxgM
GVi8kaLoyfrSzg86P1V/3xmO1DdL5YfIuN+DsMpc875aD2gpV/c2HHRHLzkSIDuC5wCuDEtdnfvo
lMloCu5twBOLD3xM3DK/E4G0+7GTpKgjCgXnopjjmHt9WdkiFFo5b+ShSLMlqB7DPCQOoiBUhnbv
5IPCO/JJtw5KeXcW5QMXmt4Lja4prRpnKmeIX6hyTFpy/IhNqjhs++NpNJz/uYyx/2ZtB2xpnSw8
CbGwK5sx7DIzEyUVD3MZplPQTVAtdvgdiMnU/1joVQBjS6Nf8j6WsNbjJKtCsh3hSmKzvFw/mErx
6mzUseoblwWiWq+x9kJ08jrpVBo05k6KF3ekd468U52W9LfIbEj6yh1xp2IFmFvQOYW7F7G8FJ3Q
eRfq/BEDf5s5KIGx/E1z8IBB3RRM+P8TwQm2/rt/NZMLdrf17aZYktNgge74R33nrlp0Lvgq6MXQ
zkDGNjHVJQ9Mdkj3+fw4DH3n87CIQ0HLNB7H39b1IBh7q/yxfvyxajn9NAD+I9xrCZK1ZsxZWKsh
Dff1nz0z8tzDOTrPPtYu5Av0Wvxg9IrPFT9icDSRMvYcaduas7viYIBrnYOq+sdthO8IUviq5HzD
DPwW3wPyIBhDoXaWZ46/rtqi96RU1h2JHQ9Wni+gwuONcY6iFZZPB/d1j8ZUWLhhq/8xjYddA5Rx
DZeKVvaLKTuICBNodOiLo1yStfPL3Jr67YbCyETy6bK58c04EXeLnhyWP4oZLk+7Lx4WDtJsj0Hj
PJq7OA8zTZshenndTBfhDYhZz8NNfeFzHI4E04LPuZxoADI1i/UufBqTB0EyqWGArBHbv5iCX+Mk
Da6GzePiPriqSDFIHnnBY8lXhOz1PktdFtUXsKQxKJ8PQzTL+WvDnxBg+9zQbGdKt1IqCFydsihC
LIXNKgia693zRNCapwDuDexdQQxCBv61gZbaVpGalQDa8oZGUlhfnrLj0aRTsoQM+KmHGtkGFtqs
paMJZvG3sAHivn/2w5m21naQEJbrdUS1/zUmpJ/lYBocqxu8eBLwEYe6Dfhw5HSR8Tvay1ryMw9C
I7S/43kAzdqLDMrHJr/jeo+N23zo0rJ7QaPqLMBBl7MMR4+3wziOQmQzcQlyKrMsiCzIuDhe/2lB
M7Fm3BvHd6HgMFgxm11Gn9TOr97zFlZscRcs0tN4Y5QQaz83r/9xeRBx5LHe0eGeW9m1Xz9ca4rm
J5UmH/CoLZSA5TBhTeg2izU3CUe+/7nWsczVHbBoZgeD3rY6aw98ceh88glFkYFr01WjNep/ZZGe
BQ0cwKrIBH3WIis8+6G2txSoG95etMyh3bMvNGmyTg9buiudx3HyShPXcwwB0xy4NbwNfJieN3HL
aGjBzQvYht3uxVkwmqz/EOyYLN7UsLx8x6Y5lr0HQgn18thxEXOwJCGVZTxjWYJRk2uCFsCOisCm
I/1+GOEuWJzh5PmmlRg0CBbAzy+CNAewNhhfOglwE0LAH2DWuhXF9n6XClDo5v0SsqIwlG+ZqkNN
JdR+nvlwq5ULx0TOrLgYJriZvC+8ZpEARDP0NsKqffDX4iX4R0ZGhqFKBihZqRv3MlvhPt5u8EeP
MZhlcEJyuc+k0nxB3Do2RDF1BPjRh2eyyDMjbUKrpPbZv8GcotFUd7yMli60fA+kcaxNOtmlSgi3
gIddcB7ahVhbGzMzBnJtszrXNx9/23xzFVXEGM9Hw/pLtvptkVEYwnwWaLBWUB9k93k46ZlQImaf
qqjxH/Ob4rXsGmNoWVWMLE++Wsqo7Nyl/q1WT1c50SDLgfbXcipIgScEEHLXlmmr9HQ+xt251hcb
E6iUDpkcecaND0rzYyCGRbGFiYTQF5fB0xbiKPuLLJffCwWc9JTxvxNCEkCIy+s2XpivFXyMwxlx
tJE0uIH5GiDji1RBe1Uk+BG3JMEcx5mF/D6680kjwNAwE+R/glMR2bgNsJyA6W710eU7TnF1Yb9B
iCfC8sr5HisT21n7D+X1ALoQSby5sSQcYDqPqtx7MLdF7d4fmpBdVAbLpMdAvwsf3tlHEh71vRg3
rhxPG2gGVSlwnwJcFb9tLrNA8Y+LRlmD+sCFlXPQyeDbqGqPgr+qwcbNZtyNrgxSRe4PAbtQg5Uw
JRXiLKZgs6zSXJ0F7/3ubbnbNXpojfAJXAHqkiC4/dG1ceZntanzmVIk3P8WnvbcKsEX97r56Ypp
IFf0W9MlLYUy5ILpJUg5zx4DyLjKKs24Fc92UN+MnEu/se6ZIXdvsv3iyYYBX2SgcMS81AR5NT3T
Fh8hbxJRVDeANuKxWaLyqwHma67pA9a1ayVfK1419b6ICfZbNX1wpUpswSRfUTynzIntX94w1+jh
6504ixp4KU3WMLwRrAQUun62cKvNWUoJFFj6pQu2c9PJKAK7/3U+IQQf2jyxqnvg6COsRkJxgRvU
d6JfW8NoCI1yfXsNVPD9D9jQQOJ6NB6jM5cUH5QrGqbg98geUcsKw7sxDgECBxq3i3bMTGG7i/ta
LXFZjIp8m79DbIvUG8ksKVZKMjsVyqMEFT07vrLqvival6MvWzWqwwIgLjNmBnTm5AyXYdtg6azk
eQWnueXm9dbwYTEfgrv2KzkIJmH2mPLYtkWjd4T4olcn96ecZX+EqEqsla8ptFPEFNXkDe5cVFOx
e4qOtqNnb7hEy2vN1siL9XI1x5Gs24dvdga/EM71cKmEJ6Rodt7c06aEDAQbwb6NEmIJYGrq2rdR
amA3sdSN9GLu8cYA2ARwM3IkZ0ASM2egpnx+ljZeE1iwjJZx1N8Wa5lksl9sue7hBIOm3W3XqpMj
EuJaNz5eNIVa6bFYVHrSsFSMuT5v89J2u87lpulL2Sho5DH5fBQNsxShoMdlUijeRpUeRhA/BC2A
2d5YGlx3x1MA+iXlQk+vGbDNJT0B01MAOLqwkI59OKtrQ3kb4cWRJ4L8vRp6U5kcrwVjmV10sv9w
XXWf7GYvO7rXxYaBDUp/ZJ/F6PliUR1TCHijwWVbzAt31AHuoUQ6MtMlBXyoxeDKiF8yOT/5bl6V
3Q49Ry841q62cvI/uOJcSfRfk9CDnOmQ+Q4UHQiCtUlYs0lX+f5/fu0doKsuXA3HjCIzN/Y9dqit
zNYZeOat/1/95qINJB7Y1qJJbAK3Qs4egSeq56GBfyxWK2qsdX/oRdZzknWy3KJEroZ1qOiUCeKj
WfgAWVDrSWhqqTH1NhwEXujm/xp1BGVnFjhzIrxxGnCAnRd7sSvfAEXd9pvZfU8IkFWpRa37b0LI
COYHFgliLiZXxv7YDgAicsx9r2iXK0ek2SzFCk9X+cLzUpNLK5rrp1jBeuu7X8MmtLCFI4X0Xsmt
51o0TJzOgnf+40lVyQHUq41z2TuJbjkAFvtc35vwZ2LFCRSwJusT4m6NJbTRTes37ZE6YmQh8b+7
GyinE76uJOE9m7+ulWlsqlZiYJIjL53A0c4ye01BrUrYNxjHhVAnmgzdsrAlm2nKHUiOSs5kcs3Q
p34XEwhSUiP2zj5J9lJl0YAw1aQ86pAFOr2TA+tcBiHnQgaOpb4BnF8SP6Og8/NSFiibUlWDQ8tH
Gos57ctZ0Rk/ejnCPmobDOmD/wfJTWhJ7yINFjpVgrUTYov/r/0UY/eMR+wnvWshXrgwCL7V7NBG
JYq2164VfVNWylJaLug7pZYiguN633DNmT8fDvBI63bXH9bCEQ0fS5ooNClL/+ZeWyMrjyNUVSE/
NDO07iSUmkCXa/LGBdmhvmNCr0oaSXNptY9K/uiPwDvT75Qp3ItmDGiZKG/l6bRKnwOxnitvC8y3
awYHwhCfgx4LUzIR4Je+RclKCTNdTWEwnxwYIBTe2PkPZwGwhU/boGeZvbfch/yQrfd3Qz1hDutI
mVBwein3mL6brdk1GUaEmZiIU5aBqDjFhRBSPxznqBHDdpezfKKwQHVG7eTDjm8rg+1mVfz6DkED
hbCJT9xxH9bBtagl1+/BTxAnTzXmJBKg/IEtA3KqPd349ip8b4pt/A9q8JlO74U7bJVECxOT6APb
CytKCmfJMmIFOSNgParcmdyHplLZcyZQhPlQ2DbggPL+nlRBjRZncGhLArZSOR6z8YNOhJccVlK1
oyP7op6MBJNvdJL5r/YRL2Sqor0P1KUFZsr5X1Pi7dQWwm2vCGOKI/h5IuymVS4xSL6kR68o3mdL
VvSNOxDwZh3/0+RwHC7M4owczZYAxd/zdSz4CCKzw8Nl5OxZ8mpAJZC/O9YbVcI/VpFdY2iDLpmy
yeq3Hh+C3vd9zB1PXCXMNj6CE7ot8BAaTeu9abWJdZ3iHXjgr3Fc6xggt4Fou15wyCQ+x6cCWbQ0
LcvvlfdEwDHcxN0iZZpfKXk/fDfSplD2+h4lcqG6/e/MOfp5/6XcZjnbtx4UJO8z3xH5dB5TQnuW
Is1p9E1Em3KhtntBbadxLS3HLGMwbCVAaDR3Mj9b+YuVq5ktLc0DNRR2xtji/BPHuK9pI8IH5hXl
RzdlsXQKBmX2wOlpG/4jfodys01CfT8Kb+Iqs3XXV3pP2b5W5Kx2eMopReDE6QSyMDkuf683zti1
ErIYODwXULFDkLAOQvyu+kEmobMwzg4B/cx7z5219CXQ0W8PZ1+sgN3qqoTx6pg8ZaXDhirKG5nD
5QUYBgBOW8rH28BaXMGovx0TVPjxd56z400xg/OhYsJJ6f1x7ZJ38lsjXqoDeWA+jfxBbcjAYAHa
RZ4oNUafYtrlcEOHzqXqoSlQtmRh8Vks1KpBn2Ma8PO53qbtFDc8YE/WgHlLfp29bhZs4p0Xia2f
jXJFYCiy6gngcRxP69BtPP9/gQ/fP1mBCq6u3gHF2gzLjG8/NBg0ayx8GNbCZLOizb0rSEv7ySQR
PIhIyzQAZYwve51A4Yjh/lNQbcDa2bBgKQPpZ9AtIQHTVQnQuHoj/zUCk/gkfmUvGYU84ly5P8T3
jQiEZyEIfxpLgyWZbeaCVuguLl+xLJnHRUQNyHjuwHguNz0MATNCsbURH6cZKU8oEPJUMTZ7iBSL
RnLU20f3tf96tKJBa2M93Oig6uz2n1Mo9xfU78a6YGac41ftahodZrmxz9ZQ2Prn8BVa6A8AhBn6
pgEataIG8pjmMOceuMIHEb/26KHf2Y9kDiptiN86e0G1G3JDI/dVrKe0Xax6MZnHcNPiDwarqwoP
Gdj12kvOhQsCQVPWiSfQYiQ5ljA32pSN7IpZMnlUe/UzUeVR8Ll1xBwFi2NEN5eauE26TddfGmjA
Wo+FI+HCGns1HrQwMJ1/joCOo4pGicBfUQp1KKJEgnJiv7y2X3mVOxO86g+uDs8G//TYif+vO4gy
aWArl7HX1JsQ++gj6RSkrKOKG02ReKTHyj1ejpEXToC8qFyUARN6zhjfeHBune+p9k8Rw3heaimk
DElq+cIUpZv8wgIcWrcj9I+zE6OlQ8oebpeWVOccWmC9d92/JmW11SrHmKoejAVYj9nprCHqbiSK
S02NmCR0GEPna032RgEx/lzrW4wcj9PQOplI4dFvgGB1f+6md7fZhngzz9KkGz6T3eSHMKi3l5o9
b5RiGFaJdTewU4HDUQpoVq4nMB3bKDYjWmBzzBWQeDQwtI53dJl4F4eXtNMrrWPOOOak4JPz2VWl
SVgbdk26fTY4aie/QVmcwhX33V608rYYK890vlMucU0w+fn84XVcX3sFVzXWlZkGwX67uy/PZhkC
CxLaiXboRFy3yROUuKNNah9IiEoK1S7iWnBHqzogWFqPpHNwGe9S+MyJJiL62DalKQfJXxfD7D4n
2udWBHUu93DyMcVWMPUOLWHzSP5R9WdEm6oXLhZi+eKMHL+0y6QVEhD5cycOSZ2YpA0j0XV8cxSc
TKEhFMFHJ+K+I/AJEqkTmMnmiVEKXI3kO9bxS/cayM5/5Wp/NBKSt/mDeHNJ0tEQ7hzKS1YwoNRN
PIWcchFOlodUFdDwsjpng5RLSM8YLCfdNfChhaBrFJ69xFY+wwleUSYZb0hFzMrRQqYllPrRZtq+
sDhDaK3fLI+RKvACla5X59nPBznn5dBN+lih7k7mztdWK4JX4xHssRw+eDsJ2m5y8E1TDzVDzqvA
4SIeKHpBITv7HRseOMNpIxFYX69nIdcjU+PsndVc7NgKTwVBV9Gs0NQdOecC9paeAKn3YbWItk9J
50T+fGQv9wXs7YmYRQA3d2M24wtIZOVINWW5l808aBWnO9GL/0y/0MBHiuWV9UK8sClITV6qW8pz
dHxo2+/6rwCED4VF3e4nq3e2Mn+87oX9GbKGsH6poADZlKA4tX0gAICK0cjKgfIsCvuP96mP/7bq
iEgPSC00CN+P/QaAHvL7H/VcdOTI+mk6xfSw/qKHDJxSA7hgNEnD+48+mJSU6Hy/fUscZy4myKSW
oDF1ZXxkGBErh5vHP6y0WR0wb+I0zxAsOqRcyiDzRwSc83YoWSt0d1H9PAaNIcCXqHR4IeD0Sep7
c8iwnRU4liX34zdKcUtXGgwAb/Sgj5xsuPKkljLnL4f+radD7BWzlqOcvzHCbLGMk+4TPJt1Yjjz
x5I6rQvKCH54MNp76/boyA4rSV2KBcv7WOhfSRO4zFiHqYC7Pk8O+qlqzmFQ5BOzbLG09Turs9Ta
mowBU7Av2ZF52ZPv1pghLLg1Yq+vfxRBRfGtybsscthIdVx8SITx/yd7YxmsHZDzfAQ6U7MhG9Tw
4059jEtrwr6kHTsDv27FOCrr1hx7h+KhoFDDmqRh2koUtacCIUOJ51W/i0CCs9RpQ61w9CBKIc7O
fDiRQxPs3pK1z+dJkMWaEed2ERPln+ttlVHhtaFFXmWaLR5KS7dTcm6YZUXXURhtbN16ykD914Kp
hGE4Dk+IHp0rpyGdZG2eQ4BXLCpzqL8H9Ijkv6x67gRRI0EWOs34IZ3Enwf0aZjj52bZ04QIMkAT
WqMOgJn5iGEFo4rBOr3djpiRvAscZfy184CmkYskiZjNmPWVBVh0SaQNbJxxBU59Pq0LazVKOuPt
NZABXkNNEhJtvjuYB4Gt6XgZDMu2F9Hw3GrAEU1kqroUpCVy0piXonA+8dZFh5wYntYi++HFZpm0
E00C1nF7EWQjuNh82+MlZkZY5uu4Xfcd8Ie5fHhsd1c4OJmuuXdUTnJcxUEAnvPzF962o8rHF8Mj
nMrz2eezDpb0KeH0953Cf6er0WCnND/IAM2KEIOb65es11FqFyqAnvIENG86+nMKDgr317mPu8Hy
4glNRzti7tXrd7wTgLsJImQo/DF5/TUFAPY0gSKe+c6UdlcmCgU2GCXQH370aEVjsRPUpCYpTPuP
UUUzHrubB4YN7+cNcEKBcx8NturMg4Ku8mBEtsp2rga3Wdn14FY3N1gieMCtuN6+C6tZCcbTFhEj
FxeurntZ/TZPHQ3ytlRwB1/3JquGBCs4g5vGNZK6EUnXtJbdMhLRROj1uUjvyG/WiQY7+vn8+Ntz
Egu5TmFx7/dJB/Nz8zpPZFUmGNFnfPACzUeKHZfun6NmIQOUXt85mnIulxsb8uCvJAyofZb0tyU7
qX1W/chKlv0NyFTYB5hDtbTemNITALbByuZWcniyk+CZkH++DBfyvV1tTYPQ+WF3oQhmyK0osXsH
AYK6l/0SJtCYjR3fbY7hPXKmePfDiSlyjkxUO0XBHoVU00il6dp6TzN7gnLEMsMTu1cJ7SVNJQ10
zK5qdWfhaamJZoHs01t0bW4R1mPJ2kRpZ33bWAMr7Hx+2Zg2+VPV+QZ1bnIFpyKQ4fdhAI94BM/x
J02q9vdMm6jSNkH1Uh2hpBsIaV1uN1gNb4l/+temgcP1+MaBsEFo69aCxX00+xsIzDO8sqy+exTa
FPxU3CBeoO5qHRYvL+yRHJw5wt2TROLxcxvyqWslGACiYTdbT4YIHWEUBfMdYLiganrloZMjds2/
j2nI8ricKvnxGI0vWISyhUhjU9bru3Ulnt/mTVGDukLijAwWlihRbYZ3hdFAX1OJ/GrukSeHkfbH
qNwyPNLXREBvzrprdvYnYiAYAUPC7LTz8k1AnIEc1xZjlVhfjUmLfbG7caCl0zoomk2yXs+FvzH6
8PgkjOVcbehBb9DB6k1pMFxlzwwh7/7wtZnP37DxXewyQKqyEqHz0zQwM6i+BjLBnG+uapjFMLMF
bquA/WNuO9XeqlzrgyeKP2raLMlTkutM17Pn2nQUZQe9U8XrkEFkIP4WaSK5lfACeBw78XI9mCHq
hMj48HGY7ZyeQ+rm18Yma44X2mrhnxdlx3AT/LIYcv//eAe/lxmCEKyeMiS6oygfjl4QuMcPvM8m
0lXWDklv2c4O7RTrioWaLj5c1O/bi1vXXJc9C/N6/1CCbPullVGZjxtN+rbJigQjsamseK83dHCn
ojZnFLtIY1RPBmBKMmAsBeaNF0r/smpaz5WOw9Aekqg2ks0Fo+cIepcBRQO/ADEdqVI/sQkqSQUo
v6oA7NBvDEVcA9Pk0QrRjNIPANsnf2N30RPuwTwsiqdqWDB73S5FmMT2Mc+nrCDzFkgBiwGYW1lu
yJ0vmz8kCdI+vHCLiw8dsCSwq5e4RTEuRgm5zwzrAHdsHDTetxxpkQXQ53vCofap5e7WAxVPT/IC
mI/aVYHq94EtSXTJ89dI1l+TYtWT5vnvCLKrpB+HB18/f9K9jJIa2xzzaA/4N4No7xOL3GKcS5Zz
ZXxQQ8aQ6eyroQa6UNT0L/fi4wZMHi/O+efcYR+UJH5oM5tatuefmT7IVgc4tUqORZFyLS4DnmQE
b+EK3kvVxRiokQq/GQKocqAOp9/AjRlZ7dvsKIxgF/xm9tEtAfo9fWfNSwQkEqa7NJ43ljT/yZpi
VPGORf86wb0XzWg5R43lnxTA5d2KT6TWGFlR+0iluRaaucjIww988JIjIhFiIqFmnfFl/mDSYiCq
hN0Xj7kD6+31+wQ/spy/fWFlirltZrTlnx2zEdR+5umSNcfJwNSJSEs2YdvQDejjTUmVetKTlqia
2kpH72njzUizYJTGg5jRJCohuG1cpgdOgS5vN+V2tZlMoYUsuPVZI68OD+m5oH1oEaD6RDghMBa9
arLnXpXfuABCirVJVQkAfzSL06ItZQJ223mXdWhQuNOM/shT0N3CrrUnaBT3CePnjT9bEmzuAavj
u+QFrvEkV9mgJMoB1XLdludk20xCknkzfmezuCUiXlLlpArX8iLbsedouHMXlodWk3C09dYyD7xx
Kv8i7zUe3ehZdyXnqZRBW8sf/YrktZ5EINplRkaBW4LBtN6Sl708l5khNjpSuKMY11P9+ZRfGvZq
Tut8nYut54971btPgDNw01loIH/mWseCSUHWZ0uJsXKTb2t99fY1pS1C5zCXIpCEbh13p6zyDiuD
8H7LeRRysZohdKEe0PvISyglKiHHd3qcnI5qtKbhuYS9VpKvaqDmkqLd402gtlqFNHvqgdOSJalN
8AjZnbYOdsFDe0OfxvzTRfBcJDUcWsfrYP2xLtY/MW5NNED1PfZ8Yp3msX2+0B3MdAZzNpLcZ/v9
UpcKDiZ92sWZUoWkx+fCN2pgTBv+zYaIsYIVJahoIX3ey5jfBiD6xKizQNNlFGbldWpKUxAgZlqe
UA4DaB9HHbuPn9weOntDtLxHg6V8Z+t8CkcKtWe7Dtot1KjCWrB88u9lc0tSHdA9wp713XswCLWr
vQppTZ8KVmOOErnTaYy41kF4IK0kX6UAGpYnF/xUz0EomawthIEhXYNr1Q8Q7Q0t04Nrx6H9w6Ye
yFRa9L/+ekvuMSfR6n0+QIrK8eJtBr6UqSLgjcq4+pNrcKNrVjWWwykJhBs/a4wVq/W+JGSGCB2E
y4t03Adw05KRZKlgmAqunqP76Y4hfBQSgNpVE272x0jTZ9dm2q55tvWCYN1yy+qx/cV7wb81C5ic
3tldvucTzfMp6H4zutmFPwvZHYYPlt5Yj5EE9iv3KdfVKeb8CyXP6i4y5uCpXXphgJDp9sVycaJ+
IU/nWnYaLBOateBod480X5mO494QxZmzTDgUney3D63IgbCrHyZjk9D8CBMcdk8RwLJDJb2ekH5P
IjwUgaNtT9WN8pu/nD8M9EjcwrLg78K6bLJxG3gPSuLo6rjbPPiCNqr2f5SAJdnuSFVEx0LmFhYk
GAbz9eR2mJssxw9/j5JgBw5IGVnPlz/byPi57FdTJroCn1rQuzQYk9cSOSTiTFf6qD5PP+9FAFqA
3SkmxunglR3LnKvsmopctu1PcPYdyfniT5xZdvI0g2gQAINtEgmE26gqy2ryaIMp4DptAB3gn1Sx
vlO+1iKPXWepzDCuavV/BhSXXHA1SBz0tT9WS84LDqlZqJrJI9Y+xAsWVE9aCtkajoIk6JlvWwIB
EKEnVCCIKJ32uhfV8VqT5LIl4BhoNuI43IJZxO7+haMxa4V/C2pavp3yckZw+9VrfuBKdS/fv9hW
sk2qtlNmiNla6mQKNq7CJtvCRmSlMvPCbF1qpgoLH9GqEaRJXknaREDJ10NiSM+JIKFN5oMaM6Wt
ZZWbrc33QAqYMhQ5IpstRugkjLy56X4RTtvVUN1ounkBhZd+drE4sM4kkMHG6Tqsc7vxYn4WPAFR
ha8+G4eZgjvBZt7dvbRZBUAcuyZ9imwFfRncFKm60WzqCU5Sf5gP9z1zeiwDx1AnCqtRBd+79M0Q
FFjtWxQH8E7DQzF8Gksn5OptW4WW6AP51AqGYYRwfR8gQIETzX9J8fjxxG6Y2WYZM/Oy33Y6psgs
zINRmRvjcJtv6A00ZIUXlUTt5TUK3iZORTzTzPD/2Js2znJyRx7+HL3JKyaxUAXID5DydzJ2trPu
qFnxXaXjeI9KOMwoJq7UAMz2Y8+uugfNI332ObvUb/CtLB3AHdAOod6u/4UbalG7WPTjEAD2jcOL
af9kSVe7dK5pb32lYPZiYr5Cfo2enMtXuo+GJDVr7rkE+nZeu2yNHareiLKCniH8+DQuX/WYfh7c
vR8OG26n1jU1CQHpNplqJt3fBgLSCeLd/+6beNS0CNqPa77s5hHCJH0bWPDpxHYtmVx8UK4sgs1I
u/4Pc0BT0VxPvw28NNuqc3aci2x77cjmELG68GBJe6e8vEMv/XZjYQDvQ0XjEG1Hhc0aK1VRoj6W
melGNPzZqtLPXuTCl6eFQiRjPg73wNQKYlGwjUvefip3L91K76+62LKMzrRk1MOW8ZCjEYfLYvHv
LIQ06Ci8793fwDOQmiRs9KP4SeFmqLUzZwlZuI2tz6BGTRnNXfmCTutq9sQLvxHcuDDZem6OYsmh
gUgn1BWM7NQgEkBG9xWZfoPhb+sg8FukeyjF3GOJj8cwYp67UWRLt5hipK62mRIMzUOVBI4CmwI5
CMHalSBE/+Fhkt3V0fbG/S1ZEJsV4+o2pYgykJiNPPtfe86a9ghhq+DsgpsoWQhafK7cBMxv780z
d2iB0f0SUMPRwkXkEWWpLRs6H0kLmQLidgC84acSjmNKJSqS1MVihxnFlBSqF5lKqsDmb/wqCw2D
njs0T0UAmh6M7xemRq2Y6MGd+O/kcmFdbcbO2oYR81CNKu0zzH4O4Yh2V73/lK8o+Cs/Me2A67oS
1GnAUzZGCSSBOrsQIeJ3ow65OLpZAyLPIOWN19DUuXf2s4NLdkGuJaD5guSAV2xmHTUlnkXUlYkj
e5aI0MBnz7C/L5Xv6CoTj6//fLwScKjEl2fogpNRmrOpjcSXISquuqdFhqVD50ONjGp3nOA86hVq
6dTjACsZyYlmxc970k9uYDgql7/Pj+RmHv/PQRx7QJOVesblg9HrA2dMZJAz1z4S96Iv3AY4SbW9
4YPXVx7f3FP503lxuIVikOT+5h6VFiGbgBSG6+pvft8MtI4SLWb9BXCaLMNu5wuLG7oueNFEJkaS
3ZaPDKJ1D/tSnu8gJurZmgtcEYLf4+YAVxuPL+G+scK87LN8RU2meipBMjneBOGMmprMa0fD81+D
6sjsSCAJ62NiDcoZEyqadWIwX2b5u80wtVqalull3ayFyBQ+jVflxHOAWYDhgCLqh6wk0GT7zkeE
WqLDxJd6wYYAR/QcWwgYjGCOAShbtf7I5M9I60VwKvMTdICss/hV1ajqK3UmNRT1OXqj8lm4ZTLP
FZEMeBr3RPzgfzFtH9XFfXljDoV8iyS6+0SaiHSFLc4bEVvkysl3kk1PXe9Aop4Rl5P/J9C7dsvU
x9IJ8Br8BPfzKe8Klkj0w0B87aNmv53vKyMyXm/sxnxLDJYddJ1v3jK2jfdxKD0DJkqmfHitTcsw
2Dz3QfB+7rzU86U5ceBN6fyfHbo+hJjXQIlEKNsXeQcz4leQdao5NCxNu7aqfAYVL1V1QI5KWxEk
dLR4DabLTKsWZ2rZtCT2I5vvNUDg1GNWpuW1bjEUJfhG/1TNXgoiKaUZ2k/ePcH4CzXnOzP3BkJW
YgZaee6qEwMWQXWdKOjkfknOCbassbkmkPbyVh1Q+t61AV9dCJiAjJbi1yQHPB/X6ikcilGxxyXK
+ATyQ0n/BRpmN8+LfJhvQqBe77jPPOM70K0l84yXCAm0zWkRLjkw0eMrmdzcJwkd7NEJoFUlcGQg
krRXvFaGPAE5DK4iQNwv7QNgIFSAhUJxawE6tUtrXKZqDytH8SCONwvZT9+mhYqLOy/6TJlLjyVp
w/k700dW9c6z/aH5hFhDiQR+clvA9VAmi6IfdFFKvAHhvmzmL6LUIgDheHEATdtYYtFZ9yOCC6Tl
uid6+3H4hvizNycE2QfxpqgHr1pLEyt5ZYbUQYRIyUbBSpJfQVHE1mP1mKfVCqH3dGUOBY1Me7cq
PtSCZS9Vy6y17TITyeAhF0dEVgXkeFaG8+8yh3o2IKFQaT3BIckE2Yps3NDSzXYPHtnPKa2CAFwl
lq9uJ7u5LGbf3nTY800FIdxOnnNOJIg4jFpUmAdVZ+ADWi+AoODRC9OLhJeOt+/0hwo+dQz8C60a
dSwerbR6auWsi5+N6gdjSH4ciZGVHOdXJENahJ3GlkvXg0LEsRZRNZC4A1sj+C+7NRKFNoCrXiNY
df6uGeINBrlpmsM1gXboc3jdOJBVLVDkZUGtuBtQ5X/LGCLUJ4m8R9N4yW92mPQ+PDXj7oH3r9Fq
PLdQ/Vy0SuzeMLaqD35qYz2wDIN0V/ZimlshQjM2Q44eej5qpnj0Q5r8ZzeYo6CeENBMTgC5G79f
rWlVjZXvE6bJttpuHs+3ZARacJ/ANs4TXN5szMpmGn11fiPA9f/d7qhBkykB7i2OmLzpeK7jAc3z
BTGvw3f+ZLA4v7BlLEWsHsl+90nSN8XKErRS+oLAQN7s//508UNE/0m3hcroXETAtN0YfPs9I8mA
vFVC112CEn34kjd5Xci/RnCIMUwwQT0c/MxEVslGkBQjHcxhPDkTC2iAY7c8wVH+A3rgEPNv9YCb
z8HsPSmeGatgMqs+nhzdOGZrN44XWZnGK/AocTj+A2EJyMruFXVhO5n6eAd7aflXMYB5pWIvvKxt
h0RpmZI4sqfOGWLBsuQC1xJ+ccYRXr2MPgcYiQziqK9BfcDPA8ERttgu9CUttuMxddBtTPoVlC6D
JB69ysG4to756BJcNRsWf2HJp0SCtvIkMbMfnYiX4AueBXZvt0KpbPYhfpyXlGngVFvbKY89Ai8P
2QNhBdr+YZ3G+Y4tO7rO1znMwA0ccqxLJKyH5cxE+9sXTDAFg8xsHF7y66D3y/X1DHTkxcXbQN83
7RLOIJSbmHNENb0nlOq2PoCCpMyxXC6TnKthnc/slzCGijod1J+R6zWN1p3IC4uaC8Xox6ryHNTD
pzsHuaF8p49LFagOzBi/O4a9T+tWiFGpf1f4ZKTbxKHN9in9g/ducbDKpfSKVHGJg5mpQx4lxSIS
SvghE2FdzvY3rwjpEGH5aOtbU8uYgkN7jJQUN5lFdSHjN5MktTLMfxlDGavB9NrEqg5leDYl+rqb
jrT2Whntx8b1QcMCI1AYVEeVJyrqWuyBxKFeCUuTRIbX2aCEaFYDg0OZxJl4sj8KzDO2gU07I1Fw
ThhNMojRRMS4UJ+1mXLn6w+9CNDkoNxjsiV+94Fnk7UWgB6ouTzKj8QrYtnSbChWiXQdd2NJ58UK
Dfe6oX109UsfVLQCANY61mEzcsJy3X67yayQgSXx1GeAyQT6fUNdCcjzFoUH8gz3Tw/chmv5urCi
5LUEJF/UxrCRNkrg8Jcg9dbZEv9v8iGX541VVOsaUb9dzDmVEQcJ9MmJWUkpaP0CfCalet1rpu0D
jneGX3APBFkuT1l4Csy/Elpist/rkEQXVR3cgYBU+KnQS25TCr6Ngzgu46+CEHpr62+aIjE0qrJI
+buIm/yFcMbiMq4Pb1Wa/4z/o+YWqq9SWRj0SSO1/Fc2bcJvKbje+l4jttnty/ywID6OI0u51Qo3
IQj4wos6JMVhumHrLQJ06GPX0/3FJxF7+Drml22g85x1EDB1k+w9bILLa9zasE6866OZjR3uWiGQ
1+8Yr/5NgCb5tCS7HiimcuNmeASVtPCEoI5b8Vodx/YSrBEkW/fs43fZIVebvQW6vpAawwLJEUWl
u/MNACsM8p8IxODpd3Ln5gZvbk7HUdBxsP2xBJKkg8uaWiDo1MzH3Lw77emgcHNHRrNwBfxDUGNI
joeybjiXU5SiDwf1qumwaOnBWXYhRBQWGcyn7rKJSjrxAR34oR5TfotMBgw9pKK8e93lGMrFoa+K
WMTD98fvNKtNQ+V3I4ilV461D0yWAdjbZ69VL7NBCu1KqcX/dKY0w3kGLRgrHHg5BR+F8y85Lca+
MUsRsvlh5ZHngYJ3G2XrHGDJhidizKrjeL8AMZSiYbOJdrZoh10C585ll/+zyDXZdwa6EyukD7Ac
Ia7soS2zrMQbCAfynggag+wV6DFCS6GqlxiAlpiI0/uP1KL8DottxYpRvzQbRGVa/CmVijxesiYa
qyh4yuLhmWe4KLxik8ULFxFqRsAxPHP4TpyxTJT+vtpVXoPT+HjIvkfLA0f4xgEl97EFugaII2T7
59r0EFPkgOpv3So4f1cXNW2kubTZRJ7/dI8COxlKHUeOfw06TjFL+azVV7IhZSr+sNyH0IeiqwMt
ZU5Miy15rMiKIQIcC31myGVMjkp4yrW/1ywueNs6uaLWqCVpxupJovMdPzJhe6gTu9RBCByWMCBo
OO91hcf20p8SaBM2BztjfWnxjI/L9yAGiewGUbdR3XBIO56m0//BFYcwzbgFOwDrOrXKDNa8cFVO
z3ap1ZVTkUJbzJQfgFPF7yqn7HdokXv/fFPnJsVmtONPS1JZYkudPVk/TXh7lXDC63xYP2Dokdem
3BwDB0iwj57ieGWJ4MUXNNmTQi1oiZe4iZcWJvS0Y//AWX0xsVQ4EESdVYFDGysX7ezv7Py0xxwK
ckXMnbuF10TqGltPdNfCKnppNfhrK4nNDqn+r6KnSZvlyBHUE5/IaR6GEyKpnycCLicb5ArNdxLV
K+TOUqC5GTkf6Mo80f5LagBPJgFZ1Uj91HjHASLhRWR1BU2oLJ/IGgHJJzIl1/7dL+kFD/ZECsL2
06ARqkRC9++jqS3jFDN0K1j7M5RBJbrYhRyS74jUl5a5QnjqlM5TR1kBzb6DH3kWtjqlsauTFhPA
wkD+WGB28zK3zxi5XhD7U6DF4JrmWB/GLvSi7a5o8nowc0g/UCuPaLAYsWOz+33F4T0vATKz/bU3
//EHtG+9NKrHB8hPtUbYC668jmfMIdzn1TSWrkEIHcitfDCE0q51BhmxgYwaCzrtAiOf+8fDdQEe
pMIJnlQYIgAE/L+142YB3Mm3WaGQbv8GBZjEpqtqIFjtHadfWVwbSJyWoCgCnkSN0HkT9SRvEmpF
957jRoUpS3+lBJYpxF+1JJJQt6gq0hzmyn7ZsS+nB8MbYtcFQebjlhChGxaYsmvsJQBMm3qkhpGU
mn9ooFnihKoYKhfRGFd6JXbK8m1iYdbuI8E/C1LVylNLiUz2nGUG1JHa3V1tPUOlX8WfkP6i6qYy
XWnSf67NEnGwyjtP8rTAh94+inzU5I89evw9CIt7Z07bBEHAf5At/mW0CCzMS//pVhG2RYb0LBPV
MAPCNjJ0uwz7H3u6SqCUzoeuN0ZzwbXkV7GzLZjw3+CYhzT1N2L5i+IFOCSNTbURMJQck07/de17
Ls6vOSOgI4hpNxB/sFGTQhGs0lUP1hDbnVpIvfZx+MacQA/nEYFgWexz4xB2aWOwbaiNkPVkW4cZ
Pq23vuP46BjvIHtFGI/p7fv2TLuLbEeJiRNofbJMx6/5wELYTV+NcGXqNyoM1+SjKpRRyquAF9Wr
bDDIRDHdvV1kDbgtQh6PKM6RtzMcFfe2taInt6JaK/H+haAoS5lOZNR/EAJxko3uUZKMHyjTtXTg
rcsqjgmlcOf0mLreNcQLyzqAuyvHAySylkNGIxZJ9/+kbvUYa1NrG/BkjyJ85Z0CYShWl4jgugfM
WPR7wdTfot3PqMOJPkBzmVXKc6ZrJBTna+u0BCHMONABHNrypD4CzftuO1JtQvsvDFKlAlSiLlRE
Anx5SVhHikKE4pcCODgR8ZyL/NjvwhO4RmwkeZ+fTQqkP5ENxo/Dgyl4Umr48AdkrlZEASScMTIL
lBo5M4OPUmD786YJp7ArSr+G7OlYYNJlm6uyLAf2SE0PJtQRwF64g2dNjMtMn4bpwzeKl2MkoW56
AABpil5taUo0GLV4edJl5ZzCYR56h1O+ZAKbU3lrD0FhbyVV445WcB16+vN0ToTjfl/DIzhwczN8
WGaX3yokGwn4bqFoqVFYy9CgljXwNMTmsSlpxwMFX+zsHHq97owFSaEKhjz3Bev9opzt/9uHxx/p
uflULhoRbxKpwNK8XMm0XSqABKISo7CgA5fFCwCmKSVbJc8IFpS7XTw8+wEmo9BbwoCa15v7Hz7h
g0OymUUjJgrNYrHdb07XcGkSV/rJ3NrYG94gs4ePjMM/8vnh6D57BeBXWpJubJSTB4Kb4zamCwJs
KcUHw8NrDqnyrCL8A/Sg5FJYEqEYzAkHDZ3EtKoZYQnbH0D3Eabxjzf5Cfdohny/hsZbPMj3F2TO
kC5Ty18ol4HGNhl50+ULfnIw6mNjbno85Id/HUsoaOvXFiDtgvr+ZWH4dT+N1o0Wv1XNfEfrFyRh
NVvAcZz8UgbghtlOlTniaEqRvVH1q4Y6Y6j7EJpG1gd1CGxR4+Lz3St/8Zpl18ldBud5DkthybTQ
qNsyeHUOIK9A1GZ1fyRdqP8BLDhHg+K0rFCVwP/gTNUXgP06MDxsl/jAA056q2MS8ta4QYKN7ZJu
JlapuBwpBgA/LCiK1HWylQW6JggCbmGqMfPuWJTW2bHTShnqMKiGz4rmhVJUzqlmqi9IDoLIyHZK
Tx7AtFVT/2JXS+CrGyKkLTFMiLMnELOwr6S7OP38Qzf82gS8M3daxvYECx6nJ9EFSjJkhZ0qb9Od
wgwUJ4W5ph2gsmeIb9K6+3DfrGg8xb2Omj94iQa/rM0eBhLUytBaCkx0f2VwZ8XyaLjb+jiTtxDj
+0/34FoGfTAu0CkmFzdaLJoX/DJMWJlLJjJ49Hm2rpqqooqEz0nk29TQShCLYe4QA/RRU1O7jUp9
L4XQ3Cu6fiU895VKVUzXE8S+LLY1UJcPE8YqFffaPMTxup3qmksQZL9y0VWghG4OnPlyI8KPY2CW
5nlW6+CpzKTEwRNiGDbe/aD8XHWw9cTdir2QurcbULBzHgUOMwab3SVonGD2oqAmxUEZxzme1CXs
Lg0IUNLkrVKwECtD9xuLAfoMBHyFAOFtN4vQZWuV8bhudxltt/dC9DCEXg09gi24Ei1TK+OyiTrD
lwcy0/cG4AVkzOe9iMxa82jxo3tZOM/Lgto4CS3SDTI/+haXiICDlYw/NRlcyJcfTxsDFcRd6byR
Fs+jLndxGCLgGOGThnmOo1SWYZeZ91dsFjYLRJbF5mK+0MFfYhn/ArT+P7x3vs0GYp2FuffnIWHm
0+0hvSTjV40gWPB0XjkEpZIjReMNySFxnKPknwb1mQPwxsWj4Mf0RVQunOAMz/mNEGDogFhzwUEg
e4ub/v5QTziMohdJYYZetItY26qfyzZQ+OX5UG3IJKL7wN5SOTDw6P42XfTI3plCOEciHnACsjy1
BPswKwRHD1fs08s40Bo+ibfrvRB49RyoSaWWkX6bvwUtZOUF9GK1ePbbw/sFUkIiVVuNRefqkeFI
4Bsz9XY85Nq2W+xB23Ozdc9Tx7sqO/kW9zRwm15I2O6gWvwzEDJfGxNl+GWxRmDy5beBDZognG9i
yQSvOT382IEKkrTLNtDY7yVgLVp9eW35S0giUsremQWGSLzXprHKbPI7Ya48zKrg+ewo001xVM6O
ipr1zmxh52z77tCy2o5ims3P6L7LoMYupVEFLikRIpKZ7kM0asSLhFjaaYlsG582Y5fC4rBCJL3q
VsY2LQ5t8e7qiECAzqehwAO/FFNVWZDllatY1iqo22CqmRWvOLZCJoHATILIjh5uAFFDHKGEiXPO
7TO6sMb0e5ZB5+tk1pd6aHT6peOpm+bykhNV8dT2kL599AEw+C+MVgynCCnBj66bfu15XRyDBKK1
xpLHjbxCWJ/sI9bZ1PH3WbmGc8eOYNy4k8rWczLT9wHE3LN0Qof3U3IuSWe468G6AO3UZAr3NLAv
Ef6ymp/EzjB6wTLxaeEWLO1LYVUDkoliZQ43bXJrbOV5SHwNy3i/+S3D1s1rMAaFFo/we9TR4zPY
t5UTRgF7pE/1iZpL2QLuOeZVl4zFTN6H9WSiLlTiz3I/Qor5m+tMeDZGy/4r5oPqFTLYGqFaic7J
LDVwsdwbMZT1Ps3ulh3/LdegOuFYZpH+1KA8Re/vThBw9l8VIdRE4DG3g42lKEu6FwFPKK5VnTwL
zMMbEwRMzjvthvXg/YSGp/EQNCZXKahAGNzK2wDTBsAzDmugLrHxmsR6FnWxfIITbXLVBPqvNxCJ
2m/t0bdzFPwSktfH9z1Dpn7a82cgF5uhGbNvr6F7w9p7NNYHpH85wbP8oiWrQ5xHwjk3zgcySyh3
Q8Y1zctkLmuF6P9NiXSKB9g53fqdI29kBtuuze7hNpuDLF056wa14yv4D81A4ZRm7xLjW8Sr0FwM
fQ1Y4C68gSKO5g6lO1Ce4wnzkvWgG0v4ICMxJJHLTs/GvKBOtTeODoZfU6r8+DZBlAfdEJkUKlZt
EPNchtzRiPgryek5+uKyZzorRQFdAFawh1BPsqsxE3Zabeban6Fw0OFakC4FoAwtrXIJ9apxYGgY
rw/KuGXczRSdO+1ZzRv1X0vUEZ207tJOMcZCUW6u8Pp9o7WGQm81HtKufqcqRKtQMEvsLXt8htbk
UMHzJTiLtGKG7ltX9Fm5zLC5Nu/b8j+E++XDnjb2pX/0QMsLpo3NTktTVomcS28rBEvLf/2ANSCB
okgRyZfgSnP7vTfBz6m/jGohf3SUKFsDI+ch+Uu65UwuGpH1TgY0CDE7lDdZzETSX181ELCJrPrM
Rhpdo5AZYwDFzFvPGX+SYabtbecGQZZDzLqcc8Wnf44LfxdyIyQ8k2LVzc4AchPRvtz4rZCUvtoa
LxMOzWJTReieGbjHvISF7yDTN6rg5WCvXYm+/YUAHcgAkSselQZBSVOLtx1FcvJpaiD7bkdzpciR
F3q63mJQDb2wU13mRZnGC6j8Yt6GFuIHHGJZGKV5m2kAQfqALv73enmc6Z3OR04ivII8kEzRxdzM
MW7bH1mVtlmHmyDlX79OqNgQD+G1yETNLUWazZlNFvOQNyVyOAoNUUzPrusrULTbZzWsyAfkXyf6
rjd4CZ2eSGGxVE3SVY+HmB0ml4kcYTZFoxmIqi6bkbQ37Qq2pd2V3pbmWDCzgn/xrZqEB+tYPZqg
Tbzyl89fzZmsdPGlDQejOg80MA8Udyijk9sdrrjZLvSVEL81KEKAzmKk1lHserllsmYFt75iXrbp
fsfFIcQZhonjrORWP3+4mriX7br+ODej3hQLh6Zwm8UwjlkY1hbW4K395qxftFYGaN/4AJUKkARU
4UfFAMlXKvFkgTBG79+NsPzIbDWs/ks3+yh8MA5xBSAeSAB6vVumxxgG5VV4OP8Y36NsaJ8Wq0ej
ZtOJEL+U7rkRckYphOUHgIeYp8k2/3J1gjikOj23pyOEdg5yMDA1RLZJ842BQe3cPAb2pUQwLXkU
Zer52KQUEgBao1nt3dkl53xOKOsWTrhu039vWzRjL/BMi+wuYKNeDHcC2Z0ax/IP1yIgYdPWRW4C
xlHOVWPNzE66DSGtfDfDr8ubFRyL8Nb5bEuJ9b2fS4Tla7V5nFyQCi+kvdt6dX/BHq5X87Kfe1Mb
vWTPwR98330JZfAgv7SoxnHtFNy+flpflejhuI+AFwFiU8QxkC/YDkk+GhYKan7yDsvONFe1VEam
1MwNCPhCyNZ4ghp5zr5N66hKWWJTaq2lkUkMaYTZKr5pc/3zvQXU2zsZT+KiE29J5sS8UJmsLQ91
3CahbTXy8GtzGyHwmLniRBUOhoGcq90CIYamNNmq2x+z/CwYmVF3eq6TQOZ0S2AwwI/OAdEgcq0K
JPpMCeQQzqFLAnMssVGJBqlkWbJXHrG02WQKfswna18o4yjJ8IoHm9I55wBxKrt3dSmj6GYc9wp+
fgPS0X9e/52tGEYVZupNTemnkwoRJwWPcr3kEuc7nyoXyRKm7rDQbGbFTZIJit3bknWpikLf72Ro
94FpExlk8iSZefd7EJgSvqnjPg4+Xeqgi1ANOKNmSCwxxbTvlhfr6/xwPYDdtHRoh1lsJ+uNriaX
Qcq7ekBErpo4hkV1V9HZLDZbTbJFJi8HaUwOyg5rZ1AjMIm2TpcbifWY1VLu5f6lqEKXR36E+nmu
yg8Q9lrVyJ4r9NJYdvUT107i+pGE0mv+7vTgHGgz6npRb6i48e+10UgdpoWLR+H6lalGkujq7E4t
GrcV4x62Umwf7JhI2vjkBoChyM3YA17nU69FzcW1otPEKZrx8feZ2Vht1GszxT28MBgLNdOsFm96
RHI93om1uIOymQqOSmH2KBzLIZiTSVLkZ94cffDhpnuwSveBSQuSuxUNoZwOtVmtLul1sQZdZq+A
Q7EpPKOy5RAwyfPZPBxZdA2lypYWIH1qF0U0qzyh8GvfwdkAU+ErOSzI6xEhZP6If/xQ/2fn4EFq
vaXCcin6SLrzZFmndaSfahwbPrRWwyPF2teFAoY9KNavfSnnE1t/UEKRBPBh4DlpnRwOLg90cEFK
Q/bniMVArfCb/1vpYwSMbTCM6+9957H3AlVCMg4nSJuic97iOCc8y5wklKIDNXWV8E5GMA4jkfE+
jhQpvyfjzC02//eN9+UEPf+HRoB6ZJKs+8betMsmUBFyHfRAHx585SPivkMAZvnpyi3R644iSDDN
C/BVW3MUvaqaQgyPUYGR31IsKjwD7FOQ4dEoQ/hv3HlUipg+YOUruiN3joy9fAftjzi52MN6Oc9w
dXDJSlaGz3WPsLlmjWZ3PEoBBo+0oGjy0nBxR9vrabiM59tVxiQl8HnvA/3J2X6xVm8uEumizW6h
FYROorXvadwUgWCjukS+mGP5lRXSPhZK2pv3o7+Ci5QiGd6RrXhOe/xMC+wmn7a9bQN2sEWdci9I
yqTqtY2AjBfEQaaqAqnzmVn+uhByA3tKUFLrJiYNEw1mMXJUnlJify+r1VlUyKLiLzAfVysLswWz
M0AfM3f+1rbEc/O//CuRsUJ52T+JYpm9sdIpLE4hYOMtiAiRIsru1DIX5HfTAUtmDZP14LIPt2rk
zR+8fxPeyz/bSoU87DaofUzcxW5SeVlMAsKBXbelM1pKMYQxB2MXb2hfhVZaDyftezmEvTQj/T60
BQ0n+EhzH0GNqErSAwTcNczQ9BIwdulCilG2U9aK27tzlnPm7Sd4ZO2XEbS2ivfEVsZa057/6oAq
bsKpHtv1eS7UVt3qy6ah52S1wIeIRfTsHVc89rjRWBMzQ1xP0KCkaZ4JI0it/jbD8cPB++SR4ecA
OKE7lmZSytpVyPOoAycw8eiLFBOvlBbsxZWIELjDfHVdCRY5ZJMKnsbG8b0fazwdg85LHiw66WlI
zXgxRS8qybc+CPfnKghPQf4qixkcaaiytJFQFrw6GYaNOrnYQGZaJROIfmKmjx0daLcVCTjAP9Af
2vVdZPibWmnBGf+3zKWTLa8CylBgQ/qZIC0iuzAL4Ij3wr4lWF8HnrleNVnL+k0tI/b0eLrkUPyl
LUeUgRE0q2+YxhhCc5xUy4zzm0/R6NcZmwWauU839O+vdIT50fYgQKcTRNTqgIdyZKX4Rm4lN8N9
i/pt637dha5o8tnHuBizu3VcEECH90DjbD4XsRLDTEBHex5L9wQ56V5CcA8mLf1dlmArMvXS6jb8
SnDBUUuTg3qvTO8uJKC38k6AOK97EDywuOMNabIRR9Wy3GvouDEuG0stbiGny++s6ZXF9Vun2O5B
aVX+ezM5ovldBgFnh0mKUtxK73pcrYKCvcOD6POVBZ18B91zoPVyccw88hATeN47jnHfgrfP3X3r
c0CrWx0eQxLyjM4Yh3w5Qd3dGwmjDMXORWRaDOi8vHAvjLc2Y9CElL7m/WdUg1xeYYFC4XTbCFeM
lmMaKfN5/uX95K6nZ/E/ZtW0Ffu0OO3xIjP+BnPhGLH6k4Qm6LtlKiCtwWBwBZ8rCXtmpU573lGg
hlxYRNqKZTZ+b5cw8IT7HUChDawEPkTbp7ZYgxl0Mj5pe2FUdlbqepzacoTWcR1MMdgbbTztnzgK
1ZrrLDLEaU2LISzI7o/AKXiB8CoqmB0M1uvvTMRJn0VwtYPgJz13Fzp4hyW6v7PLMZK0do6cLYXU
bOdJAPG/c+7sldKlspuy+Xaj7mDM06WhYkR+D/R3ijA7YZYTOYidmRj5hqEHGIZj6n7sqMLlMvir
dYPRvZTn7VBwBTtlBZePrtzAbYKxBPJccWffSzjLPaZBA/jd+PsLuB+MgXpZCagA8wje5L9QAxIC
sTBuCAsbr0gNgFHXSeA+BOHv+2mQ+HO/QJBJ1rQdvUnaJs9kLcXvVVsXTFKZHJkkxz+5mSzFmiMp
ChyZCvRazbmKgjlbOYrzMoMidUpYTFqh8vebH0MgDPtYw2MH16kFq7n/3k0H8Yw/LJbdaYGy2Lpt
z0s0TrNVneUJvQnbRZRw8pjbAm8Xs9W/8DTqNYdCpDHDRTrMgWc/QfPxi8Z3wFME5ICOAuBz2eM8
dAU/Q/JpPYtbWS4PZnNRfHxkyRFcCKwhLWSsY7LybCRFKQYczHvxjIzeIuL44/tHGsNChZy+QIme
QPdfVoAJs3Qe8Oe4xF+J9B5X9/z5iJV3fgvJV12WKbiAoP3MI17q0xqvwVe2lT2eXazmzv5gOYQf
L6wOaxNYxMCZsFO6NY16O19ovwSac5KtxUAvCvWNfMwa8c04ELbHPptb3mfIpqaQbsakAn5at8+g
GWK/vf6TpxMlTT2b+PkjFyiAGj4MEIwcWnZjAMCoDV+r8CwGeb1vs6OVE21fr25Z9tlsi3uWZ8Nz
V9Hj1JKNjhYr0ock59VWLGQ7MMu7hAIDDjAxWZbNOF/l0K2dmSPrxbgsxcbQqboT/9BjY9JUUlvM
/1qGo7GcjNAuxubYUSpMaWE6PamdwYjhBO104QmcN6AAI6FogLTT6gFmlN/OLPMbhYPhNwnxHmgL
es+uyMTKacOiiKDDxpi25jSM7D3iTYryIa7UKsoG6nOYwGtH24DaeDgwf7p73FRcpf2ArmBWZ2w/
iGea0wT0U4I3oHwP+JoaYpippSRgnsuA3XfvufPQZUR/1yBSP7SlJjbtVKyirCiCSj/zxnLygrkq
9V9GMy0bLk7E5Lvjm4dXiPuqcHfCYvgBLrgIoDhj6pPWSx5YT/FWne9Hsj5lZbUqdEN7OH0UBCJ2
NiMrSdVg5rMfzFUFH8MRwJ/JxMxaef8gy2gvPsgUFlQm57dVEFL9u6KlIkWHZbT4+sprElhXlmOA
Njluej05Dq6njY9wqIDmOCV4fYGsQ1qGTlLxENuSwC+l2eqzKtIhXeMRmgHTA8D4QHg5hjMY/R+n
sdFP4LdMOzc65XPYdEhKtQOd+MqC1CAb1Q9Y8n5zIeU/EFA2v/gxKnxqD1bTkALiU1awyzp+2MZb
O//agU5c11vABAk4g3ceEbZ/B2s+tf3F7CEGNWkoSEi2EH/ysh69pnun3T0lAk75k4j/mvQ7qg/q
DcrpGl+0GHY1ZEPBKw/KRWYIs8IfQCR2dxe2UcH09D3UGHfHuD8VHTVWRSDNgO+JfBLSlr22cmKS
eqdWfPPtTs0Lyb5z0gOSTHuAa4a7G952QYZnxTcCXHNwn9JUktH4WeFp1IlKXeSZwgpuas+R7QxM
OGMdn/RRqSQ0lTXLJXys9dsGPtVoLPHc3zeGs+QIVTBra5Zmj2bRDCWIvT7Mpy5GQI9IeW7zPPvA
sjImxxqDJLux1wOwg44WsaLOC1XTD8FHfCOGqWiRSZHxJwm0Qj5YlZRRvcHLYox6PER3gdxfo2Gm
TQ/X/JAKuaHjAQPk/EptwbbQRMk7F+9rYju/IF1nlAxdv1PKyHKYOHiD15xHBrcoMJbruV9Y8+/0
KoKTtk1Z3Doev5kmg+xWwNEGxPsxySXxU6TfXJ9FXR4AhtKaCJJdCmt+z+9dmNGD0W5XPtm0xJZn
YA8VfwLmSlNlb5wRO9gwWaP/NG0BUslM2bjpDkMgJblPV8iTXTWNGRFN8Q0vwwnrPGC2hKTX3fJ5
WkF1WF0uGoSYMLzFQn3bexccturWHlbwz2ImRI7226mbuU95ju4W3bcRmrz2ZcxKkhnkqyV+5HMf
ZPyhempc9C1JwbpIal8UA44LfJqDCIqWYtvQ7e/qB35/DsnwvqDJIYYbRKvW9Gap4W0yv1MC1Pu/
Qlc4mFxZcNPlxvu3ZjDU67EdW+nduKpYsHuug4G2uh9grkywGT0fQQ46dcpNwCrY6FACJE4hyrN1
24Cx/18GmEFwvDlIlwFsbhX7vKAm4dCiVLus5oCUceFJv9KmeSvudAB2pMzoTJSI96bNDUSBhJjC
TM9Xe/xKoEpUNYCEiQPFMottYm4bnYsrsYT6LfpSkHUs2JkfQyw+rZKC6jgB3G7VvE3l+nGPmZTG
5IahMSmBVqBnPzfq8X3HNL1tWoBOhFXH/WQNP4rn8U84wfOn03c91+fcIEJG6SlveWqmpBqFkpUJ
SLRxtKc9C8Bwzagk8+eKE3HYHU/amPLjL+a1pH2QmCePi0x4VqqPN9ERu9cTL6D+8MJ4d/KRyw+c
XjrD07+T8eoQuHMyiAIR0/bzJb0zB0f62z5r1olgXXF9/hyGjF5TGxTVUtoUGeQD0nuk+1o0LN+D
6CjJ138rQwiQJFSBozplb4NUUvDeJ77/XQHeouKpWB9TSPPDJ/JINVxe4rNR1b2KU0fqCxiwkLaK
nJsmxzwSv1f4FnFAvA1AMHb8ndwSplLzXtv07yJ6FEEHDZuAcdgawPOYEmbAoQ2saksxY7FGffPS
0FuePmJsKbMKSkux3oXVk1rzbZ6FzFsdSNxILMMOcZjwa1VhGhOYIzckBTpDLG1XG4JFbR/hY4A7
R+oy6IFJ3QJ6NmLCAvmEwarNIuGISCjwsxIUu5sapk/uojq6j8AFHL61dhkk7PUInj3qvKhxHokn
7J82PX82KwwY3TU5N8fRVipy2qEu8DjFWALFKwb6obg3At5tlSF9W5YPKV4lfg9yTE/PHImUXzYx
VmDmuNF4mH6f9jhWlVIToOGp0vcYdDw6In97IvSLgw868vSLrzKOd9GQ9I9HMgcNo1Vl5EXFAjhH
EGLFKCaJf/bcE+xJKNAye6BrHTYjbo6ox9sOhwxSMOeM3UZLn8h8ITKweHVL+dVRpGt89hmwlGm8
YGIWcBwFVDCHb705Hxbw6AoU2DkRaGrdSnJqYVK1mqBVAzpTAOSO9mpQPrI/2JfvQbVTYXlE0pnA
zzgpF22DISA4Dpan19Ws9lX9m35IC6dS2W6YfsHqwtEmOQeM7CI6u9QN8A/ehxsW2jb52+6ShSde
ZitdJFv0z8fSrJPSak3JlAYGdvO3YlEyEtmQWG/gcqWmghCG1t1MPT7SqDz5kDdS39vAiepeSNUQ
qLhQW98Ora9nepkroP9OG8kVy/VI8IONtd/9bbKNuJ+ak6hBmTh4VaoyuuGejIlAZ8gR5MjDlARu
Hz6b+Zxc3lW6XqCoMAXxCH1HE3MCMpLFlTGDQ0g9sGc0HmODg0dvhmyfWLLuMu1z7+BasUGA+khU
VorSuZq5zElX7fTOWtmTdxduClYESV2J7s38tjCjehbNIXK4QKQS01BXsPm+HZgblGMxADqUrvqs
I+L+D0fzQe/Tg+zjyhk13SASEEgU3b1r26kyeXIIxg0/BOZPLlxNy441m2vg5nrN63iFHOKaboPU
CHnaqg5jVJK2YxTYG0oqO1cfhCRnvgP0B4lLJRW6zNYzn8FeKOv+LWwGdEc6mAaglUMrk/8ZNVjp
Qh7NBVIghb6HEjWTjtPuHlr1a3G8TCmArjMyDODeIOEWRoD6AJNTTuWl60i7f3OenoW2pRWt8uEq
WMogK0VsQEksaysXYLB77PTPVf/07KERxKXVYTddVxPsw+obQ3JwaK5ahWFpX2cDCRBKPVKAKKiY
63QDxcfbq5g+a1Lm9UDUEQ45QqgrZFP+8s4AcHYBKyJrAZpU7jeaopkQqcxUnVN6rC3i1QjwDGJ6
xX5F0JEdRxD+g2Lw0E7VQOZjghUZvcmWwOp9SwOohT7s7uzR83Da3SZiz58dRVNI1oWSNebL9qSu
U1yMtctEzftf5n9LXeDouuzcJPqqjJIScQOqzGum04qfVO+6KQM5k40CeJMRavHhmIecj3U3nubK
Nk6Odrtl98IlJabonJGGRKNwqNb+/AuM/hCzmSaIhLgru0YboKDFusbOV7gsA5iPIx5Q1hOwUrSJ
BESplwKkzn+uvgPYExWaTtdj29lz8kAv99EcbgYahECdY2YXfeDxz6SB8D3iHqyxS2dOq1oLGLvd
PZ+QS81NH77Y3VSqNYI06Zs3hcAIX3TlNlocywg02zZ9NVtK1g+ddNZUJjbU1hS/OH3u3s4m5eDD
6XqXkHaCvUdSmAUZj6vvlrolIZlH4zhBwD9huGHd2ZeuzLGJqCK8BHu3A4tAitemjISXzPMsvFRT
xWvKPtxEVYumd5SR544ZronA0e9vYQOJr4Rnp6NlS70eSXVfC0zWul41bQ7FqukjxVH01NwA9IiH
SZA8E8y3/CRVP8gJPhGQy1l2iyKUlN+eK7LPwZG8oEJfYGoEDIwE4E0tys3GMa0UfBWMAIheYknR
wPnRvwPL8NtSxZGsQRTwy9vV/4vQIkyFIgzeNm8NI4k2q4IzyaK6MsTgByrH2nIjsEJT0Fv+im2i
z47mwp0IwqpFp4UDdcGMFmtWKIueoPlJBOiaprxM1aI2jdIAl6rqmLsIXsaEKJOmUu2pTgDgdwYZ
2PcCB212nJr6OU3VtOFTfhuMdZcVLl5DvCWqzpLl0X37C0CFjov6xpULod29NLGCo1AlyXS0H99n
EucyBStrq9xenDjhUel8XOPdotbM9QRIbOHHee6PQ1XQt1tUscyXP1uHPwHS7w06NVGfClT/JPMZ
nE2UGm5K70tFmdwRb3Pfm8ql/gCssXv4kkgYQWQvMHv122XKBMuGiW2X2JpG07S3WbuILReOC0LZ
3uiu2sTx+aulliu40PODuP9JQorGN9CmNRZo3BHDCtOWCqvLXM+Mp9YZYdskwz8/IzWkOSNS9p3L
3hHW5AY/Hff6NaLAChgTKArL+osiTAaacuNwWQqAN1I6SX1kSZEOgAST1KtQCJz5B62m7aLyFlR9
Q2N82sQbV0KlhPhHnYjDUqH2XWgkuMQE6wXw61lV5SweGzTwap5mpUbGrOzJ2TO8U97kUYNZcTuI
Ump/ENkIty/1RC6YXkMU49g/Jzd9CdGy7m2POEdyfo7JxddFiARPrqNWtu/OjaWk6+EcZhoayaNM
kXfnlhIId5RXUQlOW5Kdrxnv4z0DlVFmF6LLFnUwbTw8cUzzG0lF7tAE9FxXbkvxj9MuRcbOiYKs
Q5ye1rqf6dqjlgvxXwJFDhQHMZhaslONSg5RZn/jnAWrxL/xW6JgvGQi9ENuNN2RE+ff4I9YYk55
tblfsSQn7jK/bpfIOkLLbLsb8UnRs+qNL1CawCBh4aQgL6FvZNSlbWyCfSpuly3g2RTC+YqSf5ww
FPag+x6ccmCpkiGkGOp5rM9guHkSbgk4opF1GoDERwjHhAdVXg89F1OzYugTnKEOYqxx2uBP5RRA
K+dB6o8V64gicAuAq1PV/mG4BWJr+A+xDFBTSym3SDYni6uHpjialao+mH/0vB25PEMSSUZOWTNy
Sl3yGwi/bM32wNIFQxp9QvN3KHxVrAfPt0TliGOytZeCpfbd0U7ZUQitbHB20so7L7ISZigV17kN
SM6ovKGwd2vmrUwgNnKFm8pErgOI3xXhgd+xBRUs6cIxxaM19rwTgZGoh5bdZ4aHOOAyoyu3GpJy
PygrodKwIAZnJ6TmXqJH+YMh8xtcZsGTH+2fgbKqWLQlPq502nx7P+u/b7pOPtJKXsdeh59f+n09
rDjJ8QkZJ+LSskJOtZjN56sPI/usoY93yeMnvexUZnxLQh0jAVA1R4hWDc60liZ92dSeZvbf1TyW
RI3582WO4a1+HbGJb0IKUqBZyPZ4yPXRBE089eUH5pzToxnUAXm/qCu+04O1Uz8R5Q45onbVvl8n
tw7FqmBvulZKiP54aREGtWpZ74xZKf3P5wsYMvAF6dy+I+kywlDd8uQibCHhZobtaME9TjQ8xK0i
zZaHkZDN7VqTgX1BSeZcNgtofOq6o1iFz9AvdQ4akpDfRir5gb7AJfo6ZL7AhXfw9lhpoouG1vf7
oXae8uxPUKQoPqj0a3c06YDe0q95q/HyhIAQ7w8MOASv8Ry+phf72WLGzKvlAlY5ABLmo2fDZq+b
dSYsXUDcY56C8u5njPIsI7y0DZjqhK9UDHXiPV4LRxTY9HuVxDgiIQXGlOocW1xk22Y3bcvAaR20
SK5mONxqtvuhHeHTB9Lrb4xp7R2kphJ9vVzHBbUdiQuoJxA8VjFYa01I5D5pQA2IN68yFaqZ4Wow
aW90rw45y53kAXzyMLLp3rvEC9/tAzkagfdhRuI8TS5zicAMMtEKbMq4ivzxt8tti1I7lo0c3QDe
G3jnpsiZnUyUl4gc3s9gzEuNGlBt0C6stb3XX8OhavQxXBYCXyx/wbjzD5Y3JUf+8+fUjFmLBvJS
h/b8edAlZbb801KopsKJSleVc2obENL9i4iWWKWKxsK1O3+zP67rwqE1jGOL+Hwd7OQ3i19BA2V+
BJCN5J03REuNu4FOdMSAJ6xAsa1Y2b3ARxnxiq14AfHkXAyqfQEhFku5yA8noDMxoeYIzTzv0aMW
Eir3F/dgy7cTKaCgVVXO10jC1CmYwpB1wXhjFUqzI9AThvPJ57yu8PudRNtdsQyM1sKSB4D53dL8
GssSFJyXPlF8uDWWhsCXfrD+5vw32e6cYBbdfikZsAUQlRPM2tvm5TT3P6zC/f4YHRbG6tZl9JqP
fIWmU8O+14GFj42OckGPzjz/exNnw/V8wSk1B3KJiB7v2a+GAoipG2iWVp24rSIUyz+k1TRoQ/8y
Du2MgS96vlm4PmfxM3EMH2B5LTe9Nw2D+mfV8ioWYCg68HN4I9vTgj+LgFAwHkIAn3ytFLCOvlJk
Njrt/kNkW12HrR3itiK9mGafyAmd+StNY2Nkd1PMV68IUDoFWDVgoKL8dcPnRjhttIx71l3MR9kW
WPBSULkE/wDNnDmm++mmKzz16kSuKCeW37cyPRiXpo+d12TVawPD/ArE4C0Y98219ncIygqkTwUk
dhZ4COQGTscvtPEh+B5Vriy5H/XqYEGW6pgv9xzjPhtBdt3SSyYeUGCXsqe11vCyVLxe6+rlC7sp
SIRpJOARRRe3HuYbmWJPDZFLyCwCRx06Lcnpdijd79R2iy3KGqzSpN1nvpaaIwY6Zf1TA0pe4zsK
Ucn+m3JeZvORpnMH2zJXdc/e6jVTxUpn2nLUFfuV6tj8+jM8oZ0CDOrfyQ3O1vtOsogxdP1eZTAE
S8msnerB3DQp+hJB81/D0GWzpLKRih2Yi0iG2RQlmosPZAT1n6f7Tjch8JdmN8ionhLbXLpbGuTp
39ueOomFdiltLIyqfly1mbQGVGY7cdcGidkZrguJ+Tc8tckJCCXHj2R6QJZHAskW38NK+dNuF5i4
ILxMGWB1R1cuWaF5Uz0g3ouToyXiUhLKTY/5lY3G3qmxxiNXb8cywaCXqvgV0Ww6nYj9vZInNjH1
f7E3dx3MHAV4QNi7I+QclJckHaZNIQRzayrekHiFFCk9D7pzK5vZhG3WzLl0nwDw3KzwPt2u+JXS
m1vB1WjeKzdigEniXwcKj7AVa96tjKP9JS4HgghPgb00vK+jlVSI9/lQw8/mrtsCmlTmBv/Axwsu
eptAHy+TPckFQdpYdg+mldn0jC6FgByiat5zKDU4A6xToxmrKZj++QPbCO6bXkBDYmIhSfsBAy1p
0fqiOC6jZs2u7VM4wU5sSOzED39d+DwtqyPb9XFPcM+21qIYFuJZtcJJPT6d0GBJtSRdCQzx15nS
fwpYZH5VLa2ZFTYKWR3fvGVOtMHm46hGilCi65RWcdjM4exxFpdbM+XAlTWDGYrQzRC1iAvWpDFp
YIxHwkRhbWwe7XGdIcfXRNv2aprDnPOPiNLg0zPkhwOCU4bgVubjG6+EQt1TfJb2wpIxV/k1002p
WsXDkfqsuWIvfOeRDrEE5jvU4K2ujiZpDG8rrWFpuA1ACsLTAzTT7DKk8Y7u2z7zYh05A7ZNVEfJ
YbtnoYpSt46aDLbfDtii9WsFtvpaMPQ6s288vOo2RYZvuL9GGBncR1VAgzCr7jff+saNd0em5+0L
In+6DFJ7y9ftWfEc2bMD+5jiQdE5Pz2ajek/xZIehzsw8vqLuBtL7YeNeyY5wDYSY7miuCNt+TkX
Cqwo605KcZIw1V3VAIgbYSiMy5hFuYp/wUwNCBDpqqTAT/torQmQrIH1DGOaJrzZ4cTj7ZOnvj9W
jNL45RjpZNBzeDjgItpqwUAK0cldsZ7eJd2Ocn4wgbhA3bdGYBth+ghcDNVsmAiNZdCdnxhBlUyr
9EWdqUKVLb0X+S50Z6i1WbkUMe5h4lg9bdx84LP4LU9n4Mg7GGnp9JEFSpSjPxUZn65IQI/eP3s1
IPg+RuwOo2RgVBRtC0LBn2SVqpVwQW5IhbDwpsH9L/ucEe1EqBByjPEUz+odXHIsRtpK5boW1iHR
HxTp5KqMnpR4QTo/0QY7k6RQfboYl1DZl3SaLjJnHaG8U1Z5zcWkr3yQoOrOxhO2uDy6XIML7MT6
nRqtkuHfsoMOe2sd/dqhmcOHciZYztm5ujnk7Yyp4iL7yXWd3Zx+Cpx9qzB4Ngon6ENybJdCQq2O
MeHO8jLF79gRi7DJzXX73ZcAYsLkp5HaLt4h1uGA+5+C1oSVWoMrdv2V1qi7QOKZhcWBm6DtQ/o7
6tEt/k7eBfDw8oFdn1iGaUxWe4UVKygbX6FQC+KVzN4c7yn7K5KDcYH2zOoD26O6CqglpZbrJobm
QRNkG+ikvS0YXLdIrs4YVmOe2yY3bocimqQ2mx/v/NkURYcjazRzesbHU7i15hkVHtoTy+nhGzCi
bSuWucAu4OZT2o/UMlLibAGgQVa8aOelWaHpif8pBBDBie8N25YYlILdSFq2XzSnJQR/s3ykq6nd
BZ+lSGivqSYKtytqCs8xneB515UY0FTi/cdHT7NQAxIFKJnTS/W7MEyNNIWzZnPZ5UjsFyBtgAzN
xm6e/pah9b4zV+c4dbumnYcDrbTo4OM+LMS5Si3Y967vs8Dm7daXEQvKCH5JxbW8kd59qFoMxKxW
9z6mcd3azcvw0cG+97zCywrXnJK+7SH5Wyula67MI9mZxZDLDI0cQos/spc+TuuLTvgjOYwTppsm
sTOdf+AOk6gyxfcEWq9qqhfLZm/mrDcGwx2uBBCtJRov0tBag61N/+Rn4q3wIR6Vp2Ckd6K7t0D5
RJl5VyThOyE/cfpRS7mJC/TiOr2bY4TTwN+MrYRaUw+vVe2f03SnHPi7Icf5CKDiAPE/eQLiX4UZ
ajRyozOJbAbxR+pMjfiPmZKQHQyWDaDSF11NOIMdaW11h0dyv220iH3Ya6jbOVKDV5wAWXxlBEr3
gZGtXHWFjIfdhPBD7sbovvNMQWqOLOJyigPzmwE8UjGYS49PV1V22Fx7hPK/sfyPDnHE7Hy6dUhn
gKFdVJ/G5RVjye6B7ldXaOPXUSLrdj0Kjd5aOeC+4xOPGEkRpAID0kvrv5zzmU3X0Z8hOQmos/Z1
zIJH07Kj2tYkD6zVDImvLE82Y70fz6OUbNhLXJetwF/DHFXKl3oI6vOj0mjIEVbDkCbsEUsbnU73
tGK7EAeJqCQS6LPh8h2yXcJdUqeYhn2VmZhWCTaAWGqWIsOvWIAik2zI4kH6Yps2Wd4nlF5eRH55
eh3BBydXSD2ufy4IUnHD7RnOcTGsi0UVszDkd19QpVIBh94m7b6QbXXiEvvyKDbtzYIzJxdUpo07
i7Z0vB9gDiLLPOy3+Wtnaty5jn+A7Ahcle8+XXqjiHyerlNUqs68z0RXBsRAPccGqvWTBMbzu4jS
Ze9GpskQZnjwynwwzTMrBaQrMzR3EGTLJU5yEH6+D+ETD3ylfjIYKmKk4XG9Bh0Ry0+lCg6wnt2o
abGBrUdyHdcxdm0Mh5dekPFkMNHAjr3tN+g5J/9WmIEqAeUV5Fod6JbJoBOYYYLPQXJ2/g3oXbsd
nSWOpg/4tkbGngNr3c+W4z1r4Y5iuFfW2OXkPp2MvpaT5qJpHpzvHeOOfJgKxzjOznQmWsQsVVSZ
mvHHkCmts4oboLSI0p/6MXMKXWyeIGB9kKExNJUXaVnbT1JpKjQQS2dGmc7dBncihO79XeUC4ynk
aQw1PFrq/oOCKBHJn+LF3qANVXsUYWWDsxRFzn9IC3bTl+jlBaLLcWfGtrsgoc3ki5OQhXh6extG
N2dLUYQbcTtt+Ecb2rpuiXWmO07eGyVe0gKPiA3pCvd0hLW65iEeu2PHSqs3oS4O24+HzGBUbWYf
dcx2e2zfnVKl+B6erUbVf5S0PcDOxY/vPP2b9rtNu41WVG3PsfmqFRtCUp1ywmz3NPEtdU6r9W3I
pKE5TjOLHFNiSoaiFz96eAMDtAQD/R1PaEN+atm20h0WVOB638WwsGo+rbf+7I8s4Hmc6/T+7N3q
QlSBduuy7SYCEDYTFEuS+yoHM0Xcz3nOQQHmb84YB5RymMC1L4RvILTtMw31662LMh5lRN8zdifU
DL92slKx/iluDlVrS7w3kgopvWsZLvu1zyYtRd1FnOB3rz849+2OUjN0hA+yLF+anToUpmvRnsgI
2pszE4nY9MG4m2I+cl4U8l7YppS5Ff74J57ltc2B4lBA1ZtCqJZfz8WmV5nAljsm+ESywgsyrJuF
ddzwF71fMSl6BSwLVTVTw5CYirm0Kh95ig4XjboJXiKfpuS/2szsGDnhwE5KVfRTjvEbj+gjhgwp
b3sZ8vY+UzIKwv36uZnKhdO8JSwc2kQi2W66HTxh0fUbPI2YGc1bSFUzJLfQGD+yLzR6q7uV/IyT
G16cRUFSZaacvhqYRV/uQsT/ON+0mgvhM89ncTuxXnPf2WurVa4qFra1CNxjotYGL5F3q7Cm3m4/
2/BEJUR4T79MiE77bnCuVd8+qlPMMrkGCRXFHsIOAMFgYq20zVfLRtvXXB/tCuwJq/yriO/DRxjr
eWQqG78G8I677sJk9GQ/TGRWdZGRHpHt016PwkgW7tV9NizYVZx1eGVfEUdvYA05oeJDdmYMsR9E
rpDptNh9OmtOMMgg49qH+Czbsqla0v8N+maFkrB9cA1iX75OgBpKy6cS9aUS/3OcZheqkZtkWZpv
6MgQli8T+ibAEdc88tDsImxdWwGlKw9t18rD5rv1RqB634g3+GoseS+cW09nU2IR/CrccFFfO+Gc
sgBNzxLWgGc4BI6HAtwgcsYb8SeBXJ+k7AGBQeKYraS0g9qIyBdER4MRACYj2RZNvxZzvGm94APY
cQ6TAIuCHHE8nYtgPZQlyrVlvefIIscym916FYkt9ANxoMhUmB8YKiaTOaa5/Lzr9toly/bpDxdx
EBo9F4CSuzuXpXOAikypGphy5DMKOJjJxGBtlSLAlEYMMN/W24sItbnCTNNMOFui87ArePr3JQnA
N/27c/s/cBTJ79QDMThl7CkZzVUq68UxdnToU10nzEfExxxMc9T3INSSdfAWjMGexD9mzv+2xD1z
Al3Xc2G7PvHa+pXiL2Pei/4w/lPt8ZMJnHgOiAWxLeDPLNQhHjcw0wkKvDSAoTNG9ePi13Pjd5vk
2Nl+KtgMRcqqN9Ly8lfCzu4N437svtJ9we7CWzly8uBO/VPvEVcNZiDeTFjzdpjN9x3ky6Xh16Tz
63ubXxrevVdvype9o63Tt2UOs8gWICZvJ0WF4QoczNxn6VfZFUc2s+g+cEe5OpCF2ZyYpafJuhlP
gyC+EJBseWAV6AgokhAvxmpVI5cTl/nmU/vR78R18CYIg3Zv/F5EWnPs+QO9ptKmrCInFUG34l7B
UUItdpKUAYhd08TS/0C0vFv7ruw42DJLssL7AHeCyo0VqGlrLEVD38OPqoTETwBgfMwHuGAxHX3V
94mP9G/aZYwcCMu5xgxdYSEpa8ILSWZxIz4zLHo/BWFWSuIPaBS6DQQ3jFO3TxBsa9f9+EYki2rn
RFRPHBbxurd+7LVdu5Zlps4Ql/fM3Lcp1rnBWzE+Fu0yMZXcHZxdqz+d11dJ7g8J2IB3aL8LcjAC
QzlX9EioXInw+UM9MMNI60JpeW9L3V06OCHiq9DbFiXfQOCgTiZk3oRCSjMOdmOScptPBTmSKrPW
SC0cVYXAdztvtUOV4ToLH1+JpuFQBx8PP0r3mhaGXa4FPytUQwoc4C1uYiNN5l0PdhL2Aa73YRkl
Rmp4oqiUVszEfZaJiQBIBV2PjlTic5GuCvueFtVgTOlMdFRzn1fRfrK8QsN9rgBofHj/Qvs7z9z+
xrYscmU2fiywnReKPJLHe5CSDZgQtQXB4ukAozLNHHCDjxhxOFHoyGBKEcSn9sM3C+cn5S/nPdFi
IrCPciRSOAjuB/pnDKk/iLojbC/JBcDl+hzI/H3Bnh5gN1Z1GKB8Eu9hAJBNKUTJfB//1oAqgfvm
/M+RBx+vHqojYwhuQqqmx+fxJw0y5m/G6EsJbmm8uF+1IYyRbWGcU0DkNYO87iHBXCkmGBKBSy4A
IvVVZhWnDSK5MXM/P9Krwj+RkawopGXCNQXk6dpm4Ll5MO6U7vYip4DNW3IKPgGr0FloxjtI1xg2
UctQr/IEcHdF9e3PlpTcBtc0NLjgwn6HZuKasbTTTa+yLz2Xdt/VoQ6nFmzUQme2qozttnBuOi7r
sxJdrcvqqDldCwkWucXYatWqowuNaLmGXfg/NdPQHsI/+v7YWcP/qkpEY2omVXro2HrHwG6jGZZM
jEW+o6HFKLbNkKV0r/w3RUkqmmZX3qDqjkzbYCLCRn7RIRTkV3ovGfeFI39UwOj4zj0FHe76fGp9
XqkhjDHOFj4LeoH7EeUB8eYEVDUS2Ny+9v5ZIFdWE2CbYbo5TKDR0bAuyVxGTGjKRBKCYMkalUTe
e4ZpGdiQGpJJEBO37tI/BzVBOnc5Ch0R5WWQfP1I3SVRm8d0kw2yBUDILBYjudbdIaFlhHMnSXpm
hT65fYBs/fsNS7F5kikrwdXpA0/P40webzFsIDaKOuaQQzGpBnjucLzoSftEIcy/4s8W87kP4s9i
UX6+7F1cR0ajnwTFB+YITeNKj8LozAauEpCm3+Nj3/jOrIppFAUslkSnTvqC8PrqlckvUoXkDLep
cFMGNOyr27ZIGflBF45a1J9/+xFQeaPlHLaoFdxd/Y9xd8zx1QaQO1y7IEdXZ+EnBB1W2Qe7x0cE
WOL7PBWaVwvTEfV2WgVEl4UXv0tEJSZZDYhOdM0NrpgljN+20jX0YHf5R6fk/dMpPPU2xpN3Lkxn
ee7oNLVXedWEoEJsS838fXjOru5Zp9dQJqb7ymTnaLadpAhdOgO4xusWPE4m4NFnvn9p+vdj70eY
Cq20Eg0Qd5y9rUMH3NgoSK8yP93J7DBLhCa2DT6txnAQhCGFjVb47J7HthXj1pmX62c42aUqrgt9
Z4I2Vu/VrEwN3s5u72BnajGDaQN27BrbZq74k6E7GppAGvFGrqiM3RzqYJLgctd/6Yb54gMe+Uv8
XrucDlnQnxQb9RdF8ZVcdz/yOgquyh5vol9XSjz7wLilzQ/e1rv9ZLYB96b9yMRiNLjvZKbNBtqt
WPk/9DGBevdHPC6WisnwkNX+qLf2De4rWkqyBpKHZdKd9CNvwQlRS73karBSvSpbntbVZrShvfd8
a/q6RdL+mvRr9ZbKGn3SsXbiEupXlZ2su+A+PcaB/xpkV1uU/b+BHm15ZCa+Y8TB+R37FBAEKr63
TvBOMHijNbBUr47Xkdi/wDv3nec6/jAEbJL9baGDXmMc13faXZ1hiugm/AwakbhOrazjku65WxuM
W/zxW0XUoozErWR8owm1Pc5AJyoZ0hx7xeWpyaHkLMvM3cDmGLx/1k7nVTDbrXO8xeZDTSGWOszI
KsoI3l8IGwvCrFPGSv0YabfFjsEG262d8ScSdoTsPN+M9qQY0UmJp92o0m28juzo2maW811Jkfts
UHfBV/NcynwheZ1ZP4/GbBf/fE6FLhFWvb45zKXhxOMJ1hNAiVdWl1GAuJj1g0bXyBxqgMwyZsei
EhsQReU4CXNncUIrkxVUS4PJHtF5H9OPQiVwHDKXNokS97KF14tLXXU3mzMTSo8PYVb2YAXZqHJI
0FuVxMdWoqX7mO85nWbejSVE5yfqwnomixeH8n/jhhKyMidO9w0FXqQrW06kCqSrMKpurH/qi1Bp
nwNPHD2nB9wV8mP5o8d3zkcyG+DQIrYdFF/t/HhwsVXQisKH1MWxxE6T9rti4meSl5ZI/M/rEESa
tQylWjHWATxQZxIKTgyQh/XNiC/QRP89vd94zieDfrvB6bThUFisGu1D+yj080WjHpDBngmRXOht
YCFnq0jdmHt9RNSr5Vmj4lM90tF7ppMdUzBZweWqJkuD3B4X880+5m2/hU5Y1pY96vym6S3TcmF3
Sknv5K6D5+nbC+2UbUYCFOLoX59XpKEHGpoePc8unMlJ4nszWzIyZis3Le33rHHlxq1vqW+lRKiq
0Tf2UXFLyZTO08o9EifDem5dU+rJgKJP/A0K9ompjOvFvDyYu3BYfiCAZSnZUjc7Co2l/QYaLRN2
vvCGcfIQ+pbcAv0RziEyPvUeRoJtcn99SSWjsRgfPRvhHJVZz1gWXpXwpK/AxszbFGqQbzLU1xX8
nDKrq0q/IwficI5afh9MQJzhZRp68SG0Bt4J6eXslqqRM1BvDYCxq4v/cDiw66dmzKT1/uOUlzqr
GzYM87zm3H0D0Bu3HOJDeUJkgCgKCLcsqGXtxrvywg0bvtZGv598MEpKUcEPxi6N1HCXySNVpYz/
M/xJhiYCNbrv5Uo7H/7qJzLZ6HC3xVNjmw6iTs17V7cBrS/bEWvIh4nBrGgUc9ilSsONkQXR7qlW
9JmS8VxzD5/CLjOUoVNXaMQ1VKw67oh+uOMBrHmscD8coGX5O//dsuu4aiK4QupwjTt+5LKhs1Ab
IDIAivEoqF8b7oXqmf+9G2r9ajnQwkVdrgAk5RAYmb4OXCzWLxmQWBv7ojtUJF4FjzMon3j3QJbx
4h2odKTNtFqCRxBWHanjiwvWo+8YOHMej2TUHOjGIHl+tkL/fGPr2yof+uBjfx50E4qeRH3b08Mm
Ge4XF/36b59F46iEn9feDn6aK35zDSa5uvZSboaqSDsOr/P6/hnASg1Wz57BaLMWQSgd/ZVk7GGh
OU8kNr/J92PDIQXe1yf8ciDKxtQ28SQFFCIjgsADRYcdm8prqVC2IVEOWm1UqPFl1TI0qK7BfC3O
7+c2NhRoxGdHQAZswAokH7iFHkFxq2MlaWVQ3l6NXH1dZszmRata1si5xhIdxefcFbUNUlgbbUGG
AqcFj9A+KoOg1JNCGuy1xkRQ8Dkdhk9bT9U5nbP/Eqm2p7uINRsT3iJckKqpo/C99srYf4ZJwXgg
O3jvUQzImwLu9aPoNMpgVlbEj151KfGXiYDmigvefYVShJqBvTTQ47TT844vNcDXjnYynMDuypVW
iyq0ZtDmmSYctA27uIjC5g/TQilJhnMmVPMk1LDAxrFXqUxUTwUzqsV/0jJsPltFiUkIQVhd2cx5
ZKKxmvuDVquFL6LpGYnDDghrEwraipILqRu0TaIr8rNwjfo2h7I1hY0ySrC3Glk+fIzOklndGFzg
Ns2MYYz2KJaybq2L7nGIyd4ryiHaon8/4mJaKCzlj1hPGCsTzWKM0gcnPsAPcdkjY54Snk02O2mP
DfKT3kIiEzhDCL/1iPCk71f3jRuYPdq6rU9goNwslEzAEFfAm+y9CMAOGzc/qX2oJwEH5izTRaep
O419IMc5lIxxNDeNRfg3ugYkAYp1bkHqXzI+jEXBU92HmjyelmH9FvoU50aT2KqgdtdiUxfSu8+c
tDhF5TEYJP1Buqe5luTcYRWMvCH1v497VpftHt390xnyNdywlhkalgzlcwXA4RvAhwF/WcA4D/PQ
HwZcRf6BQdPeGm2ABCakiPtFo2aMvvZ+/vgQyrRGZrJ7RhMo5Vsg26NLZP4/J7k3cLOc2mmiWnlj
84Gjg70NXJjpu2muqOWdotuutHPKaNt5wrk0twbtftXm+cFr1Jd11QH7uc7SW21X+fFFq9tbdCY0
f4d+gZpXQAXk2rlfH4Fis5xisvcnEMNbhYAjY/YCyhrMRBWQ2JItasHCVFYiCnGCMjZzLOm2rulk
yfOt74l5l7Vzqh0dNhtHx26jj2BmW0ZdNN+6LyC6cfuspV0zEkgky90fzhGXwdy+Q9a5djuEM4/q
RfyX4jFOK4ZiocOEWdAtjd1fipJmmMhL5yMMgQt4L9i9wbnKMshJCGLjpz93nLczMeBLZkJfikVY
2+3w/wjm1oLqqRAFmVlqDyVAszUncTmFshUQcddJpx3WjlVihAsj55oV0RtECPmBopPwwITulATU
TbJNHKAVb75bIDPQqs5FbODr1qdndsHQ2PzQH62WY34Bh8Z0Ysh0R1QUydUoRzf+X6SM4SI+JYK9
pp5osvxfnUyU1GC/XMjmHj7HJfPCoBQWeuaSVdNNEHiH9kk/jaBPca1/95e+0umekzX7VoCH2lO8
zxmCeFhFIbbWAIzaHILEwqAh/2eDaCOuHdiU+6KvocsymChUOVamZQphOmhcvKs0Wtutda+RpsQx
OKtj2usJ6d8fECvg9czWxLZgAK4VeR6rr5biY8vBepAikku1LqnNMNevMYSw6K1U7fHktLzvsrBW
OTRUXspwrzTsX3b6iqbUh3D8L2MElzEcdcOcGOZidSk6N5CW7gsomKuruhtF+PqOj/n4ygiV/Ixh
SGLRkft929gfEgDAeSCG2FG55i7wrf8KUp8XaUHWir5Nw7f/lNnSaT2ZPxbKC7IOC4P1M2i750AZ
VKANQ72IDuwJFCh9iwU15pIPaE2SdFy822xtt2hsreZx5rGK0qCOXMktkvhkvzz9mD0yedLkCfvR
6oPqCDhjbtUmgTw7MTjLW57Kk7x/BnSSgeT5RRuZcACdHHMcgttfXopGQAuzMbU/gzR98Tqt3uFP
mzEq+aKEbjSfXcViMFRbtJHimBupK2fVuTq4Tw7D+CqMGYAmkUrAozk9JpeacFfItAgtt3NSYQnW
cZR5c4HxTZmnVFyKT7x6kGDaz9SuxbpyOHnPUm6JVAo8bKW/bgWVWnnA78CxmiWci7yrDTaxt3RN
fchIuHeEaK1yvcxXkZ+YxpY6f8ygCEYHYt0fhND+1OB5Ti6aDwcmQGmwjgIFl6JiZ3vS94Tb7yzx
ySmQGhEsbEaXfCMk+1HVbr8A+MM+kkcv8h48pXf+B/QW/gwfmMvY9H2xS4o11p5fps99uWbxvfeJ
b8ZePB6k9R/pHTDN/YEol85DgNDWUiENdgdFG3EE8oARTzu7GV+AiyMvp9liJ/AuXYcushhXnuc6
gk7bPB8R2f8lRAe4UKHAmQBPX/lprABbHYSJJ9mGKPbw+UEpeuQyVaxtjKyZE87uPmsD7CqeHmgS
7qGrC5H5vYVNamEXwDSqNYwX2Gcf4bmwHQVS9MtQbn7uxFG2eQHJrQHAn5pzRlVBckwUW3BKk3jw
4YHRi9zz2HbydM7vJpykXhz0JePKNl7rkTY+bRrFkKoOzQ3LuQ7RdM1MwACUy0xouNZJxHj1NBb+
S//c59j3bOgUbAzlOIxYxhU5wkYdsW2w+1a2tjp4HF/ArW7PKsxvmcYHTyL9EGuyIoe3mLTwyKsS
l3Dt2PG8s3OHP4UP6vwqu4OH0WhqDhH+EsvmwsFVLWoCFPS3Q8aUKhhE0ULSIKPLL9p5EDNYRj3U
JAWCwl2anO4bUG6tGuinLvoKD2t6S1wkaj/GQFtRhlTplbx6LzxjNrXFyrecFWDzWTNhhfMTdGe8
DGUArcF4fNdBI9D/DcH1B43G9BaBlLL95nJQUYKvHpv8GG/RnklDfU/CsXZh8MdiFVlchweQ9xSQ
nXslHH0fZKY0Zb3MGjyi8ELUtIlVGZyba7iTxteXTNYOSNBbrjW/+jt0csd9e4VRm3i+DQHIsveU
IMdkJptEv2RgRFxgKcyxyEAjJsHzoqdW1MDYNFeMBF3pZnlfrsWzydC2wbizT2RXqRmB166iyRL+
CCf5vjwTack2Ji//Gg/OFjWF6MuRwLhojemHBgDtoXNGzfuibnDkcwpC2ZvxxJGsIExaKXxrSGzC
4wvE5jMI5twHeVAd6b8BYzw749up8ymZCaieALZKVlwrrVopYSXwD0b55VqrdJt/x/Tbjga0IkZ8
ixpO2ojXFwfGmy6haejby7+1K7uVJglh2w6vVRpuYOgZ/REawl8OPDNYX8VyUuScV69Q8bEsxrWE
IN8mZAj1QN5qTqkyybnlhCeveBI2nU/Pxu8iv+Sk6pNoxXkomBS86iE8aouZ9pHO0LAjUPlzi3HD
/9GrZwq3pNDOWe/7ox/zCbNg0AAGM3vY6aXRd8DL/3YewCgl5obqZ1ccaRHhgxrDC58JOFGE5T9k
q776AOihgQWEZ7h6+qvMCcg7/if80MRO7bMVCoGRwHggiKditCO8DL8PJGfn/7tDqvdZk5JtAo09
BP264fUXxxRz8CTCjbYzxeRX8TxsONdJMGkqLqFXOmbLgXUfHtRWV2sBMJprseGkXmnAUJqJZQE2
Y5NB4f6jrfKX5Of2LMtH2MQ08BTmIgQX+uU1ICUVdy5CacC1JrCU/XgnmZ4tjUS1ZKB03zAHO4YD
OLnSkvPl+w+anQSEyVYGY9MXkykgUW4HEXtNv54PgAJpqWc3IBlhWb5wbYwCVjyOMf9xRBJLLOoU
wqf/sqj5oAoplzlnhjHvJcXZxJfNcYzTj2uQZrn0B9b0RM85oWqlCLqZ98ljW3qvcrsmUiahXdsS
0gVQI+2CrVrvr8nOzD1921ll0x2A9uvm1bVcTtrIy7J133B3AkchvnkmgLrHhZOFBLZWKu9e3teM
6nMLyF2W9IhCAI6jurEIj9YR9INMWkPP4qOMKsK7u1F+txw7oyWTwROkOkzSJUypvvxWnBG3e4Fl
2PG5U6uj8FmMTQhJ/V9Dg+R/wi59bH/+bJ/SrtWTIzPcTqZ3P9btManKCn7X//AwZcdLad5dXZz4
lVfRtQGFwVEeN9cXyDycdEajU82McU8QDm66ABzRyngpXwZrbRaLONS1NIK0jtqQVKh9iomTml1g
Pq4PBLO0Qlrq2SN3D7CPlMZJA7Q2ioR4oZYYs1/1/UDWqvTwsDpjWJqvgdxEY5TsZjyVpKYgMdM0
TZjJppgm0YZ7S4hRJh4hWw+nuJU7XoWe8HacqaXIXPP5k0OlSIZobm87P2RsB3OHUsfTfPghvWvp
X/jPHh16aLVeeBU1PtmWCxo3EW93nlgwx/s2AMYFMAtJznJVSIrXMabTKvLzgGLn0agHbFyy5MKw
AqLmogC8Rndi8jFRWzTwSQXJ1zED+ol/xMXYpc8TWmhhSez/wE5AwszTTIDEJ1KO+OprPoMY8iCi
K5RRuN8WkYk9RPJcApiXwbe/aHUWDdkTMOsHkkPbtb0iikTurYi2LpkWF5KirGZL9dS4ZE1fQzV3
Ph6L4LCu9e8iycoBr1ZYxOOva4iqu1lElJXkPRtIAVJ5yro5tZvFAds0IMPsucnfHuijm0NdKmYl
A8cQjVcu4HPbvB+qu4k4+B85Ky/IjkB/bEq4zDIdjkYjuEiuYxpfqZyGnw95prW560p4pQMyqnOx
B+7c/EICXjx7P4w34N+84DYPjDMGlCGAMWHgTSzSGS9kuwVqCUfBXefdWFo68G/Vtf4hM0iEKJAF
E+/ZfvPBXJKqh7skcPeH3EHOTSiaRB024/jr766+7VBLfJfIVZCqrpm0CA1xKTeG+fPaGR6gu8xp
8r0NkNjfxyHBM0ZpOkjGPZjWVTH3sWkNDkyxI/LRQFwVPYLPyGlIaDZ7/fqZOebJS98NJx97OMHD
hlTsKQ8c07yOZfmBgZOb8xtBfWPVEQRfGZbGcpQAdgOXeMwg7VfDLDgOPHULTAM02hJ8uqfYk3ff
olDi4o2TGEhqCNPqvv3Yqg5K73zxrFtixpb2hKT74D6UVculQK1ZtXwnFGUhsnTVpg640cF7UTcY
gNEYt5polqR+ic6brZjJjhvF8tgTlrWaV661bdUvRFJydq0HsHTmsmKWUelMQks5em0wyDbokZJ2
AxuwhcSudZY7tU7K1EaQ36z5xOCR1A7BUGrS2XAMygrQWJQlWvJx5kiPssBJvUCO7kv9SyWPT/IF
5lCtBsZg8U4UFc78eVJtfOGq+7AeTXM+OcZda0Jn9Cmalj465gHZA9QwbIKUFUSMKN7lsaP4v9IY
trAKehJV3+XCzAm9pY7zSs0m4MJXy+iOyCXAGr/gXBNHBoWv0Ymly5Wfbx6PMYwADjgO7PXPw9Pr
MOGdK3RNjcyB4AWoT/ttOweeaEEN7rAO+ALx76VsDh1EWQp4Rf2NJkxZz2Gf+M3bQHA7Mbit4dOZ
V+U2Vd2uIyZIlglDmiS94IOcBsRxSahYdmurxm59jN9L7ORgyRHKLKNCg5xAW8/0HrL7KNQPlF2Y
yWT3CcjZe5hJ9tLTqslW3Gqxn1NJgyNQZ0BFnwEb53K0ClZbW8roe2SArcW90iAiBum/+xP19Ksm
9Ma4jkythbkBojldkG5Xn1g1Uwhr3kd0vbI72zH7NNde/bdAPk75xdd13wIVuvVhJkiy6mkSnsGQ
FsjTtbA0wPGDLcQ43UkRuLoArcYX5Y3kaS1rM4wX7yHEjCjA6g32R5bMjbuyglJi1PlTr19wSA8Q
Xd8ORbnFaXsiHIBs0Mo66k3lEByz/wEUGEFmp7rMW20q8Dy42mq8LXIUay+zMwfYyknbfXrk3+A8
sxkfOGT/mlnp9vesKPBYlcjgkBbIYtY10SCZDjurOuBHbl961vnBj61qQy+RLAdE8km7Sip7+UEo
Op+sndaJfPWjhJSuhN8ce9f5mhV6Z00+lcQ+/1YxIbtZ7JnzPDIGxJJxKC+9zudddkxkBl/v+qn9
caf3BRfvfcAENvfj6ENLO5mtqAc60qLzagm8adGWBU3mmSB8rgh8JhowbYzhnf4cLwUFRjGjgIb4
Be7S7PHAQ0vgthIsKla2QXqvWzr/osZeHvtOjHDPtaN0KJOwg9eLi3kc5WC7VKhFF6o8dFQoB7LE
kwiI2MYXJLjvpP4m01/1ftmVAHQ1Zl1Hc8QYNs7d1swkBwjThCfG7ghdVwGscNmycVF4cHSqjrvh
skbay35UwOYKrDQntRPik3zacIdjJUbH46oRTQDHZZ9flyEH4QGGk3Ms306wHJD2rdqwrcy3a06D
uMEDSK7keUTM3KUpn5bOcveKxxZYNHTJwaCTyO9OKUedhFXiP+S0oAH2PT57pkBYDPZJMcfAawUh
iFTTPNWAmal5V0hy82a+n4YPtnsHAnZjtIR4ETgXQi9nVgjZBixw5tCXgA6SonjU/cFMn7mrWiCC
jwas+9S2JAtlm0cfcBjbk0OvBilNlQ7+RBt2j466FIRVd4vFEVKRhylcK4cTvT20pcN5wB94VN2P
9lf9Oi2ssnN6iW9F3HQZ492B6kFwGSIZwZL9kcWhWmPRTf8UK/+N2TFbDtgnhM7UGFCOKzZHP7fu
sNmjwWB3EPXyZL7VguHguKPorp/HYdyRuhq6PHSS4e/vYcWuwJ/I25bBE753EhJRzSsJnJEl7M88
RMgTBbxkiTqdwSUGu56RR2T88hbDe425NQ7LhkNRiBkUJT53vTCC5RsUNeZlge1hpG0PZ6kspxNr
rBFRRr1KcNz0P5hi70sImaxc2s0W6f9bTtBI4yq6rg2mT59wqsVHGdofv87J1+pH0gBUaIby+E0m
oghdCcrP31URNhlZcSGTJ2h4sAPKQ1xXsJyHzVmvsui1CUqqYVGpfBEjaSzt7G0nVitYy9yvXp07
IR1eqBjeUWl8WY0+y5Mq6Kb2e4lycesVQTvmxaU308u0mtQmduE1y0ir2Q3K2T/qWfcrGvSQ++tp
rJoR/XfWpnYg4Mhq4qiz4YdJlp6VP1H70G4iEHaxjvJjupsTSoX/bWDnR5x90haWAbs3wESoGeaD
aQIPMDXfIIDJQ3Ze+hEfovCGgQ4PVDQg/P5GQR+upL6MEQBZtseRm43fkAiu56jPNz0ha75SRjgn
ZOnyrXV68RXYowN5OIhGnWrvtFXliA3ELkzqI+o3rUZbUYC5S4nsO9GuJ/eqZtsYjCUpPAPFybwq
04sXiJ7zGByQobatcO/Rbqw5BHqxym7AsxlUG+CVLb5CtB+9ApD4J9dpLrmdGhR9k9mzj9UmqVSy
kSlbbg/Ft3Vyfwv7yWBeGa5yDLV1wDMXrFK+fnGaR+M4qhfIM+dp5JczVxWqNbLPIDz5WYXWBq26
9mNCiDpfNcb1RfXiQhgs+BxQ1sfJ8P0rRznTo58Nzj+FV8mg6rSUQlChlwLi093on+oRKUDK0E5r
DkO3FHOzXDYbpaNXv5tI8zsI/qBDCN68kschZ2HF+zvhQeWc7v8NwCH32KOhzoiLU9qVduBf2c/q
GZ0x/Vs9zWUOrC8h3JSkhGmRzN0+idxXqyffqiOhNqicAuXQ9DYH7F8eGi0HEZKChTLaKzW3gx0z
nGcoT4R+XpeNApEXB6RpR98/5/7IaHhNM/IC1KYPdauLo7PlHviE+rJ+ndsIuxLm04oDmAOSb+qv
9HluE5Tuj+8RpPK6Uvf6wqqypp0Kwf1WH3hBpSSuf8tdjpSDGzgK+zHpr+DRfBdxTCYwpjwadE0c
JH2ss+NgEphzky7OLa+IazPFwB1hytAiHOATxBblvgwvCfS1L3uZEzACrbVYSnMLszIvEUQgHWGw
OEeiu/d/u74LQ2ukgbBqCKRwzPrjbYMnbl/VZ/KTPrM1CNjfKHHIjLMNoyaKb976OcqvscEF2Qpn
vk0RGVnntG8UraQB4/eTvNfagS9Rex4aY3vbYuCPX+7EGYNnSgwumW7EamIwW1TSNbsMN8/+D84S
73kb967+n9lPcoBV+V/OWejWc3xH0p/4RKzpfTnESXtnUsNivGfBZs16gmrlRXhJPO3dG3EfT6O1
0TN1BxAI0bFcyY2ua/jhvJThdKMx+yeIEaiE+5mimKFbD7Cb9hnAGTOxiFLXpreJra/lIU074xOW
vA8AcTm+LB9N0h0W4I2UQ7WPygRv8T3DSkrFcZREqP5xx2Eimnirg7ZyrO5MJSz4rY4+khLWdw9d
UnPAxW6/5VQbuaIXrQdW7spawI2hAljkHFH9qq5r5EOM523Nky5kIjq+mgvQzBrdEPjVHIHDWRy1
wyVcrFPCTfvlw2FalGeWIqwOUAIskOnBC4ENPWeIiy/gPdns6K30hUzsRMGpBecPDonUxbRfmQap
raSzXLqTJ+5cNC0bpa2A5BpaQGo13QcEeAbHB4DZOgsQC36nlBLxArfqjJS0JWkKp78lemi9+eRR
H7nlW7eSI1URJHVy7VGAxRQdugZtJ/wiObbhX30NbIfZcwJQJi9WW3JwnL9fHY3lRuVquqX9Ddj3
97NNGX0JMHUeZF+itqm8chCBUBysIwAYK5kF1ut4x2MwOjjhDGViZnDgplo8CORqAYSZ8zJX2Gpx
//7RIdTDThDOawBU0q1HXxbAZYyV8X/TDVBOkH25Z3Lf9j1Dbbnj/ZtCw/Co+QWu6cd1Ceq/irX0
2Kt/HaqnC50D20V0l6wgWa6c1fnt+P9PtP9DiRPJ/LuqodrHR0mVCzVVUjiL4brJPSgCkU7jsMsY
cbH0GqCHMr2sEF62vERXYyCbubbG9chLEc1MWDCNPUq7DvRXAJXk9ZhHTBE+gDswReBzdyz6/Dab
jNtAJGIa8xeXJT/oTGLO5nJWTbBFX8Lc2iYuYuhwx5xox+hXx6nMg6pvvyMI0/ruYeV6gDBMvazH
uQVCJSJkapLjr9L/HQMZcqLE77oB3ivVQ4Bmzj0KIwdw+XbGhgrzLB59U+fZHDzf1BGHXCxaSZH5
SjwkF4yOI2O3jAkCQCE1gQmhdqx3WmHBYQ22u4ZCMU92AkGL8Y9YRNW5SUlBhNEi1Jb8n/QOkcFf
ZMkO2C6xKJj9EXKukj3HbZfpAcsGexVD9lypVHf/CJf/3wtDhEUoQZnAzUxr3im2SrZmgdrmB+e+
UjiA4OXAquUCux3lZ4bi9Vekyi58ASxXDTlLGVzDT83A4soxOZ2miH91hDJFixASWdXk4+lA/XFd
1JJrl4DlsLBD+pnnIgyJ5tAJAe4XSZ2PmvwPXE0CnZh9tfwPYv51/O8TTgpmFFSMRZ9P3do++l78
8VSIZ3zcXxdFQ+yE/cCdOHhYuNv6xqOro44FxlqsQn5K/vHBrJPH9dTWRTxCIALNCANl4aZ57VMq
dsPn2yYcBht1X+L1LqYqFahEvb6rijgwNZaMHFyk0yDv4fpPRfWVe6zCT/eTUDZALecBkzKd6V8l
ExNMqja6apNZP2Oh2RKkbLy3HCLBetpNEFtU09olZ4fXTL5rsd5599GtcQeQh525DkG5Vu+mzQJ1
SEZrbitkS3t0Ntf39q/gkrfXWhCoqQwXAB0T7ykftfE4gohfMDO/ozzvgssMqRcF3PNdeFQuaBgT
NMb1S8THEVXuUrbIc/aq0rMgn5yCGEHgiOsrIsEn1KXJ90/gq2cjqk4T2x0I8aelLPd/4FDlldaN
0V4PDRRkCwdwFdBtEZZIZ9vhzkTuFw0hHZj5U8mJGr14Ula/B4eFYxaIAoInF4EWsvv7P/d/Bft5
YHYEmqo4THiM39hDrkObrD2SHZePLREqRa+06axNkVWsXT2QLgvCxTxQsXusMNLqtsqs+CWhmaMU
sAt95u9TBI+gZ9x5bLM/r9AKG/d30LLFFFX0rZwpRQkuHJzZwuyuJ4qq4cCnWKaXgj5rKC8NdTXJ
Z9WoZbMf1+nVjihhsOTykJOHDJE21whCY+GYqgsy/CzrKxbRaQ0FwcqU3JW2tWmZIy18zGeumn3k
FY/uKZtjXz22/KSTV3nAnPlWHP2QrJid+Uc5Aw74bUxe74KN5+Mji5685IAiG459L/1H6hS7lX/5
4Mc0Mvoy5nxRD9uHG5Zyk1180EVkuVFahK+CS4ynz560B0740VrjzbuISvHs5SE0fmpn01O30191
BEnjl5ZkWSyb8NxIJpQSvyZw7xrsy3w1wn+PxgZ6DzZXNvPzIEXCPz1eDBFhn08WEqeZXNgmkIU0
BMG1JrWobA1XPKqXcwQI9kQj+QluwYKK/w2uf3iUzv2V5LYFQS9MrmPInNaPtmSl8VaBwc6OhyvA
pIFloDhk2vusyW6auE48Hik3g053wPChS8U2/AkVx/sMIsIRNe5c3bMTjEd6cUcNtWONpTtVhbLP
4KTPE2RkuIEOlyx5RJnfT0uj8IwkMXCskYhY5Jyey7THA6zv3kKYJS4iMsY5BKyXNwR2vgEZX9PT
4v9VrCrC50j+nMCV5UfEbLVFLGxDsnzrW8t7VWPrILfuYXhC90klSGFzC+lHANiZ7w+3fKN4mFda
D3GgcQz9L3PLDScbfpanOaYmxMGoyf7ueNW67WlI71NZh0/wC5mciDXTOcjRB4Y3Bpy7WNIr7pzq
8zXNBJtNwwqEBRWS8IVHYDqb2VvMTZsGYkzWThV7PsmOI/fT+YvFj1Z/HVkcRPplIyY/ogCLmHop
MhWFb+yY2h27/eBXBG4b23r10qcvVJTZtswqFe8Ob9bHd02k8bKKJ3MJjMVKJOVPLIVqgI1mG5jf
P2yD0Tig8f+6MTBGYnKWvyioyL9SZk3P2LDgZ3c00nQhzO4hyCTIesJt/+rcubUq8pG7PnyeMSQd
QXol3FOMpY80nkLtbdJPRLNn8Hictc3ojj47YXj55OiF7NWxLnywIUGEjeqcejXdWRkeivNbYX77
Xq40+to1n3DTtQKRr78k/XPSvOQZ627e21Qm8OvHe1Gi+evOniDnezPGwHzZ6F4vghq4ntkdWRmL
jP3z3Ukp/lPh9KphHVzW5M9HWdbSftjkQPME8dsHdgfDiAQUHAEK+W9NlqMX5GTJrUz/fNzTlcwx
7huLiUQIMV79UxXuquUAUhD7PmAUaQ/4Z5b7yx59LjaZnoiHSM535qEmIrcFgN0CTFHQqEVZ3qAy
uj612OfOxU7RZAHBKIiKHMSh9CJuve+DIELMPzibpveFUFLBGwz8vIW1cDwr3dRw7c/6wgYe3zDB
ic4mKClf+GlFw/f4xynKRKMQekojV1lb4lbt6lDgEW27ScIxtCmvnk9uhCPG9KvxGS13oNV6U/Hk
097uu61PmWkP+CmcUrUHJYlnfV81EljAOTMkbUYTkOM41UCQGodk2Mq1vjPVtM2+1YpjceenurGS
BmtWgdaG9IBcz9Y+79QFpIislTSyV9FF79EbKFR7/uowb4lPjpIdv1ymyGRXlgzukmYDwLkThrRK
FK7OExqDwkDKMh+Ul0QwhDmQDomgqr5VzW+pC+HKOWTUWWoFUIHAHvRxYcoPYtgAK+RumjbPSp0S
nqgJsc2PQSS5/eanRftKMtGYkt2XrutLC644skdcBKOTGvLndAT2cSaL5iiNCujm5rKygAMhu/50
OrgBVNSjZr4mmYeeKdDlmP9v9xR9HjsprkW7E07DC0tSqSpRkpU9oWHCmQOLadAH3GGzqwALrWXw
fxEM5ULrMJr2EF8Wu+W//kvNG7eUbitYY2R91lDGK4WzH21LKScXncTp8Pr+OZMbf6TGdNW90rXa
ycNo6WXWWguEXNOxhdMMl7baa4GUfNkRyriuQksqTHMYNHR8tlEyY8uWMV1nb1eyfI9x5P6Cndfs
wsNRm6H/UTuq2O4l9lxtoLRybCM+d4PtYJYfemm3p8I2Wg7ACZxSFXOG/BfjvqJwvzrs5/GT5aCR
U2iIO1J95V6yeO6xfRZ7C8Rcodzn/yqE1pAe3CtYbr/rj5jaerJz2QLZ2yJMJEHqao6nGN9OOw21
iCBcAt80KBd7E6SC6Z2pSNRXHJuggAEOVGPk3s20kq0LEjZkQwrF83/MpVCj2rjiDGhJhNklcNcm
VMze77WnREww5hEm0vyfx/wNJGrTE/cMqQ6K/CenWEUvhMl4b8vfZQlKCN03uCfv6DF3yXO9hfb/
xuK3zkA3nlm7qhuhvxBYmgkmC0oZxDzir//tT/UQvmmrkYjCoI6EKcq7tSCw790nbUeCNqSwEsi5
ROBKRIra5J+P4IHpEbS8TXeKcCOWZp0t/TNglGvd8lw4RqMgfR82SfgEF+s7J1xWberkC1nLMQfF
p2pIQPGCkfAJiFw/D0X+OKhtx5Ru8b2gRf6IFtGeds8hYGdP0OLBWSLuWAq2Xk0X1hvFXfzGTa7Z
WQ6KCtHu116xotmBapmWhLmy2BhvUf3+lCvljufQqB2QQOPa9v9aXeQEVOCnGwk+SNQG96YYF+Zb
JLkEQtLMjYw996PdobVZuA0XjJP3IIU1D3asg8P9w0Mpzp4xKOvlxQUhlsXQQ0K+9Dhto21sKzyJ
MMS+X/BI2ZkNdpKn5VFU5gtvuSXAaMYy5H64p6OuBDiCyvqhzrJAsyValh5gXqvo6FW+NysrCOdl
JfMEqjrGWKroagowx6QzyJp2zc4Y5FrFG/k+tw8BuL8GgZxPBPoL82OyoCLL5iPY6Eq/JPAFkDTk
Y+MlRVeN9tbUK3YTta9zPrdXIZMaZnszky+T9VWqntsGNUUEMbw3cHOm6wgj4MAHTjmLnK4jVyFg
G6AFqjpxJi4f1HLmfG4mz2CncAxJ1BlhT/AigVZMWgOWmHDWetQH4OLi3vHD1bbH4qjXclQcmxYy
PS5AQ4fiYVPybpvgPRVkFSQn5w5DLYrAPoKwh+SO8muxuZRCG2u9pcAvffEeAXtt5HdWXYeIz+T3
Ki3wQhiQnxsOtx4VPI+1casChloGrLmbQ4qf9i9Dp4okKgL2x5b2r1+kEI4tgksr1H3u1qizutQB
XgowhNEJ7PglUor2s0uhuzgDjF4uKz8dSmR3bmHGhvLH4sbMi1qjjmIRR8xNhe4NshrJ9V8xyxpw
t02T1IhTI0gR4Kd5oktf9sNPmQZ69MY/i7P+FRujZUV/EaX08UtLlmjEIGEQl1mOJppIDhbB0wFH
i/jVsxJN82XLrRylnN9k5Rj/NQPhjmG+4UGIBEjKjIaC0XRVBNURXYCQQSb/d9iSRfwde0ExrMM2
mbGZRiaIntaxFqbTNkWGOiLeC872tV7XPM3inNTGbZ+fLKouNnAc9lqs1LRfawwfKizST6sKrpI0
3LqTCx2rnw9Az6Gm1bhmGmis+LCWJehvbZMzkYEK5yMcGzXH6SvG+rL0Ml9eXMMMlHUbVn0b3cfO
mtgxKyHLwnlwlYJgI44aGu6WwK5DciGFpL9JOYcagrZMTZBREIj3MYEG6WlH0OLPiGMqWAHTuIST
skkvlIlqkfQ5UdgiypgE2TMVLe+qxM1y3w0hJuzDjaDeELaCC32VhoBcLWsUgilqLjzMeB7aRIrM
n4YgyDkE3Y8tkjsLPWNWm2xvPIizYGZNlHApgOvpH17osV8Kxijo5a1fVXohuAiQiKo5yjSCLKM1
nr5p/C69M5HFwHwXsm5lPF9Y+y9IMZFo6yyIxgy23tbINyo1fNGfhjMn/1KBNXMoMCZp3/iUzl3L
cC2beNJ9TqHlrdgoNL+UydepQQBiiYuJS7SmHlgN7Y4ob6sZUxsj1w0rVgADrhM5H/UnedYUb7Vo
EQQ5p2pWpDwspJAAcyjs/9p/RCP6D7Tem0S5dXbH33JNwksqOqbdmy1v66RKyn8Epe9yoNjgBiUf
lXT3pxMFWkZ88uFMHce4NdMEujFjssDVgvEKqIKkmHuyieKFGkPAK9oDt37h0j+QMpj8poeo3iTW
XVwraNVjvwjN+79QDCStgne5kVh8aSt7NotA0oi55e5LGC3dw1heEePauE3S+ed2wGeDOsL+K1+r
+f+E2tF+91UgKz1TmJ4GXjRK/SjWaBfPWW3zIY0zgcQhFrCiO4fbtuOMM1SUDdWR3FnJZZHq6wQa
srY4YVDhvKOBHWCxXXf8sCGtO/nqqLgS9dfVrPfIFuEZQn6g98VhTnWZ+ZJADRTlET0vw8uzYfNC
40Uyst1kIjSxsAj1K5iaDLWjWjiXXhGmfkh4oH0B3jV9VZn+At/7MtfDR01E3QWKzvzOMaByr6Tf
JpV/Pro3QW3j+Y/R9/csbDNjtTbJno0oAajXIXljtPmO7SPyswJB32AObUDIpjvMprL2w87b6eWi
sMmM21EQ5t9TDa8go9I4W7yNW/LlNxjFzhPwyeubiZryxcKU9d3fkS/G5pTu13nlqNe6we+mIVXo
bl/vmA2GaybP6fDdYc6NSjj5xYIfPfijjqmmKGijkwphV7nwTJlZrEG6XJRM6dTWUCJaO87shA1T
DnI/ySfsF7xBZ5tRMI1BqE1bzNeFmA74ISF5hhFUZ4rf3zx+kzubZte3LNGwuVvUZjpbvEfjOLeN
a1Dc31C+aezVGB0sna9Te2dgR2CmgkmTkPgGH3k9E7iVjcVSuRAPRQehfXXzD0unnB9b2UBcsrdr
L+zricQbpATddiujsCi3949bNVbGPHmhXnpjrDNLmw3gJY3us8gFF9DiBQt+D/L/wuv0uVeCSEy/
DqdEQqkNgmOjmiQIo0ut3VkkC3I2hWwAWy2aOd5O+IBXngI9hmZ+Uk55neMNYg7RAvFGpR+Qb87F
bLK0ioETgXLE9r+n5wCq2NotyVUnuilUBX0PFvm+FCDSMMWJAisX+ZQE3asD0OK7Xic8FDA5MRoD
ywxOqS28TXuJthPKEVt1kJiRN7VrKF8TSn1jwWDwQhRcQ5PgvkxzKOpEcYGfqtJ2d9a5JEMuQuvp
/aU9X1mAWcf/4d07H+g7WG+yJyq+rqkAjSBEXYK278OT5+zKzo6TAES0Uf0vmP/Mhi+6xYpJn2VS
c1oI5pN1OA3gKEOHDfUM9KTu93PwybyxQJrT0btE7q+3mC/E70ATC2kzfro+FK/uuKsG6afZLqoj
9eKts/2s/JsRXofRBHuPss/EUjSsCHmAnDlPbgmSG9YeuLYAa/KQ5COm5bE/PZWYLrHZhTbbmRqw
2o8uuG1b4xRHJfHvM1kPdKajgx7HLm7rW7vVQxsY/t4CO5m6hmpxM2tA+EZNLEFhNpnJpHeIK5tf
cnKPproIT5qr2f2X1DmKqUpCkz1bhBuvhYI+AqBgnusl802FnyTVw4E+1dp4NY1EFwU+pmzPwlMc
mdCFnUICSFrGLDtunNks6ziWjI/IpKUinPdqXHsLPADDZnYo+DNbZ3jURIGMa2eeu+a6aC+mx6l+
w+T67cxWqkTr145Fh53ycUyvv2mUXrT4r2+7bnu1BbrMtAIO7W7TowX3Y7WuFZQxHz/CLfDPs2o2
poh5vYoTt1JHV1KWJBgP/jz79t9d75H18J9rowkJUWP3e5AqFZ2MKitnpgfAHyBWeCqoEW/1pPib
hWF6XDdcAjuJ/cXCluH5qIP3naomYrceeIc44cK7F0DLrPVZMW8AoWD1k7PiBNsuByEgUMPT07U7
DYwst1LEK3LJJ9qjSsDqE9zuSAhuhZidD3VhLICT8QUWBsXpbblYA0JqE45f1dRzT04MXJfb2QG0
sii2azbkNuoLkzO2/HlyL5IbGaMuqp2nSkAOmOVWKX0zTYRQoPXiFFAOKtcAJppFW9wDaaQ+7lui
wB1A+v4CJKr3UIrlJ6NozryN7t4PAJ5JBURld8EpH8asT7t86ebqrH/m2eXQYsFpY43o5Y+i2zJ4
DF/1/ZwLIH2zcKQ26YRrZ/1OuOdTtqqj/4pB/K/1RIl7hKFIQ3/rB7xbAr3rG9pENgj273lmGVrL
7tWizShgTsUTktrdbBxs+6ag/EeSZgjqw5suMpe0tTmZxqD2XFwYWWCV/iHAJEWb1ycEswDpK56P
tRgwf4f0XkX+tLn8MlRx1xIj4LLr28utASNhxY08lauGO5Vzyj1hvq7M6UykpMkpjdx8fzNfUiXx
7SGHuPdjcmDQ+XSrq9YCaBMlM95KeOTcVDR1topeLx4L2yzd8zIB7hhD6d8B5AGhSg0f7Z004ffY
WcxY2v5WaJypOIUS+SLAYkJj8h1OsI+FwHaCVPgbNc1auHJK4xOl/Es81hZjlyjOePfQNiOhvFSD
wwjCLpgo7onhakPD3pVuyZSh4qKod5hWWTpvUUUeynM2DSHj4K/r4oV/Yn1rrUINvMfd7gLWwbjE
axLsFbx1Ll5CWca6+wEl4bv3FZBc/n1D4Ad006qjRjbi1CW8uwAYP1VPQ2cY8BWfKVuqbJOSLdp7
z2erK4RkO8Im/hohgQEe0FOOaIUZsyAP2huebstKWWjbVXyG608Y+ociqgs4Skml1c1UOIeao9Oj
OIuCbOofDC8BIc6eRd7YHNOt1Za8JSEKv8ZfBVHy/oO4DW6EQfWPSn3BFP29PE01o+ix2ebG6hJF
9/D4I46ZdvJBgLNHfhoy0XMu6QjoKCi77+kmT8oMZgAkWudJewisF3ynQnUQ50M83mAZdVrQ1shy
6MmE3DqCFICO8f74+XmohJweIntnQRV1W5KXDmCXW9FfvlAMKo0591k2FLNJnK6VxjO2rMr6RUwW
oi7klpQnx6gUWqxp7K2q0snak8hukGjd15kZNYyWEYDABSbn/vs/KHIHe0jU6KkQoglT3Yy8Ty7n
b4dajTGjG16lakRT6YvKACPg7ox8m64+t6ZnemD3YYzg3oZO7brf2PPv0+pPrzIZriUANBM1LpdX
NdKfPB9P7hcJFPOouomYmxZCFDAArGpC9UTsrNufGFFMoXwteI4s/I6QJY8HJRSI1D2kCp+jPRQB
VkiehY55XT13XFZKYufCZUQBYOYV6mF92uWtVJpYrSQ8Mp80jpCH0IQuM5fR1RRnWOviBYD9y3SS
2NoJVCSjCB7JkUJp6oSuQhMDi5icsGUn3PeLwahkI6oJGx2dBpRg3w8IB7eCagEt9X7XspDoMo1F
KPPY1kiu/2+SYKZZTRgRqKFju7rBmq7xkv7LGV+4K0+fE+v+XksnhbKTqKcV/WjXAoxw4nywb/v5
7vvr82IvwazONdH1tRcnJnL3gAQRo47O3cWXw6fBDg79jMzAe47jLwbKoBL73auFdj56Zrf4sawR
R78iFxUHK5mst+td+ggm2XVs9RHrVyb4LTMHiC81XWOlEPMVpoI3uoTeGwjNqYsVUHVnaJxQa1Zr
2NVyrNhbByruiJcmwJcWo2JQVBwy1EGjfNr6QVjNPxKVpGmNbbipYfolBdIgVDreS/UT/7L3qJwy
p31OTiDeqN+C6xNXtCRWFsAdcRgHUhEX4FvY6++gmZ1ma6A8RCzqaLhzreGVwT89Wo27znseHJG0
OplBk0NWVVwjNF+k/RWIP+Qka8nrvbugxB0QUXoKGN1eqMLYfZ4D51LjOoFFo1KN5u95ZtrkuWIo
wbix6TtmzHRu+P+Fs0d3ybD6eWGlhR71kMPyfPm92cdScIyfKUuhzvWRCN+TFN+X82DTY2jebFJZ
qFEdcjknUz9Ic1ILWY8qQjm7awDKbz0h8JLul0ApcIHOeQZZf3K8Rl8wdTWCc8UsUiC0+OeN6gqy
99tG92Kw7dMNzZhd422W+KHigMLE452LSvE2J6IzIgBFNtkBnFFR6PBvAAdDyINMF2ouwWcN+Xyh
V6Osipc2Oyu3NYt+1iZ25nGYyBeM+pKHmCDPZRTou4K5rtAp7L98XiZNsPr2exGt1tfzuq2qzId2
QQemxijN45oShfWeqOxtPY8mMERTcfhGHlKUnn/C3c2Ishf1tm5Ay6X1Q0R8f9GpGxpPcD4AY5kb
gpa9b+RF33GToRpi+Wh8NmkJS6eO7F0i7OpEN9RaiLF5W1xt9EptQ2bTfdbe4oxVorOxxYJ4tFBX
5VIel8qxbqRkOxQlc3lhZgu6qprEtcBHmHj9lz56SiaFTtL/Mq5/rSF2ejKRRx1zgMVVueD0OY41
9AXzSnWRQtd8AJBKDO5zkink2z98pIz60yQcF/pB1YFVuoSJBR5oQi2VFbGng/siNO+kG3+6EpFF
uTBAR5b4alYtquOHgTLl1nhFbzqpkZDgahyV/e3+ycecsV4ATi+6FpMkc1hp001usx3cHRmZ9J3L
5Sy42ZSt97V8aBw6t6HZkP/xYxHsKgfmJ5jeTEiMHtLAE5F2LhWMVc140QqQWbsdwK+z7Q7xV7Jk
ekV9PmtFKIsTN6TR0NpnY/7keY/d2dWQHd3zoq7FZSBguvNzMzrucU2urdzJaTJzGD8PF3y2Q2Af
Fpm40jcX0EhpfYs1p8q/9SX3lNIxm0b7A5frUtXV+BcH0Nb6wsJc3uYnGMPHEwPpUhHYJfd3bc5h
+hDsdlwQZ9lnOl4p3YKN3ByF/1o2NOOAMQw7QMkV4Cr6mfWZe848x1gxOvSU8PV6dlIie8UDCzu1
Gf97BAhew3/RYox4FOGEOHq9bn5RfBc6Baqga4+Qeo/xFD6fwyPyv1mwFCdWbFVgCcKFTP9OfAwc
/Fm5pBLTDZynaCwzYL529os1TU5sXKPjxlDnDRYb2JguHnwGL+eAbKRCqFoa05GM1nMcbAD1S2Fd
H8YLs1OkbHiazOSGJJuXiUMvPCkOoKTob+i9GZ9LMVoeKvEwviQrTzUgSrJIyI13ndAJCEB5m37l
K1olJlOevXTldN47kn1EWMzlDXGTQLhvsXKTXcbWKZ3JdxuQefkSz3ZGGNSuO5TTKdiUuh8WhEr1
VCfeZTNNOXlY2SbuH6jPe3P6uD2HpFWBlCOymQWMhewuOrhfWVv5z1oIQ48PGMCIMF2qNycDgq+Z
D4kfW6Kp0gBclHznzqYbTQUii/XK/okB/tAlnZwQBxwssJshNzRTHNroBNmEkbMQtMG4mRgGiA6Q
MaNyFrywwKLI+mlAANiV6KoRz8r7xkgJgjayeTv1nneZzbUMfeS4oNOgtJFm/hknAM6yrQuETWSp
k4nfmcPMY6eilo5z6ihE1XFQYPF15nsxZVtzFm+fqBpoKw+TTig63mTHcXXs9hlSWG8aUEcQ8Tk0
9Gk7jNwXKR3GOYlPo+HD13qzDr72ee8tfwaG2SVtEcUZBa3q3NaBU57zOHaMufAoaP0o/VID4VK5
kJAVuEL6O9IZ5lGNQyWDHRxjwdG4CXL8F9N1COL0x5wrmQK5LX6QHkOwqMNzCjs3Xrh23qN0CgzU
V5aLqYJdrtVTwHsakkwk41t6qid6ELiSe0NKNkMiFRL6YcOxhdjP+6luwDkNWraDMpN28qW9Viwj
x1821G9Sr9SKudsPANXNEu9tmIf5pGpy20wSKxpOOfxqxXUkZ9Ri4sHBxE1fGU/ryvfMPkplZ3/m
B7wxphqpr6PaPCuujojarxcrxbmGDraJ1qFjw6LPGlRmsjxVW/+pftcgItWl7YJZP7XRysHM8Pjg
4Lv38Syr6rhiCLojCOboHuj690U3DBn/9eUy5fk4SCwNq8F6svpp537Qy9Iqv1wlH8ZfUr8pJtIf
aj2lH5xnP3H9D2C55KorE/qCIoCVdH4dEu+KJxELBVVX3x0GU4K/vTJdL1ngCqJIzxdTA+6AfHDq
9//HC/S4ERZCae3vivQtYlU1IGfEU282zueMnMpsgTy1zcftEJ/KmJlJJ2wdmOSC9q45xK0qJIRd
0Qj4suTrzcDAcsKQalh8vXbHwhKTPWUnk166Z9Jf3F8+bpfM7vMyTMwD6rOmmXbUDccDAyugvSA5
yS/kH94+H0WQ94/iQagjFrF6d/9minIBBiizkDSiCr4zLEsJe3fguspD/SfQGa+tS46dmXfdek0k
A9T+LqHqJPoEWZXRja/jpyW2orv1ufs7+6KH88cgn9xvct29iXRxjHKxmJQ7mYIS07P86o6F0NkE
nB2+Xia6JD5L2B31cHhjixE+Jkr+SQakehF1Yu4J5m1nvzSh2Zfe/gRg51cSHLns3Y22r9h8WK+x
OroYgs2AjLzTKBiRwh1wZIiRb84LwdnPdaZmCPqjI0pe4lKcAarM/nfk5uAEnq9NG6wz+uf0qe5z
XpmonDXZ8ypeuvXKA3bTDj5qFwwIxHlpqD8kOMAorgjiFs3SvUO32zUdLbs2O/AKOOnwD0mJuz1y
txWJI734jDDFFwY0NSDpboPasVt0zyBzt+CLk6Fw54xIgOYEu39y4MYBWD+u+pRMsKEJILRf4pso
5ha9X/pQ/zD2UJUPJE02IATTEUM978n29Ls+sFYSD7oNW0HercvYPbWkAKexBUO6W8++uF+mN0Tf
S4YXNNj9x62/2+dEiH2NkEQvLeaiFmmbEXPUBRM3+k/SzV5MC17BRBpJPAv/4jpJxqwbbJAJY8EL
HM78ckkD6vD76ldG6z1aXrd1drw9mCtwoHG7obDI9fvBAxJyjU6rp80HF+3k2ObYHcfgRrcgFZkX
KWmKOWLioK+Q6GADs+7S5jP7BMpthFphV/Ejr8H1I7FkM+4zn4UYGZ6DS+J6Xs7/eDxw5EMyHI/o
qT9Xu2fq/YxTUCx6908oRuYmR/lpbK0/0ZU4hr9orUnxon2MNsupfUJwLrM+6gGIPuyeoO9YHsdW
xJbdT4EIQ70fj/yQXfdqb0/FDrNVDBgRvDKps3ov8TGpw4Dw0zOwXGVOYZB2m8I9nWii1iP+z/2U
mTCjPhzmsV88dtyozNg5rfeKVngF2lWHVPAFeclH1JahqQI6NMbBz7/2SSdJhBSS9/Xey2BhzHSE
6BDTnyVPzviNmprY/6Q7xK9PQMPKGvu38Is1VKmI3gSTWJx9KiUhxhbDlhZnNm05zISXs46ywM1/
KKAZenzdqe/mKm6GYRf5w56IhwnUYYEQxq8E83slZ4WyLaP/HoK/SUJvvWeUilqwMvXXQr7gBB9s
QwlRBUHZhhmuuWVH2DEAyf+11YWoTTUef5kh80dwuXvL5IN5TYw/qO8kHj3Rb3sXQaeqynVaWwcr
nOIQWq9lyX2NPOg/moOJ02iNqAnLEzQm/5V/H9XKr6BN3DMHR2EhmMHW9W3cIdIIz6DahZgqKAZM
I9PSNWVWu7eReSabeEQewolRc/dp6qpUOqPCsZ7GA+ME3Wyga7zUN08M0coFexliNP+0UuNE5HwN
cMXa8Dwc5BpCmIyT2mRtFBIpr9DuybOTRGGL429CSc6hep6DHJ4F2qLzAVgUsyrjjALvrpriTY7Q
+mcWx9+CaVaQa8U6fuLK0J46eQrk2i9DgJ/yAlCeNh67Iv2BK5aL1Oy69FAFUYDHnMc34Kji4suW
Swf3kbZ+Xl7/4ogVOL14R78BYgMNH7vc57frTNSLTkU4R3hVzM7B+n/kclU9G6YAA+NEygPfHGbD
rLwZMRs81ccc2Pvdrpit52U27p2AuUjmxaqJuwjmnMVcD22JrjLJdxtm8lcqNlSiRRMiQou915et
prZNn4aubLq7V8LT21eTFbU5fz73xt/0CtJUfrDO8k6TCV6v9OGk1R/wwXHf7lrtN6mXL2ULmgMu
2MfaAf6O0Jt9QtO3/ECcnhSzF/dSCiScZrLRA49NuYRp8KWFl2725uIPykQrGAlAnQWd5eLDYn0F
oySiBlCr0C9xwMB32rKlepPE/1j7JIQeLu4Zs0vVpbUSCoxlMnyxB6zUAY1N5WXImj5q8n4Y2Cet
QpA5Nbpki5qcVRVy5v24Vy7+KvXeSrsII3x+Bo9uUjRqlH87Y/5+h4j1Z2ZxS71im4NY6t6lbN2L
xRt60sk+CF6sf9hgiHVDISxURwkdQTzz8p/jnHHcfu6nAUCUjJDTcBQM+MNSBFmhQmGE1DAIFVPc
tJ+yOV1oJY+nD5mJCuJP3oynXOjcu6VM6hpWh/fNaEOMBlqpOzgrtabQJJacYcrJ5jZq0AphmGXK
+bcx692NRUOGGP0c/Sgzb86y8i5AC56F9fEUVM5wrJW+5X9ZL8CrUmbGH7XSAu67s5zZpFXd9nrZ
m3JyGsFlav7tNwj9JU5RTaeG3HXEC6ZZQHeSXb8VXajy30Ba1WIChraAPHtMRZV/G+ALiPGMMMz7
7AVfYEOc8yWHilIsoAi15P7eLQmMa3AHW9RJIsWijzhJODQUDceindelN2zps4N7z0MT+/VS8ZsR
arK9vU8i2GX1Nbyi+HTqnhPdHBRp4UyLw1ww4W/vaAXwWk8SUsvQbbsuPy/KaOW6O0l0VlfeP4YX
UTnD1d19Pr45IcgbWVHq8Q4xEwbTxcwid7t5mhIIiwVgx9PcVl5Q2+xxJhzgqC2OVGhevVR7TIEW
9WJrPr5K9yPEFcpBnmWzvVGo8vYXm/ZKdPtLlEB6EBLcfAAL3AEFz8OKTGL0VHFQtg0ZCwEBr8Lg
MgBE7u6iOPHJNKIFoi2dHd59EPZVxhcdYRwqcy9cLFrVTFyZ0PpcItEbQqplLxinCJkxkhjYOrIe
tO0z+EBUbTE5UjBA0RVC+Y2AhAQRpEeZAQf9FQb6+LcnmhqJP8E2UmhFxmKGkV7FjCZDjtB6F2Q0
X1YyXP4ZsqgMjz63R+2a7uwu02gvYzYzx7kD4fazivduHZcuvVxpM6gjOwD/vXFkhydvq1zqXmt9
F9MALFBaqAb/i1Z/hf0kaW7P87bTXQl6BxKA+VvpGiITQdekfl2+5PLm6dGcjpGK5CZsFmNFGtAc
dv4pUcxM+TIWX0oHwnWQvpF+HD0k+4slOFO/j0LY9sZC3ezdmx+KuLkbPDfjKAvRIKdmnZ/9raEY
XysULiCqghKlxEl8dIs9jNvCQ2aM18iktxMGQM8vENJ+OzdLA2Q+hes6jz52iVh/UCMBZXlv9Nqr
HJcQzEhdl84XjI1QDPwNvBp2/4641XTTFw++6vhG5GEKfP9u6dRJDfJWImxYVGvKJZoc48yfDJgS
qF/RLEpMWjl4yTdS/kOSnVv3kfkyKUTF4qHyxm82YIVHUf/Gwm3nXqUjEykf69McUuFWC/Ae0gFd
/OZCSx12KutIIbosUPpT9HIRO8w3t0fDrhMPMHZyYtEOMBFx+vJpxEtyJ6o+2XXHBgnFilowCKMW
Y3cow7DsckrulMdTcqM2edNx1FYPuJK4NPDd4MTyhaX+xAXHJ90DgJPa4N94tbmj/L7e7/pVHBNE
YeLSWacKdF8wrkKvMXWWOfirvrFCChyuDnJtVCQg82jCHEb8s1Dd7lo/6yoxxQT2sPaRl2DyGaXr
s8UOA6+sKPHZC7qa5iB6tUhPwvHvkwDDnfj8SC1F37QvJWIg7vsZt4Ls/rmCo3+PgFtzd54h6NdP
iM8ln/ZHy1yJKhywTWJ+r3vXO1jKlbGqiUB83oe7lOPzU2iixQIF91fWGqNQPr5dUsKcpZAXag+E
PlCvZEriQGtiALuas/U+h1JEJzGIbtHICkcZh+TcGljvtf1+69jOj2ZWpTIfWecn2dyZC+7zn9w8
D6cGidmuHPjGS6DDee0bPNDxS92PgFK/x5L6Q0fnR4RfmR/NC0Upl6VeYQ1H6naHLDdF2UDiyEGJ
j7UKLYkvMttU82qtBQhMRCyelpUR4qVhMakdV4q9CzbC7SunVMIi5Bwcc9wS5gznLeH4AZB37ga9
nC0ycUKWPxp4k60yR0Qf2c1w4fu0U/wz6q/PO0N9TUW3xfqe053pkeqfghhHRd81l7xz9YmLKy/M
Ow1sEyzwmi6TsK3rqwbw7XUYONNHM3XVrPPuZeS5ECoH1FAXVA75fYwalTsC2TyPoiZXE+HZWHfB
B3Wq2aPM7AQbogD+12Q/kikw3SUHH9zD3dS+yD7Y7p9KzHlh44P0vqr/+ri0t2fA8R/bfYkxQ7+r
JNhHzr0AujSM4/wXno0IoIPRtgKHgyv9tCT538asLKr57zOkd6ObiRQ178frsmfNOse5mGeH2TXX
y1xtury8wOSs9NvpjHcxU3UCL62DUc+CNp+PCmadHdMfPc8s7n3A/Te3gzYDlhdELQaGJQvT3U7V
aqKUa/3lXdLzuEy8KD9w4+19e5cxou6P7C2oOjB2iOCc5LGaKOsJPgwbpyuBqctM2v10F/U6pogR
QpAQs9VS+yLFCxGAwKvGWo3kRtlfZDyn4nn6k0W6qQfTBreVjPNZ8Fl/m+9lT/ApLoZFbgjaLz6K
zndKNvUuB4RxIY9Hf9QFnykKsbFLF4B6nqVlZer7h15+3pc4CSfKBWcRCwhXKjXottUB9Wh6aGer
bs6rFwKlHGNajkWqoM3T4la4CCr/mTL5ewk2uNNLeTm3h05GDP5u8BZxQJKnfTFN30fSzWVH1uXQ
HjecrPI3cUOU1A5q5/p0QVHdrdKbfMbtaIzNa7/7TgtynIl2OmYIHvGTGRLmHmqxS/Ydq/egV7vR
JFtJk38L9flwxAvjiF4yB5HSgTV9cthDOdy2ADXcfiFLkNJHIEnvwhgkTnKGD30V0HnNroSmWsHj
YulvUYChlWXBJN7I506ehtBb5xUbUyQIAQyKoGP1lC6UIowqd6jH1RiPW6Le6vtkhqDr+pqQG9VP
yFs7d+cpYwrbC0rh/WJFhssDEyZ3B/qeznbReLImcJzZS+Y5akWEgkD7wU1L4uHGp2oLWFu5giu3
9dbH2bymS05/NwVryuKp4AJLRc9YB689X+pnX3TxKL+1SM0xLKXFxhARyBmvtmQuANV1CgeSG8rG
QI5xtmewHxi4Cs8Inw3DmMiovVht4LmoH5EZXuUP1E5yvMe8Xc91j8o85vjCUJvYYFl6G3TUOuWd
6BuWkniadGppYmbHXxwNXSr40da1vdOOERAeM2MHB6+TfaVcXuTEIEOe3t2XKDprEfrCyYPBosWZ
j0P7zEym3MuJhPCZ6SCljqBf5+H+WR7DxGTXHS+KOjBgmOX9TIwJ7B9kdCJPO0HLf7O60/n3Dwnf
RV/6L/jMqfIx4XXrGQnyOLazyl9KxkbHIZnGt881xd1SdRJVBy6JBkz0oRMZx75fxBdvSZctoH69
0U0QbWj6mCQdUH9q2yoG5SRxieI9aDX0m8pHeV0yWoD9LNn2TWyO8CGf97o498ebktObp3zD567n
OiRNdHkOQZqlUur19qKXOLLFdBDjnhaG62fZ/dvEO2Ico9uBdIGMKvjpbB6rdo4Wxgn8t2DZYXm+
KpciRVNxaRYvLClTsWggDSw4OgIxafHaqtX9JC4/UbtquMpRqtk12Sr7SNK3FepyWf9gbmwdRLFi
Pp5z0p6kH/LxlEaQc1RlKMKISnIvfJ60t5lrWT6XTKQHgjxznSvej/Rpka3+rTwKP8VMHxbAaNBu
ZSLwg/YGa70VoZFcNq4NuobpuV6fw6ieXMqi9Xh7eKXEZU3jL/lMCX1bn7JxrEsQc28vOoGjTc+B
WBL7/+S5fVG1icNtgqV8wQpl1szeQOBWKtLOXvbztgTAqaQgpa2RIim5pZqYhy9YPOWPHMPNTmK4
mWqiHVCcvi8d3FRspADAHpdWTC87qPiRESmYU89Mb7qucOPRFnihPhyALsjhTI+l1tOWvpripJYt
9rQhz7eMlfncF0iaLwuuysQy8OhunNh8aY5GOyFBe7cRW+TCd75rGrQCiKi93ZOY1+oeDq8SloPB
53ELC1gimg5DNM6qdFiX/x6Haov7ouNWt0MmvWl7D43VL0qjZZ1fLP08UxZ0vTDjUhwSPPPX5Y70
c+5SjsxUT4dh92YwsuB/RTZTlBecyVkMwyK4wJmgNxeSEDCcmOhQDH4Z+6OisFKZuf083ZENsDAi
6sG1Wi763uswDoawcMjJkmKjJJx2djsiNyVnLDfZwp7r2y1vxNQzSWOsRm8sLU7cKPx7exqmxXPu
Q0Y5fs6cOPnElcqLzJWfAbFtszkLPgkcQq0H0WGshHO4Wn04wFbmUz9py46inZTmg+F4S0ui+RpA
w4SmPsr77U5KxZONAS7Zppu3/G/8r8Cz8kt3dM++fK2dse3CJg6wbxYREKXMngNRYSvypmkK+6qX
wRaZTm+EZqbzlmNK0oqvBFiQgZ/nqK7H/+vKN11dSLCNHl62ehKWDulVkACmtYkpkR9pgentIahU
P+3d+++SCIB7lmDV3Yqe/zGBpEm+ZtXQ5bUDKfdMYwrQwZWBMuxAqoT4rIUV+/7UXGYUz4l2ESwF
W41H41b+O8/mC99CUUz/t0tw81hpfP7NE/78lWZVkuam9yNkt9q0Y7gSlkMbMABBs7vvwUcNQKHX
uIKsRekQ1Q0+fOTik9T678/cLBdXD0l8LW+qNGkEj3HlibKJrC1nLo/NoMvDvt5uepAYdb1Ds7YN
4N3imPUo1ku69FlNqY4XDpldWz4P5mKOorKA8p9hM2ZnwbH9cVVwHCVrckWZz5bZxEl/mCSyypJr
eYW80BQj2ZW/WVpuElYV1orOT/UbN4F37iN4RTolNa7Cnb7Eig7uD3cXeSOqWIXrnehT4SYG+SLg
qm53lvqu9WGOF+UFBX+gbJpq9y+on7Cxfk0RMLFgiJK4IS1e8OKMxo2xR/k08v+V1sw4VOv9J2nB
+hNMlv+/HwFG+CLzzbYCx0VP8A8imRxMdXsJyabw4csPRALZxtXbuwFnZd0ERB7uG7MYj4cfSPAM
8xyEZSUy9DIfEXfKxIor3OnxQfZXrOnw3DCbt//ZdHeaHDBHlOFjQp2q80UPSrFucXNHDR/pgVY+
SpS9oG2mL6j+wJWPuFx4vST2JCEMrVBByJedxlpiRkd2sUtef2LrnlTMY+W4OY/LtByjJuS8SfB2
q9daoaQ5fwk8Irq0btNds0obllGm5KaIAxo8c48hrRS6gv4LoOET6liGlSwPX6WoStvlM3hJ9qkm
oE2dGSMkskb0ZI7iWCvmFlAAWKURXCgiDAsFjeHAdbkJwGFbe261+ljtzpPCw/IOQFeJszMxHAkm
N9oC0CxWQgf1rj52aG+Dcah3LXr1KUbW7qm/KZx1VTDlPOmrAQwoURvjs1RHO1J4m6ILezPGO6Yy
bI+1VK3p2YfJRZGmt/opfqkskX6pKljs45HCWucZSCyXPK1IJ+ZduLUrKJJrkvLBEIqOp/B1p9dG
/3M2SOvl/1pc4gotpyE9HZVEbbjgkCaUhRf+Gh7ZwdbbesX6lADRPO1mpECUr9Lv3QZ2cguMvgvf
zaAe8Dq96I79Gfk04AqvvumBMqdrz4IhuOhnHr0zANqAz38dPx1+Z+Jl07nk0EsUba+Fv/+Lb5OV
IYCGpfmrT7oXLCQDNxfqoKzQBIzwrCIfNlAIHlbhMzG2DMkE0gbJQ1FYskZPcnCqW0rDbtjQQyN8
D82UzC60FWmhLOSYsE4HpDBaj4jMELem5uY/pDHDpFQzyEVg4cpZJG7FfUcPHntbP17J0ibP1Gsc
46kgWPskWTD98/pZKTmBFevuxJ9I8kPdruG07SMtl3GC82/s2m+cTIt6ZzM/CCPSz7bz0K4BV5u6
9kRCaSenjSeYfz19PGv9HWhqTRM2ffOiwiA8tPcyjFp9I7kYL77MGjijQ5Exa13BcNrC2lt6cB1j
VQrqfQxRoE7+2r9qyU7v8AUvToBs6u+fYhUe4Sk4pcwv+Let2HcXIFPAua0t1tTN03eK6tBbGmS5
sHhVbTWgZeU5gTZ2QhIF8349ZHhaK7u0nheUxzQoS/WrpTXgROcuB3MB0uGMXAAmCmOxIAGSGQjM
GF9xAq5UH2WvG5nBfKFq0h/oI4Jht6KXxz4ySB8y8KleG8fqet/2Ouui8czfqIT6ekYV32eFW8RV
MQnTvzu+RVI1MQv7JWi4iZV51KyqN9EX7tff3ANNXpOAjHbdzs6DorlLb6pQFeiI8tFtm08dXJ5X
9zq4oCDzEyOcObRo37kSvCKqHA9Ml4hDLzBZ7YlgeP/ysKGdxw0jOHQCG83wwcQm5eI3XP/OWhOO
jJwMwzk8X0C+z1lG/m5RIJQpIhEJRCSv72w24PoJVN0m7M12uthytqv0uIvDu704mmPiZ3a79Hvk
1VmmPOGCSZnpArI7LweL/5Rlw1FQ8OzYGEiS1vktfsEHkppENakhNoUMsLC1C8SLR63UI0jO1KcR
aLTGaxN/8WptrMfw/miAtQsTMYh5RS/RPMqrKV1K6BIHloBebGUTsjasN3mmha/Bj7U29XBOjlsF
mvL/XzkkuOTnoRznmSpfZTGmWFbk0NHo/m17fDL90iSMZPJH+mAd0vxzRyRMAKFS8NmGdpZ3oMmA
AbnP+c5xuu2E2KgAPJSWyiXV8WNMzJC+/TM7v+0DGBEgr0S0lQxzVmk7dZJcTtOf4JIHc5bSTiHJ
NYmSNnGmVAcrBycG4Y2YCioMegvXH4mZDURn4w+c40JHxQdnwRtBexAEWuSxs8CQM6vUAtArehVx
RfJWEw6dj+hKYdNQaFlZmS0h6dCRCGIa0obT+62YA8eLjgkt6hMsJXrKzUe87ZTUrFYdqWcUCFFc
fvS/5QWW6I6XhJS63c6J+J2WmG042ja2U3ckBExNX3tT98aK86OfooAs0vrE09O7hwr+0aWDbw2g
f3oIA/dLeC9ONEQTM0sa3oFlpmP1kuAXVu/G2EBuJlgHCQsAn8rqspSyl9l7iUlU3COSZaNyNn/0
ruoCtMiGyrLRghmrfloMiiwuFk+eqW1lDHUuVB7vf18JCYbmScY2QpXW+MLYxw9ekt+bImWW8Ru2
5xOLhrFxYFFOOSQdLrXhLh3NdHtiop9ywpVR1FyDEEoY1brNBlPQIRBSau3fwAvyRAxAW265fexP
HKrjiU5uc3yzrXFhOm1PdtbBXanPWk8OcSqCPyGcqxrbX8q0KOHUSmFCLp8Nc0uuhZ0HQ9m8EKOz
S+gFUy/VuOTX83vY0VIP/RLfs3V1frGtvO1+XJcEdOjUcdlpiqvS0CLIResywDMEYgx+RO3rSYdq
XG95sLXwlP8WzulJSofxsSm5FXx8MBEjebN4JvrNnvk7zooS5Elxv99bxtcXOZjszwSpanDV/kZo
xFCK/zdb8Zh+L4YpXXRKt++AxDKO3JVEnhkQJevQnFFXrwtS9WWHpgJOKW4+b7+yAudUprAQeWe5
ulIa2T1doOS3HAX7/MtmPMDNxMEaklR1gDKcvC1mwDwu7O4rPbn4ss65brc/8GpvMY0d4Y/VPz2g
KhVbioDMEooo5katnT+jJ40Ot3iRusLPS0OL0OIVFn4HmtgeJ70VBzzbeeri473RYaiNiEQpDFbV
4o2bBxCv2MOwI4onTBfCcJbYT6o2tV0e9JxoA8i8GiRO69LaoJyJM8Z97GWXzqDEMoi8fotJEwMc
sn6CHLkL/yJmZPa8c9P9JI5ibtJ2dzr32Jy7rqrURer53Fe5bddKwdDZFTADOzaBsHGJX0cJPmXE
UyFuxW7F1TgPo1r+2FdpxvlKKjnn4f7k6ulV5RMyBo3jXOMauZ8hpkBi+XlJ0ommdBcdDScIhfxl
nbvODFDJJ2DaXn2b2tj53FxDvlmzUFSOR3OLRDdVVTFWStsyOhX4RMhdg820f30izc2/ZmNH8g5N
yjPUWk+uZT5bXxA7AmTk4Sizo67qxAVkjw3t1EGnH/GGKDplf4Sbk91LhSuaVhQYRHqNy6Zdg33v
RxQBRKroWBA5MifqCKMxIl6xg5ExCnJMi7CmFfjYT4tbXcVYrlMh7TluPM73hHexxh6Or0ruWtAK
+QFf7tvxwNYghX8KWUpsYJYEXqFtGsL9auPqwPD1hMXEzzKOpUtwVDhtfhhfhxbD4qkC7Uvtk++q
3fV4anlutG28TfBXMNAydjIyL2g84v2twKZkztuRRBC34qVRgXN06jHEM7pwRr40iAKy0tb9Nwle
Me1D+uLpPiQCREIWHA59NFyIE/Q2uoYxwzNmBlhhwRwmnlyPk7DU1V4bfPZqn3ZbrAuYIjhbYgI3
x4ZqGLMRNJWXP9kts/Mq2r9Hq1zuwqW9fxalXVuWzXKSdyRtcCfdWMbJUb48EzTbwICReCi2JW3/
u9IrFpfixk3jT439xa2CmiwX6p/MZCjMBB7LXaTN1p9RK97zKkyZXgU4zb90npipOohzbEaSTHL1
69z1oNA7lsYSBLLFH6LXW6sU7vVQaJeGlLlBPhrIMfyuyggRi3YDeM6J/vyLX6MOD1OR45cBmls9
u/d5gRVpWWaCiDQCz2ZgqfXdEj/iL7OzPqMhi675fDgguvVGKaHB2hr08HPCe41bBWmReOWtdULd
IS/kFNGGeGHVMKK93zxEI8yq9kBdb74n979MEdLVrc8bztSVX/gVOP0oX9bnrrhkLkBx3ezp08oj
0Y3JIcwRox62o6QUQyOKnsGbfxAHxPbBFW6EfiXw7FJO2oZmeShm1r8Svo9fgFJ3EqRiNJDrBEFd
nSCN0Ivdma+gtrcGNYp+G0jRRJIfBerRo5ufD6IcCirqH0zfPjRQL7UdCGueHjJS3zp3m8hmtvd0
fD5E5gPaw4nxlhDyhl9BcEDbAWzSgVU7T+zt29B7vwbyxu7v/EyiG4i7hMh/LoA9lPoMUDKmJTok
w4xWMnEJgLbevBZu9PEuG6KaQt4FyvI4Hlw5yalVM8d7TpNdV8opCc0/6LEfnwu19WyIMS7Z7iuS
FWAj2XHtXCazsIROPTZHFJbXKg3IZd86hNu7rhMuyZqVrHUzxMvTw4PDKNVMO/BrF5LoyQ19glwc
guoQYhK0+mkRZsddsNPk4G+u/LGD0ilRG+4SNWdrRFmrhqeAjlPN9PTCObagFWUP6iCpO17GmuJI
9bZO30VQvi8Z3qYfz1PlPvdpqrA0Ght2NTGv7fi88/CiQFkPN7js6TYHHt/Mv1Iwur+mgbGAvWz8
YJ5t+c63ceN/muV9MUW+cxN3Hq9Aze+X1zuxlQlCjnx4cy4Nz1wilzUoF4+WtliMEvY4Y2FIVwbF
RKQ3FK4Y7sb8hzkdpQvoTrbmGXjqp9bGvKs4UN4vHKuG6hvDO3dvYBgu89Z+ldc9ZJYAAju7kHYs
K4/kDjEY2L7gCo9gBKSyptp2EqCkeP9ML5RvC2AfHT5cIwxkG68R7ZD8g+U3VS6Nu6cKQE4d4bnR
mHnfFMe+B8D4MQd4OTKIantAiy5iXQJ335D6+9Ck+K4dOa3Jowy6QtCnZK88ikZIVduXXKJzQ1Ts
6x+oqeqc9Kb//y3aTBAYnmWz81sQQr/HCVEy4NGi1vDNugewTu18bhothfyEhbau9OnQOhUrGkCU
k9UqJeuZWU7vdLPwbz6NRcoormt8q4+hZ5p3xN+mJD6tDFDdVPWnf+mbF5cFFDVILEh7fhck0yJO
tgI8TrnAW2z9HiTiZa/XZp+gjZtTTortM1QwddEnFd5oTnHbnY8PxJ2yMITmekeLSOOZI5IStz7m
6oIjPUCmGxW/Ju6W5+sGnUDOUZC0nqLLVO0rTJgI2IYJwrMy6g0V4tmVc1bjxsjn3W2I5A27e48D
NTiLowKuOor5BIx3Qkr5yHRl/WZ0rzKP4TeGD9pKDpxiJvh16HaRQ4UARM+de/e8im7dmeJr2WGN
4zzFN/y3H+8zL/u/oem7VgZtTofOvHQ3XZGPnB+lMBFiCrbbKPQse73biFjKo+qD615nBzBYn0Qs
EzojKa+dh2qB4r5rlwtlgqsg1HbDwvn7cLWRSlnV/jppT9o+O5Rv5BBl3X9FD82I92oAsKhhNxyC
7NeWSPae6eV096w4GeQyTUrE9q6id4Oeheqrz5Kmi+8WzOq7cV3BqMs9Z7UPBG+I8TC7nbDe54Ax
zSw+GxPDQbfbycWgYx+ITsSlF7mmZ9FN93B1exur1zmdRsiTpjJirof7tbSGAVS00F7Wl+FFKXgi
BMDZfRiJf0SuOqkDUuvDxmFyoCD++CULXXTSPKhJs+mnsIKqitY461FSA4z1JJfc262r8VNQPZI3
OH1AX2K/7m1xE5uZ8ebdJ4p1c4J5wrg1if64VGZxmiJ2bTL1kzw3NXG5ML96L9KPnlA6jcftHaEG
L7A43DzCReB7of8/oxbaRhNMThuA5Ywg2LXXUkw06CYewH34lsb3htyPuejDwVy5XXo77wRWSgck
etY4i6t13hR7fBloC6NnMGWPrEjK+rEDWdd0/PlYMwpiOicJKXCLkjtu57x9ZLAti2CVeVAmno6N
3IzioFAlj8SQSxNI6a2B+hThIkUNak1sID7Xpu+yJ8Fui1etdOk1RxBufot0uynQAQ57QCvSe/9b
e4ffO7V3JcPTdQ9Ofme816GzN+a/VA2DkQ5MuWv9pLP3WNpyTG1Zqr+xxPdLFs2c0ks1XveMDYmP
4JCXsXh1WIGK/8STSWoySIc9o+OgklN7rmvl2qDc/jpk2KpLz04YPEx3VQ2s57cXNkgUnP9bLdxy
M7nH2bf8tA8Rv0T8kHlNUQFlKKc8ocfMMi0ew5tBfBC24tmBb+S5qYzFjWnlv/RbKAAskF9BsQx3
947m+68Igo9mISrTI62TivigtxyVwJiOh432RfPcZB9Mt50u4FViXZl31YgpboGUF0zNR4uDQIw8
YhPhtAqcEJYR4IhLWH6b9bxbaAPFfl940cx/wZx7Mulw0mR69C6FZEGod8GI4pns6NRjeuzhyv4X
iDTPZDM2GU/2Lr3I6tTlAVgjtED3sFJkN2zoydDAr57RJM6LTn2ws2KH2/JOa6xlq90pQBepoU3Q
cBrsilC8GB4AGiHDf6XMcyH/1zhkLbCelXr2obwe+PnusNDRKuoaBck4QC0qh9CU0VXc7Zn+CBdK
gkdh5A1k8xQVgwPMlmUnfSiLEXnT3Mvr3385aB03239o9JFlz3JyeaSOA4PljlenMwYC15hPCgkP
h8IsLmaoKknfLe4YFEIhZAfe2vHwRklzsif+3k4IYi1M5pRkq+/UZhabvLkDHQbhZuPjeedNYqZ6
7HNZZsWv1kA+hMEy0NBJ1qqWr9NvpQNjxbxaZ8oUXRzFfaGc5+KweXJlPxg+jXHxLwimiQcX+ZuO
o8QPs04xxeIA4VBNYayqXivmCI62Mqk2FPCC/8RsN/5JX6P2/QACjaU69NxsZzMr2NEwZV6+Iiws
WaqLl6naAnLq+kjJV3i25SkzRQyJh1gg6m30rfHHdiWfVvRsymvyUSrpCfzglw01dV1Uai1UNYba
IxkJNfoMhMdKE7MBBmEj6Wz+9QN0uOxTisSqJRCzTXbDVm5tSFtkq4XWLqq2e85r8yNYaOYzO/5Q
YeQMMapfz6oJeEK+BLAmG2lRzDFCZRVdXVSGkv96glFN2BFV+eM7CovIg9rvOe3Py4qAU7AcUoDy
2aRzw+ENOtDwmGKiRL5fTtSy9qm2WCZ1d+UAzqdffQjueYx9Z6zBIMfIYk3HF/fxXRc3QIrc3igJ
WbH0TgwFY93/+jg0nupB9AyhqmNNQEem2K2lwbFyjZWdfkBB3z54guboW0mtFc8ZdpKKfUhJ13tG
s0YXmVHjr5S/j3Y40fVcJTNKzs4ZKFENTj5PwTw16v6Q+Kl/DCOpNwI+bKljDJef/W7+Dp3sWdQ7
WCLrltem6N4EPVOaNb87d2Xc35nYBwJRY4YnyofSrmLny4DPdHTtKbXKC1DJQmK8W6V/8zfUioMi
Akyi9UStAILWIFDeKzc76Hi9uZuJBmT7EAMXgeQDRy1eNQKR7ZpQaz691d94IfTOsd6KnmAUR+NV
Yy5ztg5vzJZeTNsxo0677VVoVQFTmOpqjmKD2e2g30RnXzOb5aExXBb1bPRRoqzaFhjkonGf+zOh
QZsEbNGTjEwaF7n6r1dOc/8WkiDxiNkKe+eINAiJ+aNNtd4adoF8UPqMm+FJbXeiiii0KNF7AYd6
yVtO/rhsCyCb6mn0eNiKbCt7/p6pSIBE1mc0ErXL7e9XDnCecxxN/5TQ1WnPDFja5uHP+HFVy0QS
gYbhbJumAhrFjD+93fjTVmUkR12jiQJXC05/6sqSSv7Ii8AjR4K57wIlE8ddOclsUCf2MQFhyyTX
b6xsDi5JGMkeLx/UNLJ26xcrxk9ltjbgNVeXEd7i6ryU0qyjceW0oKoLRjUoJEGMEJIKhnIItj8b
wtRgNhfGpdq3MVqdEO8Fzpd4wTw4htAv34XZxqkNhAiRLnLJ0QDQPgnUuw4lza34G6GFyepiX87N
Eph5BKThu1jUReWRVU0dRSBDIvX16Xp4oqi0+AaDGnGGVFiUkHnj/W1lPMC0i7+90FzTgY8dKnSh
xiyw8INrTDGrPtSL4i6yra+GZuJfdWrTcJFSkBit6hSC8JpeURNmlE0YQKU904nAyH6hwybUDYOP
zxreJuVeWteDDGSHMml8rY6kLNZaVrxOB48VJAgRpfFqAoPURmpstpEYtLhiE0xKJT3ihw6HY0Ck
td0ZyFZjyE6vg7kfiZJGtzyrDAlq2L/2FGKJ9Sp5iT5TPldxAqFAEqEUlk28JwKLobzFJWG2xt2X
el2Mc1/l6dFAG4dpKhAfyxvGSoxJm3NpWJUaxCbYYMDVphiOVfpsfgYeYzJpvlGuz1pO3H3uCLFA
tLX6e+cVCDOGmgFYj8hwlRTDP2Rdf0UQvU/GyJvZGEh01SHCO5rWBhDtQZPJbKzMLNfc6ajTAAO9
1gYwoJp1EbXQPpmfHqx8NSaqlPbUDQWPf/cE44TGLBwAxc7Trbzw1HFcBIBZZGQdgZrQjPydIu2b
imVfR4oZV7HDtTQj4kGDeVyO/SH/HZVHxlxSo+p1plUu5LBOfHK/4NnkMHoV7+tzUYBU9Bbl2qmv
OdaXwSk1U2kocRsVrA9Akidz6dD3M8o84i4EMYlchNZA2nqIxDL0N9bgOvi+H5XBh27wwg+CeYvL
p1NnN8np107Ko1N07Uo0aQNgM+2fMQG8TPM5iRFa5njwR2ZWXBcTety/vmkDczTQpNy953VoA9uv
gaQsOtNxK+lBn2/+ig+yb8U5e3qzZ27bUyQXp2R8s2Sy4u7uh8DKGL/xKr359m8LRBSxmSdnVd34
3PFYBIeNGrTissRHV8+5jvK4nufBnlSqth5kji1yjmB8Sm26QthhbL/LUYvQ6cCMvNnza+eeSClt
lmGwXZKDHWQpvsFqq7C4vSoo+dNhH/rG63lR/8rPAU43VpCx2/qB5rtrNgBD9DuhLQgdyyiN8t+d
rWknRs8UOo6LDVuNthQKNOQQDf+GKbWart7UFd0b1+7UP4PPDPGsjoBuUj7QCUmZ3sesJs+Ka6xC
l0NkhuYZBhCeDC2Mzb21U1C18sUoTHEayIh18iDUM+gFa8wCiSXAUyBm8l5js4cmRcZVoF/T9fpZ
d0z9eZFeo4F6SpyhEAu3CAfcp9tj2tOWCUdt7BrytN5fCZbxMJ9+GaehCHzZyYeoZy4AI2ytY0BJ
3twcFEK7VO08V8LKMlFSkcxwgg6HwOrmJI3Tu799J2d24AuyBJqd/lY5y3hl9OtC3ezM2aqGfvBo
FfxXBS9eKYz1dZLjxhJ9lO8QRUXFYSoRvtZb2OObqIAkalep72t/vmH++9ht5f+vSNZHp6AGYf+y
EUVfncNVOKYjvnszZywKn84aaTGvuGc+XD58e4JoopC77O3KznTBr3mQ51VL1QpoE+xL31sjgGth
qj2U7n7OkebobjbdqWdnJ311Cq66mHP5S7NBBMGEW3rF46d0/bmaBe5v9B6PYzT26RacXydtQoY7
x3aCwZphNpltW8Riuox6H2cFjNDMKVU2orw8KqQmrULtxu26bQVyHSs04mxN24uS4j8qJwnaCoY1
wSVc6GbufpZbylzBE5WZ4vKMkAZwQEQoBr0BKCUlkYybEWPWqctmL8AI3M3qIf82pfgkGbigHp+d
VWPkX8j55wZeIp5LDHagDIjmmaFqRohYsDmsZ3yslk4+Nd/lGgwXgwxr+taVN9qQbddP3DIbl+E8
d+k4YjfMqDS9fJPF2e+/JMfigsbNb1B0jkdePX/3LzPC0SwfGzduIEK9otN0OXXDptldyOMv1vyt
YR/TcdMIpjNIqKIP2FIerBbpvykU84MZnT0yeS8GztAutHuujp5nSH3oNALVh0d/JjkHKc/L0ADB
GZe4O5AyfM08pvNhQ3eyIGdrr4808M0j3cAoC5jqdAH6cD1h3W1lhyriG/TlxMCXU8Z8c0mhX8Fj
7t59CC7Q6bT50WiEwJeDab6aeUuByfCmVK19Yzp4I7mW7ApQOwXiE9yRRwz4B4NFFEh2CV6IIhwd
kGnhc5IZb8EkOhcmePvy4IYBP6rh1zN/rwGOFhU1zNQ1f+ef/CB/MoyRFHOvfWvEiSQj8Cxs2k0x
eegnXx8e+FZ0U5EYLS3uy9kUdmGSKXitn518//VLNBja8Yeyt9rgpwbHRA0LU1ZqhRG/ceMcXSpW
V5QWWoGosZBtjb0KlbwCBITThAQFzkgNXmBIGy8lD0PNiV2jIA2mJAJ7lMIjdizcJw/KhDWev3uT
laLJzqEQJrc+QNnnlBd/Ct25gDeuDSy5Tdw+fnCoUjIgHznv1eLaJAy3+IKxHcXFrTxeXjNauTvM
9jUmMw7zC4vOYmt4bu9cYy3ZurQpgXIC3jUInc97CEV9yq9oAIJfME25sJM5fqrBpGBEmbay1CyZ
CL0bgQhEcXkAZPNytRKXXGBp4B2eeUBSPLQ+OhsCzsb7FlQRfV3iXwBNjdMovtZ1EllkqMsUOZ9k
I+YvXHDFcd+h4mUC8yyIa4+f4gAL6GSjRmtss1cnUbt4BZRunqckGlv/XyLnVwpKZQGmkfdOwWj/
kWziXKDqb8QVmvqh08a7epqrRg4LotNsWwgUpBRX9GF47QbvXzSNfhiWlJCDNU0vseG78b2t1NOo
s8DdUU+eWXOpGvW8Lk8BQ3eLNVtlIgQiXGx0z1RAIzJotLPuedO/8J661szY+wLCJuMRNeFCAsy4
Me2HVZrDq6wGPciCvO3VVptfBnTonk8aJGjOyull6JkZGGTjbb1/moP1P1VXFZRtZr3r67MySaTk
XQ/YQCRYAOEk7WVsnjs8VCHwQUie6aY7bQYVDRga7OnUgPE4W4wsKMm4zplSququougq79+Ob03S
ROatpaD2yOrTB/982tUKqRpf9pLtAdPYfOSp2yMZvhqa5BJIbLOhNDL3Sqm/Vaaf6DfiBooRrJGU
SngbSjGQ0v9ztoZ+MxVpk4kmELwA6EwSZVIIvDDdCnjYNezi2YZNSs0yO5AneCwLFXARFG8eYDjR
PzU+Vq/ZXbAagtBBbkW30YaslPuxty+NgrjqWl9pWqVzfHDXAQuUY1tj25aZ98RbHuEc0dnG1PnR
CyWnWPIHVmU8ahtikzP6OJxoLg8JxhVTJZehUXFISdMTfJhjY1mAhU+JaMlIEiKO+LwIN8Px/Ao6
7Soe054yLj99IOwRrL29W5AqONHU/TRmydqDHAMQuYMgaYgAlFK4NsZ4m4wG1zEh3OEMUE7/Cq48
VsYgJ3XL6vEwll7v2NTkp1cXvlESBDUNakso85bWD7PivYQwYVF/lraMa6sQ+//v2DsoIH28Z8Ue
Q/FimY4eWbbkMNumwF4Yjh+7Yi/PckCCesaZKADo/WxdAvcw9NeYRLoDl5o/F04GATC/pIqVpMMa
8VMze38Bs0ckNGhLWyRLkeicKvjLYVmZD5GMboQca4Lqtco10mOsSh67OjNfGwJxAk9hXb7oUIik
jROSIJ1pjL88rJWu6fJTyyQCilIS/qorptmxU7BFnBdbVPmgZjWx1Wdh6/VL22EyZ78cZJ2HtzwB
9P8g+LG0PhxW//jtUe+Fjg21b/PxwI/wsiu9Dl6561vm5gSy7EaGEtZPiSw3CXRfl1dunrEaMiuU
wtUzdTbchHENSHsll8pJF8WiH1iIT7o0yFVGDrWnbcyi/Z5vw8ymBI4DlbejzPZLLPJbIZk26DyS
acV2hZNxkvkd8/lbWv7Lc4rUkAkTQMaTc5YbxZFuWXADq+Eq3dLvnwMUzMHFVC0muipqI0kI1c1I
XvK6cDq6r9sZZulp7Trqideireo27V0fXVe+0/cF+IPwunqneJ6jQR0frIVOQuEWQtzKk9b+GxQz
+Wwma94AYi83ByACJLxvvd4AR3XmIiJYLdOctzXN2TcA8WylMPFrbZ/vnBC44UqcIDGrHcerEB9A
R0R2XKTTpuP5kIgUvdhACEzNLKw1v1rCOgg/BkL3aYi5/p4AB5aCap08zVxjQ6HBjqx8D2a1kd8X
lADh4H38iowzza2GDLChsy+5/IAVqr2R1KxJEw1R6LJKOAJpc4WM07QegkMfyp48Aiu66DEjjo14
lv/s7LaqvvJJZXSiFq0y3I2cgdcOyENxkYyMbg8lZOuwH8MPgUloDPOxzQkmBLgREIrT0phL+qi6
PVULSj1A9hVPvb+jOoUfY+B+sTLTqnU/AZHKIghrGH30fNRZ779T1nliU7/WxHUjDJoIkqpYEI3t
fUC7canQ+24KP+/cXq5O/PjLAqQ8S4dBvQMNCffOHjBbT9LCEcacYAR5TwN32hNrcWnjpq/Guoru
QPdU0sQ+dLPpUH5tGotK1N8CHtCsPDkMFxaEVWYmYiebO9PYkLbYMiodV5y/MLmT3R3G+pNJZJ3U
lmeGhGDxmlINrMVGhw6hfdtFXwZvNQ9OTYZ4j7hUZq+0QJ2r5aVcUzkXUV9hKnVp3jjN3k8Koy0N
UFvl8CgQ3X8D0/d9jmCnn3w9844+Tf0UkgXJnHhFiE5kyNe7hrtJK1Kz709tdePDvXrvcmwePfiT
FJJYgSlsk5h0FKX2gR1bYsvt7FX32eIX3373UiXgLDgBJ0ty+qWj2jb4ezHLTODEtCIoXhsE2rU+
doY7GE9d15PdZpJU+7G78YOA7aHMG7+L0TFinUI/o0V+/oYAX4LVQ/1HgKlrFY8sKjMpZOrTsNtJ
XeXSu+KUcSRBFOG87zQVECCkqeSIb3aNpz7M1sz8hfTwW1IJJEELAiiuW96Ke/cl/hfGSO5NQkPG
3tCYqQc4fv/i9Bkhr2az1BBqpEs2YFnwCnSfA0sO13pn41foDTbMI2Mmw1CcLLf50tAE0uElh0aF
ZtKMG4w/4yUJJaGl1Um1XWrO0M0x22a5tob1BRX7rM7BJjJW2H05qI9UxyIa9sg/kLjs2jOZR48G
9cQegLfDiQVTZTH8b+S3nL4IxCD9sDJqzJyy9pXSWdVbh2U++kOdySDQx4AysS6O552gAlPp1Q1K
N6Ao3lLPDBtE9SoZ/6gcAnAzbvXXyC8niLUIBWZ4q/oX1Hia5pCHEQScXjcboAAdrhT7onBYE8k7
UjCLFY/A4+3LT+jNRatvPUduJJ6cZu0IEt3jhLY3h42335y71J6WOtdtWraN+GvY77ERWPyK5fRe
/nsDKxmu7M/olXKtQ6CYV0mzO3LxxCCzDs5wCcc2xBDU8lFSSncbt+1ucmAdotcHoXGul0wEOOuy
etx8zCroLBt3NhK7OnkzqFRzuucAReWjLLpf5Mk64cVGvRDoBKja4DG45047XdXlkdceHZctMVGY
ZSEOKQcGHAio80JCHDjxH8FU9XkW6LRps4wyOPykJcZQPsyB2wnM79Ay22fsmH851i0sNfvLnteK
ZZ5Njb4sRWjMs2Fu3OFkn37FJlB5VuEKarDIi17fkGdOQNcI8sw5+hYO0RkWVFM5ItVaIVoDBho8
jNV6aIvD8orR2zS8Tvskgp/QfvqfSxP/f+hqBZWlcgI6TL7jkoU3kI96+mh7Nu88Atp6sUdWUg1U
tJPAakgS+fz2DoH6hrb5cR+JEmxE423Sl39hubGRLvg4/KVicHBnSWoD/Ffq0o+QGaKAMKhOtCLo
vzB5kVE4dqCAYe8s/p0FJmDqV3DqwRX1OC4U1bp8EMiDk+Q0oxcn2kcPD+i6RhXPVAAFH4WksH2U
d/sv0PoQpGDi49JSQksbOoZv6m8i/GrD67nPCbjYEt/S020FFrdQMGw/yBeZ4ITKpvYBBvVDZGD8
VlBhoUlEf9sprKVeCMyCsKH/hbh1cRUNCew9D6ZSOP1uY4TpmlIE748FrvBmX0xUrkEz/pd96FKI
g0hEOu8ONvYEF6yRMJV9zvcQrfWhnpAXzw+lm2YRicZ6HGY+h8YOmK7CjnkMmFeEDIZ4xST5wEhW
X8P+4i96JTk65eJIuMoJwfeQ8dEm+onhHSb+LQixI+XJe6uneO8TQEddS79v20MZ9xUzFSNwcqZr
6LjI3n4l4ZIxYqKtAVqj2zzjuBAo9+fK4jzLt+FSIG3+L0dEhPe/iEzsXF+SwSSLNVfXw/LI5aGG
xzu/R0uPp9n4nh6TP8aNqu+XjSXB8zwsRh6M1gqpPZk4alQcVMEeNMYGDmo18y2nPpoFHONSwJAa
tL9h8YePjHXAhyE8JV/thxCqhYfy1hJ5cceDbrq6F/bwxqVJh/2VrY4wxOsrFOp4n1CX3fzyC0Pe
RXAB/YWWDpBZmNbhhpvfN7P6VD4sR19xpfx7bOBvUjT+NTM7+/5Ir+FZYk3sypWm+XQGAqR/n5SY
kwE/duvYPqayG7Xrsmflq5q0s5QNqy4EsYqQXBGHcsfyXXI0RLBNV7WfhLAnnypiRNGuJG63isA2
wK9SyxoLFRRkeIEIAQc9cHxpnv4A8W9LgntJ3RoRVipC4BynCxVwNl4klClkI02DeIt+3i1Dhzb9
LdkchjNMemy2DvpyxgrRoSIcumlDd/5s5qMWeoG3//6LRkPUJ6hVDIjrbiMrnSIBsU+NB0JNPuf7
ti4hvecT+QlPAaPUfsKV7a7ypm1uYwpdC22gfBSCaE0WqD8DFP7X9RHCMezu+cL5XndQSXa9IXAC
r4zMNTRVgO/nQnXxa2oItQ9F8bxDTcQJDiRXyjO7LMqlg/dcLKpt9KxrB6+564X+6rVNHnUdLpfB
Ye2OLEJufG4qIfEK2hXWU0GAoIbKWtTvKS/t8eGm+P07FUS8voCFctz+wJBLRNt0e/BeBrmlTTFV
Ewvd/FPL2rE6FHrNqqhsS3H+VI7SNoXFYS48rwHU7YheA+kg+NHI1uX+BsbgFdC5Al7B7cJpZ9vu
+7H2JhhHBhn+pFs2P5bRD3fmqTOHzSeG/GPjIzQt2dQWId6dLZpTbyWvSKNsG7cqHDzraleP2CtO
FFPIvoNzWt+zJLuKMRmcM767vXusEzEb9XmiG07csiBQ+edS/wVE5pV0tZub1XsPDtrqScv+/VIG
PIIHtCSURvHmG/jAx77SjwURGGko7Gd7yJfOpAUh8RgjFF0Yxxn8JVpD0oiVfRkAJ9K8xiby7IIm
BvgljrbUW16ZvV49mzdayytSeHuUSQffnzz2iXu66tL8bPLJS69E8VHjM5vLvihOHUP6b1wIMwwM
crQDlIFGPMxtw7kGJid1FM6konlAMyEIbGzE7hYoREW2sY9lMOu+kBiEEI0H1vG4AXvTjdd1tFbh
ncAacEQbtV3b0dyXQqanmtTCgxOgfyrbYag4c8Kk6+dlskCi2yNY9FBgzQDov7cIDC8vOGHJ3O4C
4C4eG35/cPW28MlEU/LXKOxzPCNG8rGl4gTN1eYmq7PzfFB2y2ZOVekidAYVmMN+6hVT7oYHFM0w
P2R0ez7tC2Vsn88N7VFKg56KzlpYZHxzNseaVPUJ+wXFBf+P1X7sOQQOJDvqfUn2cdqzFQdZSNOP
t+DsLoDrhiroPmZHCxJCmlV+VEW1nRzEraxVZVvXc34beVopgzJIKPTsVAL9xn4660zz8TMChWyE
NT4x6JHFW5DMQZVKOuNmhyQRsyOwX79dCbaYEDVs1sT9+FzVk6WHD0gp+PIs6oU6n59oW+ZYeHnC
ewigToBw7X5bdxROpjZ/5eJDLfdgBxlYuDfKfQO9iGJBHP2Om0HJOH1u7QyxvoU5l87lCfgSgumj
slV61qTYjGbESkl64VZ5dH0v5GwFI/2RwLbDyXFfPi58PUFexn4i7c9V0YwAP0uuYWMMdp0UF4jA
06L/5R7vTz9vaQAs6lNfYSBe//BQYSpwuoJ9Y73zT/cX05+eEt/x/wRwXlIvv5KNigb13USEOw63
bxYsC2mP8/MsMwIO2geMPeX0VTZ3/t/Hl8233puS0fJbmZpoVw1ePSgC0jR+nEydqbJ7EXxqHmpR
UTpFfD9pZ7jsitqkZpZx6bJzB5j6WdDkvjEHXAYSc4ONyv9ZpGqt6bsgExMkH4iZJ6INCQNQzMW5
X499fyIuWHn5lvFDvEaKQpyaTyZ7W/CKFE8RUHWYC9waE7B/X8/5SEXGEJAYZuPxORx/k2kHqKvi
jdT5hi+ohjy2QWnIsO8lywUm7uQ0xEJcRV1OrfcwBOMA17hT5QfRbb9BKWhAoxleREn14Gjtaz9L
J+ez0rYFuFwuJZ9lTVszO0yfBLbimkTjjudAcMd33vs6fgY2SD7oF+NPpPkeDOUkDe7+p5kMdrJR
pBbK8wpE0FIhyGmB51fhL0GyLcmj9MdI6RcrzX7X1VSdLLIrfEvNACi3VlbdyLiHudIxdEIRAXj9
6ajGm91KTR1N2s2vUUZgloga3lLPIacoXJiN9k0B7UitawZd2BIfzBe/CbMF7PxW4HUgmgGOUUzH
A5mY2B6dXw0xIJst8bczdKjXizbNq1WeD4LaVOAfF+vPbbfRLGJELh0kwer/sY6P0LhFQsXgRFM6
QhjMzl0YhcMmmudzb2FphWH/PmZK2Hc7N+8hdtK/hrD+kJpA1KeSs/3ISeYvkZGTizvFIKjGFmDY
7dTUzi9031i7Q1USh3nrVU3bSG7/5607/3WPU17CMAea3f8zv97NAHVNwMy1USBeQuslFDI4Zeok
OUYTLRQT0aXzsGRrxI3puJEOB1anqGXezsVfqbzIZ+ierA8K0YeN2O0fyq4nlCMQM5tBEXX45KXK
FnPSJxe/luqph3mVYYluFPlOHA62gcA+/lihAkG2nvZGNZ6TTBp7kDYsNe7aNr9Wh2fFjRTj7lkl
tIaj1YFzSfa/105WhBSi3Tcc1+oqPnz3n4nCf/0WXS/I8iqLaH66NqJM2Cjn7w2x4VX/JAKEk9xR
l6q3U2DstRReexqZNmZhBO7slSx/+oIfnoMjaRkAJQJba/yowxZdOsTBQqpTfXCL8aqJSGoBxRpC
FPigkDk5JyGgv7muIBdbSuEKe0uQ4JeF1MhXvZO4It7sVcVc6GRHeqN30o9QlK6rPzxqpKF+uLxE
ZTibVC+QxiP77m9x/Bx7DkraUFITIx4IvP81dnLWl3FW1EbH6yXlLV9Q/aPWrzsU5BjmGDqrMYzB
l0ZfCAU+bLIlRT6ZZCnS+szbpYq6oS+1UXvWgp8UedBkBpqURcZGqedzY+8CYMRO0G8Qz3vtontV
tKmV1F5kFANpgimbBlrWzewDIZ6Mc1EewAjiNcTazTLzaK2Qu6qvZYAlq5jJkamPjcIDy4w3Ohao
wXcx5AXAPPV5pFjMeYdK/bq4Nq4Gamy+LDdASJSgTUjPdV5v+/31uwAZ0vijMdhBrMScdeUNXK88
9AWhQcxsV/zDLynDJ6HXkYzxKL+uEjSOjY5pxrJ5BfDCY48/+3U0L/LiPVDk5I4T/vcFCDLaoQYT
gWqUXUvkT3hgUpHOc4wCb2r2y6/fAPlExyv7tXhw2PdJf65xeREJfs8UOcn+bYMTGLKB5fBaEAEB
kKWPMdKnBF+Ss5vpQrRdkruE1voTaWQh34wgbA5N7J0/d+xlxs1vzwXbx3AkGGN2WW74mWvCx6Mh
ow7nXcy5JvgklXfIscolM8lauOoFPy0r9cq5J3A0Y8bwQqyYpentIpbI2d+V8216LWHjItQYKil/
3br4vXHl9/2Zr06y81J02OeEorj3lHDra7CtBzstk3zYfBh+Ob3ULvs0EgiSoouk76vg6H5+K42b
T2BCe3LXo7hxQXYOrW4adP/5ki2jba8e8aKN8AP0JGYgCHBGpGsznrR55kFXZhWPQTDtWqcJCTse
OwcVqTaC/LMCT3nt+rX9alfb54mR6OO7pi8r/4ZM3aC41OFVrNqNRgQxICc2Runxz5sKv7EwQXhf
n+pfz++zx1cUZYg/ayse7LT9BFisPM7tUuLmvSEkVMq0Ksu44KwBsUVciwwuoxEm0/i50sJjM0Jc
TzIpBgR8idvBZXs/eXIQ2NWO3xyKCAO0PV32uC+hKGwt3ykrQevgTcw2uepLH8TV6ZZ8h8vPydMz
9Kqup6RGqJpUONa7WyHzvy4MQglTi9R2XUsSoMQphS2tZa7nIzLoH7K1QjizXlL/HSQo1GFTY14y
1dWHF9AeVrNXjxHy6AUhcEf+AbhbwXquhW1SfJnv4WELKTunY8UEfXobxyRAzmTyIhVeVusV4Aa2
smPWIn1+0ycruj0fBb8EqdVSktgV24al/GnjKuU4OTFKEC66uegS36y2rd6fR8YWZyFIBhbqw2sG
zGgTKWgQRCVcXgzyTYoHcnHnt+0WqCn7awGx2rXy/IyQOCdSqTaamBwQ9msgJd8gP3r4dbvpeTPu
wKtD4vWFqhq/qRGdNYgXxjguloAIA3mrflDOoFuzHRvmbYRHAokIG4Qdyhj94KUrdTGjT6p9yVD2
cESHLCjfqYd6CeUWFSVD3F4oPEaE2lGC+2LVWZMSEhFSA4j4C0KM9AHaQxv+ZSihIOnLuw9RgdZn
X2nhsiPFlW3xNUhrWlnkei1COr7HvYlyJFQnZyAfET3K4RzDTQoHo3refzJxpguZN6XnMbyhAQvA
xbwm2k+HJJG00Tr+4YF4wadyV8DnPO0NvpPiAWncbtQjOcDevLL1l6Zhmi3UQoJgZxlOblOO+pUQ
1pB4dRc7e5cWJUqIHEexmE+Yy655U8n7GM8bXbjw4PUrql5RT07MeTJ7+4cSrhnOjszGutHnsHK3
ci/sTzFzJVarnjQM0KDQ5a3XP+DZ/eqzPSZgzeQxsrUPECwMDc5CPpMN9RUv4b5SPcfeCTLCPsTW
RTkCQq/8IoX+SRbO4uj9Pr18nbXNSmbbsYDgpCahFoHAL74N78epq+u0ePuK1IvHIJKCx89dDg7A
c9AwTSGeF+jKBgvSoT5giFSCU2hoQsCLdQXUn1lz3/W+NCsu9l1pO4SCkVtb8PCKO5xRCSk20LBI
h8Rt7qp3VE5D/S/5I+qwrv3MOKcl8bU3t7hLM1TV5bqTi0o7L/HMQJGi5F1e985/raDOZgv5SARJ
VRdZhvQxysQq5oEVmd/JH/1DEE8oKsXZOTD4UZM2Co1GG4ZGzbTqs4enDZjEXq3fN3mcW7CPl5Jq
68SufX6/q0xTiQK2KdYe6+HP5Sm0a1d/QCdQqPvMeIdemEuSh27J5yJWxx3yeDmEnn8TpwJqLw0A
yBMK9oJlVAniEEHPOntOwGIPslX5jSq/b3j1p5o7p88c2KRe8S1Gyc7Gwc7jqn9Af5qp0129882X
+YkhEFaxH8Da2jYNRy3IyfklSKQDA3pZNyikvRFg3OcGBWkdkWGVhJ2qwC5fG3c6bouy83/3cB0N
i2D9mJgOlvlZS4c4ezQpSfuCm7dr0KOQAXK2jP9Hj6Y9lB3BnkdQrYUOlzv9ZXN2lx2P1nnFUwao
tJ6Tx5XWlYTKrihqLcsz+5iCJPl4llA1CEtRRxvNzbOXwxDKmOg7ZMvdSRTF6AWupk3tCLXQcrWF
6p/MyJgzkdVXdhm8BOXJlNcvqoRsN/jban+zT/1D3cmPUNtFp1PbyF5lMSKBt/0ulF4UT7NM/eVi
DBK4PouvAywf7pluLMfS6WbMgkr/y2wqPhUbvYz+cjOF1T7K6pRGSbTB3Il4ku6jU0thdJvOnXSG
VVHtMxivP7P8NutFTnuHj1lwuOPQWh7GOHJOffx/sjg9656m+XlMSWD0Cdjj6chuJZbgqsSpGon5
cLt9HW+b62s93IYxN8/5F0jqSv4708VXBVfmQiHKGmx3PWUjzA1G847+WtVnz83UKGC9MPy8A9p2
d7E14/xBlg2Q9/pA2WSYMZ1Kj7ysGM7zvM5nqc53hU8SQA49OFIuwuu16Qn1+Ouud0sR9q42Q4bb
x2r+r4Pfqa7ss2WqROF43D0Uqc11dnIPH7kNaYeO+s3L/UWuU690KfTppvxmxHmuKLw0wJnQ7W13
ThojwhK4jboh/KGiwQVJF4JTpM9cj16xR8TWqGyvQPbruhux+AMqd0LbtKFSCg39hartifI0qbo1
3SHf88qhD5zFFeEy1MUGIFYMuZ8JOOFFB5qTE7pjsvUTaC571OQg0PzZx/wOIPwZ9eKvdYweaAwK
GLnRsmz8MLkj+W6F8wnsY90y9xycwkCofedkwTtFUs8iKZiQ4ddqn8fbX2Y6dDjAAwhZlbAhutko
/cvzxjsoiuKYYCIznCJabzymexAu7Rn+iPxGBVVIjnWyL3RzRFP1znues2jzQSyVOz/VwN1wF6c/
eNhhW2YcT17cHuSBEXyZcYREdw0bsGH6ZtpbF4yzTaOruXy39S2zgIIOkC0+DZgiVxjqm9UtIPoM
5BgFCTRBT8BAQ2bqx65ELeGzpt7uTv2/AM9rwYyYViGXPKtOoS02WAlDOwBb+SuYvUvxfwzAL2XR
UA5UEyXwVvT4T/rSWBfTGNEaAV5A490EuyoaNdb4HleZUlKcb9V9SVFkTOjxVrPG3QSmh8oLi1GT
P7w4QC+nboc2cAfjj1B2tyED72txxqWMybB7nJnqe/1XLZBnd+UKJdcDIe7OE+qAmIdD9qqfi+sY
tZWNd6eVgVl726reD2xuma5CMTsKF6csEdPSt4llEM/xTh9hqTN+Tf4xp6QVYltjwMLEIt33NDSv
jG1L/sr4o/U7e5pa5sbCGBCgKlLrffbOOeQoZRKLoCrK88zAPixO7ZzDYKc4Ek8yNobvq0BRC7dC
KJ+tlezws2ogcZi1lwM9LBb6hIomwmOezmr+GJBh5nb3xk6GTWwiNFevKkXFCIw+m0RiJ7J3fUbV
GFhDiKgF4vXuigntnh3kLL8pzSD0SDNkLDZBrJsSdSgAovk8XSJ0kgmuKDGCZNrmKg+uqXCvZnjR
xo+4x08cjm+IiGZ5v4yHfjvZofYMLzvNO/829CEDiNz+Q8OOqHZ6dAllL7XGS/MKPDhmIcwgmpnW
sEA5M3MpcwOwyGatsKj0bneFI7kcNiH603eb5Xm0UYRto55AJITg13Fhw71y4Nc1suFw9TblVs7w
89fRt/oHMSNk3kLBIojQClEI8+dthVM+/mnrt1RuNxDmjud04HmswiCeTpvuPIhEfC/IBsUV52Ti
WvKRhf7+vUBI82ygcUdk4KfK7i0bnsH/Z7fhSyH0zb1oOyiURrKfG/uy+qfVa+C559j/XYqRUZYu
MDdPdmqpKCkb/8bQDh3gZIRtr4nlgvIPvyOrYHe5aLT3coxtMYIwbU6JAljC/3joWNQmh7JdzMEU
INPdBfJqosjrwx76c8vMud1q54xmH8b0aZoFbORRDEbRUKa+PHoGN0UCk0gGfjVg6jmENLUPqBBw
ef01ym2/sO6tCmNqsXvV0Q0M0j3zEldUznLGtWIurx7cAhiUQPbsKcLhG+7DQoBvvgeKT+L3g0Ta
k64IYKbOeL2LVEFxkFBwqkUpB8Oxjlmy8jUXhYNnrcIy3DjFDiXg7EBjx0M7YwWEWw9Cz+wX2OxJ
eXsAoZruOQ1OK+7kI35sgbz6evp0eEmzWPUdcNaRy6bvfCYDaEYO6qMEBgl06Obus7q1IqHVLxif
AAYQ1mT+N4XQK3Xw1hC74bLam8YwbOLAyC4y1IDtRV6LO0vA0iS3mDbHvjUL7Yezpz9d5aBuNWAu
ILpPIK/srO8XJhhmkYPA7E/RydEJaioQCN0ouYMI4b/Kb4YyO1MoT9/FCwDywGllNcMwZr8pBWZp
0skHqV/POtUAqlqRiIH99Mi84MVxbGwZ34x8F+sDjA5s4HqFmo9AJKChQBW/vkAKMODG78/WNlvF
a7pHYAhmWV3rgnMEf7EOHvQa5HYWmrSbT1mInhkitVCVHi1L/ZN54F0bg62O7VweC7TJ12LxvZlj
iqVO30qx0VYuMhmw+Jt0riMMQ3bSDDV+4+ey7WEja7KHEXJrKzPSH7cVAs5H9wyxszL4yzaayJA3
Liocm9Gi+7WgePnzNOD5vpenf3xhaUsgCe+yMAhekdyYR6K4nfCxo1xaECPIgWGwcdxM4Ipn4sok
wWOtSwkHNPjGIiaM7/tKN8i9P4dKSal/rbdSUhKvasp+iCfSgtGpZIgIunXDWs4EcuDg2ZLipZX+
1O3YIp3MAbW9F6JOJqvmXTPbjCqcuMP9TXmlJMnAc6tmWxItuLADM0Ywe5OTjaD+DwDEhaRTHsw4
5KY1eVwAlWOhZGhawq7EPS9b137HNjH2RmcbY0GJFrpkFl7GhIrZdpxeh2MV+MfecgHwVb5Wuyto
p3N2JJKD+44qyRMsO/+mnESgl0t7h2FE/8s/yM9LeNnx0DPw/AWvvhZbNuBfTHHNy3jGdSJKd40n
fkoOQIczTC93pPzBXr2HgoA91sg58quOhgeAb4f/q3KduTFRAeu1CYD82tTPOnMCMiMRCfpS+hlt
rES1QXSlrm29JWrNtDRDhlsvyjxddTc5w8bxMeHur4bpOP9+aOTwl2m3OaWaTTS1YeMw4HZ7aQHi
/Omn5cVoimuvuNj10uHXjPK+qqOEutpGJaZ4BZPy5KhNLIYoL7V5xGoUR1MStJTYb3FfQoz+k/1/
bVrIvgDCIDP+a/z+JOru2HYXroqy7YwkZ8Rq6Pwy0EklKUPS31bbri/JIDZEvQDL/s7Xkq0ZLtr0
SxF6jkNCalIGpJHxWtxSOtNhZZOJ0SeRLGdjHLS6O2UsIWncLC9yRTFgTgdsRelr1ErzLpN8EQHK
BT/eca5/SVyu3cPsv5slj/l4xGwby5QwHokI3uRG6idrGvqrAk4jJjtidzb3u2GSjHEgkH4TN6FE
8E3KCvfcF1dGt8Px4vB0MAQZVRNBguC4FDvdAlIsiYePO2BXlAIJArgSV83w7bEnOq5794G03iT/
hNTUgTWtOtZLsJZpKLjxJJL0Ws6Zlt3n1vtni7r3ffQWAQMcxcQpm9xPLrmhHLAV59zXqaiBWc28
7+RMpNvHelo2hjuQao8B4uK4N9UlcN2uFqKufiUtvouiPFT4vw2mXIYYXqOnXmZIlIjDO1kVmxfS
cD1UDG3qTMXfWBVyY8qubchYhp6ogpdfSh3b0FFLWF+RQBy7mQ57jDaTxXITRwLNS/mIfrZtwiq6
/zDBIYRc44wBDNLnn5Bc8IFOJOP6oHHOioYD+YIJ7y8nE2ffYOWgdyDqorvJcZRGRBCnpa5gsQws
WSVWfXyt9PfR0Yjg7rnhNoVGaI2X9LrVH3Y0S0f0S4W8kTO34RgUsbm+lKnuHYQ/KSuCaonQbQUA
xniGACl7qBiLoN8KrbmcrQCS0f/fDmZnAtURN/Hb7lRlucxzCsPvX13bTKFFYTMZORuc+/DX6ous
419SxM9U0alWCcMs8XPA4afV0D3W3DMg934dQZvU7rXsqgGhSe0b5C+oDUeuW4HVHZX3gruk7Klf
doeQKLjiXkUy7foeazrZaL8plcSnwTiEtKsghkfHa87+DF0qUtdxpBwdgxcggJTW2J5hlRvqUl6f
8bpwTKCYPbZBmp2XNkIE5g2zKVhhPrevQhlX3qDSgNfa5D/8BVtWXnk+6ZBGa6E4zNmuj7UKbHew
Kcvt8IxHZF6OCiu2iIMzlca8y7VH+Ka2n47BDAq+BAFPsd+1clgiCA9hcf5g6ZOpGJH/LxMNdYcp
oEM5WxcrkR/a/EJWSfZjdR0Ga+GZDUrmBme9xoAf+MNYlIh3eWKZvE3c35SvqoxBwhGjk15xJjNn
QnK563iPvwsC6SN52apAoabKjCl9Y1aL6CBnygoUuF1nA2Y43JtfyK9esV5EgsCk50mhGkoPKLXr
8+Kf+QKUA2AD5RJcERdkvdZndKLXKFHoQlsqYni3EMehdgNrm7NAu4dKADRYL67CP8U2KmTLQa7H
h5WZP7ww2ffaSVdVke7afDtXgl/oYqCStpUgiauP9Lo8eJB6rQivXoSXvEaZYu5nfwb58RLbblZW
yOdcg5Gzs0PibqU7rSJ23Wj1Z3+nMJJBOvtoKKTC/tH6IEfklmjGYIcgqpyMsUB1yGehSQuvF2gh
ppb3614i89Sx9fLZRgnmUKXn4K+Q0HToCpuKOHuns3d47eHLjYS2uqNb5kiJvX5xnTeXvwo3oO9B
60Q69mI4gOYnBRmFNlO2zDo2PNhCMjBsqMrH8lWwpARLgQu2EewCqPtY9q6j8XpJMED1i4VOMU+x
FG9ujjLTh4mAvJ+Hr6Z1HEVMf5ZLkCYzRn63WJ+vWxWcaU+jFrZQeQV7EBRj3Yq1ZeOCZhKgTC3U
X3A5yPA1LPeCytDQJL1kXusrQnin0U8lxtZFPLFyiZAwarbJ/f/Q1O1OxkR54yHjejaE+7L9aCw7
3FdbhfzPcECn0MY+KpqrNwY10KH7NfkbG9CRxWakDpyK68deRIpDdLNLpwG49N9Old3mK6rZwYP4
9RtvfNgeOZBQ7+obD4MFXR4pQHYvH6Kj2HWsCf9mYwwl1GPKODyK3hgWE5sb0EOsseMHzrIMKkDe
RZH4uUgLVS3UfMV9wwGBWRAONs60neC0UTBXhmsUcB/X6iAmy3qiepe5czhLS3X99EpP9ETqLlbN
EQn9nsURH/rEH5Cl9d+OJDzg+6McthqXeY8CK2hcxN2Uhp7VHWgsze1lzt7mUMFhDQ8QebSIErKa
qrQs1eOt3Tdxq7o3CJisrmiqegV8EQOgCMoXX4ozcpV8N4xvtlC5O6+oz9nfRW4xLuAaNTb/8mc1
VxjfnUHsRH/DcrZMH6UfUdpBRQIXpyzvmqBeIJyK0b0dSfKi47GSvw2KptpG7XtO8VubaeEMNJve
mU9LPqgqycqowSWAUrHaUIQU0LWJxOt4OAgQhkXM3vu+kZrSCELohO2CF/3OGegiXqa3u1btG8wZ
e/ru2KlaT0SbPf9lE/gB6iUh8V4tO7DuSAaqlkY2zAh0l61myqLMFjOw3x/rEodJWPD0xlxM9xj6
gv1TlUeUxq+7dwRdigSo81PZ6fbN/dXvL4YHrC/le7giTEVFfBpXsnVCAzsPSuyWCOQC8Ub5mk1s
FJT0cgDYyklqFik+b+ccNLdYP0xMSo89wBXNiEiSQaIg+XA272SJau4y+EZnnMlRdzITb876Oqjz
n/vxsECqQNj7xLwqE4WMcMOlQ6ZEF0waklQRgqoq78LwAnKpucWp+RLVBVwNE3WL1YpHiRtjVkY8
S0k0Dmormc03GLHEEomaFfufCQBwhZN7ZL3AIlYhoD+CBxV5sLThILBpsEyIvgKa3lY8HA/oKVNb
PZUbus0Jxcs/LIl7OEuEXcCZZpf/+Lk8SZi05o7EYyx1prpyHC3xlYo9iQUNW3YmbMIcd4tLNd88
O7Kl9LSRI/wets5WM96aia9ZqZ4XQTCC2iJy3FJAHIKxv0Zti6D+Ihr1qA3chnhszUnKZaE1Kw4+
momEH8vh8FBiPK+u7fhFaIHjCDHhp+oW94s3xWOMS1Ms9YwuxXJcMCHzfcqDEbOA2LUDQZruhndq
yOE3mtjuOCMS0lvQgDt+5axC5X4h9irr3dPOfghiJk2PXbzEtgyb491+GaZzHD+7mRSweR3JQn0I
R1E4rg4VxEWhV4I9uf5HFqne+XaRbo+IOTxkMpvCQJ8mqxmpxcnrj6/TzldxbOTrLvBTE+6fxrL+
5JAVc5ph+nQMJxepDt+VA+l3ufsC0YjZTNRDz4zC3d6IA2ZVGAoP+0Ed8fYTe1N3ouiq1wRdp86r
aGoq4MNtRBuMc7ZmlsK7h3VsZVR0mL7Tn3mVWN1ir1bpl900or99BT9h5xjsOuGZsd3osqlQ9LXR
AWKCdfZRRXnsfNg7QZGV8pxSz0AKb/r52VoGjlzVw8soVKndg0cikrdbIIu/5Ny3EA/P83wMujqz
gZKeuFAUBKLtuC1YsO/tDlM7GSR9ys8IJELFGiLysO8n2cZ763oimeF4igj/kUM8bXjD4t4lWJFA
oQhhqiz2jCMYYC83Wuzji/lnaQC0T79Dqsj+B1p7AxBMhLdttM3T3cWNZ+i8/ryIbczAER5rdkat
HubOK6RwmdqEWXj4lTyNhvNnboK/n2hOaoP1SH9QFtGAtZMO2t9elZmiq4SW21ZZkT+kZ4BSSgFw
nnaLuDY4rrHho7DD0w054nb4qxOhx9mAmoCQwuLT4qT/nCm/MarInE0rX4ZPyONLSYVDRhbnMSsI
BdRYAD3xSzm6b3lTlMhf5czwCrZgBBibuuNqXXb8VVGmsG1q2oxZa9gdkPxcRmg8foNUeOgAOQZy
XCFcIlsQMAcCTISxBABDGfXBjLJmtbTqMrGkP9GTOsCX54aJTbCHZdFEoWX43jqvX2w4yKsGBsGS
zF0t7oFEFRwqxpUeTKHudi89YJ2V+f1zNgaWINKwQhtMkXRyuKg+HdpKDQ9uD3Dj4k7JYZWvevnb
XZbTkuV8+ysUvvfn8FqC6MqcMDKXIW1vZzmFcdfiGl1mKRFJ/L4zQ7jYIBexbGgvAoTQK5G3BWFk
q7eQH50W5phhrv1tMQ+sMqDLt905gd8rpOtuE3WIjZZsijCWHMxQb7xBnbN3RMRJVpVcazGJYLhW
JZxflDewUOVaKLfboZv/G1dPrsN76N+rSK8l+fqK474XXQf0kv5IA5v3BHQdXTojnX+pAnBhaZ9p
e7Sf4WNatPZdm3pNF+RU3VOWQ+aVKC3Rt19gSKwG+1mWv6EYgN4AWUAh4yYVHN7mK73HM4/7lDin
SgleTrXqmtxE4tYnpU/JwiRFUxy4oMUYYRk06XWFfszEstvncoxgA6E2dbpD5foGsgyLR6/LZill
zjgFWdFsufvWXVDODl6vfbwcoIn6fYqB4aTOLkYzY8ZwthIT2RLFj/5GCK9wxB0fYFPrg4W4Fm7q
3T2zMTiuZ9O0JeoxRtP+wcRIJ54Vb6keS+MUtlYitaJea2iC3ql104TJTAIZRXE+WUVZ0bT840sr
EEmnjyIzQ67zbA1D3MBYyQ7sAQBImpSOtOJkhkAKieYYFpGU9ma2p7JAhuvF5HXfs52azoHB6loU
EkCWU9hTj7TunxmZB3ylxwR8Q9epEDp+wNGWk1dDAdlAoVV7ISFdYofOSGuFdrJDsD2jqUMVqR/h
hj/VpYt7FbYCfVMLYYpBot0DLAq60tlsusRYJ6JAuv/XrAJvOOyzUP5FRwbsc3LmYsLWYTWq15Di
zLo4B/94x1kUsKz22JfLrBruhxaOlX5Ns2vFptfEJqgUmY2NuMa2e61Q1VAGgyASizHLESPfQGDn
XCYapfPXbo42Gw0TBIRRTMV5sHFfs1ImKO6a0nwHEnvrpM0jFnTXIYoYmkqOTzhdchK5R9zagsBg
HPIZIbcdQIcFBTlwtK41HhV3ADBTC/T+5L7H0O46eqtlsfSgjYPIWatBs/mZAGI0t3ED7ONAkk1H
tlm7svyiKwNUvNXZaG4OOq2JbMQVR3cUOmD6wdWLzsnrJ4CYIkFrIMTYmPFeiKB5A7AXkLdMqQjs
4R/C4Mla9FqSWbEcnSPDeM3mQ7cXDu18RzBo2WQt/ZVCwrk8wZMjMBFLp8Y3hdRg5h7f8Ncoi8ec
SydL9CBli7ErZh4d1HC3u/wpA2hMHJFNqrLn/i53yQlbUS0RayFVZwh6ySbZf8fOPPDF85yeLLlM
2DR6sZDRDF6qo3Czezjcf/65ryNC8rCd+1ECycCRfsmBK1SYVOt26hmxatemtpqxcAhQGkZSM51r
7KHwtfCnQNyUK2WX+c0iMiqNsFZWt1w+Cm+WqukbHbjce68yWv6V15Uknkt6sgYBU5wevQdo2tsM
/zAJgj6k+n5MJ1VETVV/t/N6A39zNeSL6x11YsQUctcf627jFhPsNIG+neHf7HuyX6VfXicP9h5O
hY3YeqbW+f0IiLj+/yfViaM0B7m79bw43CTdLmUiEz4IyiVI/KurtAAsk8+/veATRK59mYYITuTr
KF/Z7Ju1oCcuMW3uGhP4CL5JdFZad70BmyjQaQ36UvRppNk1rDK7ZZCJVLaHlB5BxjxHfqGiy4RX
1TWBDYBXjATBb1PeOH0Iwmpxt9bal7GzTuF+DO95aYOtCM0+dHRU6DvjrQgy2V5YfyJhWTWGWChj
5I33/g6u1K2zRyvLIw4nQhEfRyOEzs81V3/J0nL7voAsnVTBjDIaJymT4dHYKGCycyi2uTjesfNZ
BHpMmSn+dBvMaGGV/HbMCr7laaes6IeIeaTn3+o4AuKsRYgnUaYkv34foe1aioZ5EZckGzVXf9tW
xNGAlQv5y3fvieVwpYx+Px+gdPdmXSZHnkg0hLlB4DXp7CpuvEc9tt5Qxiw1cL34h15zz56TFAB4
LypBXjl1QhsD0BQLyWNoaKseP4DZNww1lfZ8Xvn1r5zc4+uFGq/7vvPYwG8zXPmxDUpqn/VOxIzc
bLJjvMPbwqmzSas5ZGiMnqjpbx7X+T9b9tiK1Dmd0Xs56QHO9CNp3jhBIDicmurwA95BjqXxlBbV
+R/M1RlXAi7vSAM5uJZNQmFWT3Idcgn95KhyQmYRy2CUMHxRgtJfBJI0lxP8DSDQB6X2dflIMu2b
yeFlgdixSt+hI3x8AKQXMKzp/Vf17KzizAr8o/uy1GGh8oS9sSCE6z8iO6Ko1qRr1RKPW04SeLNI
zlo3Hc7vnvVCMj0HFoeOcV34V4wMJSkG0AHgD4nHCFF3qV/zXIK+NJfbbPch+K0HB/wPX70Ood3t
xbVBvCp2PkwrtCH+RqOhhUqXRqD6Kvp6JkT+pntNIkL+nJhNpbbH+vwPcGiW2nODki7nv9Vat0sj
kql1HbJkABIil/H1uzqS+QAR0vsh9/AJviPwbVJDNP83KVt6uAKJmGuk3dj69eUeapb/pmWWnAcu
A0f93L0abOGBsiS6ZRIq4zIp0st5liigG+/9sOJZYg0lDZIz/NzdW4Sk7CSUh+BDPO6YKfn/MevK
7S3+0dkgYjWQey6iq1VeyWEJ0/1w0tcsXYxhd8fMayWJSB8uSJ968XtblwncyCFFZkRt5JtshZKM
B3j0Bu65fx7Mt/pIRfc4Cb3kfKMco/nayC0GvbINmAWaF0aHCYXs0Z9wAIcRy0bp0vUWFWRYlbq3
U5pryDlwxwMwyHj7iuabWWSlPkwLdShjwtqjIx+0Mg9tYQqY+adMsk5oQjdoXOY0jZpTQ+xu/n7a
wEwwWxjLA5KyrUuXNUtFaUdw83aVz0JBXB4H+im1svHg/FpL8c8GSpoNoO68qWwXV1A1vaND8xc7
Z2HhciyNp1P5IQ0zOuIZZWLMMQdlrSMBI41+FkxdKHlJuXA4epG2XGrcg7taeWeZw5nsvlYo0PnW
DZbk7H1Zkl1I/5oE8Jdv/beWNioVRg2f2U9LjiEOk1gQ1byWxKp3ICTLohqffExgDj8nKuKUrO8b
G4MLdrDmIJVGgIChN0pF4i/m/kvML/ZHBz2Wx0DUKa7mXqjYI7AgA4c6MfRrP6kj44eP9r3dcwZq
8bNxtK3/3FEPWHivYXdJUhxIUOADcp45j96Lcmv298CJN38FqP7k4juHblGt/f/Vtmw/udIfdIe2
ppRQo0hCLkSfUWfLgVLJjIu11qQdCUDlo781PXKYKy6iK4L98gnyDVUwH2GiA5SQjevlFzanwxAD
S+moovfxJfPGmuFk/1EvQGlQo7Ib/EyYqurvqcU0szEBXh+IxhIFsSsPZ5miIPLg/u+VlnyfLwpC
SEQ+jiYakAzY0M73sFjeIMvlwsbmM7qiIIxVyDI8BjUgkXNWXujHOek+YjDiK6zw6uzIHo2+44QA
6qAvVmABmZmwxNVUEygYtku7ufPZu1GTBomdPjaPYA6w9pGZk1yLNe/LjAf2ZS/jxUNiE8HRh1Fb
h8pHh+0Bb9ehdK0yHuS1bkOpucGMMmeeToVnAyfArsuHbK4d+EgJA6Mq+d0Q/Kg3mHt8Hj1wuOx/
4gfk9bdp/8w9zElyrJ7xAgKvpsbro4Ju8qnrslA3y71Sx2evUw/rZR/s1DR8pWP0kJdT6aDKvDH+
D5Vx9FNXkRZGDZgXaXIuPoumjXY/j8mGvWhLS7cbSI6GAXexdvb01QLJbYbXzVdCpn2COKfXbu2D
XQfRfVRML6T5vfUHtf+g7dSXc95zO04wRooj/49unLSVrXHXyaYqKITBW4xSimXIY3IaiiquRLnX
o0lHoj/VWPmZQN1D6XGWzGxn6RFXvK76GurMRAZIK4PkD3Cb4Kb+Gp+yVoWwQW7gMixezA25bBiB
9WgvysaFRjfUu9hc83h+VfSKYt5VmOSqk5/MrfuXcNxPXO79qGlNthJRTR8V3YFhI15rwEOG2zRv
hdJEFl6dz6jUWy78Kp+sd7J0HKAX2YlRwv17qg53ywEstSFHj/N3fGSzzsEtjtzPwHFTX3UIMiuJ
v1gyB3f6HzCOY4gxo7fXjpJmT34AmKRej/jolehkT+OMHMESOYQleH6W+ki6CxKfqVnKiH78bD4O
DveIQp0CvT/0nwbQB7gsGqUSy81FMIol7yS1vGT9sy7W5IirmJf2rcoJ/HF46y8jdsligLjNsWEL
q28eWI7TiiQICmneGj5rVU4C1A8jjUCC5dP5BCW3gYSHAsOOUwEbn/Pl1Ir96jjJfU+BXKx9KWPD
y/MYKxg4OHfzqUByqcdR12igYqWFFX6kMGlqVlbSf1eUliGdnghNw6IiK/ue4/VjxYmBStsrnN0o
XliqS/chDDt2+/mGIrd0mqTY29FRtTWEU2OQVglZkN4DFn14ZTo6wb7YCRTEtIJge5PsDb6pyUxq
48ZXQhO/Cr8FJrOvsluQWkRaIl+CuESVAMw8pcpPzbspFkYEraYm2Ajsy3KRkr8rbiEbn+P+VcOW
HIofKRr8O23SI2SC1C+Wi/09ObMv0dCI98Cslp7a+gzp0XxhSx0dqMh1ynbIYIU0gL8Cx6oE5Yqg
FkXSQdOC/vy7KxGbS+lCSykJ8+ILAjuY3pQVK/ubH4+P46u8i3jMK74mlCSzrqnVYixlJXoa/fp5
s9mqgRbsKwt4A6hRGEOlwN9GOqlfH3nHjhagfIk2EJt//bq+vYLIDidhl64Ljh5EUMGxUaxAa+ej
gp6Rg3ZBlvd3N5860tfqz8HowisJqf5SEBgCfNi9mMrSdQXJYb8dBo0eU5MdoS6ZMhloGQdB0a+B
9z8aByITk5xnTdoq5FYCwZapqYxTfOHr1+948R71FRgSLf2CCzUVq45e40VpsMyKFXKdGBwMvmr/
huEvYfz+jPdf25qcY1ZvoCz316t/kWL6cvM5lZ5K/qlniC1Dmhqtwblom6SvI6sISk9fV0vObZJ1
8t8/EDOdR195i9RmG4mvC2Oqpa/kSztIIfHU5nn49Ol+FNdxlHetn/GUXzFYwevBoNWXr0ks4VKt
vvzdxaOE1xjDF5i5/EQQXao8XOEbPnI63SiKiGC2zXB0re4VrfKxVarEUpG/eRUMJjywksypWxEr
JOgqFPjwEBsYJAgmXCHUV1DKVQX9hK9oZ462wNBOUMHSXGgwCccREW10Z77C1MW0D4MKrMnno2Xx
SujBfFilswIotvqNbmvwVnVIvK+/39DKip3SG5fFDKpvkhaVaUQ4k1AtCuIWjGGw8BOhm3Uv+7GX
7fNTZlRXMK6WegCDOVcb1DT4cb9jaoxcMpLURbtr9bakKFA0PfEWLmZo+LavmT12Vp5aOUlJPTyQ
n9MsfErPuuU/zP6A/eyoQI3qzUw1yXIuEf5X/TvLTGJNlQ+NXjGoaa4OJR3a+msmsUbpudhy3JF5
3grnJ0luG31Aj1xFJqKG5IlOlDOAKBosX0ZZDNdsIg4IFwLxk6juDy3j7gmkv+YlO5AYESIG1MEN
WU+TQu5AXnwzcd4vj16Yhpu5+XGxSml82XdHkpv4SaomY0SMP65vfY1DqZn006Wnh9P0pANK7maK
4MKfzN5GW8RS91X4ox1lV5eb1NY8Y4wBkVhgj+81FmtLm/fR8GA93LLijY/Ey+P4zi7PUi/BLJJf
GeMZOMEw5AEDcSaXeqW6NNinvwfFKuerYOYQYLDWagiiuwFOG0u+HK1WAVz+TZOeuc0k6+8V/Ec0
1/QQgbfvZthPFDYIC5LSYcy3RkvTtzQ5ofYYGxVuhV37ZYNNg2/y6E1vciEd5Y5J0XdBupTPNYZl
QToIuLj2FoNFdivAgTZPW0Ej0AlkKDR3WjUyuR7nPd+9MZn0dTMSdKjDooFdoEe0uty1FpWThjhm
7cjxRHCSum2TQDlfWXlooWedCknzo4L0cKi2yjj7o9Vz5UJftCwYrKpgfCu4vrREL2wLWX3eLfte
kgap2V2417fQxqhgIGq/fkoqtSuyacIWC5ZpACe1UgoylS0vo4gu4oALBL7JWQ7hgn5cS6VV6lom
jGIot3bnX7GufmkJRpQRh0VxhJ1rdDfHGJOC/6nCeBxdZLnrkc8Lw7gngR8wuVxq+/ar2OwEPIMR
Jww16xYsc2xIYt4cnrOTOalrlngcGml2ZEJIseJZjUjV3lANriPSowqeHBFCZrJ7U98i4nhLJwDT
6gMcGNNqW0Ubb/wwdE3a1ZQvAGx+Nifg4z/KpMCOmT9AMjGZOxhExZZwDf9/8ROo26+NcJdS+gRV
Eo5A60hAARlvPYAGE2LD7khjC3/BY6XWtjzyNsNXLQ61dA5xXhzdslRF3N9SayCt5guWA+kj43Qe
Ks62f2TMtRVhLv2Bb8+dP8601cHI8Lp1swLQinrlrlLorKby6BFQn02D0V6lg5XRcf9P8Tcrn7Y+
povb2P+NE/8gXzAcrGGgOAfDFb6QwKSuH6Rt9yFCl/roj/fU9Sf5vzzh/bZDUfl4arvIZLLM1IPK
6hBV5uEgFMropzx9MCL8NZdLZD3ENpHo8d2hqVa//aFNA/CP91KYAyUYlTpKt8bUEp21ZOMGwkN7
OPiOmlD75j5Snv0fnmrYErrG46Vm/PiXaBXI1m63LSmkZ8ikO7VDRCzrs7h4BmT80uaSZkXa61fg
LXPNyTcsKum+vMr5HRmfzBtYH2WkMlwU7qCdg6FLG2z47uWOsWXCT8ZdMU5Fz2vJmUEBfRajFNE0
XkX5fEbYsBKcJvkdTTL4utF4yu5y/2+B49q0Nsh+a0h/GXxkXt4BbB8iajrmrzI3solgSS3ZqWTw
zoWHGla9+YshA5A3vDSAaq3qpvA8iGWb2TQxGKW5IWbm9hzPYB95sU6HWDSl9+5deswDao49BiZD
wSpBtDAGN/3GO/B95l6jegsj0imtgh99mYnUjXJh29yxMbCfNXKZRJGC22SEuOqikcrtDhzRu639
z71aLqBugDTHH1KwG5BxPd9jm0sfea1sVP2DlKUVOqPOSSt9dK5cL2jGfUpWc7g8T3C4OebwxW63
9O073cTLQuoNARQHVGV0GUsWnNswJaKXj6Zpjhds2yomXBblXvOeCL8Aj7YZDvroRFWSLFne0zOc
tyu1Ycim0O6LylVqK3JU9L06VKaoDlp6PyGsrtsXoY0Tc2RDkWV7Ols1fW6ppBf1rHNVKW0Ms0UB
VoHD58ej+T82lmZdj8BxUg/OWh97LRA0OoCmcCCHIXhKhDx7RiK6FebvQ2xmmlg+l0tKNR+YOVd9
pGaMUPWrNd2jfwB7pUqs6CnE4Vk7iY6ZIAiYLCBT7bN3GgXYTSnaR7q6wjNILE0iClw1R9KeHEWF
CigRzQE2J2OsUjN3keqoC6h/dUpwCuQFJUZO0JX/OC/ZaqA67GnignMmFCt50PW98AzT8L9veQqW
4IYypXKBvzS+QkNCovjAj+St/Yi9C/NVtm+DN9P9vtZ7RZ6MnKv8FhlmRWJtdZjULmue4BoRz5wa
K4JgQ/G1OYJMTpRuPMLKjevkc1ZReoY/a9bgtxqubB8fAuNgkEHPIydx4yG2m3lVC1Fef2e/wguz
N14V92fiuEPIxJ45ZRBgw+jVUapvdKTwxwR5T/SZDNJcdxQ70kjLKUe9/CnS0QDs3iXSuYTTdhf1
oDpjR1qNIk5zr/uFY6CIUbfBXchQA/VZR8doQsKsmoE5RswA9lkDR8iwqd71D0IN3DkPo+X1RH97
9/2EfdPFYlEG5fxkm6wyEbj978gSS5fS9LI0HBVdOoznuJFFGULs1b46p/M6biq8cdspt9b9X71y
0C1sVH6MVI0CjlYgjBn9IiBDNBCvrMMyn7efNsf+i9BOM3lqey9zqqigZYFqHlsugur6KDPex15F
Ta57rFxj1uuDO1rOnVFtO0vyA2GNem/mXCVTVE7BdoEIj5lm8DRKcrdh0YGlfaMfqSZTNSzh2MdR
UphCuoqmkYV8SkDbz7NJCYYdMlyEAMWKNCU4hDB5mOiTHc3r4HKZxn5AAAI8Tf/Qyd5pywdGZEcA
8wCrbx4Va6MBMOlP7haFhYdLAWbsks4Ia5sIdAqhekvjOWeuBmPzrYqj1gCBEY4YSrHpBi++GVM+
2Zj5Gj5j9P3DeEqzKUFp0K80s0Z4AUlDZ3v79UsoLiv9iZQV83VIGOzoySUKphxDuY8K8WYIoIK3
GILuiw7Z1SVCtsVRjpJ7E07FcCBjlM8a/cL4iKkyXIha4+xJ+MS/ukITAL77Vt69yolcb2VfTxN+
IOYJdw11VCCGrByKvf1TmRL4HTqxybQWLVM/7CFe2p02ZfVAZlp9lyCs3cSA8YGN2B202uBEyjYU
i1sZRPseyL78lcuQYHzW6ur3hkuur1enc1NxUqobMsz8X2RdB+MATbRmZZMjclHl8feweR5/0kBC
OMhKBaCCl1d6w0jqaYqkQaCPXl021EAyDyxHMNtqctOy8LLWfSfvoAMgr4GaYhWONIl19G4Ekz6q
MuNR+j9If6zTY2OteLSV9ladZMRD2UN9d2xNU+ZznFycu1SS3Qnycz9sL5V8wIbudqwFPqI65CGO
FgZGzhEAyEvJVVPwkyEdV50IMGfeFtqrnuOLbuIE8a5bNhj3p9R66anDttNdtz6tny9YTPSYSZsB
LT+mBZBj1bb12Djd/+yff79WaBgtl8QzQvu/tgJ1Y6o5qmFJzxsxtGGYm23vOjk1LYKR/nsfVLQw
vj470ysaLoGNZwKoucqn0suTpQuCAWKu1feEDx+1ak+sJLjn2xB15k9cF1+0DPGUBcvkYs5yvbYY
WlXGARgrmG6BzFeShh+KyeTP6JOdBlWV1NF+e7MZL2Pj9/lVbqBUf+SO2ll7ACutp7MpRqgSKwNU
8zep0rq/E8u66cukXhwyHoDkHFX5KUnneBk8C3IhIaDfT+brucPLi4VlK0+NVNxpScMoCIZDmO6j
BUtBG938NO7kTSH5b2NWpsFzQr+YbR0GHUaz1GZqRHXiWdh+f5aNayl+FqvgJylga/FxhR3JbxFI
6jlHhHqyjwq7KtlhYrpVryq/zRhBBML9rwvg1xzBlAgsSf3yJV5jEdwyIDoykDW4MP6cc2RXPBtr
Uus4LYfDJ928c3gttVD4CghC3NzFVfzbRfEbHQsZ4tSGVM80F5vdvEN7XkiABrjaN6Cp2TPm/jTh
ClqpbTBxFExIrZRf1bOyY8CBptfDlMkGCLcbv7ET1ASLoqVWqiJEdREi0JJJrIO/I3P60zEdYXJB
fK7arcsK1cmIyRYgAjPsWySg4wmmePBEkldsegE/ylfnZXxv3SkjLgN6k/A1Q137O55LETWTpAke
sDpwISVLj9+xN4FHtnuF8o0OUYhKE8/ixB3fAgTOV/Wzl917JIWWi2nVxRRW7aI0799jR+gsCTV0
owS6UyO8Nh0HVHRDmtzC0jkk+ZsziDWTfJD8Gi6Bz5Kdq98FIap7KzdxSe1CpgjoingD9PsYMmBc
FV7cb1qgy+S8DFhbLgRc7t5TeqYUJHZ3xSytKpyH6t0CBUH+hHAS1eFzGa1brNOlCxC1VOzBwgMx
+Knp49cD+FGoB9O/xee3Tz/5DMw/myIxsU1oYOaHv3aZdJ/kB/sefKFaFgiQ4qhTvwlrk1sakp20
d6tN68Y3SEF7pOlBIYlV8mj0BAGmCVDQb/oGU8gNw9iA/nsD/fq0rRoZgURjjtYD+iuqCG/XVZmX
VQvCJK8HpMD9mJyh54frgEromwPaS8jzwhMtJW2dIxSssgdwR8iTRpC4T0ohiWp/JJ+PqRxnKmFr
+PqgaiFgnmYC9Tc6lT/FgjBcSi+nxo3tWVDuc902RUfFE+KspYAIqC9oQ1bophYNf9xyJ2MvBdGJ
h6vF7w1Jf0DNKn7FnGhDz4fgReoppqLil7U+lULI9yFCAgk9l1QG3LFP0M+ju8juRUmynpRFWISW
e9UyNHlKwsKarMX5qNQvuShmvQomZSwjW7biZ1JDb5jiJxzDLhnH9soAaIWbjbRn0E0nU89SHABI
0LEqudib1mS9jSrEFiJYqtloziwzo7NS68LoF39AoaBobs0CFfnXY7cO1uRWkZmfLjXX/FZpStjr
OoLXTfOgtgNfK42BUPainD0Ca2h2UHDDGpPevp74cOrllhf6cNcMX1wgykx0YSX1fCKbFpmMnFbl
ZSV9z7kVUvPI3iJOh2yFVwEHdPq8scgc/F1vd+lR26aAbF0V9yl9PcL2UEmEDgx6z5pMJ3SLnx+F
Kd8ve/XPdxcHCTXCp5c8VsNSpbnmyajoN/JQRTADj4defg7Ipw3pkRsWG6JXLA4qgYJe+V3rUjGN
8qjK37hGSTrDYXkfs4G/8iTcMASpibEhtzrDXevFRMB3USotIKhvX9H551ussT6S3I2Dt5sDct0N
OfftpR/TGKSK9GXDZcrPgU2RfGnVbfi6YZ3xqCteIrOJuinneA5yOAERQk+4GIXAZg2+7idNkbwx
YaZ/g3AJBAcUj1xbuB6abFv/JT0MoeMHqJiMqD06XYwxUEESRz3tZaB9wyIlF7GgnfIH2OjWgs2o
hkCkMHDGpAjNapVduyr7jsCVej03ASPOFDrq+0AQsCKFfAnCm5IJAX2CBGO+YcvWRA1jDpBMsEVZ
KgGOlPDQBxpAJ/X+A5iRudEyy2o8e12l6VvIM7esDdU60UbkhuKFGWahHROXGuPtC+BmhNK7LYpL
zRca+g6ToA+j9SXgXIfT/fW+lPP4/sTv1WK2WgaCvl/70DdpYJFZEVtnCG56PCBP/fue18tBUqw7
ditPp8aD8j1ODGNz27br3QuRlk5mdj5BseXnglfVfIx+IiuEjLY8QFs/dONTfuPec62PP2wW/EoB
SZow/F3XydDZxaV+VKQGeBQSMImSoBotMOi8FHxWoICVB6EH3Gx0k9+BRDUuP0mIk+bKG4K5nwxj
qrlrBWusdqtY8MycnBX8tcLVG64wY12Bypla/Eb8PS+JGPkU0h7BkrT0gZx+UFtI0UAciJx1Bcse
GExJl1074Fh4RH/6Pe0EQQZipD81nMh+HIB6IHj5XRxPZYKQ1gpeZ4igfDfcUf1nbcczue5bRV9F
WNyIEmRXlK6u3R1nr3XXDV3ZvrcKgGIgwNlxhZSy5UjdIZ5/gqiuiZpOvKlkT5V3m2FUYqn2RxNH
OvXMPhH6V+2fBP/sOnW7Q4tjjeNkekLFhsy9U3VdD0ymAIbMpARgFmJqETx0duilRdmfqB14un+O
y9T4agO0NsuapIrJOAWTrXU3H7q/dzpu5TH5U8x3AzDCojOGSyT2WTnrpC9pjgUez6t2WJgHzk3U
KdflgUdrEpxPGkoa9+HYX6cGJuuLraYeKfPy8pjV4xEyWAGETw/OdwjBYIXNeEGioNlXsnUrZeSo
SodwyvhSTMFY10MW62aJzOtHXXi/GAbyd4PPwd+7w/q1Ju+3BJKL8W42QknFXWljOxG2XXY/1MQR
F3kGXDOPjIbQ35oayrRVPm7FKBiEZp6mxfgsG/F7JhL74Wt0VTRLmOo197ERTSc+XR+9UmEi3oi2
MgEAypaHvw6Cnj+eSduD+LHGqMiTWkn331annYCXHqYXAiOw9C8PpJ4KbjHN7MqvGqRVtlWbcAt+
UWdwSQhhVM18Y7l4nlNA47YxlhkgNKBdj/rZFJFJSrsmgwVCcJohIRxfug2N8FZGOtjH2i1tLp/s
6dQk9u4EOSB12onqrCelGoxejEPFxoV8idQumEVzN3aLw90dzIFcTTWO/4pEkUQgDP0MZH/x3v6w
0OcbW/740qAubTouUWYBxh3mQ2HMguofKb+mcZvFST5FAvoAHI149ijHZ2Z2G6mzaZAidfO4hARX
L28apPG+R+3l5XVZgKOzPhTwWA/4q0jZh4jR5hB4Ib6ny3qegm0L6txrF2wvUS/3YMI2QRz1GNqn
3nu9NrQk6XX4DZPwaS0dqGfb96traw9eqnTx2aO7d+BHP+rtDans8OIqVkLp6oUrtn/allBUf/Eq
Kalolw7Ud7WMB9lTqWBZpLgRGJHAXHGXVMNRkKG8Q78vb8z+++5BzmZYnOmKP8gTtlhQPWEI1P7F
vY1idbAh0tfHvEtZCbD6tvAfiMU+jT0oylcExw6KyPfr+Yt/7GduSwHstivIp7/PGCNQx3VhMxm9
OfnbFhRhcNqdWLTTg/hKSVqRxJnItcxhRa7l8Ugz22gwQ93hkjVrdjJBRCfkxDYkB87xmdUw4V9Z
HSy56AQB07KH4lf4NaTsgXuWiVYD9g0wCmps5GabTSEitMUtagodnIcbEWOo67MLemw1s9I+ez6G
MwqbWH7tkKG8HR1f6yeTmWOLYqIiuUyVyjQvsEcdwi+rDZY29nua/BKpzcame6nBmxsdlkcbuSEs
ZlYMB6gjUYfBfzsUfkLWiZ/YGkSetRwRVFgIRXxI+A0ID7bks/f2oQQyvCVn+Ylt7ngH+yhY5buv
HCUBDoxZhP7HSid9h6w3Mq0q7s3V6+wQpaFqTQCRCw7WT30EwoInVFxfMOVYdZKQbIYc82wnZpnP
RBJO2HjdtVdCe/RRWY8JJO1K0qff54EjkEKSzlJVEpumjaZba8U+dbvDIDqRKMWWX6zYjjDdfI0a
/IVes8GycdHDDpVTrNjikIfRnyBQa2IGXvhN6aNmBEdMt5Gl/DHsb1q8ZcboogUFRJzLnflS1BOz
TzsrClYXgKV0Sgl4PDeEBQjz4AB3ssma63EmUzMn6gQAAO1jRVJ8ZcJZPbbMNoJyvl1Ypgodo4uO
5N7Z5BAHupCLsDtiwdoAtD3WnxnGdNc46svBhpKN5vxzIRQDczzfAZc48Q9GMrbyNLFee3TQmlfv
7IQjNzlerWr4lsAhH5bolYU5MAy1iDl61/2/Kq0EVTp5xjiWC1fYWFN4R4tHo+q+6hFn/2CRXpg2
tSIB3+MjPUSNbhL0PBMfdpJLgcoC7rFz4MM6JOttQytGvyyKz8nFYMYp+qpseWF6QMj3vekLe68z
RHpvtFgSmh/QxOsJz7pnC3OXSly9EPvdM727KNK8hJVdaHTv25Ma3MJ8u26PILKrtoGoI8IM6H4s
tEq7YUjLODr4h4BO3zWOF3vd8srDb+Dnav/OTMZ6jQ+cDCDLa/gPbktDKuj7Af36NObHeVTsnkKw
YjXcnC0Yd7s2Se+T83jVrtvWreXqKF0QRPLenS3jmoC0b/R8Nkl4XP+Cni6uKN+1F6w/Nhb8aYDz
R8BDn0xiFLnkLV15wth8BST2ZMmJz9DYWh/E0TUEvV6DUB+6HbBnUloQMWr5SieTRyXzP33t6V9f
ZIp9QwLNZKa+97WtyqGqEs0+rYFe0+E/KM/0TS7xa1sez8wfZv4u/V+MJ8L3YvNiH3bKB2BU6IOS
oac67ED0Of+VAk3o6a+UX5ch5h3OcMaRRC7kOQqe86Z9nprkCm5LU7ObdS7egTQn364H3bBGTOBk
XpgPCZU38E3qMG024rjHWlKO1VLUBHRDy/qB0dlwY9qUmvSgCXGP8+wHAwMOvl7q33DvVmBT7F/G
fP/kpfkqKS4NpKFdbNg4rZE6TLspjvly1aINMtU0LbzTU+nE6rbBofHmTV95nNy5/92arBG7Anzm
UafxIPbmDua/p5AmYtoTdSqIqKpV8v089XZUFcJAcihHN2TNETQoHnoJytWhdnMlKaPfdvCtnVXa
7WBj31ZBMuP2r9SmZ4++Pr483jWJzAYvUl0nghe5FB0NUGm+P5dvVQoHUnswg63YuGdGpN8HvhH7
bbzgDYtHnP1qYmgfGCHxMgYZ9GNgktnIoRk1MX1SGho47Bofok65B5U7UMmXCsIZ8eDvo9Q9iX4Q
NmufAgp1DvqsNvyvBYQ+d+S4EEykL8DzsfO/PQIzKX0tDvPIrln9BxiFkvqyOR8pNzvvILEVlsA+
vpruUAAR3HpA5OqC4L/YtnP2FSlA26aRmPrFjLjqEPb/udsk6qbblg7YhQDv20wK9Ep5hQynKxZG
Hs+zxhg1Z5RNa9CnnY4fwDn144RZLL/yK+3HwO37tm+y9H1Ae03Bz/JVVN0XYfm6tPReRYrO0rGj
U4R1hsJWPhdVt9hsVjVeF4n9BmtmS7heO4QiH8cpUnMQUtyoWkn/xzqNt2nMvjKbBLKFJ6AIfmmM
dMtCuO+NikCpIZkV04jragsABoNt9sL1jH8Y59Z97bCGbHGCrZUM7lDcqFGG8271BbtQDgfwbS89
tU8TZ2zH2p4c9l1N+M18mB7vrHkCqOHlDwXfdJsTPKZefRDQJb2X40WDCEdjXMK/0Qne0s9ygUHG
OxAHkQGOsb3C6RieXoiHaMEMb3z4rA4y9I1G9p7FPtzkf2pemlGqb9Sf5GjWNR742g2u05Fh3H8p
4pP8aXdtK6aHE5ICpLbowesWgD98tYDvzT/0gfg1hOnYzWfhpdWmznAZAYzaKiWvCWPy5e8urrQp
vd6VWtxVnhWeeDm8bDBi5wyFUcGhV43yRB385QXq1LKQCNR0Q7rcabv61DjZbHm1KpPTqjQdYWdI
ffOcyhEmk0y0Wx8zfjR/Enr9hVlww+B6ztzkU7AzGwB5dPTpDk6vSf388jWT40/PSrraIYyLO6za
G8Y2NMozDQRapHSpBf/vg+ASf8XbY8PpsGA1K+7sK9S/TmUvVMD//RIMGo58pnZO4EqHJAer3c+T
vih3inf53VYC1GnzwaV5xnbdfrre1KLcNbO/uRS79x1tlYf9mCr0CJR0M6vUjOLZKPzaXLIAhiKT
+WgfaeK0EtULdlMDczGlT84Cd1kmgvxLeGUslLZ3mmypFWcRc7Geh+2UpAMHtpVL7xikJGqxsxBk
mAZn3jxR4/n6DAQc/Qh0FUZnDaAczHW69ae3GHN6XXdP4TJm4aUpAAuNy5GvJThla+nxvpsbbg8t
8zvb7IFZBRQcduDWtlO05ltFWaMf26paSwgeNj5YScUMwCf8ulvWu9ADgpqXBiIXeMIev+CxrEN0
N/Hnx9Ga7hWResV+i/OFEm+RfnSKqzkbAZw0nLRAZ9gfyyXcmGzI7XLhOSXbd4PbATGnBnQ0ZfZL
Litfhn/id8IXXEUkEB7MJDAb+meEp6cEiueifkN5JgmPuUIFrLJpIaq7bKzR+RFJsoOJirsk2TpT
4E+h8QQ8Ghkr9pIdLSb7pr/pUnmWnTNukwOTUSdUOIlMmC0Oc8KgKkOzY7sgzEWnHNyVdX6U3JEi
Ghwj/KVK4CTXg+0i5KsZAZ+kT3afDLSwGICFnOSz6xZ5S3pG4dww7oeXLmDP4yOahw4j9GvlTSTq
nzz4CJpGzJcGE14xU95i8HDolWt4ZJitxSQ5nMEWa3KUHwuVkJnupCY8ME8smAwA3IxbijvkfoG2
rMo8I5u58Cin/uom5wvpuf5FJOMkuRkmTBgmZOcZG4fcxjAkernBGI/Hr65MLOkmoExoYAoCD8xq
I9hqSEgcZdYnwGNHVV/eI62ZXV1NsGTduvVs667La31ArmkT8BRo8AatkXOL3Gue66/awHeP8+ub
A2x7Sma8LkeCmkMHkexNzZpuV+JHvzIcomKMqtJdsU0AxeA0x9IccvdHALmMn/r+DiW1rcV8c9KP
A3gCPjDsZ+5p7qVaPrK5u1lyDEw76Raze2vP9Z4FQZH0X/n9f+1L3LVbaqRuJgY+jYAxrzuDrn6I
FwvYrLGg1rE5FMsorIZHafaVPkJkBwtUw3tbiOJspk0UcWHNYvXTL/xJFUkcQgSCe/i7xfCXm4U5
gRYJw/3Snm9Gq3BD/JARmw67Y/m6vpJNy7wlXOwlFTV8v3KnldRYneFdIaiUkYj8/tegBsH6sYda
FYowgK+5dyNJQJbJcUxitliz6CPBkTSt5iv4qD4Uae2X4Yabw5/bTirpucEUO9a5n4zNXbQprbme
AG8332pLpRkc30Sbz5QTF8UNBgzF4a+sj1M1p/rgO5b2zemqjPgqiD0GVmf1MjWaeU/vcKdFJoNs
FPDXdQHuFmlGdaA0/89xAE7NfuvXsW8MvZPifHZ1Q0Cof/R99IQNyUgfi6YtG0DDfOtYZAk89UPH
OMDoqeaTsiHb7gr2DfG3VgON40jNt7KmCqOzOzAWIfViR8Gq/bSDDyjwEfGw5awzGNsO6NX+WfgY
0Cy6QYWW81DHnelZ0czkWcLqic7zHZYfiyuNG2JFKvRT8XWtm1ULM8hyJqWoplM9JD5r8wo3qgbk
p6Idjn5/qEp9KrBRIFRAx3m2B6LE0Z64makkMtEY2rCXCkTZdKBiBG7O60m+uejCz5hLZgZNQ5QD
Xs4EXnq92fcAgxbEO+YBKsrZhUGsXbdf0FlnsUG5ojLVuk3eY5tL2NKf/bySJLDmzZBedWTAc/LY
8Nvogx/9KvcQoH0SB8vJHvMtYpwKSaUuY1jPrPP+TsadeN+8iVCUo/0HmhL/vOfU+xIyyAzGFQAI
QdaPfEzmA9Asixz0i3sZpCtTKuLISLlKyJMvBPZZz2Wgun6Y8x/Trh0MWqI8cZI+OyAkYfh07Tjb
H/dGKp7v/BHtdnx+gA0MWssyJhdQQIIv2NgEj1FkvI+QXKiRTv8rL6ernjQ3AITWWuf+nPAyf/6U
YZs/ZAA4vqXfJ8aVZDnatgrSateQ+iQT6uwU3iH1x+QzOGeWqQSc/SoRvjMTP+HYikJpx3hqS7Sa
Sf35RLzmykSmf8IT36rDY/gaYn/d/bzXBy19oqSW2L6fLC3RpIhYFF1aiZV18GY8mKdDGVewJK5r
BlWp8ePY48jv3CjGWFerI85LzBw5CkKGnxS2PS9bMoBbCWmnTvWIhUH/CIcBuKcCfdb6hJhkWmyZ
K2T/Z1mglCVauP0BOpDr65LDxsoyH3Pg+7VgrFcgX9bIu56EMvR5yubmkUm8HqNex91btGHjdLDL
x2g2fK2d0ObrtAjIZoArSI/XE0cszigq9bJOM9N3luuG7xWtzG+io0kmQ/sWyavQnW+EUInMkczF
kzl8UxYHDmaZufkk4tIYjXT9iUIYBrLNd6L504xIL/vTE7rYiPO5J2j+422iPUnLgzOHD2l0bNzb
jiRp9zWIPaI+HjZ/5Px0uE+N/Rfl4qExSkXFooTCq1yqvZ+LCIef8+3KioT27tyOP/XM+hh9VBKL
JJj9BYMeHGGU1BsEzgNpSK2XS76VNVD5iJWFig6WCACAa95a2XwzqfSbUXz0smCjuBUFsxcAEHUV
+LX8uNguuftCSDC8hgkijCRb8n2SgAsGdUGYiSMJ9bc/kICHUUu/13P2Unr8quhmSKHG0s8Y1pPK
dBQtaIgnxoRGrVqcsnBKo/QF6cRxdNbe8iuPn5IqyuFaXxB8FgvDirxQ8jM7lTUXC+o1P1u9TO2Z
gU9N356RuLXI5+iwrKZxyi+Eq3vLxlfPY1591Zg5XeAnoq2bXy8Nstqqxgm7z0HGtj2xtWoltrTa
qJIoI5p/sX6wKrWLTBb5bmFflcz8eEldNe02RGSu3JCu16ucL2S985vbp+HjR6fNk76YEbvOFXd7
SUVm2JBD9YYSsyfKBO/cI1wt+1XxAk7ocpqSLlU5vcYIrlL9TJFPwJfh4XPZdV5uCox31AAf4gEj
4lUVjymkGpb9mVc/Ah1QzOP7bsBfsLPoBIf/2we1f+/KQRTmxjEQ5DblPjcahzOsW0vELfjsh5cv
7RoLquAk2A5iLPvrW4OUITbZJsLRZpKtCKXTiuwBWvJ6mAWeyTE21ocwLM2ZixhJbZfJxYDFVS38
Qnhvdr8apUDHJidaTV6XJE2ZpwLqgaWGTsXtzUQmljrMffyFXpuPrDkb8QPdTMrIJKAJM5yY3tW9
FpEqnou5jtzI0DP/bsCtDDvSnLLU6gxtEgLh2MPBJ1DkjMzmHXDjKejcpsvxEmlhWbX4Ii3xz2aD
l1D4lB4wrQTU0gAok2iGPpnvoa+fpeUZXK4Tmc6HrR/UgyzF1jwhJggeUYxfcofLHI83wVFAah7v
W32ASvqgDQccf3FCV77/AkyaYQlEFtDrkhzst4CrPgbKOGm0i7RM2uQoCTMBZyX0pFLlhpkQbU+G
xEhFAyby/QX+hYrtsZeRNyADua1eXR2Br7UtI3AI6UqqrDwYIGvFAifjR8WOdglWx9CeSR1WwWzB
KmaXwdmIfPjvCUhk0nNEbi6HyXVSXzSu/VMx9FZEldSqchmTGO8bbJGUe3I3XZ3RhqsmBRRyYQia
QIzC4OmjSKuLtY/SRfAqeZ/F+iQMIwPj26XAGguwWeWhzRV7SFA4nx5am4L/xHLUPUEhO5CeBFQV
ZW/8vK2Q6iW8rESiqw7FzezZ9nko6G9hnKa+E8Gb+JNli2cdInFZj+51gsA2ZLldJT5w5BnpZ6U6
fi1IsG1yZbc8OLCd/YuRJt6utMtKSOrRgQVKTlL5cK5nlSr0t1CHzPO/1avZEdAr/Lcp1WPbWfK+
txvEJ6duVEYbmOVxDoGxm/rB1NeixeSHNbGlcEFz64OSK2kP07trduVRQsQgh4kJvXTokp3LQJO7
Jn/en9y6tYc8P5PnInFX1wgmwbLF8gSSc5nNFZu5sW5KI1331VeknlePiZ44jk2Pt1HFp+DRT6jQ
k0M31I0ja9mi1cEczSFxJzKLHX0F4mTvkXtZuPddMpdCfV0V8KZl2BkOdxMr3jVwp34gDU+E/T1K
CYN8lPp4EQ6jATfDNb3FF+KW3N9etyfeHH3xHkcb223zmfFDauhALeDfel0hKIDxlpdgvyEzG5iV
REKfO/laqicM9OiGupCjkftkwelmg1DrXp0hAd/leu/daqnwq5SyT/V5M6qtH6DrczfyIPHTMEfZ
KmhsumIdVJLDRARPmOCUJAbEqkT7G48v58Jh7oBe2if27MFmc0mICu9VfXH9Y91WHxCSDDcEFOjx
RD1ULuJTtIo9TEP/Mh36mg+A+ISo3zKC98xlmHQLzwyycS1v/jRodNFphx9Hbg7Pk4XXGer5QyDU
oi9jLjcZw957AFYYGf+q6yA45Ih9+lWT5c1E/MhvKYCZot48Rlx/vgXpRl5K8rgvcPsjukbB/GjW
AgkHVORj4vN+Jlsdu7heHjmrX/jvwHyhAT3qGnK7WVI5p+JfXJPd94ldTo99gTpL5WAFpTB15UyU
IH7FcSEniLG8ZgEUYmuFrN6CiRt+w/wpqg8HEFt8t0vUY8HdmFqrnxR2p93DwNcAGbO7pzwqWvLn
LMx7qmafCFdFhk5mUNcEhn2aymUw9FBZlCkJld4vZcIoD6xdr00cXUnMBh0jdf8JMgKEzvaFTnCw
RQEmRXPkfOABF9iW5f+KrI5bRApVWzfV4bZeVeXADCYJmWbRWwFrshDcbDlL9nFkaNX3Q/6c/PvP
ZFC91T+rTDuCEFMvEFImKnJIwSmHWxjPYr3BVvQc8n6ZdeKWfX/Uw0Qskln7JQoXBSmd4dcxQTrs
Gh7eB5bVpDvoIcPb+9NDlS2I90kxmPgVxKfArhkZf90vaCUM50O3K3Ab1Nc0ydKSELP2eHMoJYAp
2ROg6Q7JwzvnPi5pxr7wGw5nCSkCcuQ2tl5ork8ZISlvuQCmX4aNzV6rltf+s8cgWbmoOaHHJQJ+
FURNXTUf0aXAb/NcjnmW2VkpPnM989BVrMG3D66mxub71/bkvNTf/2RvdNEgESiBQ5tzwpwDxJwS
77HiHqjUyZ/t1LlGe83vLXvMjFmA34w37nkrIB4LLYFxmkIut/GJp4TVuhvlQ/xog3SAE/qUTVnF
KCsgkmC4qP4cpMazfWe6uTAnmrTc0nrFiogafHv9NsCX22qDZIiDsdgJxrYav3gZMN8whSe5BseJ
xc5GPiIz6YRJqFXC4yFkC1jXiRWQ7oyoA78uder+2AoP2oV20akNBYn8npFMaRE/yKdBsc54UiSb
bsJv82HWJroP9bWD9mr5VXdr1cjfozOqyVPPaN5dgsl5EZTe96n0VSs04QYI1XIaXP8NobXIG2LW
gBiuOoa6Lp6P3B67406+2rGBkfOhELNbmBH2CE8n9+BGxfiz5fhr+mfTHOz3tKUmBaq5jwJRJjEV
kRDkoZOuoNJCqFIW8ybisIGFfJePLwUQcN/eY8dwu8+lh6qCXCLZz3E7WPIUQk7/fQrNrmhrnRzD
rAg927NOfhOi7GJAep15btNl9/ZKDEI/iULWL3dzLJ/h/50Nvlo10hHA1XmrWNRRZx7/LsxqcwBW
gj7DQNftm9wwmBT0b/ULN++d8R/UividaPdIUfYGwRS896sCSWnku1FWHzHCBD9L/J+UNqOr2J+V
o87muwenBQMDLZ6bBilctbFi+1MGTozKEp44kuf8z3YK4gI8k19aLSI65/iJbOVbQuIkw8wTe1ea
FQdo/S1FYgasTuo3r4YyGG3jxaZcNO0gisVrF8TkQYE2JecObtEnPWb2CVs24++t0oMdI1zp9sUs
+PQ3l1rtzQ20q776gBDK2wmnaqIMNiR7cZsKI7m+4JKZC+2QbLZyzjs7s8M/MNkBAUUhBk1zu1el
FuRTcz4o0MPhrcQGIzBO+8+im6n4K6sRtdD28HMnTdsaIvQc00RxOjgH2mXlNUHD+lSrxL8z8GFZ
52mblA296u1ZRJMFk6lHJzf0IF7bru94/o6sAJdrhByU4H889tO1j8OZYfyi4xxoZnwSQTWMGX2l
QitOM6JfuA6KXIWluePkogi6rjqFh6QwbIr6HBPfZ/PQuhdXRIwTxmHupLUmYAE6EStM+DSdcmqT
mc3930rBgdi1ueYTo02HUufOJ2bUUJdzf30vnU3VaDSJNkgy/gjlRD0axT5phukcVd3HTV8YpzEV
VoaKvLSWU6MbucD+KUjZ7EJvVznr4f/K2FtW3DtrE+RfT/vq6NLfIe4bQ/fG0uYuEWUWZGERKYZl
t+f0P25HAy6BuCpJKaWY5PPKN+ekupym52ca1jcBCGKMpO1oOk+KRwCYWfP0vk7RSw7qJ/0cou7A
QdWvOu9O5Ue4iXjcTp3+Zf6xNe45ZrNFxIVPtopJT8R8CSde0BmazwJz8fvoUaPb37NdDo/T+iIC
9Sk51JhXJp6aJQJWcwK0afp4BM00gjxdJ324sLkbmSjh/1KgFEzQgrYAgzMwvwegyGnapznglSCx
t4pHXoSGtrplrXUl5cimMWHnbhPQTfzoWt/yxHw1j5zYBvMg2twgXhNUFmurCMmnZQwDDaTfgzOe
Fgx0mvigKarMSWukF156dOWpq5ts5vIUW3vFUKlGCZS575fVbrCe10oUhTQMIYb1hRTgvF4as4Ma
T3tWpphyT0FXGc3DDJsaGaxjxdz5SzsWfojp5Xa7NLVXrjV8b9wFX45lHx8GjyRPO/6tgnSLlK4S
XId4D9WqvVaSiL3ShnTULNYpFhTxws7R+DXUDhNtCqzk3IRoGNXH5MHVyZDkoZ45z5+lol0u1FAE
iHLezDuYJ3gOyXr4uJHXFt9z6veaNVs0dCuwL5eQg7K39lQAwSm1xj1vhLWqQ+dSUb7oIxoxTFoG
NvFr5QUHKbUxdf99HB3YCtECckFX7yPTlNKvOTfpuOn2ZvbXiCdoX9WCwh7Co8axyjU2jDjWpi3/
ZzmKdB4+46mB0ciBRLEzwdlNXgWQle2SN5gacPH6mMTaiIbvtaCkI+oS/D2OFhO6UDliEPCtqUe5
xWGZICLZiiFzc7fytPkvn3krzlaGAR/IzARvUHBoDRbO9zfsvXa5tgNfreA82ljuE6AclxMOotPV
cUG1vDl+ITG8GWbWeB5XBXstWih7uIUTaARZ2+cwn7eq+7ybBYMcnKMQwvj/FboSg93pq83IScUr
+0Ln3bUD/T249FG3p5alWTjkdAzlCG8GzumubC/yR1/I6DQ4Al/8dmyGq6NE5BgA2vvEnf1jIbXa
bVSjemZ5vOBX4wXOZX/iErPz/rkwvX2PM3fn+p3M53FATG5WxESwg477Gh/yrHLS8iyWhEnXx5Tx
+3mHzWmB4jJkq5pZ6iQbvGVcu79L4FFFcdhf33XIXU0IH/QMvXEEN3LdTdnL5SqAof1jCttnQd/3
GBN7wgUlDODHI90Pkj5W0/PCopVnZK3t9dA0XCFs6YrJau1Os9hupUg1jYhA5AuFBnVpfhNdD2pt
au+pqP5MzcM/v0tQnYIgvqejCzzfePzDVR7fjqG6gANhjJvYtq49BDXygjDmpzkctfZtwOcBP2cB
ZyiTWTat3kAV8YQWw9KX8nboGaxydSmfX8O2so/z8DJqi06Pvru8kimW2TuRBXxEp+glDRF0Ezfc
vDdAEuJQE5dtp9CS5WCe8QRS7/0F5G1hbL+FVLm205YRPfTeQxyHaSrHIdMeLSyP7bQ5fHtHldC4
Z4gwVLmShpbmosjQQHbiT9AyHmtESA+WI0oupFKBykBDXM5dh9nsp1Lnj3mBz8G2p2KXCiIwhjqC
erQX2Q/u1VjsQttfJsUkjAymw1pDYt5fO3Sd72d+S4CIvdBZm5kabm0OYlwcPBMWeUJ+Dqf5D9ZY
gEtqrxgWYtBoA3F2gDQXEDOwh0waHaS29hDXH0HA7mEW7C/2hlPkzNuWZiTk+bf+BGkwJklUeqXh
gGnc6lFP+lTgZzH8fwhgskCa9E2wrYV+p9z/0GMyofixrM0DvbV6Yi6F6pmdyqsG2R6i43VSUq0V
zz15v8l4pFSD+lHz/ocSvL5XvnVXVc8vOnvMn6CjjUW42DccO3vN6Ul9iViGMrS1S4PI3ZFOdrs/
kDePr33Sop91kSm4NSby1Z0QowVlFHXo+Z2/hxSrKi3bigGZAzIS6DpdC0FBYmSk2Zc8lP0l/mIF
btEDAulRDxexONvFq6aJeODTVrJj3rarfVTl5fMp2poAceArF3yV6oGAM+DJUp8P7pUceBBCJLYJ
0F0x3LiXRs1u1ljWeDzFy/YgLqVurrHzpFIdHmwaZr0KvrQgRrxyf2ZdqAFCqK0gQATOFTRjWNrL
yV1m3DiiuzV0tzJHI+99eNqkpsAjjobtiiViFhJPK0rjTzxQrxct78DFP+INlURGTQNKB0VM9nd2
AYtAiWRX7WSSYeQeEiI2JIjDdu1hSvcM+GoT8L9SoEiA66DS/HIc9uWNY1lESuKZxb7YY/TNUOSG
QS6T34+M+iTiivUUmGhPF/5OAIo9KI3OoA/pMdNycdZf8fXKIL0to0BYjlLyktcQ2Naj4TJZuA4l
sbzJHDxDAUkRxHAq1curh6sKKQTBGsHC+ECej9jlpqmaGWM0oOJyP6Cd6TQ6OxTL8kWMy76c2b2y
xNQpD/tfL1R+EIbdE4xoLKoYHw7gTnUGv9gSgoS8U6zZyVxFuXw/k/XfTImIKVzCkgCp5h/NJ/49
cfHenMmfkkOcYgwGDVu0LGXcZIbxLXPLF1ZHcy+bXSMqxvGgrml2fRUUm2t5+fElOrQ4fY+rc7wN
TX+Hu2tj2olbpzIyQ3z+HvtEhOvGs+AkOqEutXBuJ6/K0lr+iUICXyL2k5FnO5OYcSwlDaCppnPY
TKCp3CBkja02jhmRatdUZPshIm2SzxxGKPM0U4eNcWALfSLRx37a0Xd3fhRAFcwe0kRJa/9mn2AJ
3XwjrqmvWpP7egQuVGPSZZjYuMbI5fvo8AzbkGW1I8FMJzb0JeJ3YFRrTmkcIlH2Te6yHXQ447ca
Gb7Z3uBgAzw8+OeVYizF3czv1RsrhILMmp8UenLTfKBlUqg2bThLf83UDT+/RYzWdIJSfJsdTQCE
j9xcZfuP/4N1IQGHfl5lSheUsqsZg2LBemydK1O0kmfSlJ/iS4wzKXP8HpCOB8s2umY4YSfpORj2
+kYHcfbLnSedAWQ/8kT/Vt3LwtbwXu3UF6qGCrlk/aBr01SEIjVaulzNqBlg7kaiaSIBISzA+RxI
MKaQbw4GvHcEHGyMUWykmV0sye/SwjNHLoTOAWBGAJDDNSdZ4ChYly41trKAstX36j5M4jvsqZLJ
9yCNqqPhA1R9R6Kd9WuCe+AaYw0vNXmaxcHogqWbsLi5PfyMEeETl8nr/v6HMRzLfmaXu5o58YVc
H944VbsIDN8yilG4z12W4dOetGT/8q3ON5/SUbAnpFggviqEBwrm2iKGnzHar5M1unDR4UxufSvk
wh0aFacQ3Y+84+QEdpa5BY0QVUKgKFD4BBKpNrrjg5+6MOU5j9lYIiSeX7Xg2uIkStJU+L8BAV2c
Y4yncs8oNeD65f2F2236cw2JvKHP75i+P5UYal7l2Gwrie4bd9hPZ5xtiJRa6PiJKv784IZwM9SZ
iPevCbF7lnpm4ERpDk695tQP6H3AS4rv3A4gWjaQIM1WY6cK75uluSeG5mTY+oaSJcv/ijhmLKCS
q/HxANEBeYYNZoD0vuUl8IjRWxy+3zq1ONcHiwdNiS3s3bumyhO6GBVXkg3y9FMnF8BPY/j8wfnb
Yz8JRAxSIU4Ui7/Q5QL3CRlaO6Hfohrr1OLLSbsVp/zNPc9V0joButS5a8s+6XhsFuyBZTsdlug4
vVJkZK4znOHTr/wMIuW9k4IdSjHBh2qBLr8qFHSu22rdwwdn6UY9uDooJgmgLXNhyXAOzQQ7XhxB
bLBuZuVt230QvHTzV3Mq3uDmE9APXsmOKB7j+p94C63iHmgF0gyo45YU9XO3OfmOGDX6qIo8fskm
9u8heZsLBWq6oVhyA7SHvSijg5/8UmbdvIITn8aY6Kjbf6Hli102aCJEcAlcpn4qjolYpqp0GGpg
KM8QSHuGhNcfCbPfQ9euaM9La4z8IoQUdXYr7n+s8vC1BR2nrWQYpYxN1OugAPU6H0EtuAHqziAO
vNLT+xFL9B+P/S3MB/dxYR/l+AV316nGRbstxlTczlNdxeEKNE8QWEPOwiqnze6HCfG94Pf8LgZh
RfFCS8dE2Mfwo6I3nt2k+PGFyk2J0x4n5txK7sJ+Is8unYyEoVEDWs5k4zfgFdvHKktZVay4VMac
kW7D54R4qGJJBhcmp8QiuIkYRoODhWgN3q6z58rVBxlkejU2E/5UK6VX7vN3mGAmxdcE5AcxjraE
eX+Uy0lC2ax5kleSilRXMezHJu1u/8FV3focDZdpPsKS7LqhVyqu8xxaGbgstc1ZGZDNnBAfl16B
lGUTRtsk3PY7VoGFyz5SXKbCPySmDJJITrg84WdNRyh73L3AWg1TY7BT+T9Gpaeq+vGTUtt/FxYs
ysNWP0KwcQF8jxpQaSf0vvHTC/ntwNJVZ4fGDcP1xjM0EfWNMJxFfH93IM9FFPTteoTGCNJejjlB
RJ3LjCIOckEzPya6kmaLaLYQNaVvtnFhhg4dsk4yUR1RyqyCbnrfSuwSqtVQTE2BmOgjVsLqNqrx
U8ZG0LdMriBw6uZLgZnoq0RsFzqawU/QmGFhxx1sJK2wrulnffVJ+rj+nntRS4TCyjZfAIBx2b+o
sydc6XIbslWjnA7I1Dt7EvBOH+gvm6ZNkZXxfWHg3L/BXdHeVN/BIL5R+slDpuJSUAUkc+Pqp+ub
OAMjmdzfCUw64VM4FzHHh8D0/FP3v545k6hO+ElpRnGhTblWhc1VGEYBjrnQIMp3oFJ/3juAmmKh
waU6dfge/7DqdLY+TbCHoQ5S8e6NRkXrIDfGtyTjP08FK0+9rgNgNjpf2IKX8HEKvbx9p3zODwgF
UmkV4eQrwNtGWio/JsxlYNLco9iZ6MJColAR+JYygIesG6McdoNCsN56kSdbPQa/fBIXKelq/Oi9
M9IwRSatTzgSEfiEYu4ZRtzca/NR341OL3q4yEGWHdLFsPlqnxNXgLsGRfhhrn5IYKy+sMEcMUqo
JYHOhAcsaL1u0gYJUzzBoojdCOt17pganbMplDFECQqFvPOVW+g8E9ijDhY56Gns4ATQ/kshrnnz
/kuQMWDp1rIRonbaQ7BYWCB6wtGCeKpB3n9o1wlbk8V1wNoZ6xcuQFIb+IyMd3ENODKF34XGZ8Ej
D8pjxwRIy7Sm4hbfBNNRKSX9VpNgeHDwaqIjHdTJL3Fhp+n6BaR5yKV6faqcHczdY8VKI6C/Xx4K
IGOTWMxCx2GcftZ2s3l0169h+s3QUfHLhFRxYYJ+bQJIsrdKbbY43aFGvZa97QXL1EiwDDGWg3Ic
Wza74vQ7Y6LFRzKNBoR2amqdYB+3gt9yWP4pAW7bPLthyX/FRLJgnXXr6gH3VMa1ODj3rnvUS58b
g1J64I/b+Jn2FKBYxkE8KP3yuhQF+vmEH26lyEiQ2egF7Z4lUJ3ORdT8n2CDENer1uYmlWLJ9ynU
Ng5TIBZkbgc3DAiWfFxpRsybHuwZesTBn9Ajf0/EMNL6iZEnEDws8gSfskWMSAqp0Q0VDMRn3YKE
z06eT9v2jlGRW8iBbeHjB/Zxd8Zx6QVcKw7zC9oe99+XRAdYM9ZYisrtNvWTtzppq/pzvK3XDNBU
Ke5VhvKPSVZzizAoXghGAkDE7wrHpMALMffNnDQg9MH5i98EAgrEtqa9TinXtcFKP7z/XTkQ6b4E
MkK149RTLHMEbtyPV8stXS/1i3MapD1fmWIReCiVQy1z8V1kytclpCMVO0xGsUr/9/4Oy1/kyoA5
W9EXYM8wxlyrkHjY7vwIylRoPTYUH+jMLYADt0dL4TOl6YmEa7aCZJcatvTRhTqSax5X4qmJg/Zk
uIZ8jUpEU4ZSCa8PaPAWu9YN8zpa9+qZr1tk3BS9m9n7mlv8EkOse93NsJCWWYcN5Wfm0I3LXRJT
HL1eR65vRi28jEAuM20Yx09X1jPW1eJIucTbhTXudmjHrV8HJAhMqH+zKwJP7y64+Px25AriKpeA
yMjOBYwTbHtUJIs7B2CsicG0tj8b3faGfnuSfe3MOtVh581i9qpIw4C/N8eG9K21ro43rLdSNYGy
1E3/ijO3JxUOHL0Km7aMMKMm08GSAUbomWav99yCCHGHos8AWurHCd02SdXVe8bc2LFxWCAamcDg
yi9gGwOpLT9Sa1/McEMo7d08atAJe2SYky7ZABbmqRSzqw36gQLLoAEdo5wbFt8Mhb1/tuzybQdR
kIzUMDt61gmsrd9RF62M3dOHG2ICxuFgmZ3mqVn/MH4whKpWB0WvTwJ0jchhYGt1g6mA2LQPqWcU
VV0RAFKpWNSwUvj+uPC4IDu9kSkZT/QVKKr+bhUU9NZC+1foUyMtT6h5nXOtGsomst0beo1MkP2g
Wy7sGru3qN4im7w9pw63Q4MREb5TvveZmF5lPucmRiuHlaPkUI+J+xf5rSWkhkhu+uNf+MEmJ2N7
sJrf5Idj55fjWK8hegqeZe5ezP2SiQQUV4oeqqbHXkW6hidmvFZoLLBvrgx3fOB6l93VRmTagOkF
T3fMlv7iqSMkashz+Sjd1iM5Az1Ged0iadAz//F699RpN6NnbujhO631O7SeXLvtFRbjd6tCnKz+
JBi8sM12d5uUJP7YYv0mqy/ECF3ZXrMZwp+Vccno+WRRqBc36QfIqUPN6JMi43y+eFomCu6xgNX5
lkdmKmJ0j4sSq7GpaZKFHH6O60C0bJVDsX2NviR+y8PvWUuDaMyJW4OsMcOltqb5Y+0obp5p4bUU
0z7uSuvTo5YA+tI7oIdzjaRn8l9yzqL5xxSa0yrdB4ni9WlkgRBbcyHNTj6Kg2lwLgH5UpLhBs5d
vWN0wbZZxAF3IkBKBTFV330ZBIXv6K7C1D70cMrWfw2ti8sA9ZAISHceP3NIGiQX5aavybHrKy5R
KPnsQLn8yWOy8hVsNponDa7854lpeIHD4o/hdkdCW4+twfECVG4gUCr4MslRnUmcZzpYiVUknAjG
tunSm8PfmxmNzAaJMZ3Lhw9XHo3AdUgjQ2wGcmTPBlWB46Mz3b+QeRdWwEJM2gbaIxO/DHcOC/IL
KSP8cjiHTRP34wInO03qcv2D8HaVZw+D2A8+0d41Szl7E7JxBhD5C6PO5Wuw+QKn8eEQ7hF4sfu/
r4l0L0OeAG/yyvVBpBT5wUSk3l9LW1XT3UonYiYlALYYvvv0+kJOr5gRlBbISIPVlTbyL4lHs/Lz
bP/8KfPpL8mJzlc8KYCHeVQi1Y5WwDDlnTwYsGEozzjYsqECVTFpj1ZUJsrvHuqVYDRzPcZEbjwF
2gSQxpnezyHIjgyhEfTi3EATGguXPx/zL1sKopNSsEINFTMaNrohl923JLTcVngu13AyikX1BVXf
eKCgZWamMIxoNvYWDhLnqhZHvu65g3s+N+43vME9bEbwrk8+rgxcobIcx6PIaPPTheonDwf7Xjnu
f9sCrq6A+N+vgA2rlWlcOZJeTCgWtUbcRuhs5CsmnAV5KcDEhNHAMQSuAuhXI6ge6rrNMuLy+kyR
wkqynzDcds0gk84DxhOEPhE8h2yPCFb7pEwtlu1ywn/fN3NZ2Cghc2Kd7GXrgnMkq5jDfDE9m+T9
PPHb6Bu0H7CDPxYARtsX3EZkudKLfXnznBo6zmIlaHcAdSt6FUp33aS+2HA/+bQaJfe4p7txC+S3
g1fl6UySozcYlPPCRRPvtAixVexeQT/45KVurTjahSBBqezp8dcETttM3mzw/1VF2y9uBxX16iOW
CCRu2muF/VrFC28C0pLbYPoM08eOagti/GM65XdlPavl3jlsfWBYQKFhEHAkuIiJLHPtzyGQGv5L
8uPpvpaAmqknRdliGXa/KehI5ElLW+IdRdPFvDNSuUijqeDf0zJUgcLB5mjh+61n91RYM6GXPltX
Q5/hmtiRJPh+XGFl/oXmNsrHwF7+ulRuzuDbyCVrVwenmSP9/XUl4/yJZFGtX8L0B2sufqWRudxl
QBw4EphCJLfAq5cUMX1wPmxBC6tK0ehq5g0+AMfDgjkDn8Fz3PGgkaDz6w+og6fs706bOw0QZoZv
r2aTpQN6GFCsgwiHZ0us6c2V008rhPT+9/XSpMXF8l6WfJVt9sTmWko2d5WmVi2uBfPcSOH6J7C5
3VYofXMzLAxHt3lKnBC4kRkzKFHhuhnuycMszQrMdLdZ9O0HL2xpOaODRw/vvhihu26P+MClqv7R
jjzBNEPU/W5K/tfgbkbKI/+Yt2dQ/GhJoiE8dbTtW6X1F9AgYveIzCCzOXcGr5ke32c8RJv8VH6G
3RPgc1W+vw6uMTPC5JNZp0erraVB9I7xcMsGEKQo9BEZ9QXhSkvlFK51zNc3Fp9HhBhjakxSl9Ek
vdJ6f3bdxdF0Wi+Pb5O44D3FWvt4Dn/8eQw1EFzc5Eu5uuDDG7ceh/7E5WaxdBJCU/H0ttj69S7j
PI6fCpTPxy7gIrTErYQkGJhBTnsOcQocZ0vcEcWzdt9Dd4M1rzF1zPSI+RwWs7zJotF7ldY1/e/j
hrqV1kAyivCLk8+exPhPswmTm2E77h1vYTrrBtoToQ3sHBB2OdAe7N4ZfxH7VxtWnlwy+ijLaR9o
eOl+hTCCLMGI8LniO32s/vUITNiBKvCkOz1Fnmxp2slJORcJvbNxjJbCY9mraPvxUUuI9N1vzljd
kqUbP/DCW0rije1tY0iMe3pEUPIbuYYyHZc29xVqCGXs/n0pbD6pvYrQT95oOIAlc5S2v76P7M9z
qqeJKQglkoFTXHfztgcSwnNTiHNPcNHDM0u4GKWFi2tpBFqJ08qAK6orSHzYSRv1lkpkpGY9rNTy
pCnDJ95sViWOsZiR7i68M4/oEJZbK0sFr07GbNghfUq1PFa294Vj0PsMbykPstpmcDatkoHXkg3x
FMQMxon3Xpu1zoaDeKgnC6Z8xMXbIXtLKwF8NLoAUdObkZcRb/L3ZoHl0hcUq7g2i2dHnx/fENX5
wX2PVfF33LSQF+WE5VAz1a+6gzH2kmo69xYFfXVC/mxfs4FiaCpUsvd1O7mJtMZt2L330eps2G90
xWdA8obZlFrwajnO4qZULpHa5aAk+9X5hvyIXo9MpJT6u7He61QjeYFePDGqNMX7+Y+KVZqEOLaY
0mWPM83uR5WRTF4JnHvHm3BZVEISxPbUKCzcagunSzyH5YmwYBuUoI3bFNA7hRZrHvtCg7Ue8SyN
RZNCej/iMeJexghn+n7+R/Hq6jeVeSeA4Y04OnPy7iV9m3R7WAmuhBdhEgW5vdamFlPljDB2rRmQ
SM8z5NF7GwMuUC/cecDm1lyCgINnTkxmXEtiUCaztZfgtI1WvVfmAsG+mNa+zs+W7031kV/Pbzqj
yXptFetsDlTibzalLBkNzvB1SJxcwq4p5Ur05jm4GApKWi9P2qehkY6jU+ZyNxVRFHFlbPNKf4C+
d72rzvu+LY/zBEuUNeG3EkeCrhkX3ZTsjSZRrrqOdqh26CmaUXXIudhK/sXM/RVnC087D5xicZyh
QhwzzbAOLPT+IqZHl9pDSpWzkUPtbkqvpJrOnh/KwP8b6+B8yXfrR3KKJAy0qKhyZxxiyYjZ4pYO
M1P/8+uElyNWyHMP3oizpjRwFvbD+uFKMpW4HsypzY8zwrFa6IgF5w3dmBKa6sAdzsXlJjg1PFzw
TjeP21AnmgxPLoKiNFCDOqykZDQGclHW/5Z+7L3FeaXRE3aiTLyb0UlRb0MEP/t8g2Q4gvua0Usi
hQFYjrdNcZvNSflC8iIS2YzrgJN5vnzQzmEwKjS3JKtIk/+l5+kUT6N8gfRA6ZJ9ya1tzNM28ZH2
50PbPXSfwzuPSMbG4dB6n/tivNI3vaLhc9zqbWL4Vd7zaSuDf8DJhfYUNjocOn8dhuJqag6SAvQ/
wOBfwX8vuga4f0iXwwLv0hk9pVFqsswtN28p9nvsbIOx7YXptP08jLcQ17Aw6B8zGhyAntUT9sFa
L1iOyJy4tQrnaLzE9Hdxp7jC2ke1it/pCEP5YEEWwNXNDjlgXkRiwvFH6tLgKBj3R3NLoPqSHxou
h0PO4ZNQm7TvFAfggvbpcT5VkwuybRVqyX45xU0/a6MmaBndrjRp58vmnrdUVsu7pA38G+6e3LDc
HB79411aW8Irn356cjdBhgxBXrlICG9mSkOEX7GtqoW19Mf/7X35cx6NTsjNfKagFTw642a3w9Qs
rnPVctmPM1R+3mfBO8c2aHJ/NZLTjgrB0x+U1J7c4R9ufB3gslUl8VYXacMbdeo/N/1DMgh2WiWM
NAhQ47iGU6rc66vqFhDNDN5ePjtpgaRdUnxLwnbeGSvdO3ufaxGr+szdhrForqR6Wm5JlglhGZC+
yo4dHMMtCMLZsEzimy1mzfkySWxmxk+F+GHN0WgxdRMsaofMFfO5KlY4zoRlmox6YwfPW/5nAeSS
s6un1UAzJmrn6eBvQzO2eUiv+GUs2sEPSlPeyfsHrZOMDFwi6CVMMMzccJnpsbz82FbDyO7ajCUa
wigzto3/aUvuRatPTw+iT2JeXwiXgdaiiUIIiI0zrOE6ZqOPGAa3hCTjqwsXSKScdMlMcpjFCW/7
8ll69KNzeYM24VRjTOr1sqLDb0wX+IVaY7mMW3s+Edetckm5r8+sycRge6lDCO/8dJS6k0n108fP
4mGER3ftfVn+upTJrtaAjdfqtN29OJHZX+SpQ+WhUn9pTVvrjppJ3rE60q7N2TFon2yRdNRIkVvG
++BXpXw9o49R6i7yyADvKOywRfMZdryuJVN20jd3Bu1YqT88qghcYkxuaa3e7GxIlea1VjPabP93
muVv9Tr7Q2qjMhDiBtegq+7GR1LtSKNmXZJ8qpcK28HGf+z0aimRc5NdqWjT/PN1nwfbvOgIvOMe
VuXm7urjjFc6BeZbATZZKua6hzX4kpiKqdFOADsEZwHUU4q/dg5ZNFHFbhe/Ph7K9E1/9I2oBojZ
wKIbosKCZ+fG9sIcfS8943rCttXYZbjwG0qQuCFRskGxi+EpWWGDhNHqvlyZiRILTBDS2XLej3mQ
aVEiCBgLXo4jqSM8gr7sklQIaQt+PCGOEDi3GTouSDjfoo5mKw/+gBB10EwID9XlgFuAmzoqJIfY
mxLrArvb1J2mLykJS2J8MNfGAuz7tvVTNoNWtjY9hOGB7uMbuRMMUzv9Y9JX2fV4M6t59Nv7uVvI
BMW1u8hFe7UIOWFGhqbWg8SuL7U66pgwcKw0QFAgu9zys2GVSfDReKRcto+JJDYdwwILewkDfiLQ
gZ1VdcW7mH3JlReBy6ihBZ6dgpA4kk55r0t01glWVB3oNjpba3sE7kBNeMBkg0CMhW+vqM6f/Q4D
I2BOHCM6rza+QyOGf2V7ManHlZ21f3NHuzBOSPRTP75X9a69fC7KZaT+13UYi9tNFMxpL+2HDazD
EXG08Z1cmWRkjGK+S/T5aV+b82ITF1QmxOqsSv3WmM3HiNzZleNo6gvMicTyPqQ/ofJkToL6hN0/
2+fUZgBwOchKh5GzkEf+Qy3j6cU8jbI4EJiOtP6vosrdOZ1n4JBG4/s/QBzqj7M3uXrK95258tWp
B3I3H0wLgcYRM3R82kXc8wpMI4hjEXYozxt72GRNlHX3zh0fa5kFqXW03FG6fZ0ngLlhmgvHzwSI
MvdQ/G9aa9ziL5Xqut08ojYGq0plhj3wh0Z60zxD/39zIiYDSsMonsq8b7tTGklVuTqPJG/kaEIL
DH6YEgCR04GyN+GIsCs5l4yif+7e4NklkF9U9nMc2dwUCwy/3aCdeizrqB/DPuOF+Yoznu1Xr8Au
wdTI/dpoFfh4/e2NDvGAujatEP58ECj0tcImtfH4qqLGDihJ7zt4us7mVcaS3Zhbup0DfOqr3CoE
eatT6vDJkBqp7+AideZltruJhD65fetqb7wP1LgnYGjspBVC3/X4At1WFduikj6a6E9VQIDRu+iD
IHmnYwgguTdpN+bOk2qFlsLAOO9CtrLLgJaPDTmeyVZ3LaWU1Vmi1atMybqsLGQEx3/Gjw5GCFPc
uNCxVTIbPvlIho55uVO/x+kbssIzgcDcURPCzmfHorDDgnx/V/b7JASFcRIBcJrbOaG0x8lunDQW
kE4tlgjC5isINgFLQ7ySzbdHMUWUjBOS1NBVZHdwMP79wz+K5w706Nbu9fxuDJpaAI6B1GhlvrYO
5NZ1fE3tVFQPprdrRWAc6RBWXiJ7p2MLlezWCnMfKBXrmpQAluwtoD+UW4MMRge6L1yF3RwXIxiC
3txySUuDgKRpRc+YFRFAjHNhWiF7hMxXmQd0KlK4gxPs8woFPIUjsrER0sP0r6ZSJqG3OObn0o2B
Im6F3J7P9Uor4AA4OT3AR3d8xCH1RRDRjPLermYQnoFrtN6iXH1HtnK7NKeMYPVEaooS2YbM6TdE
UFvNzAwQsF0HD8F9ZdXOVIsxpVbw5aqwvljIz292c+AQ7QhL6iAWn2J2VGwDRdZQEC8FAc9lkcsN
puTIX38OyGYFTMqnn+oNINPHzafuymaz0+dv5FHu44m5uB85XuJhjmK+iiEuddP/agezGOkIv6kn
a5IOCx7wUvpczm54ilpiq3T10Zu5uSJtQnd+vE58K+TxuOmBecEoLgPJYeO1gmh2wIxftL3LFt1x
lNK0vpswq2t9P4M4U9GzysogwIC+oL6n7109uHB0QRiULm2HyXjU+xPEz/TCNgd2WGLWCZ5p2mpz
qIrL0bgOQDdEryjt+maF6xrehKTt9pbb22AjyeEPD6LqFgLesPtGS30hrXDmTzNckkOm7N0WtoxA
zgb4mbbUg0CZtp7E6Zln1iLeZG8J9s81Kjg2JdUu8moi4kF6YQkYvGGNk0oVPLupgV3dn+Afkx55
ORqSiTbx6CXbuwzrV/nOWQTbocnkNzY7ovo9JYvb1eYUMY8RgF60G2seCIKkHRbnT1qxrpuX1X2g
ArMPYt/2k2avh/vm+r1J4p1KggEWAZhiKUw7IzUhClEgWTpC8wmYPleFjN4THYNhCzptG9JClTKV
fr7QKRHAjnxZ6ihLqD/2I2wKM8PzGIP5VgdNrCWvv4R3Z29uLE3xaTyYUl4ui+Zbgx2GuoFTFh3h
N9U0Z+Awp5q7b3EV8Hw1E+NxeEtFmFi+z5mHjcwlptqZhJH1iGtpXrsoien+IQ1qPuO5KmddMcgy
8DTpfQv+d/hk2bfX2TAZb5KWlyD5I97b96gbB+Bs+jZ5MzUjam2Vpd8G8rplGuM1zeKf7jtaLAYL
wAiKW4ZDqQOo81JVNHlYM+MOJhtRh05T/+RWBxgweCNBqPV3n8BWpTViBOoYYfO7lsYeuttLO/kx
/pVffeNtPaeo0kAWeYCKM6j7SsNAtotdKFMaczTIr1zd21cwiwpN1Pz4mjhD1mKNtlDSiWf+KuQ7
XO+K/w52tHn6kC8o0eggibYhsk3GACyUPgM0FiZ0rCAICImgd+S9gy0Uya6keR71b/s12RYI3n+s
+IwGvYNYfPuDrkMAgrn37966rkkhyGGwzxzl6Hcqy/x97Gf5umEwjnhVMO2a8Zpk0mqOAEKLU4lJ
mmm0cN6lIH57kLBrieELLuNo5rXZQZerRxsrh89ZyReydztwdMpfF0DsxzrDISuh2xixPYtBtCmH
jJprasvy92qGOmmVuE7uG9ED6gaZfoUxGPyFH6nEwJDff9vUYliesgsNUrAsC6npIaIXWLD6DTG5
uZ7gRAvYM1BC48P/R2onqylLa3vjlxPRv5C+PGOxfUX9sUIT+liq+mEwfu6Pgrnlc9Yqb3BsHdsq
gPmPVisccS/1/B+ApXl6I2s/Xw6NVWfAqSQhdP8hWaNQ/T67OvPsBDfhAZpoHm6HtVi1kCqcOc/K
iutWTUiA3vTO3EOg1AZU4rfoAm5DMmPzzHSpaROaJeAofPgLLZstliJN2ohsQQNGbpMTdWnGafaf
SWaB43s0nPOk8evhS5mun6uh+KVenOBy8HUYnMnRtp36Msd/3uwkeTdS44T0XomQuvb/z+h1u6Np
nCwCJKvMm7cyoy2fBDcgb7+r/lVlTk0mj7JE+xZZZs5yh0HF12XJjrLtS+TbeuqrMvfcVex32bzf
1pRb7U3StlOkE6ZliCR6SWERbh+8o1HwqiLNvxKFZyOg/XOGrcv6T9HQw1n0HTewYW5yFQO3fLqc
ihNxHcZcdIvtOuzSFzsD3WFf62+ou1ZTPojSo8b+Jv/YnmCuDXT08YIIbKgM8iet2YiE9OyEtL5w
lBP/gbb6xggsm5ywO9pUQO3m3xxAqpqMojLpvQoq60FpOF3WcwJtswWsv/MVgQNMsHerqJLUp7sr
D/aCK04YP8EHa8FDdZkyJ0b3QbrYXQESXf9gzMAvOKLJlilyIVolMnozcd9xdQDF3XKRYQEdVT7z
PZyHykIi6BaRjW8BbL9ljWUS3qPjYtn11JLj35G3eVzJ3qnPbpoGzTZxAGY20UpInHO/VTBLEGrb
+99usto8VVgAcq3Bdg3AHksxnk2HOz70jRIQq6Tp9ffd/90BbuW3eq5BydALIc5ZLgyMHbDMlmlh
jHgs8vBcF+cEaKgF7DETVCSkwuYiXSE4Hf2vh1PECxKBlDmIX23KPvwrGCP6h+6J4kXzZuL2Kvn4
2kqtfPrAz85/hw65mxPevAt0vLGJ7pj9XtZK5yWjEKBT7IHA5yxqOts7heITAJublmPXqSH07qyK
CJoVcnPBCh+QdCZYXyFnwdNzQDDQET9GF/NWDpqsZQGrN8ajThMhzuyUwxcJsIu1Wde90rb2XBd7
dowLoKQkgNfTRfxKt3+A3O3NtEjClZRE0gOx6oaVLRLRrJbSsMT8zCyTALVTS3ZFnF8NpSudCeAG
uiGrvLm1u57iFE6EZQ14Y8eKLddyuO8Ud1hrDYJBnIYj33QGCfc+q0UpXTXstEZf6VHtRuuIL8cz
GFZeUt8WYdRVJdv1HrTdt3DsnxEROACtV/lsRDlxXeyXPNsasKn8+aArJGjl2L4nBhmvErsvDKgZ
fplyzMFFb8sG+7uxlERMsv9/K2juH4PnU0SPK2iXti9qzlrbMa62mBSYGwMk044IDfn7hgOHQbYz
wMT8o9tay8DSPRrvJL1oTsnrpWr45IzwDzgW+a6cRFjA/RPDi8yM8IICvvpNf7UyJFnNwGzBOilc
05L3opjzp7S2OHj8dwBb+0tCwx/+B1U2wYVjb2Y0OG3mfTrvm9/NS6v21t2/xpcTNc2gsCqBvF/n
cVrmauFuNkNoqcNJvntF8eSsX8CMKXndzt2NUXkcv8M41ukn5nrVgm/M+o1Ditn6CtADQfwqPitP
d5eQk+sb+hD/q/8S4/FC4nqfi3KIsgvfYzCtihDocT/vwMiwUodpQWGyurbULWbRhB5WFq0DQXa2
4cwd69PANIaI8OY1TUWokh66rYcaeAprDAjJ7//OAc7u0vgnf0DAlvOWm2SAFNp1WmZvH+IcTX1W
zYNKZ4/uO1HVlnRL5/Kmc9wp+dhcckUl0wnK71RaCu4OtB9FJbT/UX59LzRBlntW+szHUod84rDR
El0SSFRqpTkIksYIhaieXtYEDCOowmmuB0h/gf4Khd0O89MBNARh4elCbrvFPjczC6ms2oAFTiQe
J3PtiUJBRUFDr1HoHeai3TI8rQWUdjAoJC+iQZ2GLT+bynTNO8Qblv2+w5X0VsedQA41kN4sFuB1
nn9KaIXsXzirkORvw47X8/0qE/po7KzoWQGF2rGKrqddU1sheFDiw06LJuxUvxbdHdcLe1r100Fp
L+WOLUgWhseGzUUVIpDG2L4IvfCu1KiCly9D6k+d5JmF+82cuFuVHyDdt/3mJBq4oziGu2jeKEUw
Ebcm/dqFUr98qlahDNkUh2aK2OSxnOo8lJq7RTsZ5dd2btfItt/5A6q3ni3GcVfAOTwLwmI2u6I/
1+L/kS0nWxRlZaRrE2lBA3Wx8ipEVczUQvg8mrfNWs1E7HmaYaJ4xtfZHCYak5tJ40t9h4F3Hn2M
fIl6Clxe3jZ2Z3GStZlXo+l4ZUs5+y2sh23tlvkhf7GHlqvWRvNK0dqlzIhz0d+PLdz8d6Nin8nl
eU81YXm4nas5q9jsFzwgom5L4m6+bkNwxqyG43BTXVhpvaA6NGtzXQ1++wxJfRywCP4E6RBoXfsK
YER37CEpB2CiV1qkntMf3GFpQogqhmkbEbf3o0Sg6NIzt61fX8F+EORse2nw0YyKpjsrYfn950v3
sco295TZldvLppZtH5ILQ92fniAI0ifdMt6b4DSJtVvnveQI33ko0Ok6GQ5CB24rC9iAYiP1iWi3
AL/0UAOo8rjI9OGIZNfN6mkqQzNLJwShLosQgRBo1lWSxEMKyH8APT3HkdHxRtrWwtm/RqDlIvZS
E+OTI5i5q4hVCGxK2JxHbmlMUHDO6UQIFrUpxT0hpvEBsOEzPeUfoZTRBexdcdxIAMbUqor8C1gn
gp9NoJWk3+5t0VCF2RJweE5CSdG5XxKyLRik5Hn9OZxty1OszRXhy6LsU1mmyuZtzVYKqWtUXwq5
qpOQ00cEXgXMcian7bpOmk2fPoXck9q6vPMjiSyYxUHZRL84QR/6WRNx+KwrMQtZ8UHh4zyDjMOt
nTS5KY0XvU+a28aVDZNisZeXMpyNKNg4ax7iTisvMSn2td49YGK4eS3wdOmuY2EgL4tmHU7yDfqn
XI+8SuJw5xQDuQRgLVArRGb0N0nmeB4xTzwDVpJ9V+irtja/ieHU/0Fh4msvojugQzkCtyUULYBp
Mjuxkj3Z/xiVbMxbNQDGcq0z6Z+tjLorYjrV+AiAjtUVHYoDIC4mxZQqvj8ujQ7WVnCtxrr1djDk
o/T0u+o+BIxmah9Qpnr65VVYcG4giToUIF4kM1MZJl17odlFlmJ0qi9pLKjOAg+Uqd2rsX/Y4vtG
RUXiGjra4GBt0mE0K0AnlAC1VymWzyBb8P4hDj4xfG+P5CZG/C2xJsDHrRZJjiMYO22C+OOMhi0d
igj+YsXbvIunKuLOdyNIEVCH2lDM1LMZXfKsifej41jt5YX7Y2jTGOMy0XelYUL0sVQ605y8fgZ0
lnKpHPtzpNgvK+VhW/zUFu1q+nP/6E5vJ+nnlFV0XgpGd1vLzi2UwKqQV4htlVLzEJRmpN3iFG1A
qIHLoyEMlP5NS5mzeTVrBEsePTjEhJamKnnhu3ZIpwqFKFHmasG5j2xj3hmZo4ND+NqewwFuR5uH
I460LmX8J3y6PN4EAsmIDKRd29kzSakBZ37ZywQmig4cikJEwpaJQv36h9xpRXfMCRB6XZBuYIcW
RV6IiS9NsxB9+QZyMiBr5xbTZWBZ2bzc4BJg/DIO67qFgnfRFyiUAeXNFnSkRMTzW+6KwMjmbVK1
gVxw+HiN5FgsazCzCqqQBIn39Y+yiB4Q53pbm9ZbCmLTkZwxedxsdyHBlwQQbyuSguKaq+FqJZSR
hpeioVa+lt09guDTKjBnrz1Jybkx6cRyBOr2+uruN1OBwU0zagrN0q8EepLlRW7Oj/QveMzdb6FI
mwNd4q+F4VVKQtWgroTfkCBHxCnkJpxEIajhuUtFwnEbCZpCawubYXiROTtecwaOhToUDqILAA/q
KC2YX9ZUqXVPDAniClI902dI6TP7R83Gx6b4x248NsmN5BGx1v73yVLkTI5e462E9YBMAy7tZk3m
JwsYAG7GoNRjE+wMyf+3xG3J5fL8fL9C9I78T7h3fts79hoNu21Upk2UJ+x0VgR8NFkZ8qy75ZOP
rtoByCf2MXIwR3JSBdfBmSBGCDDLsvMJMD1GggcPIawgGi6ldnRvfb3c3dTOsuMYfeS1fDdpIx9S
gueIb2wyOcSBOWwZJrsvPXnRSFcppOr2i59zKlhguBOF2n6bd2MSvEsYOe/c3rDbGox3PleM3JY9
7goZd6P5sAaTNHBBp8OWpXORs7CN5ET3aijtkaNfq61PMq66TyebUvGFCuY/sLrK+ZR5X9xuzoLf
Ws7QfywGRBxD25AtryVcvubI3lWm9n5Uf6t/eVtevbEHUxB9BbaSLq4c6IyG4d21TPFhNgtSKrJX
ZxSeS4FAkB5wlD8ev4m8XszU7QY+FQwAgKjnpGgsehaHeY5HlQNmuA4Pap9qLxAxE00b9hJX9je+
aiOko6wQi006jcMV23PBdsapOq/kthbXoFWkIOjcwjo1eVMJYO1T8LPZ/URoEqu0SRyWFdKx4pka
948Rw41J4a5cwSVreotp7ORLJRzQ+7+sZ0dAmGM2Hb6y0nkBbJo6rLLxhfro2PCMjYB3H2iYrHB3
CaRmX1eshqksCt9eF4+a5DKRYGCo0mvaee8ALLt+ajma6CGxIjGUk7GcvuZgQ2geVQK02o+iVfY3
YFRet1wsKj6CFIAaRlF0quP2CVpNisd0XoZ32Gdty08y8JeuXsYIUAvIbfpRNJqT0OiDz6gZB98w
64LCX1XKFanytO7E6GuL4HGqWS4PpMvfodYFh2JxaWQU3PscpStBsKY9mivS9kr7LbgzLWWi2ZYM
vdr7wujTTZCjGqp+camIT0Cj77xtWYlsE4ERwB7PFK6+XBMQVUnJCMc6YnBV3mBYKCXwonKl74fz
1PzSzWcwBcVDq7OptndQLEjgGrXhdBH87TKM9HnRZPF1L/jMQ55Hk6T/0wxV1MqgZtkz7gKbPUZD
E09ZlssPYeVHyX8ZJx7JVXSHDnO3PNXkNslSSH19XP3wWyySYmUX2LgYvKePMHNG9tIgks9E4DNR
8g1yxJolPgT+2LR+S3d1AIH6D6oDfHsaybCxwhO+iudoyR52IiLQ5ufjs9qVS3HytVnGHiYFQy1Z
IT/a/cFkPd8VBB+jKEeYEAEs3nR3fIaZAxqoOFtI+cI0NPocruUFhobHA3MJsgPexJQO8u4ECe0g
3ZXJ6WXAfGUJcUZVpFGaJenj4jbSy4ycYO+FKoQzgY5G7bm8GLTSNRdWgMqtfxhumEX1etlmcPpz
+wKAbtlg3WenM+KnWpub9fk+tVu7PUZ260rhBrbCmZODRRTqvlZymDLJpf4asst5/aU5juLCtenY
GX9HScFlOxDRWX+iBTP73pQK2pTbTqWiC/aTDFhK6VTwHhLJ5yVo4P2rEOEbsZwLGYRCWLn1VcUx
+c029uW11lPo8V0SuKAhx/I2YcIZHB8YONOmmf5hRTJD6lgmW4I8Du+TThv4xCaPlcuB3vw3B1Ea
RxK+AvEj46aYQREw2Ag8ueP/sAuMxJTOnsD9gJYhz8e6OHFEpiDEn2umIYl6tZ5eQ6/crLISRTNl
xWNOP1eHD5ENReEK7Q3xFFQYA3k+wVUwqbSN1DBDE1CJqcVoiHl2RzruZH939LmoypIldokpGtcA
q5pXE9diinpq886tvLlBqbPVjCsusc4D/gkYxZsHtXbCUe9JwuigZvjCOvWn0B9u5/mZdtvsW1ZH
psizaX6hmX1cSJP6umUXbyhJa92x2BlwZsb8UtwrFPD9ku+QmWou310Jj5AYfCDJiHUGaci/Kcav
wKueWyhBvo4ut5HrA0fFHyxK73hvX2aYvTGsguKyj6TdaAf8wZiwKkm1KtmNVxn/xv2yxeu6eLDD
MxXo5e7x1jFA76/uKXaEm08d41xqOtVWbfljs6YoWN5GjQW204BczBB/el03FwUORLjomrKYt3pf
6dwV0OgRPiDtnLf1uockHEfn10X4hBFIZ8r0L9M6fAEG6eEuO7HZ1LznbBMYC775w6dcJ6iRnbVE
BWQCI2vCi+sy7CeoY2ga4Kcd9lUA/8VkX2l5ExL2QEKGkMI6Zms8JtOqzGzYXenRNbt62Nli7ONF
BJTo7gsovymGLgyCH1rMiSqtJwDZX3tqmwtnn+glqsbrF/XoAOHjPdu3eDDdkrAVIQd+A1DqXD37
wmjF/MAPD4DlWoLy7Cn3lwfCOJ/75WD+9cRqRsyJJv6zNpPTjUfnW5NWgvBOuyWwI9fp5RNLXwY7
bv4mbIWpUSOzP8PfwBGSJK22PVwFhFxsomsrtloC0T8KP8IXRPA752e8hNGYOLVGPy/GjE3uyPzM
YrJo75nNiBe9DoMiohK37fii09PTdfT75by3vT2GzXzr3TGttz+4K9kHMlAYtHlotmmL0PNHKbYV
wkw0PyxUEB8I0VGwp7HvGGks/5lSl67j/7TI7e3uxPqosN2y87TKY9uPK20JkN34NrJuMyd1b1Qp
8M5JNxIK/SDJ/7iZQ5U2LdEWAM2X48D+xugkEzdZF9Qfr1R2DKt8Zb/NHbX8MRrnLpGENwifURgH
gihaKLWzG75q+hA+gKj1LsPhywI2N3xr6kUiXsQ5Ceggvdh39PMRQek3gJ4WXO5h1E8exyiEgLu0
RW3rzsoyWKqYTqx3fw7zKoHQEkxxPXAagAnvADMMomKZqPC3HrkMpZzY6JamaonNYzLLXev/C1HE
rNGNZ6XFCcb9v0EAsYkyHyv8rnmWTKysAr19YGIkSMUQfBT8o9hhawRawZ9AJYZrM9knAFaSlisD
yoM0CNrZp4WjkEtbr2k7JHIHgNoQVraqTWiatNXiIJOND2+8SBe0mjiYM77rtIKQMSUa9cJbPWao
1kB3EMxaLmEtSb8E9TYZOJ9349wxGn5XC8br/rziYwOrHU7gAltKloQgv2rcSJVxHtA91y6xhIc9
gf2Fpy66vobkVK/xP1BebooY78xMvCr+aQFdqPRAq9K+SwT8OOrhhyHN6Rtu7oiGNvcXMz4qlI6h
cJ4rJFq1QgwECF/JqUhZUccW3OTnPg82cLSSYhj5YOL0ewHKqQKRWCsZhqmISaSzoVUPw4AT78nc
l0GJhkcHm3ad69GbPszuNBjgCRpFtjfNHMV9/wQA4lcb9yHDrkBS4WeNuCgni8yPpQOwiNiMRS6j
rihqzVhKKlTJBjeeHi7dfvu6OBzyFsJDJxRarc5MOxYR+ABVbDGpDKOqP8QzwGMTUejBw6KFDbDb
q5lQdx78+iq5oCGC+ny6sYKcEd+aIHKzlOBhOhyrdn5ktF7ChH0PQS7Vdqvlpwz/f72ufKoRnS+G
aiSsufdll4/lhEDnrXxP6tv9pUJn7CSc1C3+tU0c+++hPZr7+fCgnzTRFvmxe6ce9J8UOLFvE6TO
OPMOG2r8KG3e/X0XBW3eagWWEKpFhTnKuDRZVO/qLEVipu32gsUmcEdCssLUST83hqNLIi6s4Y67
b63BW5KwZIIVFthjM8WiWq/P01IbQu5PcFfR8GLEF6eOxoqdATtU8D4unugkpEVvJCQgpXa2QdQf
u/jtDFn+SR/C83PWVKzAYPAWx4R4f4g4Y90RwGgprC2Kk0j9dOLspqnwZKIW8d32frrYq1qr/o/h
iKVzUxKk3z84XwRLzIT+jG67WxKbPZYEI2M3ScLQvM1an0+iCXw/pA4CMXrKWXV7B4ETIsRdmUc6
eSN5GlYKBscCF7C8w4m+rFDtC66D4DNROHDSXVzOZROpUztYHR+/9SGUmlnqlbQkxJVnFmBg4ryn
bA7tmKvQV3htWyMbVKSLErkDmoPNU/g0uQqGnMYeLU875Yjpr9KKZmUktFUS35hcHyTX+y0E1zOF
jFxYa0zdWCi/ImOlTQX2yAAXwyDlEw6JtVfVIPXSm3ENM74LV0D1otLL2BPS7Ezv7lMWcwFKcquS
zrPegc29FBZr7sAro4n15CN4dCDctf7g5HeQ3Klelgq4Rzjl/5rFbdwytOvYiguItqjzW/xntNYf
zKes9/EnYJiqNjpPjPO6V0Q+yJ87blLDPN17PFMDd9KSf0dGAshuhUedvwbHUbWSgWmpvNQVqqJZ
zu1fTAyN6xC4n5FJtv1N+TJnrrdjZeY1Ij0rJLUW5xqFsUohWEuOQ6jyZXUyvHpih7hR10sCOJV1
TBzyf5/WlP/rUrNtjaHw7cS3/XJ/dThaD6tw+8pczzWXkUaVNhyc1FhpSXbVp38WUFn1XeMB+yfU
CiAuGNzFfOAHjJwI6Rsa76izuzXf8Mmsy+WkRv99v/70dkFkxQZtjAx9M9AwBQU9kpj2AOgxN8Hw
cSEJEh46izLOlJ4Z9Cy5C/AMhuij3E0hOXhrf4Q2E+c2SVEbRJ5FIX4OhokPB9kxOoEM1XX6pYOv
ieBRizCAG8afkh1vkCBb2j0E7yMxFYJvTWhRHaujlioorc4ygQfiyM8/isBtZDXZM8l/SDOsLH4P
ghlyM9QlFbE2Qc25efYyfTqlGzEkdAulZS8WuVtaf8YccQwzTMoNMs8/ZOSTl74Qiz7hUOZUA+Id
RSy4nRqGIfBdam8+zo35FEX+b8oSRIL5g+dozoZefIMTEHpC87PtdOvtEnmvCIso+IWI3b9tJhQK
cG4aho9Bkd6Ow9NJ64l7EV9A0HHB9IRWoGdm22H7ajMUgbG3BNLf59tSwmeiEI4pCSjQo/KSWtqU
Bu8/Dzr/Td4g425YXdLz2C3CFaDUVWgn/qWT9CuNSj2KVH9QWLOEzp0EdYKxwww6tOu/GtXjXeqU
AeA3J7WULlVq0uvZBQ6GWTDDhJKyqwfrgtTcDdPfeaA0cFtjJZDM+veYy46t7fDXzBYjAGsYHZoN
p6CQqqc0IVh25OIWl0g+Gi4iAAiY2v6mdyHjUD0LYFmpdVuoAbWGzDQ+wsss5kHX4XyI6EzOidGR
4Y6/o0GwmPvdpGkXm5Zx5IWpo7WF+1Mvi/jFR3SMQN2HG6HhEKXx+e+tz50zXA5Kgrvj4h6Kw+5v
Enx/Dgu7brWx358y+BzqsndJ0hmA1ekSjhgbyyuBs+f8xNL3Oz4tHOwPRuGKq2dSAORZ+wrEpN32
MzIjRywa8PxDqA5gc13/azxIcdcIclQxKryHbyZxVdF5VeMC/7q7B+upYulSSlvDcqUKbfeP3qa4
fTklPjYDtKbbZM+YeE19IinO3yqxoPCgdDFbJk8toTHTceeaXEVSgu9PuBzCGQFO+R5f6zvsD8Mh
zRjBf1sDlqJ4IpHYXzoK7eQbY64M13xgI1vY1WJ9gxewIqJjsoUMgXJ92/b/TdYEN6G9NXPSYi+/
/NqjbITZSXEhBE9DnsY8EpgH0hwOhQZGqoCmbKJ8CWkeewtmQLvhWTdKwfQnfbX0YQ283MwHR/+Z
rQ4vtVJ8nZqC8G2q0DSXq6nnNqbHRuCKHXXpmXer08BMzDxWlInGT8IJlpwRzPI/gSzULlifQyO2
RXYrabhLa5EWjlUDcQnQeVhxbWZRja/1G9+PYGO8nIF6SqCSx2WfsFqe/XZiumbq8Ub0Z0k2iXWQ
F1IEMlc0bZmt6kgq4eovZzujVbWwp+KXbdHP71Qg0bPH9Qu946PmFmdTYPTc2S5yzkDggguGt48l
4idojA9WQx5Qm+AyzWKKsYEwQNNNDlNnCQ7lTZqRv+stglKtYsfITu9g/Sn4YaP8B2+W5wLX1Uah
MKS5v3YSTeR8Oa/3BKloXJ0R39szvQYIpVW7Qz1J0fCtaMSYdMOD5QCfOzMj+e6FXUu6qlkODsIB
/t4EMcBl2SgrhBXhZrSV2VeZ4aZU8TFyUP8celwU9Dnu7hH5RM59/Z7Q5yVcTdRC8x10p84nKu9Y
XUaalT9P6pCJh5VhTn6iLxz299uwbLzrsR60TjqblKLhbmQgBi2wgr3JkM3FQQNAe3U6DS1ZZzo8
xKGlO9gguuZvv4ggz5Z6aKM2dnBvrwj8RhC3QO+PT1DAphC/+K3j63T8X9AwlcCYCaKnj1EZo5/m
kVkn+4Yn8OaCccQ7ToNY1lmywt689+D5yfwOxK1rNzU8raRIYHl+9wHfphykrGgESETm4+pe2Jb7
B6Ly2kVPRjVauefqX7Yxz8l7MkypkkU3Ix4YEMIBdQoQW6VU3J0ee/vuNBtn7mvulIo4hjYwxcyJ
muppz3dnkrwYUBoOTb4GFidgOGwy284lD6GsInMXsS3IlsjdIMgJk0kflwBwSAS+lBFFdxqkJkY3
p0Pk3eQpqjhvTSKJAAaOYnoKXtlf6YA270+kLV1eIY2mdlhAujd1h6H72bRsuCS5pnogYqT+yXnR
eKX5yzz2NC6gGfE7AJ/0m6ucH48kvQrPzqv6JfuAfoGM3SMiZoFKO14ERstoCCxtetZP6ymfEeQ8
O2MKmaZFJTyMvV7ZK6f56bWIfQVOr9aRvTZrk1AuHM3gE21PFrNPRLi8MrzBG7tHjiBsLmzimx/2
3iRXOuskfHtELJEdfNL7ecvG2blQARcrGu9BQWuzlXLRPPvlK5/w0xUTHOvA+XP1QZaM33vC11AF
6j0IKQATvb6Ahin8O4mgt8bXDWletHb77tXYlK92weaKk+v0Z4o/SiIW8jqqqpBFKNcCpy2fD7If
yYxJJ8ilWckvR/uONAjV//Y21fgxHNuWO0MH9utk2MUXDhhyJXqa5Ts3whFBOmgPO5X+Wu2JPOi2
35fY/Tu6rvMsWBmrQMJgdJRXOQIJuVgNN/EWhKRvHaOPcqDrsw6HZ08fTAiIbJ6TDVrFurrjmgzq
uVU6X4Aqkd3asAmBzbO9nnHW35LaxQzd19F/LNl6LnDg+K2su/NBPP+YO35JE0PWrnDb+K5//wRd
Jig/aLgzJJDREdQKuwoN8Im3qbfAf6FdA/k9qgFQNpB/VN/h7faxJDlMhJ9eiY4KOat5VRxdnBbs
5fwEdoU95XRJnSwYsI3VTRardFEdX7aFO0/Pye69/BJpGzZzxgCepiwSsEBScXCaWNQjsncvPzb/
fhTFvEWK3uzzp1Tx5xibWm5FHK8eHHHtO9IZVwZyNJqXo/2/mMEOU31ZuiqgqlU9BUJOjtMIy8Cb
6IigRKTzgDQsKhnNZ2/wNoRtc111PVR+u5rnH5TpN6dBkbAtBDGhAnVEy02lxw+So3jPdcDTOqwI
0EjlXD+5TKxVW6IL14h8QjrJreWGb5l16Zb1EjYLEYhfUeceytO5VxWKDUod9TzFuOQm9GUqOB/b
BNub7y/+pGPxZflCQlGB2YadPhDO3Ji1n04fwG4rIYmaF2XT4R1wJr3r8DNTlS4NgR7yohJzO7Vr
JrGrddeK0TIRGnvIcFxihP57ZWZQtkFge0HPpGVZR/6SXuL8qr23VniSyXImFdRmClHQnKtm35jB
sM6dEKe1FctBU2H/9Kw9YkzrvMLiq4IXuU4OWjlUvE2p4zp7I00G7KQeo9aa+Uw418SX+TwDAl7C
i8wrhDjzwX9paFQyd1GrNZrin+aBkiUxO03jCjSPgaeRCmyv5/8LFkjuwp68MCq34pU1koS3pVB/
8zvfKUrKVSL+li9vWwnPYLvAqh4ldOphuREh2reumIUmCcUamqxxzy5BrUYLnVZa0Nod+DeG64lJ
4KZXEwBeXm0N26N3+Tb736cunzA3hjq+SlPsHqHnEz+wBme7VmoiFC71lp9KWAOLF33wY488uAlD
T6MOkQltirSBxQsVO1SmashNAz1fBitYCc7/CTDgKf0zH/k9g+MrI4a6HUtyfL5DAfOC/gzsGxF8
+lkmo1SM3DcYWbqA8GJh/UIlPqy6iL8IJRDOwB3IsjeiKV85GMfnmERehDolf3vgSaHeG0LMslU5
2MdfhhDOzVDUPX+y+r4o74mQ38To0VZ9Xo0ccJVRCG5Jydq46OV3TvmfhEbJnKzA/lsH51SfOD5S
e/ExHRHsQG1rm0ckmgckpNxkI9/9CMqam7xfTxo+Z8JUDdLQiNcyFEghPvFm3ko2MmWnixra9s4n
d3WvlWKBAujefdxbMIuIClMzi9EC7PUu7Vs05Aska31BZH7wHd9GCFXp/cxdHQsKq1vZoTqi5ZmE
D2528TFZNI9bAqMPQsm8uWdMwmgXw5CFuttIRasVZfAAK1xFnwOxz+C8UQGUHH/YziZLY3hruzz3
gdXnpNfcxDHGJM86rQFqHQtz36OF7EP9kmYCPJy5HT6pzehzPoknBbZofvLAEOUJcZUgftShOHY/
/air5bcHX8AH2xmxQZDVcAEts7gOGb0XbPyoqZOXkLpOD+D6+HR4F0ZE62K1yIdIOVsHuhJzMhRr
8kMCti1cJ14bUMP5AIaD/tol9gbh4BZ7oYun1IfPbIrs4NAy2j7qYkUczB0WBd0ocgs7sTH4Esum
wuWD+ny24Gy0ai5p6yznW82aRHzPlDeGFOTSTe0rjgCefgwunTlVfqF/E5Z7QX18hazuJPqdd+EE
0qFsTAcJ5TGiUz/X9DyfnKDcuPfXkrVLL01kMsbGDq2Qg7tfEbmeVbY2DhQ2u4KlPc80P1TsWTg4
d3+OGdyxMDlp+nolEHmSrY4D76dSmpszNK4HMRBkjH9LlJDqwqn5QQ7TuyGTYjyPVtY0R5zW3E16
nmDCFyz48cIt0k2oSXWmRPw8PvSgvaAXl+/CTUolXRPK0/vo6uOp/ooSAQUPt3QSxckM9YRr7flw
nqd1aMjEDsFLGtu7JsuN4QDRJokwCA9aJVA+FYTFjmr/iDGT5BhXCSRTSf8iIRM+5VpZhAXX/LuT
rumOghMmA9tt0h/xuYnYvPmDLBz13UUjAEZ2iIBpjDXDmBQwM0klIAPT2CFyqJdl7g0SomN3EY8N
Dsc4RNunj0ASQ0Qzrfps9TMUS/SzbSimysSFd8drWXocD3g7VZwfoiXj8s5XX+sh/y5qxNsfpkvC
5npJtRRpJ7FP+OW29kqNJptz+I0vN/VKlCscaIx7I8cV1Ya5l3V+N2pprfA9IQZI2xVEXJ78vhQL
vnwtTBPdUxv8wh53qi/Z4dx0icUiaCZ3+BuCWSMrOPe76EzpNgiQpsAECiUfny4CZWxg7e6eICrM
ZMEdot4etLsKDIlzNP3XBUgCY/189pmJbCdVKXnLTpBDdGaNeRRqH6lvC6qOVFfF4ZHzFJIGkv0t
7aypCFhWMCpsFRDwHbFAeIFOw8WJ8Mi+wCsF5JPds2ao3GZOCDAnnkOGphZSi0rnWVHS+eVWQzgn
/6jt4DbxZynmURlUqyer+g3hifSzibGE1GNk58WczGYlRZRJWjY8cfVCIuKMIEsGrVbuYT4JaaU/
VQ9Ahj4eq6RZvx9FV0b+ZKhpukuI+pWVosERpNhNZIUwSxllQXhnhfZK4f00Q7ulqG91gNg+4+Lu
kq/bugFsPH769vxiW0NCMGbRXA10RImVmagpy32szmLJXqYrVZYn0RfS5NebfYby5O2KmKfT30wE
hw8ETBihVO+FgB6Z9Q4skshew08GO8LCUbM4UaMAIva+xPL8Z4+/ezd6ddn2X0GmSzZf1cnNpjwv
R8mlY8s1Jcax/2tNiXJFFHqYVGCb4xdeQvR3QCUXlBuAj1e5yi/FKZ73yHv4rf7aNcMyl0CROp1E
uPefQa200RQNiXinQiKX1+DcMWUGsNFUPzY18AgJFD5trjzjfU3oFUwyoiiLXUSSx6DNRh8pO/IF
2pAu49HlCf6N8qNUY5Ff8rojSghso+gXQ2C5RuoLCGVrQ7tiMkJnmrFopMgOmr3VCKYbM01EQ9ZE
K/LQwSvdfNpN1oNUIy+bOb/GhasCFXg63Y5nq+TQAoIrJcQvQkK7abpcoLK/KM4Ti390x+FOh/qT
aW0OzWi3IvQbKQzPZ7JEWf4bSJlUaRXn/c0y4T3KJageK1HZA0ZfI1w3JK0Urx6IY5FqmM/HxJ0c
f4k97ZRx5lmAWhFa/JeCuO17Lo6NMEzQD3OLITFhnk8RH7MWvscAGYuqFYRA79zdj0qR2VAu2hoP
hmXzY9++oHAx+2ehPdr52L7+rZz7w1/k6gvAiXZbr8+x1MADgJFlEFSIQvWN8whG6TT8pnxC8uIe
I7jZwYLbw+MI71cc2gnVHrQ+WY9RX89P1iEMw4a/XzqUYfbtAbB/8/wQH2a7BWhe9nUDkMZTzwhD
IDmvt6aWY50MbaHdPZJntjBzVwztt0GN07pBjL4Mi5Rn+gjrilr/VxDVLqWY/xB2PmWQx9L6+6qr
5SBnH61o6Rhi5SL12+COJU8U8e5kjYOAPn08hHaTx10SLjFJfuV+7cZtwMRCln6Y3X6Y2mlExUNi
i41gKp5kQiuwISfWm9WHiOAqFEJUIW8BcVyP31ljQQecJhK0cPwlxGo5I1ryEGbKhpgTIV5ew36D
aqKMjFcOfBYrXysRT67NRnRQ68ibWWnGYf6i8vxPQgXQR+qRmw5gkww8sO+a9LtNpKt9ZYVnRkux
gPI4cW+VJCGLq75tkRJM9gxbRgJLH6tpGiMrBVPJp5ru2P98m08CbHi5laWbHwilAhyjVDGtuLPm
EQjt36QJoTFMTJeSieugkVk9m27i+a8jDScZeI8O9QdvNPeSPgLtHO1lxxGv4yKx7LS7YpeYbJq6
A4/zbZhIMsy0cxhiVxuLmlwM2aKmVF6Ky9tmikGluX7Xcj+r0iAEtAmjNA18LR9yLJN9DehRDHKJ
jNgZOhTlcEwY/WDoAQj+XlF0nupDD7XmSqxiuEwrhj4BTGVCuhixFgHW4XzMyCZVtJ/b0ta9zLSL
S3SFKPt6rm8b2x5KrBH0XFSi7E1BjaH65jcLFBrzYcctgnDUy7WtfopSM/33mdrnfPnzb92QOG0S
uVsQ1Yxv6GdTxpjpJTpf6+8Npxoq5xwBLOdIVefSOWtenpUgkoLXoPw12kEZZJHj+5g2hC/C7TQk
DnNnMjA+dPtEflDe5KqsH54CT8tIzBjDLNlS3OMObrJwbbGQwUHo6xMQ8x9Biok6jZSa56cGDRuR
RsFZpDms0CGmpY543DKbGTpgoOUOwdfr2B5lUZZlK12C9c3gONw9LV6CL8e7ikr5Fh4PP1rxPdbG
M2aPKy7C88S6iO+JrQM4cxzGkM8FDd6b/bmtSUT+znGbVmqa9fuP3/RJ8NEzBycSbuhougKj/RdU
wUpJf6ewn08gAzzFBOHLP5beUm64Y3CgZ/P0Ogaq/Gu9YBx9GayEOFfGN7+/CZy6BIihAKqB1TsG
raNKFN6Z9OH4cu5V1i5c1YhcQUcvim6bI1iy7tdX4b1ACPkSBysmdN/vOPYERg74q6LvGbhxb2F+
wixG7Sb4lb1vCOUGs+XTkcMyAhskJ8KsNuYMluOeHDqzLQHi8j8APMSFiuOG2lk5QwRviGp2X61g
EjOs6HyynhvtZZi2OqEutKhDhiIUEvTGC+aaurK/8m/yedqHpOp+RwOgvrhjvuk58PQy7pwoEtWs
9h1FAI3DeXUmeVGXgJy9DNINMFQTPPRJW1mImFqMKBNo+182je5y04FJwL7QLAU9RZpZEU7GEU/V
y8mLYfQ6CmwmMWzQsqh12iZs0jdgk2sxPVVjqMPZladgk8w7geCXg9XaFI9mfTJMKn62KevlS6c9
Wmzal+XNCLCi23XBsH6ySvbcggEutYCvFRKtCYp+CvMdj0iSpJql7hRXFhuCztZk10zDboMLYo0D
Yty5/xBhIb5MQHlPSVONDI53naooC+Mh8HEd+eH0ZIe+H88aFlOzgKPQUyXAHy9rjuwAoqf5e95d
D7f+mENhxWjhTUpSX9n5DuYcX7N4kgfDHxb+Na5d+u1wPvrjARFfAOaCP8fNBLpI8b1YBiz+cTs2
P3v+eS+st7j+v9NDCghmcQrw00cncyHyfoBBzZNwvhaaREPRDXdPYUMYixOsd086BXs9dZ2nmv+J
/MKymmY1QqQ2dWuvStLUKBNcj+C9tL+3F421dmJ/cziyVH3R9ekiwI2iEhn7RB7M/vKk5r3oz2jD
+ziR4tbnNBSza9sOEB2RCK6rE7VsLWNdiYSsz2vGCjmdwN1cRZgUBOOF+DSIX3Sk4gpnYLR8g1zf
CMUOZQKh5HvBS6x70xKc2wVzDAh10uNuZ/Xz73KXH0U1prro3pqqvdBPDpZs4/RTIL2jniw2vNA5
vewTa2UD8+sS1mB9KQQzCZRdBxhC0abo+VaPKgw0zCDZQ0OW/twURPyDiKjNJPvmMBNhXflUVEnP
3ZZX7o1D6YU2ua61H6HvjCdAnQ8gpV2x5/Pdq1v7A2Ue5ek7Y2owCmhslBzL77ogp+dzZ6sgxhON
elOW7PKJVT2xdT5kXjbXoNerW7or13/eG8xumWsrgJ/1oGCD+n8mEkl30u9E4EmElZXuaacghMCt
RDLCiUc+34u9404WCR14BDB+3Vmirk3dZ8zDPGX5TjAcBfC5aAJSN7eUBjCVPBnFpVvMznaP84QJ
lePiq1xjm3Dlt1FjwEnPtypDHeinxycRbBecq/Ukk/0gMCnZuUy4+2Ksz7VcyMI+Wc4NEyZloO1F
EGN23vytbHcxbt90EgCPoHiEQZsg3Cj5lgSTjdWRLrBKt3+KoAqLGMU9fTE4GYgnhi9MhxbvskbY
BEGKk5r9ujLFWYMPGxkzfHxn0htDg5SHC5Scq8/Fxb5mcgWTjbVAPtVIxInupakkcBdIcEKgWaB3
Gab+F7NdvZhgo6cmFrM44ggP6VjS/po0SMxAMtdkNVuqyqs1sZOhmvVwVf1SOGQl7axA04l57sdM
26oHwoAs2opyIUNSUIlQdoVR9D2Iwgx9muXDnEGCAJLd2UaUbIaDekGWNV9uxCIar4XnLqIsbY07
hAvzBUiYjSfoDuRU9EX8a4BYum2mQbrl639M955cylED5DmjRTGMJc8Z/Rf7MIvkYiO20fTeHwfa
oBIePMVTtxRru3Sn+xpU8rqcY9WqYy4uYqi17VoGaoWRx/FoFeM16dX67HM1byMp4QBG/PejPmvQ
p5CBQpVaNb4DhGrrucIQWcSswIqHKidH/XFkeyjWQpvMryNOBAfsfphgowW6yx09Iv3gXt7Xga/r
Y6MXXnLSXSgSYutimauS1/96Q6b2rSgd2wGxrxb0LVKyOVBecJXNAK6e0SS2WXDXAE4BbtSvKfWg
gQYMyQEYh9r0CwodhaQ9PPfo5WtPBvGcLDDCJwK5iQ5QwOV7vzCwIyk2b9Vi/bTBp8Dk0dQ77bA2
kAkGcZUJI0kyw3ViR/mh5YjVlig/Hejqq5i1DJf+pCICGT8/8dyyYwN4SPvlBHKIECJROSp58STP
eqsDk62H0YFNRWeY8YE6318Uk3VmBJMnsDU3ugdC+C+Pc42w97pJssJS7i6M4uuJAbOBCG9g/L1R
8RVpQ+kajf65rrSA0qDzF7M9B2OAZvVFFAeODfDcpT9dug3IeA2ExWUmv4J/wrrzB3fMo1vOshzc
3gzm7F8Zpy/vJSNjYF7R2FvYvAkPEpQFHfSWtwEw1lQ/nCjVWmuest7VdCRFcda4NP/rgg4gndGe
kOrjemuXPU0zNUtrNd82Tiz0Txrl6V+FVpgv7pzdNKTpMG0lXVc085uzOSNDQijCs/Y+x0HlBHZp
aBloFamgqcmZmtCWwChayY5ZkdI9wFgpS5LFsUsUhEwBkxLne5jRxZvkzuHi21qm1KZaksKvf9e2
+U04JWC3P1iHWpeU7iWQpkJO6F1os44afX0jtQsCT7XTBjj0x/5PUxGgGZnKuqBurUYd7rytjMKH
kM7h8OQd+bA8FT/KB5GHiqjgoDDz9A/ngdZHskU9gdorR0Ht62V1uF/Sa2aGi5QohQ/5ODr6i0G/
xVPkUKZY+4ZHfv8DUM046vI8zbVlaico06rtcQ8/pJLZ+6eoccAUkREPsR/+i7cTmGh0jjT8/19N
WjzdydpjNoCsyKZu/9SVtAYzn2N0ezGpmQm2B8B3Sv49MSw/FVVAG8BLE1vpr3zsvrczTpE69YII
/KiHm8TR5XqQmREb2eQEjGJJ14j9/Obfw1EV4RTMAA/mE2gb4Rfz7J5C1U7+zaNA6Fn1mEdWe7du
49m6ZdUN7ugyJ7QWlCOcK/MKmueP4DXh0zd7jy6XufRxoEXBSCQ7hzbG1nu1tPFLcA4KzqJGst7T
L4rWov/oZGR2InWQdc6XpjkWJdjBsrri4QRQM5ewAKUrMBzEp2AVh8zqH9/l9K2RPOA2v7VB84Fe
JWtubcLzXMifSAiZlZKME3DBTCtty1xm/1tJb1ORdODm4W25Dg5rbZ8ZAHCXdIsKXQ2liO7ITDjV
Uh2xbaKbmCvIIX/xwQcuwHW6hJ1IRYcLFAHmKu0NYKV27epfer9zPdYFm3NmmiZd0xo/8Y9JXApi
4WlVCCQvHFqk8hNsGf8xyADaYE4SdJKmzRBOKT9X4UybCSUjNyPgFGAwJw7KMrBuymIg2Rcm6Kmg
+aeBVJU5nUCkGDRiM54VLYFtGAjnhJrc+NRopD5vh2+oI+iS/OiFmGKhouYUVAHviduEd4qILWtg
X37z2DdNgtJoBjaabGQUFpNw246RQmz1uVAGG1UWEDiTYMnaKJINzjzCi3Q86MO3QiBilHWhFkZQ
Tb2I0yp0DJwZnyU3Ui2m3U+i/qHNSBcXF36RapAdQumpTkWGfQakqvUZLGmoMfRRjTFJkVS8Vr9H
lMX+G+iyiuwMRDtuShQcEv99OyNGPE1rumPNv+iQ3PfIZzQlI5jPFbWPlYzAj/jAgnILLugm/o5y
gtoIwnsLYDDQWNXlXSki+i9iDaOi7RW++p9w1wdxyoNiZ9PPiczoj0xWG0bw5z4cPnsVSZbkX/M6
mN/CsTxRp7xgDzRUXllE07fksTzL2B4aWb0AvUqGBPoTDyDtGETpEKMnSrExfjTsZ+1FJmvIDzOX
9va8kjENftvb/SlGdOEtx99EWLUxw/gETWx8hdxX5NBR5JHb2JpEpCKkKCeUPJN5fAW+flawbFdH
eMywsTwi/BlDVPTm1n6/im1jpclCltHx2R8j+XlG0Q8aTdvrSngRd5Nblo0QyVg7pzgaXWGX8whz
oj6aIpee/4CY+sKU8P8ybbz6dNdP5/XQMu+61byL7tlA1XY94uhEyPzbIvrfzzqSGk/QYiu0T45M
RoJX29L3b80fcJwN07bUaAlL1Jy7mTKecKLeTqoPnqLXuKZ1whjWiDohhj+MY4JeRsntuaWW0KgK
s+lyH01eJu+iBlilIIBWtGZrucIEai3HNaalNenGqCONrm6wKDoZidwx2fiDoJxIJzHESn4MTtOh
494KSz2nRLiVKKdCJkd/pjrGP0ewpXBVCbUE+2p7Tae2fVQOWa5D8hnfD4akpBK3xL9F3WZ0rxIX
seYdbEWmsxjmMRc/0i+l4Yb8pu3q3Da7t9FEtSvjZTAHVkWweHmuy+yH3/9oPe7z2hd7Bp1/dJlx
F3xHrggePZ6mem1NGfpkjLG7fpXQ7G0JRZIImyGRM7zDA+FvubdcK7cVPbrkiMlae68N8HX7kcwp
Pin/AOs+yIpW4OrrB4j3pQU+ahEZFyWNaZJnVG7s6rbpJNIwBq2nsZoYM7pm1Hr+VlcQiqGKhwxb
EpsAztUi33ne0B1N0yCbhFn5avNohxVVXBnigvM+kgUW0tF+b/E61qwDw1HKbWdsD7i/3n6SSoJj
+g0h5FP+BlU/ET9pOzVXSx4+Nfs/Ay5Bxnnyj1XXCi2RsKNE+qQMyPGNXV8d/vOxeOzlPEtnj2rq
snuYDrVKxI6kY0rWmnwYCBuoaxe+SJpHJXlGaF+pZr0s99tEXAVzXxsF5n1SmW35uA/IU2243g/3
xQiyveYXhKtuohWt4qqEmQA71bf0leNznBEAk78q2OMLapsChbtImxvq+vx64AnBNnmNF26MIERa
t7AEPcraHx6eQ2VnYc2D+0otavbt63KZWM1ryauvwyh7eqRQJdSCU6/nOhUmRBH1zGtDO4CGlteS
uedQpeEuc4FcXRMUsr6Tqt65AI/zU279ScRSAUiMFf+7Gl75RtnNPXYkEBBOw9+oaJhGt/DJQKBV
pEeHPuhFopZODdhOaXDSDJ9hqs4+gD3wZ95VgTQFRGU2so4xyRoCQi20z3GV3pbxs/cWF8k1f+Zy
xuXl3XWlAN17oejV4pAYeOiWOgVt2e/Bp1670Hrxm43RJULwLJCr9T08grBDUBsQldqAjocKPxD/
3oDq+rPSuvmWFoGCDS0YwEXzxWMvLDH1ARbyD6Sel3Ue+pc1GXi/th6e3y/8cE6BC/iKQZkjuD3r
lZ+yrCj8DkuezjL47ypF99BgF3ItwHXCZKEjVmhzVAqAeg+3ZrtWZGZanTY+AocDHNqX8QhhAMrN
KHC/IQLqMfRBVxHrHb+IYeaPERIxE6BpDRV74ZpoXCnxcBLjC/E+4yorPCxNqtv1ZnQ8Z1vCUw3C
3opu5c78Xubp+6tMl9Pu56GzQSS/dKXlIi4mWUOxGlq7AATZXsjxyfUW9hiQ5JnwFMfViKhnOYjf
6IJ6JeH3/9Ku09uU8tLWc2lqffpxeLX0vmMggN266etvlPaxuBrlfOl7K/5PwjC/5T8SkjpNsnkZ
UJ8BDcl/ca8+UqiDcV1UPRdqllngbhCXLd+80mp5etBreGYL9GtHe9BU2KjthUyJoiac0iVEX/D2
iAn1cbda68zZCnNi2b7jtJLWWSFlBEzxIkSGZfiRIuUzDWTJgnajUtFSgZL836F8vjJRMVG30OLV
AQf33z6vkuvq+A65n/lzLgiE0Uttjv+CYWDvJiJXd4j28WukEu2e4NrWjw8b58PP7qqBCcKalWuy
/yKEIYbaAhbcVypWUgj82W2wKDoLKuuLKn6lmjOOO0FxtE/PjTarAd2HiyruGU9lFg9Bn+pqqI/O
Xzif5QuZDJumCYx/sCHyNAtyrY0B5n87D164aDF51tmSiT9q1dCISSXyo9GnLVFOQMCv3WymFvfC
Q8KVqW2PWy2Cgb0LGxvsdESblHPRvPc/qCiLUSm2KapOVpm5/uy9F/uJQ3r5FRuQLiCj5pz+lRui
MZs/2IKXxHdq6HqdjDnU5mDrTi7vT0waNarmo1diPxrFnQvF4iPA6rjzWSAkUvwt+i1dxt/zLd5q
uoujFVQGILH1Zbr+Qhko0CDY9J49AZBH35cymqc+0SCd1J+/UitkvDpar8Z8E2/3/4bpkG+7RWw7
R2zaQtWIHh7WMR9j5u3hppcaeXOP+xzY4skq7Sy7NkZ6TMGQpVPp8baoQbB6/fNcMB/J2R13fX4i
PMuQ0lc46k5yMat6pUQgu854ICF+5e8IpZck7lS3V/5LODn/soxdkmvnMjhqyZw7jvVjaF0fCv+C
9jKf9z08jOf3N/tyQlqL+3Mdn0STV3hdBv9oySCjHGkEllbQv9YayS1E/seFKgWi+nXvdChfnef8
WbgQMGB7uJ1X0yE5PpEALcfWK+E7pMYdmtXHaR5lwLA1hC9hNRTrZm1vWbaTNU8w+KYKEtUnS6vS
q9mwUjQRbQ+NG78fSqB9gFY/UqVKfAjykRAo2zDJHZlBQz5uo+GRfcYsYy5XlwUuxm3BGrQrI4tG
nVkFQ0RxVz2/+OrlFUUsefcvyDpYCYoRlumzHLeC4ejG5RgoyoL/BRHeWri566d/cH7M3pcWdh2R
CJ75XVDxMnKUvP2YoBOALZSwOpu5orbjKWfLauMda/YbJAxxEjP9ePRPcxgF4CvxmvslsbzfI5S0
jqvAnT6w8iHNHO2NJ1be9lmDiLNJXACU0EmZI60LiGVpZ5gb+y8SKLimQPSieoIfdKzDcsn7QrO5
EBR2/+eHRlOq6cMh79umw5OlmJuAk9tezS+DzfN2dkstbRZkwLsQ8bVZySiT8sbqzqw+kHD6sxI8
YyuCK5XJg2FnbaJ1ZEDzhpWu3WgzkodmuEU4YQkwxNZNO4mP0WzR1uB6pydlje14sb/7xQZAWLbp
KktVlaKr6AlkRDWHOuSF2sj1Z0lhaeaPBlfGRYI8QIUAwN6Pph21S1tK5H1MPMWduvjLEXl831D7
g1NF5NmH5Owd8yRqdTF2k8NKSfjI3ui+KPgClUe0KJT2JOcXzkc4+NeUkGQBO0YisEMa0kHStJsS
lahfi71KHlfboGVfWhFfkTlxgcruuyMdcK4WyMNvkocFVejxD44JemINY4LeyWQZVyYxNY+v+GQi
i+Ub041mrLpMuWXQwrLw6h47Nt5QXQjhdIgYkUFwez4I5DsdKnHLvmDuTJk0z6fHgPGse2xktGw1
AhR0QdzNOU/TmizPfqPrng39UivNAcA4nyRt8S1m/+yCDrLDmkTC0i6xlhWvBe7dQP9QV8iQuBzA
aZzEHnWP7yOqtiINYf9JerEBZQ9bBkuDmDoTm3bCRSDwlu37AXBvVoqScEUaPG0JLM6xyHKfy3dM
bLPWPnZJ7W87hOVLoNg6TvfabfoWAfBjX30+9wqD3OA7Bmr8QePaOWiElBXMdfkpemJlq80ysuM/
9xjnXkekcxH4UG8C1cGXo6AEMW1ho8BHSV6BBi/bXsk8UUhUYCIz+GOgJv0Vm24YcPK25SU6jJ5J
IHr09vFdV5mfqerfwwGhc0IeP3wWWA6tE01ZpKig0+gP93AGPuLOGxeuknRxhn+AuCujDEHH2Bef
VyGMTrviJqRqKTA2Ak2bACXu7ekf9KV0gJcsKIasKF4rTGV/UqdaQS3XIz9Auax/cqGlw5GZ7NYw
USn1Atnu8kC9ZUsJFthubf3kRg0QGDyIbCK+8fykPpfq7of9xdkkSqmxRd4IVf1jIVjPUc3G+Fx8
BJq17C/rZzlXaD9c/HjR3odD8faF6Z13Q2BD6KoUt/VBR4ClSuzJmQ8OOASz6/dWSy7Tn6WDuE/0
o1H6eCwq0iOIISpk6Uat1ZGoeTif8LzAMiRLU1nZqU9NGFkba7dl4o2WeJBljTVrXgnqny4J2XQ9
y1tjH8L2mJqObxE+AyiJ9YyFfMMwaecvXmF38wmR+7sD+H/teeM08Q9a+Ht2O4mNLCg+1UA5veCn
8yodqQFhBtzwp4UcYYXPcnR9DiIadyyOzgnbvJTAWAdoLGzxS7XKlDsraDCyNgJOc/01eCAiggTI
tFA4Ax9NU8S/+zE2dQhOAXM3B+6HyTHdvvLZm+bhuB2ql8I/DgvFg9mKii8GXiABudBolT2I1MXb
Oag/R46n9j2ShQd+pB847NGxJzIuS06ejRLmKAxJ+DUBoXQTrfaGPGj4/m97A5hXJIrkv23tDBC8
aqaV4Nm6sMdObdlYSE/BR0k8p78WY81r0HiksDLEOszyiw51eozOC7MdQNYpmrLT8i18F/+nlRuY
6OrxsvMYKIO7+I+fQzMGiNbl8nRi+Z8U8Yhb0eTUVRLqMRjqoEY6TNzJhk0CcPzTjNeokoNwpey0
YYzZq82tKwZ5LbOL6pphOpzGDkowpNOPee6kTw4/DixU2HWFjU4gVoNF6D80rFHNjaec+PeCn/Il
5BKCaY4GTY+bKEEl5NYAYoRiLrsgNmBfrZK79ngCRFJofdUq3i/xiASjm5tTmZOVR0G2+wDwjhB0
zN2ycVBXF0VvJlxS/f9Rik8teOtui2pLRY4qPHU3F/sOUnAvtR93hM0277U8yGId7t27aM53fHZV
ql+tV71MtkJ66w/EfsIX4R/8th6b9ZF28gfr/LXdbJUGBaignR8TgPq9G44XhTT1uQBjGHbYWVpy
S0YJ9Fesx4hYSKMWzFt7jBmII6zRFZR84gUVFYZeI8uoF3nOEFGw3eM2QxLyWjQ8rmtyzB4I4e+c
Tdp9gESYHDfvg6rGUiCd0uFXs3OUPww0hiqYBfS9TXo67lC76E0guik3FWTayBBDj4HrrDTIv/4S
eXjB1u8LWlWPx7xn/2tDyVfCnvn5NFN1yt6vVbSVWwS5CZ4FfYV26Zqj4Kit8oYl1ILYrpHETdem
95bZZIytGmyFYROHLB8DUyOxBM7aPTc4oZ7eRGGP80c4WR0HmWoJUxRhJUgQJsgMHYLX0vdBEpYC
ZxeHszhL5OAGUMIbq6EfrQ5/8VM1W2pXXP458cxXjFCoeGx+RMyx/HQrVpAWqX7NRpADvhbvlYDC
uMCVVnmQ5UfY2HybCec/qJZ8JGGnVbO3zX/no9PXfbIn5AkgNtCQ1gKfbxrPhTOptDngx8kE2kCL
3nQuktQqMnFreBNRuAvp/uwCKEXNIlAnwnQYeuCaJ8YQwdbG8fl6ncWZxkXb/Kda1lT8Y+wQU/YX
PeLv6ZkGdGOgSnlDhvGSIt4bnDwb0+PuBM2n0J5vTiqJRduFJq+O/dE5irhVU56Dl7YdZZr5W1nB
OTESttTF3ktZynwmNsw+vvh2AEVADgDbRjyACnnIceldvU6vOuQM6LVX/B801f9bOLZ7AuzUVksV
7fc1AzfP5tp2e+FVE6+dXC+bn79A14hruQ6iLGQ0jDZmvvFWpzep4RzFeTnvDEmQvbKJ3Qvx0rXt
6d6CIMmp6Edd7yULy8i0hovHYIzlRggiA7IVB+b0MVPPDdLjUY1UjD+omiPe4VGBJDHP7Bqyj459
qpDlQr1+Y9wyQaqb6o+Vo3xHlxkhaefESNIIdjLR6SYfDdXaVuo462Zgh9P/IsE2Jgk0CyKvskOE
ceQkPIaGoBcyzDlTNS0y5amU5nm+68wpJqgCJx2s5Kd8c1od35QgZl2LcDfQHHeNkgfpUZdFrtgb
XoXNJUxKN3Fsfer9ZhgqHG64mrWHI+h6KX6MaxOI38AMUttzjHvmLs5qoFMMuW4e/nX8deZ453Ey
7g1oEbdyk3pfvyGD5ZXGODiV4HBvp5sWC43+PyoRSO70uaWjmbeDab++LW7vduXMZSbGA1Ou9JvX
NteQt3Y74NzaPdyn7+jMXjlVsS+oYviYtqEpKim7T636M9Qrt/yMG8SO8+0l8t4LVnc5nQnmtbOr
08ZnAkg3Yd/nTnnuoSO+qc+MfW4LgRLHFjfG5KksD+wBvfGaEGcVD64DeMICM/vODOhuihsK+sQA
bmlNbRzxwPPQlaXbI/hcrYVqgH8OP/3Lebq31d2JxD1AE3s6BtR628wJzvSL8J6ztCXuVIqfemE8
URJG9JOPf1uC57NR44tePGHWjIUfzkjp8doF9VeBagUKqx6dInHSNyfd2fAvYTeLyASQ9FvWwmXO
WWTHC3zRwe1FPtRX67sTTZedMOO1ml2Ndy3LkBfWtQmX6JNgwfO65InYFG1rkiu6N8d7mHAFNNDg
`protect end_protected
