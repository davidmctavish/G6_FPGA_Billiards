`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVxyk7XRM4VsQcD0QPYws4xsTeDPKdwWYfreQJ7l1z8C+G+JAKZ2psrNI+b5ecZ2ziPH9MBGr/oY
8XtzCKmjJw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VO3Jpo4aYF9TyVwyAUb3a/oDy8Yhm9ea/9mAjNtuOBRL0qoy0/CWzL7D+bc1SnZvEP4BG903Ildl
dM2y4TNyVTBUaU7Cz+LzZfu9kCPWnmttlx92LcMKLNuvGUMPXmV5jr3PzSFEvoDuCinMqNc8uKFO
Ux/aX6fmBD8AbQfpK30=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qOkimDe0rSU5f1zKvoE8a4lZw1WOOUxh8wtTIN0ys09AXuQuNNCdfu6VL2Xuj0Xus09sBU1FazgW
XpQHuw7XcozHRlnUFKPJg2P12yPJsLRkOqUWtHTUXmH/8s2RglOoEcmFeX9FVh1IRMdnp+D/F4GX
/80OwH0Jtm4eUDa5EFkNoIfhlOG4JOG/JCsYRnsAoZAbyHMEk6qPxdOGDrYzkbA3CMCikTuE6wOm
0j69ZgENzpWR5aludQDu44oKZqgkdMKNm6Mvk//s2aUOTBYWabbSKe/I/+cEp1tWS7+9AAmaVwO+
KwmsZsNR4Ztb6OH4hCq0936o+bycwR0b+Wr1VA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4df1QYXbx3PmA5i1scwSy/ZAJgZ0wNtl21eeCeUI5h4IQD2UalJOUkc5a5UR/j7lX9ToyF2yFHzK
L4EoH+xXm54bGihfoaTvocQQsWhCDObbmBOtqB6WS1/bog7FNgoEObi/E19vJsjPSd6nCCdhglZ1
j33mJRkZed+lVziTR/s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rtu5N6w0tnewss9ZQUyM3gMzu1D5Ba/+qJO2rdGgk0QN5Nm+4TaVyiEXzVM5DP8z3mycaRD+z4HG
QXarW6RH4GHKahoLlSY8cryjSJRWS6D7/Z1joY2fgJb8apydMguGWjRZ/uW6R7BEimGxB3Xuon63
ZdpcvKZmoyvfg0kjAjor/DxtP3SP6DKxH3BeegGQKpP/+5EmCrAhhPu+NA21340wcbghotvyYusJ
ErSZhtj+1FLwV2sO7TUt1etBG8nf/yETDQPE7Q+zX+BzOktmY3tIKds/9qdyDt6Qb5WIxLMyaMa3
eyi0SGAuZdeDtK8Os3w2ajEZI+VjufruVqtCCw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17760)
`protect data_block
yvvRtu+tA91Rtyv3I35O4K6BiUlBjs7LTFLRc9twWgYZkATXrSpXZut2NlvE8mcC7mB31ueT2vlU
P9hzhGYaJ5GcmScpsC1FKNndMfl3Ug9Pqiw49YT0Xp/AQWIr+q38Pu2DmkLm87YVBi0HN6JMSu6G
rwJt5qvXJYVA5oSnqcy27I93z0KCdBaCW4BhEaXbMLEY+qzcYsWxGhgjRzVfC2OhOSpdpDr2MKHw
1YDri1cTZAVy/b3L8VUTlyQx4YRG+qS3u0Cz3dOLm9nglzh9Pa9XJC4+Lnpli7w7vpvakaXaH9W9
I9Xs/9ShuVul4UrHUMsoz9V5jcPh1iHPT9m0ZTeLUdfod7NEEFDW47vWU8XjL6iEqBvA/DrJKrri
hjJ//n7fbl9gjxGZT+IKqHleRVz+dRiS/uTuRo22UsAcWrLoCdroE0x4MAJ9vC0vScZa86PQBj0m
ixJFhU15XHesAUmaWmkIVFZdUdZL6n63C2nZpQmpBX8G1td46ib/xrjcP1HPzbr1hPb30S/GA95D
4e3ICss1yPb8NZCwvzZHNKYRJlVJ6EOWwDxLeBOjWmUySMUcywo+toi8FWztPmB/Fzs/gyRSBxsb
FBe82kj2NTjDK0dD4XCcU8bGjVOKNJ3KoJmC+0UD0jihX5N1CdPg7+/bvmP+MCdk3ondXZKJzYI3
9YFYkr0RM2BhF57jZwHcHHmFJrakmG38Lap7lsdonuIO5mfOOuicr4JGW8Qijs1+c7VMc6LUwGDt
YKznnHTq75vwwVLxmtGYpW4RTIuqlZmOJwC34kp9oVx0+wFtUxMvQgXry9FwUwb2gSWRseSfbmMB
auDz+22lW+enEoOu3PzG3plNq4oQP2K2H++ZU7HNTNGSA6VpJWDQ1c8o+i7+XEkyIqt9DZHUxb+3
HlbwgxRkMYX88B7lb3GnNDLF2YzkJMgQjpyPi+t3N2MtquCFuqNuaKv0LoD6+mwRceg/hAylp3x1
m9DKQ0DcKuhctFlcx3aOGMXc0mzgjh9Umxn2Ng7JEliL6/L086w36Jar0AAtsKsXZ1NsDDBpiIeT
c9pWEQj9ud2144CtZKOT9/hr1wy8/jpi1lQaHanlWWtc/eb1aDpSY58hPbltVjUTyizUFFWsqQAC
PGoqDXF3N036pR2Ipsz0lKGQE6qHOZ9IQByoJkJfVJQFD7arWnGsW4G4I9tdTj8LBH1I0/XQKvur
lSNx9C6iPx8J8GemXPHqEIipG+GgoeMURYc7ft3GzrBdwbTFPm/qrxT/0vdju3tRDBl4JSzWO+do
z/s/CD6wNYNcDBCSDKcprRdML0+tkUYr6Jexl5rxIe2GBG2XGRgBDqc+wBSNJY7VVfutmSr3NjPK
RJK5NldZFn8fT/rjewbLV4flhMn1tgsE6HhNm8GuRS52PpzP+BK3fCtYvb1mnkFy+e3mwc3RgZ45
5iaZGmsBwnJwI9GcgMGoWSDkSaL/1PrI03WtUczFAidTPvIY08FA8CTdX8Bo/j1vK5yj8spVzrNq
2YNw08dzyQOA6p4yaEO8Raki3qlKk9oCGUe72zvHFj8EIo6DPYz7MTOBMZh7qLr1JDqBA+iyQCSU
UO9dElHR49OYArhLqejxnXEbJqi2McLLRKhJoiH7B/feWKz5mjNEjtWpHgiwx6VhyEKkL6UZ1Rib
ZtiEI9gtUbhZ6XzaYm3TiIRoYgTzxH0j8bAv7Zy61YnOi5ds35hrlF48AdxPXK/eT9RxLQ9JC4D+
xhLyqoQdstrt5DgaM3NxG2mKEJVH9uc9wj8j/rmn9YrBedhVek2F8Uvojvb9UP2S80Gz13xgD5DT
uHlDBG0pjratONtNE06BnMLwZRtD8fOAmitaJqr+uurpGUSmFSP1C9+FHTWgzBTdRwxLO8vYdEOz
WFiLspZhFCxJpRdUt6N09XI21qtC+0+ZgVoJcuL102pig2HCGw+mVSkibp2ZzBHApj3TyyQWeR0T
soE6qVGrU0cCA6w+mgSp/LpLjFALA+nFAG3lXPvfyzy3nWkgcWbCXiItZJY+SdblaE3tEF0j7zRy
QEv4a8Rg+L6tHbS4IhpoHW2u/3VbDszbEYb4sRKfYUA0hAwJaM8jOAxyu4YRtJsjn94Jek1Taiie
hp0Ndlnhy5vlx4q5I6i8Nc99UyR9uhRu8iqRtT7nCYuJSAzDby3Uxqh6srwmKPrb31KF5pRhTgEE
hoDR5pRAhvr+p6GEHRm1IAJTB/vA3Cmck+beIM8DaYRIdaZnzC9N04oH+sWVHExAUc9WW2ZHotPC
yowKFvokfu+7look6EHxqKtkI6qUIsFrQgy755fSnh7+GR8EVZFKqkRCDv0zQz3m3MIaUQ9GzxNA
nVZg02l+SgGZHXvy8wOZE4ONpWcUccgX9k8Mqf2VrJEhn7FTdwr/L68VLWlWyJ51gTID4qsEbmQR
eUcVhXwZ8J6/Jr+tfQkihSE/r9/FrMS9DtCeXZFSTXFkRXX3jwy08FYzVkX1AU3nfi5uob/pWe44
jJ4c+H4TgTK/YFd0U9+b9+hcQ/PKCmyuUWlZMD2jh2m6YaM0tRHT7pTE3k+5NorK0KIzBPhuhR0P
kwadh+BfDa9Ed/g8FI4r9aO+bzUYkbubz1m2BkiyrHNUN4b/jhDQyeuJYsvVZmik7vXZ6GcS1rnC
ZJpUE1bWR8FcYhqQoncmXGI126qn791BoIP3g9UyBSGDJ/hK/eFW6lylhaaJjjVsKepmxGzcVN1B
mCwVpKVdTSGBmK72htH5om7KKA2S1rC5U1UUj3MbiW7ZNwfDd0USkl8imBDLwgYFtoEE1ko8C7Jc
eUprl5A05bpIwcNw4M1zuvcSJzD1rtWdZQl2vo3uekE+ox++ptfYE1O4Xj/2TqSRnKWmvElAWcGk
d1P93oZ45PNjviXZ8GjPM3O0qWdvlgjvAq0xdzA6x0TysB9PpseLW+g8nB6svNvi0GhK/LLkeLYg
V+VOQradYifDOr8PNb0cqid1ncvsR8+c0tlZfcJr23pLfcE3Vqz5wPmHYoK484/vAUmQUEHiXjLv
MiKyjk8ywnYHQ/TOYWuO5OiF3b4XtDucLmEyRzxNB7rY1i7qaj6wGs15PP5RLOMaDOI9Kg6163IT
YHmjt12E1isvBtgqS4df/zN19hcUsAr+Hd+fpoCiaRD8qfZT7eD2F7aDUpS5tVOH7gVSyJWqzQ5q
Obv9Yhw7rja/O45RtfCLUeQNveIdOxbYJdxtkbtNUL4THMOaUooUKNDHf2XRJ/IU29P3yYsch8DL
w6GDueFKcmhtTaLLsoIw5tztfz1OnR/Ji8//265ufazAczEkWZEuwDJ820UjB8sYf6rqgnsGaFMq
k4/RqF2vivZ5ejxFZq4j5HxYIkrT0dvfR14iHiz1gFBjRkaPy0KB92AudlRi5GguJSj9i9apnV0C
9Q8mNjw2IhqKOYuyV9e6QbBpKJ96If+glayPM19wkoNu3wYrQpc35Fto6fYKFdY6dhE8nKPhcitV
/uItKlA/SbBd82Zd2+R5YPNcmQq0sWFXHgntGjncAGogKw7gdfoVMOM8623k3ZSxgx+hl1hERb55
2VAlad1Z2TVWotbB4SU6fYbYbkgvMzH5sJuCqbAAKfcoPFz1nWbbyWa08tpLEd7dFgSfxRMD6emG
vbRwvFQQjTUHayp8X4YhTp75/cn7s7BNav/nMANVwbzv+7PlcCBDE/FAkBmre/mWCARVoeNQi9yk
Lmy+/QFbBCSDmgH9dT+J0qyptUReayys26DpOx3zpnRbUVqoevpDLpdsoEIttEWQIhHlgFCwxqwE
aRk/jq630RhYJrspYYhMKJx7vBModJIEGer5px3GFiyOMr4+4I2Loz4N0yOCB4NxzVtMSM+DMFzb
Yqmp3TY7W03MSy4BUlptWvy4cfrCDCrea8duJ43frMTKFTfbW+IerIgRfu6o1EW2xXm1cTpBK1C5
GDw5N3ENOo9k6+Og7Rv6BqrZrvmt4KofAZpoRQwtrvIUEswUfZzexMH0dWDua0IDEUztjkju9U3k
MYVajimuyW6IXCYU0qQCvsz9sBM2LLZ1x1Vup7fB1Ec5aPwU/UHatOkTm3aX0ZLYdmaCrVM88w9G
XHeo1x2sSQwb3bclHeYGqJ5KFtGY8NkrjA2kOqD+X2jo651hd0o8X/ii6dRA1MaQa3XRL48KOtEM
HH0PUmnhNz19o5YiXS60R4NMyF8DBJ2arUQqgtrBdHpYd+zsNwOO4FJe/HVkB0g9fp75mEMH5PiJ
iCp8PJo1jsqW1yWtRGUFGwq3z88uUmySC3W8F4jZcCA/IVM3H1z/nL/Xi6GkPU3ho614p2M5bRq2
14TEYUDIUMMz5OS3VFeKp3NLgKmCpVj7tbmiZi9T8Yde5BbWfETD2YjKPY4NPYiw4TNz+908oHc2
yTbewFueWvL/NaEUrh1xMwQw0DRkd8xsxovrukJPMeMMIOpJVuHAqxeQFIhjwyO05shLRO+8ICOY
lVC8RDu4KIeHaBIdj78ETsgHAau5157cMpNdCv1z6u/eAEhsPNaTpoYf5z4Ulz5+vbrw+Ig6ywPW
AC3chkAwdqF9uooKaqUaS0uaMYKHDaK2y5UfVCBUcfko4mCk+jjZbqPR4oE/RY4mRKF+S5KVRb51
goeafsPpARmOwOZcbpLNMXGonqOUJEFV7nFBn0sn+mMycGAzE+JXd2B03sI8g6vqICD4805s8/Q7
Q9RvYQCBXt2A6pU5gu9eZBujlJ5yteDEmqSPNTNLHzUtnYMoAcOjjRN+mnEfti3CP2YaqZYc7AEK
EmGhccCK28g3Iq3fyEIwqSG5ZMQqTqoqd2RXD5hdEa8/QoSw8h+tBDysQ5iCskiecYnVoVm2sJ9g
EiFptSQHJIy0hyW5bqu4IBzo173gYuxltoA/x0vJsCyFYs77QhbyJAFsJLmGHqO3cT9lndY5RmIe
G2IsYZVzwYIn/hCH0vy7GSobNYDvEMIvGBaU5p1UTsf1zLoaBwNW5il64Rmt8mWVqr6Q4Cv07zk7
YKXZHTXhEeAgsPcWekKsDPhosTQ1OG/Lbmqe6Xtt932gr1mKpZC9HDG0zXIrXY+2oSE8WilO1BRy
J88nrrr7Yu0oYnF4wZWHuAWIyjgLKyWWX4IP/WRaze8T+DWjRzYC+x719Lw3Own8W4ws2iTfKhys
/AoSQctmniBEUleebvUzkP/54oUfgrmlSFnT+LQI1wpo2T+VfQtutqXZD+Q9onWKVVV4HeEbkZlD
NiZEFqgI7BCHMNKvyQsr+gN3d1+ljxpDWwjLTifh1kNDK1FTX628L7Esv/ze15vf2ojo/9c1/gl/
t1SV+B85OJEVM2ghrmoVc/L4ECZPJK0ZQo5F/4K6TFqIGKCvu6JvWCTXCXXQuvIJWVCf3yQ+xB28
CnIRjnpjYhPYNojhQfb5Zv+GZ7LFqZZ1/o78veE9yuWl0lUlNLkf7AciAMp2qc67QqLSzbmp+IIZ
GRPGcMLDzgqZMu5UoNLRtDcIK4IdO68RfVU+DfGj7azU8UasdLC7EXFxENSmQ/djh/0I4Ci41R+q
wsa+kmx3eYs+rFXPF/gpMof9+m7gcNIlaKRiKrmGwaefZwbiLS2b5ZrIZ6dIXfBst6s3VP1CYaaa
+z49NTCU0GqV80EBrXnRQ63CMSRECEHoQlN/WGzyaldjxjHPYO9Hmx4A4l37hy0X4CBEgwcgcLmn
2IaYATXcAYJj2x+86KLB5ybH7SyK4Ew14BYjahhIhbE/HpiaKw6srEVCnQJsybU/L8kpmLrJFJJB
A7L0H6rsyqypQ0Gw1vYRNT/Iq1SfeeCbJucKyPaC8FIIMxhLscoBs871BAGV6PnoCQwWlPdh7wt/
cV+rFe76p7fOp7y/iWBGEIZ3hi+nWA/1wg/Gwy2n5z+TL5zSsOLvSN/UaFnaFFlJfzsshhbbzRjm
u8HmR4iISYlZfg+PuCGg4qWDzTm+W3rHe0IKKFdTl4GXGM1/EpTtOAqbIDIWKEIZkJ5l8b15nkSy
kXA7m+xG+B2kCr6obeLcnH/Kll+3TvkRO20Bb17nVNUb9o9OAtuAZf0dsN0dkMWVbDBmARX5RrB8
Xaso0jhmy2GD0839FOGPRmjq0itlZIHy9gyGxFuelbdXGBP7YJlreCebt5nS69xLW/ntBMeaobHB
+fuRF9ZeLz6NIAjircenBW7v07uWGziq8CV4rmH/bVbBQVpgNLXkN8+irSvzIih6+uQU+4qnhkGf
6DPM1CIN42m9ynyzhboG0MwLmsmxfHNu6W7pdDbuQK0nD+bziOLzzqrXLBnyPXGnwpO2QuvUEpHz
JbvGAC0fH3+ZHVgO2K75xWmD0ckLOS8k2Z5yXiDsc+mex5g46t0h1hrH4Yyvs+xHhn22sZ5vmAd9
z+TAxX31wRoiRQvb/b9h8k+DfNRbYFTRb2ARM5f0wglZ2CBCHU3UDca46UnCcX0s2i8dCJiik+U8
1YIMvzM1YeyL3p4mMj0N+JIFkUtiWw2Iimbj4Zp6ofh5N27FA2Lw2SNpuIQppGII0um+Cd8fl8LJ
wmvWzSxiUir0Ax11Yq2EPE4jm3nKtv2sY0E6lx8WJYJydjXzqOwe7I/q8cblI4Vw7LJj+vuX/Vac
5mEUxAfQSPmHwmPnz7dWxElLo7zN511DK5ZEC8GBtiK9/m3RoIfI1+3Csl/GLaL5uWLV5jg3nmav
Y0x1hldBRI4gGM/8vCOKB1q8BY8TbeB6wETtrgJDpKK2w6lzrgVWA5wHTPjCuFeJZQKurXZeL80g
JJpIX8UxxYd+U6Gg7ji8gqW9cjciYoznCFRSJAcwiV6/RLQ7TMkMWTU2UPbgRRUhP5AJaTlsHLBG
kDpRv5sUys85ONbc5+pksLhtG+6Vd/mWvnomEBms1/e+jX8+Af6n98WPo67PSdCntlBBB0GpSw77
A58uptTtJh3ZnWGQRMSuQLMvad/WJZKosSXA1e4gAi8brVgIYmbIc2kzpFVAw8CT8ZJVQt0dh7lh
8tVc9ifnMjHMk7eBB/kSfTmYqiH66g/FPPIMThz2zJc8uB+JcA65L3cTruK5TAIZfFjQsRhDD+jo
+IQSPEMe5sSQGn6lLvuEYseLQbSEswNwE1xM0mWOmQTgipmdzDR1ApQU7CJ3glXHI7CVSZ+Ptc0x
tMhQKU+3nMUBMdbrbWczDZr8+LtuVq79gy6RjWSEvDiU8k/C2jfU7gvAAhYeQmEWA2ZDfrBZGMUe
ctwS4RKrBsgrdotouRos6i7rnUYet3BfSROrkb0kSdMZRGxAyAEEU/HXaAAC8PBph61GdBPOjY2o
ucgy4/5j59ePvr2AHV13YPvzcUThetgzbOE/iQtfdAyChyoVx/t7MUXlzDXK9YyFeO5akcWlv5cV
/tZmdn+0Ip2LqVVRXFEBSoKdQdXJdPtlxjfAelCI04ov4YoJ58o+t0nhwgO7bkbIx87oHNgrzQ2M
F9Nx7WUW7kGIwr83dm82aDD3MxmSYxoppKine4XFBSQuB5OgrdtAHhsoSTFIgdLrqVtjPempXbGk
sAGCyeTTFU5G+XjRzr/5F6bDtFizNprxJBKDaht1ZHz7ETvgFDqUE1wXMVV/4EQdWo3mWO3IzFHy
MHtIRlXUch3GQNXGHB3VG9FfABO63ISUv+i8letcphRuJGaIqd6D140yb1j9b65V/pllsmcXjxZI
Ah43oD+OViZ853FMzqnn1m6QUPSsMZIRyqrAz1NPtluN+CJrw1FCZVpiTakwpdxU24wYPLdzkJVt
MpfNjTp4CfPgAm7JSZ8uNwQriV6W+lMhO/nOlWDmWdpkvsTuaEmfMCDUgnSLOZS+lGvmuwQqc4c7
zpaP6+TmfafMbg199BGBGKHnAzZYORNMzqGduqQH2rfIjXYsYhgEvrviZ02MrjLaQZP6+Ut5Alf8
E/kL+HVFFRph1szoSkmJ7EBXybrGUR5qMCQirKzjN+9O+mZGlpjLRjEm9OvwEI2YBAdnbEy2PUIS
EppQU9iHilUApIhfes6nYf+wBw90smvQ+ggytyPZpyUuHI4qtFg7oOfeQJsHmMUTERb3j27kJedP
2tYr9qiiRWvUkdwJ4KJwqWf4pQgGognpwYEamf+1nPv2wTMMQK8Xx/yjdn10Y0/KWTAYXLQMmYjz
1frZ7sNr9m2G1bncTeAGzAAYatbj5nvolqrKxgG3z0xhGVUVc40Ki2Nepm+7jD8G0IY0ml5LLddn
YbZpN/8M3Qhx3Xq5oGiH/2TnC8sMX0iYn2UCyLxrWczitSRdquyZOivyQrbiaox+Q14RjH2RZNd5
aQF0j+++AlFnkxA005oCTlPjkpfMTIc4RxeeLQJ/tOK503oFkgsrCogo+yF12lnKy6igucSzbMPn
3Wor45sypUNSbvvkuBCYT1dqOqZXmmu2OwrJxxib2arzDMD+Od3/2YCFIL50cnXvoIjhEB0DXR9K
/K7a88aV7qbJ4DHBzJ3f0XIdiFQ8SQgz7J1rbVBgheu6FymoZephdjJLqZb90iDDQWVJmojtbzXg
gFOUIz5M7rwsn1szvg6OQvvyk2BO7F4pzU/gosxylIy+ZgksSmVFg/qaV20rZ1k+aSKwrFaoQyeZ
RFL+1rHpj+IbGKJ0T6azxeZPrSBdULXO4GIJdvr3Qb7m1uZp95FUpJBDu9qVsBeW+e88fCT6V8gX
VS6NTuR49358rzHdu4P84iHiJvQ86U9hTj3lb3jjwQAZN8p0kHLIhJ/OK3HNXw+RTjLj3vFhUR/i
IRh025GWPgCvLKW/Fcjs6l17Yf4iBubssKiYf8wlCs3fcp9iubVKMP7pRHwefSdGrCymu6kYmLgw
mqeCa1xHRtdyJWo9Qe40/RZF/z5wrG4kAL6/QY4JsNK5IuaqdL11AZL2SCSWi+If9d6xMChOcgdO
Kz8rL/ul1zVN4v9usZdnQoWuT37LkO/XTV67Fotcg6wt/2SklpnESLjZ8scuc4uMPNBaKqJxjusu
l1vSBAc0RfX+94qdKAB1kZkl5L/0wR4MeVpy7u7MCHssLTOzpzCO9upNisBXiFFPDC00CfVouYZN
XXF0RkU9ILKEeChv27SW6Gi7Qy+jku7OC4OkwVTtOeSe3uN21fa0MxUAVDqDcSYih33eUdQ2UgQt
L6AkF4QraqjCQmkNLaNY6/FADaaIph2sC0y2v4R6EliBhBDUC/ueMaaLEicWDYdky6CenbfyuZOC
Uvu3Y/IwIV5G1ioj22TVv+/LM2NMXlM3efeBXVFLlpk0glMoySXNMXgPIwpcUbWKr9MvEuUqvHfU
Ua+EPFCKPWY+MPtNhxODgEaf5SD42ilmAXixVxbfQgZT8KDy5ESHSevUnG4beDCiUOx2OxSZYEd2
WecJ3ZL6564z/G4fc7Om0ZIOU9ng5EgK5ufct/8wDhJxhrKfWKF8oGMAz/NIeDg+KDpnnOd9TWC8
m1C/nAlPRFVJESuKzp85N/iFta4ERlbMXC3KbBhJx19efD9AzC6BaiST96FqCaEQ0gbAZg+5M0vd
sd4uARkYKVZ+saEmK10NttpOf8+fMTy+o11z0fGYxK7evc99er/Gbpf39qG9yEfmAEVRfphmZPIn
SQf7u15eABhrE65ulYC9cW/1kD9cckhW3Ca6Fmggjt0dr5f0xyY9FGPQPcKlXF41lN5BHyQxsQIA
iGo9RSECpzORa/a8M6ZNFsEFb1RNk7PIJWUUTwA3yGJ86kp56QxDSwHJ3pphqBtvncSbkJA4qxYe
VYFrqoPM2y9CnuLtBx77VYq0P4lNlDZj2jk3mHJrjUoyGQJcNWMrbXeusyvrDBumKKKJuoCp8Ji0
/RMJ+8HFg8+R4uKqYvpIJg8NyYQ8vYA5vtYccRW0jvZP/i0U6PWDFr9Jttd7mvkTVOZWVQzQwIa1
CX0sZXUqWjeUdWRk0PgpbprIfHUzRGF/71Zzu1yRW2GCnx767EQ5qKMpDIk0GPjYaqO4xoSoi9aM
1yz/MP17scsZFRtDTEX3mlGXuzvOXzoZuF1pv+cx/HZyvxTWVigsZvXDBZjLh/wgy0creA+fBV1k
8fkV6zAuCk5dk5WqKFfYd+1UeCPMcZKIBp4CT4CSOy97C7PdZOfTtjBE2N1HOoaQ2ZxOQQfwlT7T
fBNkY0FZvjuckL0I+G/gCuS39PwVULFYbFIzpXBM1Nbej2d5BRC9Qd2AZu9sxMPtcZKUu95Tnwhz
RLTAtWmI3jpVmutYnGnpM5mKwhhOdMO3VOC5v3YpF592DzT+6/6Acs5ks+nnzpA1Us36PVKcWGkE
M1WjUqhQAuy5AFtL3rF2Roudc62UHxBXUcrRUznmTU0m6HWy5ij6umKW8aSGQEAuTFkgHG+/QK3t
lkny9IyYFmqLI8pYvOJTBRa/mUHj/dj/6NbKzslOo2YhiygO1nVPUAcgCQY4cgBaV1HZAFPnSrue
xDDcyoDCQ9XAq7HtK2PK5zi3RkeZ2APBYNWexQi62G+cTV00wfk/mJEXllv7M1McZl6EYNB7w7Wy
NSFsKlLu8YEu9N+Kz6RKVjxTNxRK8PL4e5PF+lnFbOzA7pjA2WZ8s4rN/GBsDQxj+iRTW9eFFwkI
55pwh0HyA5SIW3FjpJUf7cIrlGZ4oEXT7+1t1T2BK+cZECsvU3yQPWI0wujjI3BHqX2Avcr6Gfjj
Zt/BOCeLm3WPYbVnr5JtETvK2x7GxSyH+9LMO852zV25Cd+48P/c6S2Kw0ca728Ny1Y6KGbL3qlP
4EvN/TZ7etw5UKea706IUXwIQVwpP5jQ938y0oHDYwffAWQlBszHIVreDFPDhRH7grduFfXwkAZq
Xg1+sBIztw+hxqlMs53QCz42G+g9RWycycylepEsvcSk9fVNm6VmgeZfgi6X66giRnNJpU2PIBAF
TmbPAcrMrGqiw6Igp/NT9dLv+HdaubjRbMktYivcwKhtfvRJxOMuhYot4wWlUUavaDQbJmW24VmJ
ZwCVPPi6rQ4Nhst/OnX8HNiq2U/gTHWXorogGqfyr8Y6nwQ1i/rMdmxoA7b/GE1m9P5/B6xamFQg
EwXo+CxJrOCPsGlEdrtI/EomayDvxVj5CfvkkF3AfbS1sQsfyGGG1tUvsuzyG6HbCWTS0DgHLYKw
mLw/kac2HudY+pRGugwjN7CsZhMmmjhzcrMq0IOLuASVzEQ07NRtu7qYo3gXq8qnNgGi3DQKDYrw
SYfT6Pwt/XDOLV/1Nwm7lrkBfprfCHgW0qbPVabJczWZCD+LcxtBQw3gU2094NvU7pb7yPhlgrq0
cS5wrnWHRgkSVTP2nTdECUOf2uvdv6UAYuKZB+WHxfuNgMuJy+NNx5KfDuofgKn+lYGw6REYH3Ka
ZOfYztF8bAdIPEvwSawpzhGQAiNBWeC79fEj8BBPy695w6r/wK/tqaFZeWkyTtf0I3GsKFAFjoZf
KzKY+NxdAAJi0qPk4lVk75CJ8kptfpPfFywJQmfyBb975TcM5vpsuS0OLQ7PPrjlQ3gHCKvA+H4n
QPQpKtQRoRv3axSt2d5bX+nHX7sDe0XLK+YohWnf6W2r8ED9onbhdOXu/KX2OHKoCbv/dCpO3JIs
yPgJIlcsES6Z7VNPf7AG2iCOhM8IJc2rkfWNF05kCosrhh9zj72ovE8RIohjbE6NHLiuUlA8oede
e6MJsIbj7L6BcoK50YtZJ47mkqQ53XN8aAc4J/rI7owAq6S9g50tYefm3L0nPbuCGWHERzd2gjBj
eixz+xrcNM7tnJIQKf3BHG5GEXQzMr8loXRSFArDmZxS3+X0oRJlIt5ZBx6wPaJLw/47C403FaVO
IQ7rKIj1J78aFfPu3+RUWyAxXdSUla9IOrNugivXxl+/pixnEdfqFhdGh7sINrMDr3Gva7MydLld
aT6Xxy2ZXoCIrn3QUJYKAx8iSWuYEwP4DqSnDEcIzqyptarJmsEalMCp9GrYMqhCwNqKhm7QFRVH
EJZYkgW+8UMhys0ogbrtFGbOrQzAPtBJbeUFIniW3mJQMXc79i1yiE21ixQ8ixak+mrYSNslA3e6
hUZFTZJoh5xpuHQYY1nBk5twjasanafpLNUSwBeNbZ44LL0/WMXxVmEI+OffB5P3t3OhAtcLuUmq
dmfqUu5wfet7GcTzjZMame10OMV+omk6zhW4JKpGLlaOc5wx6/zoGhGWuaT+cWFv7j06y/IK1Ge5
VwYmkjNekZd73ikRPgWbiiTGW9uE4WwlB6bawr+FtFUk26pt7kv3iGZfcaexkYk3gFuoCjMatcxm
5iJBYNcSz8AWR2X2L+XKSxtSf0hQgxgqoTL2UfsFHmKChrS4gCUThdVlzTQXUx4eyHaIJJH9DnFE
M5L/7tl89MeROUUOeAtes3QIlHeFFHBL/Ji3cfap8ryGMN1/gtgWdRFkXnoX+G6hQhXwma8qXikA
LWFDlKPRFEnz45o+6OCrGzLwe/otDBFLGfQ+GWVpN0kV/uZQ75Sf0e/PsUXpFnaLewiSKank6gwi
8yF+WH1FQE9YQ18xUl4fwH8mizCAxcpFYsA0t+RbSUT3n/4OMU5Qp9o7PN7lBGRIO5p6cMtXRnXC
JfW5MAwmEbuYLebmtXFTuJDEJn0GyquYWPiwpRZnv1ziMZpHifvHl8+OztIxJd2mYoB0qILovXrv
p+sSoT6d+Qt2nOaFyPi/m6CB3U6EZTDb/lY9CEtizEw/HAA/6VwkE8uIX7K7vI/hr2H0tduoiiNC
Z7Qlv61NGDw+Zsk5lf/EB3d4KiMTGGR+U3OwHtOnm6VYC8rcu1iaHeniGKq68Pd4RNabdW0SEWBG
SCsEB5twlwDDXXKD7ZjGPdrzFL4xeUQOh7FvLbwmC9sr/yhddMvrFkA2V9wW905QTisuA8OW3JSB
AUh4iRU5p3eIXnK4bV5DGLg5qrBMXKp7ITgTUsrz1GkN0djgyFC0XYoOcjI7B/yHlOip+3I0y4mv
lvXPbxrefN6gyKaXEaeKqc8lkTrapgWmcul9IqE2dc62oipP4yfF9dyU9mxlW10geK1g24KEyzGo
BeRphtKG4Qmo+nfR7liloRHvowONq++DWCDl7U64lFtPGM8DVJ8L3f2O4dZ63W280QNqOHfM+D3v
oYV1BCKRuIDzGPh+aSQpVALS7SpCpa9vz5n7NadTJvhdFlHr4KfuJX3Dh2oImi+n71N0Qn84euc1
fOD4vRyV2dyrbvpf8ZyzqYuhxBpx4gleNeoUIVPfagb2FoQQ+bskrJ9Fzaop3uYeyYjVHHz9Hn/v
kD96iS4c3YZAm2tkHGVHg07+rB7CjCZASOlDUuBZBYy/Vf49Oo6ZIbyPX6zKW1HIZX6TCXgL2RMD
Z18i6bS4dVWdamjHoVM2FEWy0zWmP48ZzqIofGQ35eZ/S/W7DX9ElshVXWSoz2DnttgcYeQP85Uy
g9m+ziCUZIcadRW964AoRUA3+eqQFMd4s3bDuqBW3XcuFpHSRPXh6t0Fs16Zxakn48FFt53gPuPn
kWccmrUbXLvLcqhA8NtpSsiryUclKgessi+7wqGZwaOZ/56iVBpZqOJwABqb37gDS4naRX5Lhm3s
m3HaTaYcXMsCHqn0auTQIir/uX4q5UPZFQ8Bz8UC3UKxfj5ULvWsnpZTirNjNzizmAgQT8RVbgzU
2G5ppcdSvbuZsNpQGRd4Pb6lyI9TgsK+1nbLlHGhemrdiL/34MiuObwmSLc73QRRBxNgFET6e1Lv
o6xWN/l6TErNc+6EiEwrxgHsEDYFHeG6qnW1ueS9Lpmo4/z7e+6wy6Tl/b5WouFHRr5e9BLEbuxz
42BX4dBB1w/PfHqyvQ9VWKQ2jLS19zH4agGu55yMenuP9MgLtErIMJT+Bl4ELPGwB6MlUUqTZB3t
VQC2OppjbtSjETZroDDv09xkwKjiHqEFViOwEy3sF9EdAetnX005D6kuc/K3fTbQi+m6fMRiKN2Z
BiUYhf8XENvED3ZMQxboABD11DmJ1e9Fs74DiyxWCij5drQwOkqqstt1vqKAB5y7Yfz7BEDaiFt4
N/hwftM3GyDIag16EDHX9KUEehn7+WAQVjm8M9q3X05bEsi+YJzDYvQ1YUMmCywjgkrU+we6Zlfj
jwHfaDlARpdR7SkNfEHejmsi+v6oKmporsGFi/PV6Zto0tsGqVmsM4rG7ACZ9Rr67LZv2ZBYmau9
YMgEVa7MgE7o+XRH98+6g76U+vPo8sDSXBzjLxrUWj7LbaLAwHwCiaHAk2NE6S11a38XlxU9q4Rc
V/ZeXX8H7FNqwpWafLtSUSFGjVEl2UPuR+LqiFTtg5pDbXTI3RUZ/1FTQXdKgs8mgkiZobQpzFE/
rrjhpfu5U2VFgUt175KUgZwXZkH/mSNkaexiOIwbfcsZBAy/tKw0ZMHpRgmxVxs6aDNEnWMppYML
mirp99KtxeiB4YkVvhoCIgRH9rd9f8SjF4hpmqeG33F+I/8aGa/B9TDn9mIOB0MkA9G27OhNWHti
BhiDpachcuiKHNRXtROW2tZ6QSKltulLhEE2tKS5ySwwxUggM23fjcafEriJsOg/75JPoP0f7KSD
GKya9azUZuLQNLPDToOlCvYyOgxC7DwAJSzAineFxmxudrjNaala4ME5f7ber08k0H7a98KpnWhr
7Wj2/ZJ+vEdRg5LF5JobYzKvmpaM7hGgOO0Y0TDtIOO7HUt3HbEwZQnXW67gaNwbS1SMvRGswaYx
K6wkNU8q8NKtgBuc+BLolYfLBZRJcyR4yNDpU2ZjHuWIT4ts/OFFXInD84SDkSXjHApALHfZxsnt
cTfPbSH8fDmCJm8Vuoqw1xgU6RGcrAVPTlI/Bq6t7tCPO+YaS7Zc7owdZvEsNMbqoZsmDCFe8doV
8cVthfoNVR0f3SFwHIhWyLqcudCO3w5Kbmclzjof/qugz7XI3W4up1D76MJKqi3dcnruoFlabFxm
tSwx3GSlL+5B2O2YixhTq2xSfw1sszftRCihJ0NMSoRqkcjUCZWV/isTBo0MmbQfNmdasTOjZ7ew
2BGPXSHQT6V3s6XY14QEqIGMHPF5erZNNQZhY8yMaHagYfd2U+nuwBd7aS4EyGQFpNTw3QcKE37V
hGX17EZiG8Wq6MY/44BXOfTCtCeKo/byhuif/pVMsu+ca4R5zGuY3CiVWYEsPvzxF/qKifpxZi51
XRmtFk0dvxCb9LZijwdOxnyH8ZiWDHs7mJnDVpcWUMPZU8IvqumksK95mbWFPl5LqmMFM0jEs8PD
mTfV2GTjPFDNIyUlS5wgr5mAkFV9aGhFTJyxgym8HJTFTPnH5yHrrcc8JJLtN4hU1di3Xn1fE3uT
opoRvS0bdUapON9OlwVhd26jM7wCZBYB6trMJ8Mp76myBkkv39NINwvcNz0C9PjTC2KxxPuukWtR
w/yhSCjv3HZENtmeUszZgrIUGEER9oAiD+owYoWYlewK0ILXabNAqrhmEBqBHrr9oqgbcYRDzuYy
tXp0TFqhsCtk673OJdQGB6Oio70EYcvfK2+/+lQbm8RY3MMrGTIdFT56B/KY7jNhS0GK2TQxwqhs
TRZFKV/ZJk4siqHTytH15d/JDe5gR0ZT6YLiWctRZ0o7rDFAuWGOts2T5plZkYkKlicuij/brRUE
VoPwjXc21Asul2nGZ4oqWITvNNvqsSj3pZcib/NkEb/ywxjqeutPrWHdY2z9bYYV0afl6iN+OJPF
mRYM7kLjlkifzhHkjMHeNI/3PFm0mygSZsjtHDrFRcYjNY27pFqwHt2ydv+Y8I0N1SDHvn9BLNJu
oFVKeuo90KYeeut8r9DrRTYqFOonG2OEQDDLAFRufZ3qQCoZzCVAz2808ZTxpmyZlUrqqRB5eNoR
fjg1JW2zKpsRpYXTmNQeMRdldk+Feri5oq9cGD5YRVbI8qXrgCFVgnHaSb6bgNKjoxu7ljGDhDlA
fyljqWnwjpwLnJrnLEEPxCA0T5/et2QButOgW3nnwmS1l46RTyIuJvDC37QKPJAoZiXW3NONxQ4S
VMkIxUni4WFNp61+I8ALmhKWYBMnSF2olRUJgjx/5EoFbnaRnuG71h4SLeOPIDGWQZc0jBwrQoy/
p39/L/g1wLZ3FqNDV7qggQZ0GMY0PqS78funhvJ8e59DeuguR3c8Qw2C0tcThu571K4wpX/OFbnY
beeizjT0zdkHhRSex+8gBUGhTbaSXFA+qwXR9xCY+C7zYRTKO8Nx+cPPqtw9pP9PxBswmjqhEKt6
3Ck/ADyCLZdGREp/A68XVGVvHb/JvfOg35vhDTnY5YS2yaSxtOlTrfweIjcpHNm/KYIfyfc8tE37
vQgFgsHKTN1WfK5wTNKf7aRiY0HC8102JHI+A45viX2RWjDbdLJq2Y7F5ppx0BUGXajkekHFHtTP
zGH4mWnc+ZM9cxpDbZHg9CWY03g1SIePCaPv+IQWravG0Y5/FjoT60o3H5FyFBudgMVZ3cp8VzJe
LvD1NXLx34aC55OogymYf2wimfHqDswutWmnj+tuNMEDOInqQNq9UcHM/OyxxtX8wTTT/NRUFeVm
VeKtfofxOPU4GgEr7q/dgpmmyUwpJdTmUIWgEo/EFBgHOpfX6wnVmKNZLK/35u6h5zONTzL/dQna
H6zFQ6I+cQKT5ug+al7l3k03OO7iBB2zXBSdPjOWpTtDodnsbHMw86WcpUsjoqFkiDJh0K9pAiTs
yu0YtLXYhpLRc8vLx+nlNPLnBlewheD6Rsel2vUITR+Y0R+LTIVcFizL3RkCWpgT8Mv7GFBus0bs
tXa7x74NoVvDOv16dK5Bp6co4kem5MjsBMqulNnb5qAiSRSAHjJVEcbgiN/ejphUzKhhnQ2rLlmR
J0srKz5SDkt9GoLIIQYs5LiQz7IybWCgpgj6AsAgzJv8o1wGzGOJFcuutKhU3byY8gX4mvT1mcoL
+oV0fltqMUZ5+7fYGYXRzx+IoKYTulFlekV7KaIy6pn9anlT85vVRhfq3tNZZRGuUALVSiHKp1Bv
hSH5jlo6taMLCDODPF39Tqvftq6OemOjXklUiPQyYpE3hA7qrG4TTmxYZzDSMPUrCpTcgg6vjYA+
icfYFMU1pgr4fLmYJ0fROfPHuGJh8j+aeRnjdDL1S9T5mRS4VQFv2nBpMet9lpa4++KbevKGFfwJ
BO0QF4h8xYmLMoxmJE4LfilYtw9dGxV5baelDnfq58HheZD2ds1QdE7sNtEpXV6y/daqe+F0IrwO
EggItvtulBViDAFHzzEs4Ors+9e3U7TiRkh+FQouUA4zwFshY6xGA6Dbnol3ZBzdaBUiUM72DESu
4f8i55WEiA1ksZPV3YoWd/4fFxoy40yp+YAThVsC3PUgYwIJd+HeGGy4QmzfwbeK+mDAR9fhkgPx
nzDL3LV2Gv3HmCCLPBRF3HWk89YHpBOvD6r+uOVfqkM48561HfV7l3A6apzVHxEOEh1IyTyiN4f6
3KVzCDqCvavPKeaSnkFs20XLbL+sYELy1lix4/B4BOvvSBa6muSI5EwkO9IYHRp4SldDU/BoT6Cf
qRS1nv1bScZ42MttKPlYo5C+D45g6wpNReoA61TtaIEPBZNYtLw4TsZyYTF8v5ZzdClRynhRzcCS
TDxMcqXxYDSNoJqUrB7zcYe4AU3uO+Tj6wXoA39LLbsKtK1EY16dK5eicLPwSoFRhW+yHzcF2R0r
WPJGyuHI7ddZdu81doAYgdtje29f2PoQ7UdSTUx5TaBtDIJ3Rj9hzUirGokvUqbl7/aQny41+3XL
F7yI+f+1hfB0KztcysNAoH/Ef6mEeMnfNIZ1MWfgKXi2mHySkygQ6NWZ6vvA1E4qyMJXH6Ff48/K
gOLCxf9q2hiWqZQnp6Xn75CfUcw3BVuhzDPyLdr0RuUnInmBo6zzYXmuhUgWD3UZOwbOLMbQde1E
4+ppigWbA6D8yjjDH5d///Ez3Ge5UANdGKtn5+zwt6sVz/UnNbLaIxHavGC/XYYHjVzK8UBa1goj
rRjxZYq+/vP9jTUVM/We05Tuu6Vhr8Xqgqbs4LxdLvSY5ZRtfkiZ4ZCcUX6PAd4EH3/mr2iiXXwk
MaHxtETB5c92jL0MYVhAngHcoQp4PXcVgMM53uyhUPz7f2ILQV2YDlsJucEYfDq13cpM0FlEQd0h
5mhrSC7d1cT9pzwN/S9h7Qh/HzA8ELwUmuPuJDo2/TpqVz3rFrdQd6zrjucPEC8bNXyMJ4KKbI8D
jSOb8qPFWrNmF54vmxSvOh/OuuWoD9f3nVoFgkV+u9aHOriGCvKVf9fo+9RKQjPtDXcFXUfhU3Cv
MzmWBqGndqHMPSFCJwZft7uzO4LOPPH0VfFoxWhRynQwCPBocMx6x0YUJV+M3EFU6Vu7E3kJrFsl
y1fn4yO53dC25b8g4zcCCiBPZyfjr/dEPpI56AfsYVso/JiXvsCGk4Q44hgxk7E2o05UqQCMycBS
ygQjxTdflOik9YO+XOKbMzwwOKB9IrJf7iEl2lQF2K+TkGRUH4+zgS1JhcVqHPMQR+DJxVpWfM0M
H47wPKt6giCxmkkimy+FeHTdZ6hz+24lzsFu3UbXHAwWbAtim+kz7tWoUwDCuWtRez90LMVibV03
s9OTE0S01WDnqkPCfv23N97xtDZeKpUclYjzfg8WN4IphB+xKA760It6EE+vAg6sslhPeEtILCY4
Uo32QdRhD4sEjjub54P8JzSNxRxNbgJXU+8ynehszPSEyuxl5dDi1AscV5lkhXQ99VE3kbMI8ilh
QVUy1qYXE9K5fiRAV0MgOjL6GGRYoTf4n43A3FTs90xm2IHT/tG6dfy45aY7VCkDyOLAsNg6qbjb
S+am1g2mbZSI1nM9RhmFc/sBTe78Kgm7HWfCi6EV9WsWjqKGa5AaRsASsm7bd1npnUKXCxM53zTI
77Gkmb968Gfj1eaXjJQdf892eoN9RwJPsCC18O81xXkHoHW9rpUzV/NkTfGJToNKY6n8O/U/gp3y
AG4NmQb+ohRjIbQrMorHExbrqsFGL4eC3yc69mOV+v1CTYsqda7U3Kustm/djGTSpFqDUaNUmNv7
s59H+WB4s7H0P4v0ac2cjyGb2JiekKYXjqytCQsMiVJwOtyNM7tOjPKEr5DFyVazHv2pRLOhaGVG
87WLyoRqDpuHLeZLjrkoa33bl1FYrCa3J6+jJ7/V3xNnIZQChJxZvKwYAjZaE4fMV2ZZJnThqFaV
jzThXMsUKhts7V+pxPK+9zyGMAfbJb+gqTodEbZFGJ3uAmuFe4/D7u5r4ULee1EtBh9bcw2j+Ola
cNtHZu9ufBxtKXSETdazieWpvDhS+w9bsCl/1kwyTaNvigZTEXWAX7zN8t/Lv3wG6d57wx/BxB+E
F8OAUdaEA/l/kXOG0XbxRG2wQEbzuLgDFSmrE62VEjJinXmf1q7lMpmlsJOGH0t6Vpx6OC8xz8e0
9F6q/ODk0dxRYn1TlLWz5oHLnk5CLNiWA8DqRrYx16q9uzU6zk/7a2dB6MGsTzhiIU00omSXkLY3
uhJSd6oKTQspc9w3uPCrB095lhsz+vGhD4iM4/CS2HsS0zXvKKDnVX6r6sYwhAYS1txJn8cHejTS
33a3FzrLh/Lr8tihbnmzdHQJtk+sq7tZb72rWrEbk48sbF9yJahsTCRqNmxxIiHoM81CkKoI+Lxh
cfc0D5Yp/MomiNvkLGAQL9gJNP3W0OyucO7MynZvbq3xjQW7UGuTkM+U7elqqbUSHoc+YvoRMbS0
Wra3OUa9vgiPvfWOPUXkCzQ+GZz5oh+zUdgV9KFSEg78gDsnyyeW/ilBD6TtAk9pe6QKH83lGlA/
2bWItSalCQk+8HJxYzEowKqYFGa6IaIc9tMb8mXj8fSJrYpmGSaaPDJJbiFsHkgzUgKFO56A6/eF
ldbJbZmhU48DLTEq3y10q679uNFxpRjMbj1VLTSaUJ5hhfLgA9jgL7ku8ypfmsyML/AFtmtYlAYS
x/hfNfqd/HxrFDj4suOVtrsEgFli/p8rQFuk8bUKKi+qMACYCmucfH6KPKuWAuxGCuqam7J+SLhy
F6DV5jjns6q2TiCqwQ/SFDGGwNWkiXwsljkpcugaJxrggWO350nMbF0QYxh1wDeVmRmPTvIktQeN
C2vym6ToRxoNYTF2Tp4Y99bkBeDapsuHhs2C3sEBcQs8X6JL4hEvCnkrhPhAFYDvUWiWd97v1xEF
JXyVXUJkVG9BXgkFfhxRC6VBtIUPWaRXjsqkEhgA4GfNh9Ato1kt2NsNy0Yk0TuxhhyZVCo9JfjN
xOUbhJqEzzlTH8+IdmNPKx43EGDT0Lrsk/UOaUPBvFWdb3GqIMg4TchPjXgWpuyR85DLNpqWKB3K
K2K8dzks0hfLCIP0o1ZrJyaV6vTRLX6GDJX6JZRDQIcYVYCtM38a642Um1FZz9czprkChHqQfL3B
NzQrdtyK7LIW3fUDo5pKTkFMk/BrlxVPsmRbDFKf4rxCbgZA+dTNUmlpBauC7VYTM5YFkM6wgAQf
kvhXW9lkApSLz8wKN03C6wRC66r8yh/YqKG+OjTUsFovJrTDokQK8MgWGIzpNPRCNORK91DK5GNY
HEXIaZzdLIwnRbeaVleFh1M2/3aFZkINsBeVqebQim1r/XodkwvYfRJymSowdoWJn6/gXjWYYZGh
nHpo+U87TYAoe/0bNSftOYIRvEYmlBQPHk/YuQ7Jdb5hXqiv8iaBtaRv3kWfgGc6JF0PyuLIJmQz
sePGBoxGEAi/gTPFAp5q7bYdVvVh+ebZ1KPCkgVP67PIAZMIBdM7ytHOVT5vyhBUSnzHGj7tsaK/
AqD6UoWrkSts4FsZnh9O4M8pkE8Vm26V8YWdgHnDnz87zqQ/CBdX9Nf6pLsk7Gm/k4IQqgnaYV3Q
djGKNtk3QKG8x7u/AfFVjfC3uxos9Lej1HjxSt7yMGU5UStm3a89d3ADmdllSmHXG8oaJwgC5yD+
6ZyoV+S6O/inHAAITWTqNss+CZq3wQ2fSPRm3iMIYujSFh49ZWF6Y5hhATGZ7puV05IkX1gc8Ela
qcxST2cD5iqJ2QwgOpu3pXIdq8sop2UlJ2ii2/Ct6PF84r15S+LX3gLwJ/KnCGF+GUwOWmRkx3Hu
v4EWljx5OFiNNQjpL6/VF8J8mZgV0Yatyn1p4Zb53UROPaTcM7aRopMguRKwhgpbxYt/+eTJW6XO
DU2onCq+kdiW47TN2oEGrRxvPPPOq8/oSOfJtP28+4j2QIWKpNEEkyM1waSHRIK9ySAFcsxROSmZ
y5VUaZHpge4mjt4o3wek/wS6MwWVPMsAu3hEPxAU1KQr/u9URt3MMa2fLlo4iYegrEEYe2yLrrAN
jfOlfFl2WAfnBn0q9dqaZPhtJGkjLcv87aMFcrI8E5sRxgPWXNHe5E3yM7fFaxtQ9czAwy5HBQ7T
gJgBJSPfEfU8e3x0JPGyrdeTDJ3A7ttFutTZr1mNDvkDS1bKipmWU7JPSOW9iMIXgy8z3KaMV17o
y3aq0spIkFtfHwEMlx5tdEz8T/iwPwSqX7cnQdq/VsqDUNNb4SVzr+cYcHaGI1VbX/0HzDuMomQP
8bBDfD6NPr3YWlufkhrsbQfYW7WwfFtn5mraBA8+uYpAnFvNL1nN6ushsbMR1N+vSXjcYN5NACl/
H2124SzQrgKMKsLqQRU44LOU1vbHbBKDecnaquvebNH7p2feemLLqYcfbhQerM8RTzfGlW92BjUa
pGu7s0UvPCSvVvGLI6kKWChXl/Ug0dnDJutwDJbPGIIKIcK+2NPBDWx7NvZcgk1vLArNWzWWN5i0
Z8dDhZ6CzgsX9JZYvHPLyXwjLrgSDXp6EkJ3xaVltlxsSPjIWuSJ5UR2t3a5j70+y53DA5hawRIJ
BflpJHyKmzPzoIY+XozhC5geLbq+MLSTkXTA+Md2N7j1po0WdpbtlNFxKyHKeOmAG5tXoFNxuonX
NfKY106GmQh1ErXt/sv1FnwsfMlB1zi1P2UI7BNRKZFKqOrCBbJHJCnZXGXx5HE1jHd9qZY8pcf/
raU+1iunjRWFwqi0m4Q/8gbHQTiFqXI0Vta3iD7PfOvOLzc9cuejpa4JY/ddtS3kX2TIpZRySbii
XgeFxsoRZG/o05PSNLi9egYTmlUgVS8d+uK+3hIvzh7l7GM7KBHA/q9Nsn2MXkbuM26NH3qxiAea
Dn32PsY77N/kRaam/N0h1Zw1y+Yze0k6Xo7SvXAa3PeIHINvxYjsqA0DUbJAr2qJQ9ez9vPSqTOB
Dhbd/08MfHVAhXHpF3fM+00YOk9kcYkG9Ri/eeixt2oEDZaKzJLnnoqvFxeWkGjVuZfdk5dOu9v7
ExEKEHZo+ZvJiEXLjjzmDtZFould5AIW+q3ME1xdRFAo48yScl3GdhltW7oIIwCbxONHp6pPH1DB
UKn3Dh2Z6TWDBMdTMe2/L9TS7lojLF/dKkQy/l5IxcOXSsyxUWAVpL5ZrB9DtijZUUpLiHlAFei9
Y9Z+k80OmqZhY2yO5s8R0ALs1Ft48o5GjKhCgHF72iPb/y0d1jf95FfmUoxwezzrhskMaOCfFgg8
AphxbFX/k+52qiLuQkjtJScwGnNfZDEzWfMjSThKXVI/arwQ7Tn55JqubDkyP18b3uYJ3czC/KiX
yv+ED9+8d35HV+DzUtygwZY7rrisICcU3NFk7cc8i1jdolvkOva04x34YiSWT+zjbKj39iDgMJfP
nq1M1Ah0h3m9u3TgvvOjbzfU5dUNe5/RyIdK0LTLLKGFZO1jZL2P6ntEgfg507gCdVHVavN3mTHX
IPwxe6Y6aJ52LnrwSvqTlTplUK3PXqyywVm3ukSQ8najZI5ITtibqu8sJzJxPESP1h/CGEy2irf0
tKuFjzq4iUmlE08KwGR6AdQ90uUyDZ7BInDpap0TUFE2yqj+Cmg/RLdONz44miMbIJ+DAxSUi2MS
CVoaEGRDgZX7L+1GCwlSyMt9OauSexn2E56pMGI/A/PNjcGrIdxkutQoK2YRlg7i6f+wNb9Y2gcM
YzNWLYz5uyo3rNjHRcKm7HEbiWcCdoOlOc1k1c55wLySin4bgMGuA9UXa2pj15QXYNFMeJbtfhwm
ar4+eZn5WyZ6Q7DhbN8CKPpHO9TyDPvVgQmrAQcWSBAx1hC6wirnvf7ATJlrz+DmfHI9E026mId6
KH40lG9jMqfrWu7g7s8wz6nIBiamEhcd5objUHUEmMKbsASQjGVhZA6QbCbgAukMJWUtjQs3kGXc
FgiOMoJpGeYNPE8MJgGTMl4eB3OVuQh36cD5wqXzYC8GP17NZ/0WINIk6TBXOsOpv1WCDSwhzshP
zuOsK8lBIWHJFZMEZp1ygQP/cGs0RyCqkD8ulUBTV+K+EZcy6DXjw67oee/ALKZrhgkjW/cAGZxd
eGZowjoQwZjMCPMMu4WX0cMnUwzIo4hU1IQi+ktIpNRZkliY3/li31LBpNye1mMA1I1p7/jq9Rb+
No3LbhHCont+fMEy734+6OiLsjBXts+/ro+qRqYFtjyT+k0RFo619T77Yp2untdxkjuR6be0s93j
vPwKi2VrjYaTCJbKSM0oj0YtWmM4nSWlNLkS2h2rjbGdujgcDPlU8I44Bo2G1oMGiCui9FodkZtG
kOBqtjbv1R/z+321jpGACzq25FPJUSd1xst7U+0GLp/EzuEpptq4ISk5nnvG8OpY7afVlV5aPFsj
MBQKt8uSzd/dHgxVjmPeqp1cV0WABPcaLzC/ehxbi04Q
`protect end_protected
