`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
G8uxspDV0QwwRW+WGxQnGX/V1RIlMY83W8ZpGvNjJU7ZtYxlCV6wsCwRGM6KBDcABFjtUhtQZBtw
TfvfPMUsHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FdtIfJb83WHUVyDW7s3GfYhhyG0I7+alF4iW/EbCZN6MyNVYb3FTXHuxUUXTRcCywHUTfZqQX+6f
Neu7MprLT/oDxJLJwIG64izJ850V5rdnChFxLzlYp4FTrLDja17rmOJyJUKN9UZdeexhGmSrfGz7
JWWv0omEHHnGrWXQlAo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
puC1CYhlmGtTfG0QTveyvf9qnpE5W5/vmW1lJi1Rc4U/U6uWMh2fqt3e4uV0q7R2zg0p8AN54vhR
bBz0L9+zGhVVWD28rQxcrkI77TkJaRZ7DQBrr4RTEC5LEQLZA1rIvxpEUAhvHtQPTbKrERYeRX2x
cN2upOsM7sd6M2/91HZycOkX3qSsklP+r3Bly58PIuXfgLtCRL2HxNon5IHjrvbVlai1YZXoGcRQ
9jfSv6OkB5hfTSyCuup2dawjsaFnZTCNwwq0Ler1n7y7CK+3pAhaIvddt83WRt1KFZ88yzJVygzl
aG8ro7vmAiVkPMfaHhDY8irAzj6O056E8bBWJA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a3gRbf/0Snz6XCo5YMy8/MwXnPA7qth5ds+2CJuY9iYvS5NBXAxy0MgCeCPz2lBiGpOFVF7qGtg9
9vfZDAEH29pdWsonq5T6PGvDhHKrElPj9Yn1ERGQ1oYXdSSJVBG0+II4fF0R+zU88gz/A5xVQauy
nlrSTf9SLbJEKCiTqAM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A1/WQyDB+nvLV0GZzluskGhX7ioyVR3UZoadrJW+8ZIoleHGDE1EPsai7mYH1h4c7Ni7DzIg7it3
3PPrg1D9uinkZxHKRSBY0PF0YOwXtctlJYsQbezgpUWzRbUVDDr+1RKgaEZdwnfS2kz1eF0icLgW
aY6OweOsRP8CD6cNkSVdGsQjbjFucX+kQ2+Zi8cCJlqmMZuRkILoIuKlgxqKtUNrOALtXIM5GmNV
yk3kbRdDsNk6wSt36JpHZZaVK4i3TRzWjfLl00nF85QW0mKUwrZZvcdjyFM1ZKO0wQdxlpLKYZuo
qPfSml7T8Fui4NjLa6Vt0suXRICMJF4VLEvzOg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17456)
`protect data_block
ZF8uZHL5Rb9nKP63ZOgLsxlSsAl0ILe37VLGiUBbMNz9REQwi07nU37lYYh6kzwIewiXMgWhrnpg
Ux21OdDK1R/sKU9oj+CTDtrTZ2x5622OS8xP3cY1azpNQeHrFOtJ/aTpfgDlRsQgV5T1lpe5Dqsm
JHIXgFBAkkWCsevSrF34L+Wl/m8aiuF32qqPr9xPbFkZbz3cQEnfNFGBqtSbQDYkTGVLnBrl/qXt
p/z7KeGkNc8v+2U0N75M+7GVaP3tRLY8QY8XF4FE0YU1ulrSGCBWES8w5Y7O5yzeOvLOGAt+WECG
PH/rM+8r2cr5Ef5svtv6A/xFVJPXjXu7NtaZzB9Ds3m8EUgRvlW4vfEVitxUk8PWc4p15xUh/MZQ
KgikIn+FeaYNL5oVacuj34vi4n2TCikDXImEbMkhpgMyh/aExt05L30ADN6Js+73YBEKLeyVwR2/
ScF3xoq9KQNG7IpHw71/FBruDftGOkcj16xx3MLzWOW1B2EWj+8bBd3LwH3QS7kYr/u+9ZG72N6n
WYMNbmpmlRq52f3AAzLs6zFMycpQqbAbxjq+memcTr2xNepMO+KBdeUGECLYu2PPRKAr+9QCPRK+
dTWOc/kdwDbF315Nvy7lqBmgPj9Yn/tFotQiCQ8buTTbrbDsKoCsB0N0IrkCAKXUHNvOmFoIklxh
OTn+MCQ6X15LWtrwqVMbTP56h7lqLCeUUB9bNen4Wk2buhRMuztERE8Nze5t/+n9JDkni3TG3+r3
6+2kpa06dmxPrXoSkFN58nflFd3r3W7l4KHztpq5DImQHazGMO5l8r141LtJMoYA/aQfppKuNLax
CspwcN642Wu9nvk+Ha6jCt9EZff71loacbFFSjoeMYLXt2O/trAengWIp/Fh/UXyUAuev9AEP1S+
RA+2TxWH0r90RzpbX8WRyT1QaYpatVtqkJawz8bckuLQNQczzahpe3ejrjm7/7OYZFqoGIrSxbiP
/XxiWo85IN1vEy0tqOWq+9Mq+DpXUGadvyFWHQtlbjKy7jHACNOHO1S9t/Ni0BOAy+RsaB7lqdYU
UdgoDjpgthURLYst6B6P85c1NC9XutIg4H/4Ki43Fo/MuqZ2qo9Bp4387o6CunkiRIZS9QB1NYiY
wPHbh+LgYDnPb+GM5Gce2lb4qKliJOxekmzm/E2B2wtR7V9xTmYT9ju3rsuDRdIBuz3xse8X+nVP
6U2S/4L12EHuRzRRlt46QfKs5y0KFgI0Bk5+CBKpX1DkUSM1C36uQdh1Hw2ugrWSTlv0cBZqpHJF
Sdrl5xR6Y0a1ttD2X/QghQ8CCWELwLw5nlohkxKCKo5hZL8gQo8bfg1LReY7eeYZ3/VTLdfNK24k
/RyR9XZoULBbqGgyWhgbqKQ/cc2OOVW3TdNNwebG6+rhQWrTAWCk/hdcSwv0MeIHahdPynOVeZHK
ZdlL7jWMnHd4X5YdCSac+ltbeY+j85jgYedXq1v294DqMxmJlCEcaRs8At2NrvMVwB9F+CJxJUFF
7Jn3ch9EIG2evLnrNOcqDjNA3CG2kJjgTQpNi30UCS6IRGDfJfUrnfe7wta0RtXOrLidunoO+QN6
45yVQ0W9mlMeemiVy8ToFqGLWHsrT6c+EImfzLl14xYcxiXkAGijEzoNnYEBTqQtozbLA7wZ/53W
SU0EMvhQmNRcuL4xNFq1JoX1o1/UdWqeTlPF08QTKFXFo7csAFGSNFKC0gKbGZZOul0OMtMnjehV
KndR4ee6lzalOIgU8f+gCYc/MgpeysjS6uq6DfckkKENLgXl6PfZEwUDbsdJ65+gcccnWkFOMbCY
WBXnlmTsbG0TVjhWm3cLIE6nxLKPmQNVrNh4tujNgLjm+q/EzB5rPTimaioCzX8fWJ2fbbSx4Xt2
JXG1aAZ7irNXMM32t04Qfa0DXgJ3vgSUn05fc0w9DMq5d74fWtTOfssQAIs2Hn7Yovz424oPQNvo
VthBAUr9I/S2+fg6u56jYKu2P5OXbwilRxoksLEDcAijp7iL5JV9hgjec1kr8xfUdos0g71CxrXo
ZbTcOPCIhTO/L6OWbaGhRmq+7yYFrxWg/J9iHFoliQ4N1Zl8MXmM7MpH+otB2WooUJN+HKxLFBwq
HRJQBOmzCSurb9Ebj+suGtC1iAV6PhVArgA/O6BWTiqaR1vRhoGEApmr99hF8vJ8WSkjZaPhKOUm
7GGR/WlVghZNM9RxXbtDxfsITfPSTwgXl7oeRr3T5kQAF6aXzYlMRYCN/gP4nNDEUEQzf+7Vdl0e
fBmJa2aDswIwy2aU2wHdgr4tIZUqg2jgCgtJ6Pf4R0/RYJgdGFHIA/cPKrkbR9uDFqcHcSnYvt6y
niAC/IPGmzVe/DI0SpUY+Z968qY/pxofZdlI5CXkyZ4m/gm8FY0ysqlPb/C1w+hLVWJVOMb6PbH9
TxUCQnhvoeM+YVXTtul/pfMhC8eSB4fVuwrjQfXfKneYl59SipoUwqdznLgycCBt3a2kgkciMCak
i2h+/qqAuFN5gJXWyMGZg/ujXPW9UGKl3pNqdnj74jBvbTjgcFiE3wEYZudUgM602M5mNx91yb8y
d6til/fBtvJo8dgGEYm28efeiu7juehEvZ2an8erPJx6qYTqqn1+leD6D/V8oTtiWN4XxgX8NKWR
gfQQVu2vQA4N2HZ/mT6pEAMLBtPVnDiFa+ZuB+8ivS8Go+9x/IyMTMAE12b9Rqp0pGpTNrUWM9LQ
6LahjjbMlBT++X0ZNb0RPQD8aQk/CoHo5zAwMpTbdBWTEJ6SR40BFHIpgLQ77IvWrIGUz+IopbPd
VeAQBnKdNDAcsyqwDLcOKtPyBlYyh5QU+pxkdmwWHiE8R4/Z1Y+STYtoU7KLu1vj7E0J6CG+JvsE
JCnO7acAfJ0GQJg3s+zlZSmX7A3KKzj5fPCBVkZ7hDHrAjDNkMUDnfCGkmeuEIoKQm0TXSOJ1bU9
UjZ9r+wB5CwBlbK5bmWAdQj6QwhBdMJKm4aZ6bh6uGS6ovBoFPK6AW6wugSoyjUFd5vzTiI3mblw
y1t6etROgFZYsZlpRae7Lbe3S7n/1Ol75yuxDsAc+KK82sMbPS7DudAbDm6niI0EkQfGE6dehNQI
4E7Imc8v2cr04yZ8kB+Knfgw8iUvlf2Y5PTj2PUwuXteLxWzqkprC8UZ2blbjhZAaE06DMpnp+hb
HCW4qbZyCF8rNpXhqOvO1LxFzVM5OvRvvzftOnkipvkQMby9Vs/+p9iXS4PQjnCfYcixs7saKrUn
x5c2cmAKs9rt9wsOqQzMHXjtbRYWO8cJUWrirATB37fBfUCJAK/k+Jj16wEwROW6tDxIOe0XbzfY
b0uYNN73rC3vDkeeMjPkolpPwv+VrFyHAQoTRyYS8/BT+IQtnx2Lwb4drRsGdlVt2TMVSACUUnLH
OPm7KApDOxVoezYwLiFYUijbXs5jam4UHl29k09zb9LNX6Li22MGYo384bI/8xbZf5X/K8G80Kvd
2HS5GPEsIPExxnCzt0XMOpxTLOygE14CmJRb5RDcsBZpWJu8X6jY8qV22Pf/mpcunytoIx3TTd8v
p6BF6OHDjKo7/7p3N16HgtxUHJ0NJU0u6+Z4/0LSEGMkczOPCbngBReDXsdRC9Fm6OlOXDAtYr5K
8GWRXGV48l0sB7j+hp00U9iI9dPukr5AxfxDVwyWIHhvKg8V+1+w7mvNdN2BSnskubxTiEf7zk5o
XHHfVFC+CZfXRHLsZ87zXvLc8F/wvhcHl7lCLuXM1f/lqLLlUoY3Kul4b3xyf43paWD0RlULbpRV
xNM1FQeBWiYacLmHLk91uxhz8f9rI38J8O4f6d0Gtf+DE4lyJj4H7uTO8zgXZa8nTfJ0cy+EYFhb
eeIIDd1H51RIsFT+BWABcVwPQSrS050IpL8OGi2oAUKAYDsp6UjMgca4IQjJfBZYQyQ7VYoiZxTx
YFw/I2PfAz6TbnJkkhcv6FWFdwHjPJ/0K7v12t1Buv3hAyIdZyibnaljAC9SMNN3YqbEIhXjV/dQ
2199BtwPkhJprapDw/5ceBBLcTDcDo/gp1nAVN3fWVGD6K6acJmK2OZ2HT6BoOC91eQ0Bb/Vro+T
4VehAjlxJP3zpKWZKykyFGHIlz9VT0nJ3xT1GNi9nE2RHJUAlMM2Iz7eBzG1x1fJJBEss5i0TmJS
OcAqyKS4aVNS1UR0nEdpSw/lGNH6ZFOUveJGgwq4Ia8n/Ls1Yc8L+wLeXvCte/d071OjUQiunfHq
rp8od0chGIpsVIWiw60yDo+DjdV+p9rlOcFcqvk7SeD+2kirAId2wUtcV838e9vPVTEQp46z0Tld
U12y25E9tGLg8mY5hpHjLe0CZGZzQJc30GOjp9gPjPX5UL82AxhhLVw7enzx5wDtu/EOxDlbJPnA
lwTv7p34LunhkAKA58I6G9IxQc/xU9iOCCUGZBFgDfvSoYP2CgUMBctctd9Yjs1CVSjUOuMh8D9t
0//BCzox5oxJIwWmKUHnH2wTuVuUEgs6DkuOGWnRhxWNHeVmUofMZMDTiX3g75xDMzeZ+YN6YcS0
PkX9y55Gcc91DZM3YkAuHpmX5EBKy561w09jJ/0B5isgHvNLww3CqSsbiIp29G4aTJOO5EhDC2E8
HTxGvNou2AL5zTcD21FgkrCvExylqRQKYl3ynWhZKZESYWbq4BPi2RDFElLElWv6osQnOFUaDG1/
dVIVU0Qo+sIFyHylwmVKn8AwLePlbjWK7chuB4TzE/v+NGzbNj2KNx5J7Zh8mOTHq2RFg68NuCsP
EdT3Ge2ChcKDXdCZufsUCvPZ4xjchIy5RqfpBxOvyVXV/q1x62f5MeLhykwlrx3H/TH7msOLbf6G
x+qhVBYQHcWUX8+P0CqiMjNHT77mt97jR9oYmPNBSYWGAbsLrpw45ChCl8Um9RJVgjOImy+wKeAe
0r9EGzFSoViBrezOeY5b/nBrEwqy7EcENRAdZQIOl0Bk6OmZa2qrkTUbXUL/dCykTaadg0N6x20M
fQmaY1g17Ftrnzdnr65NJbjmTEK2p1eafExCqcUxXzd3ZoWZakC4LThB5pUzxtgX2v7GOcXpdyCI
EvC24h/ADhY1LrMJS4lvkuqww+BYSsoi2ZvYVqldpG0bL8AFAI2GTe9DBRtPjAUkeBRiAL+tuSyz
/7Kav+u4koE7B6JCbntCw8rISVhEvvOIP4xb/IGUZdNTWhRsLgYl8sULpBZ33GslXsfN3AgDmsWr
bK/EGJjORsdJ+KhTJePA/5FnSChA6lzcdhQcfR3DiYt9gps89yD2wD+FEdTsohJkjfH/3rX9i+SH
p1sqSkxYTsD3dnl+NAyWmu0j8jD77vUJ+vT947n2Z3X7LRWmgeZsnita4OTEnk6h9WMqpzn3+OgY
+Bxeyxcv7d+vgcfTrmUSwNHrRs+ffi026m6Frj/eC+9VVET+MDjBKko0JHYSgbho0cFwlteQrmry
QeiHlk106+ZmJf1f1lMGBzibgi03QfChEhyj+mqsQp7/IwylA6L7y6FYeafXJ4TuB5kr/YV7OG6v
ejI6nne7NBTCLDTZu9Tc01kOuU51d8emK4dt9h2gbge3f+nUqyGuw6861r0SOlbSNZjDFSG8mlrS
z78zTdibaP8BdFYmZTTZgFLxadQSTry+Ymw6OrHy3GA3y0Wo2QI/kGZ9+LBML4+sY4VCTS7p0kJ7
WtkEOUzENNWeaV9vMZL8B0eP9ZI13uICsM4FPeNX6D6Xvm51Od8mqYTYVCvadJhGzW7OuX7JvDs7
MWnWm15usCHdqRvkFX96/xdNx7kB2tGYFj6Z8kchsnkC3tTlrZ4bse1WTRGUcGG8Wlzbpb/H9AI7
bo2Z1TcGvSA9HHGjCa5Tq2OQEvjzd6DPBsLyCLckfXP4CDlHHbpYNlylSwp/72MFMGiVgt5u3sRb
CstDm0KvQt2LMKnFzVd4wl4AvPrLuulcQsWQ1+d+AduKi8CaZVmzNnlTK3eS4HcjoXljSdEwax72
jyfCil9zcIGSmUb7sgmliZowfxYhaSwg0D0IC5hj+yl1V9JszVf21q4RiQCwV2lZ9FMaa87Ob2K+
ytZ752ei6dGLX2ijDYQnAuMd+MHpEaJE/Wq1+YpyXHO1ZaFvdFNebOIL3sAEGrQLn7TSCGWLRkcC
tDWWpjK0rrOlrd1IqfgjwJU6EJPiUWPveVXDkc5az/5lMpU/qebfqOVp3Qf+8bDTmumv4FXnool4
JGkxkOyfcQLXJfMHsteFSdGib2Hjg5pfGKCDSz+gMqN85Liv41mWtjrW7bboxz4RnK7subKDw1Jj
9asE/gikQa5P1cGl2eLL66gRnGuGzN90Wb1TJcKRUKYow5O3xSykFV1AnOirSDnAImnqv3qT0Sqj
jXEIb+ORYoVHNkKZSo5M0aT0qCNIqwjrZv+ywOkAeYV77Nnu87cBXcOcA46q6z5pOhHxoYn0MaXz
q2AoTX//lzugC6kPe07t1A/2KSx5bOf8Zn8AWPMqnar87dC4D9ndOPO0Zes0C/v7BCprN/PMMSu5
hwNKYieHarly9bO8BOdFmv4yT62v4crCSaETiWdn0ZHTCvCb4XaBvxK93IGnhtsVL7N36VhUgeJg
YD8ope9woshls9+shz9QxRsQYGcw1YnC/snFYeZHCayZ8cJhNGgKFej7RwVEyMOc7qX3cHT/12Xm
10ztJwGt8SJWcQWlwANkje2uCGZ8Bs9fB0inBuWVmc5pkD27hdms4hrA2802ZPrlDNeh7s2d00HK
TzaQd4Qx1ztsSsIZKCQruG9yb0qqv5wlyz8yB7RFQIJbyXIJAhbwVCyUYczW4TsRsmN01hvP68N5
5wTei+SGxBoKm7Q908qlzjOeT8WrpGYlxJmYtBoEzzpMTnwDE6CQ8ZRt8/aQJ0aVgzHE0DuK1RPW
xvcyeCyzmOKBTWcfBI6akgLzV1wySc78eglk6YKRc3zZH6ybG+gX8XT5CfuC48FGEPDi9zrNcTV0
oyiwB1FnsrrugTUNV+YGB+RhVQaQ5h8HJthygDFNSnJUIe7jKMGtVqS918X9gPHmzP0Xluw2Gh/v
X0yozT/AbWkVHAecB3IBhgaxyjqwGtOPWb9ibTKhpqILakwDx531Kc+zKRdJjKAwfDdpE8rA7EOv
1mevnXd7l1+o5EN0q3ON2HKmSQcu4v0//0O782VfNO6ELyGVhwuu3wfwciFRxLl/f3YSFitCQRIm
ToDJAKd/HjUdkQyFEd6gmf3BJ7GzuU4UZXyMOZYJFKcaUoeboFCCLslEz6bd6f3ZkqFMTV5y5VQ/
RVSTm+FJYmkeL4l3Inod6YAJvtOwo2VaohhWBn+v5GIH+gBhotkWyhmK/Qr3BpNX8kNILbzyoon9
xDEHMX8JfIL1wldNPl/WbMwtC4ZgfFg/YGdVTmu8Wtp0Og1DsFmaPAzvMtHu4Z94pAfDLwZflgQk
vEmbZx6bHun8b4pTztCJ2TPTVd/2m7vPoqgG4yu7Md5F4EX2O2SAT7UugtoO760ngLkPJVHyFk0d
BaC7/W370ptutUGX7zVJK2vyyuDQ3cJv/YlvyMsHKrxnEdOekj4DbEIORFAZYIoWcCsYsvC6IZFK
oSgUaaG9BCyVdjc50LeSI5dDBZ2Hqop2dySW/ijhH3TgQ/jUh/OZuq9dNahBHc6PVKlcJP6V3tOY
IqWrnWj588LI9BF6hJrkrX6OY32t+1xbt76dSj7OV1yw/hxBkiv4akD1rPV4xmp4thJiItVycWtf
Ldzc8zU4FQYGo81elfd0Oll7xDJMz9Aa9YaxU477U9SBXTtlgjJ1gMkVl8S9OUItiM29KoJ/agWY
6K4xpNdBk1/KBKc2maUAA3GOYzLVi7FldlcyftQB1gOLKtpl2ggQ1hlNyd4m/9Zk98jVxbzI0z9t
QWaE4RfZAtHtJTz95A6sz/FdpZqjd2CU73JW55MOjQjB3gQ+/pU16teWIzOQdcQFcJeUNglUV9A0
WzK2T1ctgl/36YgcQjaMQMg73wJAIFvThQNBGnRqoc1gZ1AWQfc4DDS1EZ6n3wCsvIggeab2qvxz
SQ+0/VF2pYOEQXgQdD3ZQZ71TrAgjt7v8iVFjwrBi/o0hmzZ1iiOPa2SqwlSbPugkjedUAUMF4yA
dn4qbSnb19QMe/1phK+CfjHkaJ4AlW3FQNJDZv6pOTNqmQ52QJn3V7cHhM/HmWq2Fthl7FAMjS9Q
Z6eoetpQ7q71AGT1dH3O9gehPKclz8ZHQqR3WOJ/Zwu5cDoVeGO/dOuLAMO1VwpYB6jldpThHK+Q
RGuvqBVg94GQ6G6wsSDmnlcDlTcflMLBN3pkvKPLoGxtvE+sdlRV6+4ancz99mqqqosRTahVkoy8
3WtJyRov713NFOxNImg8yffGj4ulyFXiWgr+LGJe1+ZKaovQ8sjgD5uTZ0R8htnBrnVpfdfjTPim
kcspySYuTCzmy8gdOhodcpa/QpZlwlfd/9Tr5V9Zdvku4BtmS/WmeT+VeHgdrre0TNy6o44sGtjF
YtkjsAHzTZBUIMStK6mYnEJN8u5x4CrJZdmChZHdmsLB9NBMOM80zvNB5RGsz0+YRUrOiwtIG+uZ
SqK3BJ8oJT026pJj8PeDnF5qkFNROBWn6lRAK668G89THwKZviPOu9nPqOmnaVy5t6b77iRMUEQl
G+lOwdywqFHDIk92ErWWX5JIxu+b4tua7EgKqCzotluaEiLJYIVkF6lz8Ob6ixHQh435rMjuAsBM
OtS6gA65iLtutaS/PGnJsKJemKCal2VB3ruKVWapsJFNBSTsw9QwT0Llg0i9zMXUySjhGlq2HUZ4
Uu4Uj5T1kH2nYXtrCjv6XmLdtG/xVrIaauZCBTIaIkmzMWzsRCjwNheslQ3IPhuNlSupl51SYNuB
ejiixfi8YyXvkSgkCiD+vZVGkj90uZrtE21NwKYj2jL30Vxr/eECpV1oN89fVwJwAIySKcRwvzxC
s6S++i7jUxFR8IyU877Dc7jXkMjb9T8KJ38odcbxgtZjLoh4vFQcjFaF37OTPaDYPhj6bchMk3MO
Vn6OvPLqykRM53p5A/3R695XBhIhh8hIu7VLBR/XeCNd4e6+UR6r2E3cSmpmXOjYtl5kAMxwfpad
f1gqER1dk2jNl5g2PabQ4gj7q4C3MhH5ZIhA+NF9moZw5ofzEn0qv687bkAVX02FMRcrK6xnGTMV
j2K9i5Sj9xAmuJFyF/cny0Dukqh6UEKEcM+JO8eDeJ21xYMeb2DLs7Tw+lRzvBFO1UMNhZbDttrZ
WIUkBDJGCZtM7kZLckNsYci5L1R+gCaRVaC2CYcHBzhyV+xFeaUMhY4SI0f5o0A3yPNlMd3O/Y9z
iJ9MHlDIx9NT+TXZQ+QEEPJBB00a72NFAyYsibqm7g0+Zv8ku+wNR9buzQgGaxiLUgFNPfc9V2M8
DAguLaoSzF1cVM1xkbl4ISkq4N/rGri9CMAtwoW6W+m6C/oQosPBuR3atVASjVO2B9kh8uepvBZ1
opso0dNNGahQpichYcNepF82LdvLTfoJRw5cqITA1Sr6eNmZFgXhTxhurKH6weqY7SUcXg/E9wtj
8lfILbcyNcenMGbMkInmKXIu36J2Dl3y5OnscTQcEjYZTycaanPT5yxfsFyX6GPmEn7kOAx8ufwf
L6gsct/FsnQkQWB1N1/BnVIdrQeV4b+5mVl+X2/Lv/EyjxXt/nx0eU2+3cfDkKjSc6RiacZupw8V
L9vzGlqw2XbVxbFXFwovOxzqiUhn7J1YTG5Qrsl6oAz3YqZsLQqoDtbSn0dOfq6irFszVx5gIvA/
07nvv627L7kzg6TehQEG/PLUAP42UKh2MXWtmWSU3XZYvu1asGLPENZRL/vbjnClPiIh1H+/ZVeJ
sfVxrJqe1o2gisb17Nzw8yB1fRk3Orudz+F+M1p4fd+PyPMqG8OOmFd78n1TVQriXW8W/F/Sy1xt
wQ47CLEogMP1s6RIGceHtw+dkvYRFo3p0B7C58j+0KSDJSyefDfTlpE7ujwlj/f0JiERWT+W7DXB
e+6z4zB8M1kKyxNvUqWJYURyoj0TDZ3I1Oc5Vwfu4ml9o/sgqZOG47ddOU58MYO6S00QbaVkX8qD
vVse94gQ/zFek8a0S6vXZnSu+Y2Xd3YMSS6spCoe6tXsCGhtYtwJw4M1sZCAnHSllTt1xopNdQS0
IijJFSWBghV4uSD41ik4+yo/NfKcZ1fLfMjOBQXrj7jqiUr4Kk28Pw+DgBKpaQ/Ln7E+nfAazCGn
GT9hCahtYNVLVn3nzHKHHJVwQDGFu5FTQLXJU9iZCRv83FYDyNw7xh9x9y1xbPlAcdPCTJbP5i/k
U/dm1/xvrCe6clrza+7hdaJoMwdZs3jE9C1Td6eQJJ/TEw73rdPdOom4O2WxRmuPX4W6hTu5Mjoi
MRuq/PDAky5Dw11Z7/w820C6YwofYwyTq4nG3vKFsT30gRxgzSSqvY0gMJtCtB3Ggc44xy21nO8U
M7yeAoiXd9fQxw/8bTAZGMB84ZVxitdhxbvU/x2VRmG3+H6GXPh3F4/Kjn2f2IXDnbr2eo5OwXDd
fPjyFxb3Ui4bgn/D36FT5YkTvz6g6dTUrogOgeb+UdY7GS79pgdwUPeJ8jbRueg8ynQxQ7Uv8Gxp
WTgPAwSitflNO5wn2xWhD71oHM5qZyvUtT7eFvEE8TjzNFRuGLJkhGTK6LSCfKUoJWB9trbjUBiW
5xQdX330XRZ9u6DRYqkDy18U3psoyWTxZeQG+h8FPYVHsfUApK6XRaO7IbauQGYzVRjuDSBLOySX
DZT+QW5scVfMimpYsMz7Nr3wJyEIDt/UZVJo3DL9CdG7cID2o2CZrLmh5u9sevWOV/L8J+PgvJcS
CMRUdEo4XghNzdYvdFlvu70opeDJMOgcxmD4CHuWxxhyEub5msHJheczA9OdD7rb5bpqjIk+3Jx/
q6z3maxyXCas1PIZ2bsFFwKs+mBaoptMNbvpLpjmnoL6Ek5YxdEhTsewRIVS8sG6XRHiA1dqQmp0
cxyjhU0iUOqQuRn6ZI5iwV/jAhBBKeLUkgcCBsAyNBmpEMUxwhcitwqFpGFpEsM6ZKs/svFp9VHI
FmdUvFXjYYEC7JIxpmvrQlq/h6a66jgmy4MHikqRSpWowf1Oa1NgSPz6/QtrEUpPBy4Gun3GWvw5
+GlkaR8XgDDEUS0kgTby0A2C8XMdsV1gIHEp59HNOJdy2sllnDjggMpxyz1XetpiAW6CjeYH42m5
3ocwaqxkLWhQPMRc4/lWfHJFbogv/ADHrU75FMVoztr9JxuniYqTpefyAHTVCJXh7fTzKhLXs0C/
BnlgfLoB8w5L7E9LXEwD+aSiFvolNm8t7TqsY3XxCk24aMA5MmH4LEmqxSCaqjfVT33mM78CCQS0
5Fe0K9ph671geFVNqXHnOUqu+qxkkq9ww6aaMWFGdXzLth1lixYxUVkEoRy77zoRaHSNfyz1AD3f
eghrRnB/dsVodtvc59lGcWGSLnKbW+ygI58qNKv717RboTFwSoDfeMYaWRR5VbXLDMphhDaTYVar
fM9SBWmcG+6tfcdLyzXWhxvR7gVdv42piQX3GcIi1XFzN1FRHpTBlHZWALC1Dl2GhVsSpRFxkemQ
Xo+5rp2lo0jwFQc8Q+h9IzIly8TM8Rw71bw77LBvDUWCpErhJz1Yta7u/pnk58rr0r+/4vJP1ijb
rxJxlPJtHJRRfg+PxuqbGPgw5/O4A87Oefn93zC0+UbIx1P/D2By++/La9JZ8TUKpsFKmaBkloMx
vlC3HhDqAWxIk//kHJFBRTkJX7Tc8CZlF1PBjrB067JQICo9hUC9AuvpQ5fO/PGY4N/jChCX+gD+
rvjQCwzOgC0RQaniuYc86ZCouAaAV6uuRYnboY6lQsgNo/t7rbUq3TmF6rNzxKlD96pLiug7Jv93
reK9VXFUu9+iTdcx5qX3WJR0Q0egZQo0FkI7JwdK2nU7XX15wMh/aDKfz9O/BtghK7y8qmCjbNUU
1B/ALFHcXEyno74GQvphg5z+cKxUTnF2bgQDc86ZYRoCni3wlzwHvkGPzZ2fLnS83Xfd70+NfTyu
inrnw+ITmtb794w1uynT4mx+7LeMAYHlOf+efof70cCkKLa0UhZeU0ni2uMKfrDaKChj+upGanoL
klllkZt4SHaeZemh60IUA0nVjleYPxaebgBLg+Cf7J7X/fX0dWgyV1fCB044DUn25JDXRFQ5ne5d
upyG977aAT5uqBzjwMIG1XDWq7svPB5A8G5oBXvJj1eEOwfOYEqyEIKg6AIuuVuPsbHPBwq9auWd
S02WnANOahLIGlr4qxRa0gnHQ27ya/N9+BXiO9wHtYClUwgerlX/kCxq0gqcNoyRDz3wHRliBIWf
+Vl5aRmDz0054hWISMqks+EWhr86P5tmcLiL7NyGZw3JtG6EEcNoz7oHGjuyxz7+sKjv3v3+PJ3I
qhsXZ3819OMoG0vbYcelme6pzs3EGEU7En2txEeMV0b1dBtCr/dyyYlV0cEjlDWqmD/EN9SOeu61
YBZIJPMyr3XJ+IVHm8w108wMV1KxOz+1P4iwQLJ3oSzeJ5MIjqTR0rSd6iahxcAe1dmSSKHoNmIg
OsLpFly2ELttfFToBK7YLN1SaOgXtonzvPELvannsGe1cBFJRWOXtg/bhiYaum2H672iqi7RyQYV
qKdrjRNoIquwF1/gl3yyGbwDfhx+GydSCo2QAQ2HZwQOcOX0YFVPOECytZRZ07hc6eE8m8mX6d9o
cUJWZHJY6tbDdHX7e7N4gZVvo3a31tu/AHK3HwiIm+WmlPOcunb0wKlimd9Q5CLFnpIAKC48lu2J
Ougc7ux9pn1QH6ljmQiaDhgHK2HNAu+Ziqk4B6YaIfgEX1TpgWthp374D1R8/X44d8Bmx7Rz5UOX
qYdJG+sv0PlPwVZnZkLcbaz33zEE43fSyOxt8TTE5pNTnm2LFY2Dr64WcKPvCgLSYFSqksuRNW5B
6863X7eDLAJTOS9TCm8Uc2QCiJWzXxAbBnbGKilDbTgingFoqQxKkms3Tzkxi3wYrQkDJzFQV/El
x5qDnnlpYcBQaYf8foYsexZsCHi1VZFKebHCvY5TcFBuSw5f/64pZz91/igyN+qa1IaogkMs7+d6
/bH3eGZ/3Z+0OGMg5Fs8S7dfXwp4rDWJqApwd6lB9UMZl4k/BulqnPjzEtVqOIN9j3mWXDtxI+63
OaPZOnm46mq/Ytk4vBX47yqkUCstyXxLEVMCCtDtoBsTIBIwmJMlmM07V90QNS5b7/NsbtUMveE3
R/HnAN1jqhdNipxKqDzsf2c7TGtu31Pb6yYA3AD6bk+VNtzCCjb5Y6xboPY1dj9ti6cdZQyU6s08
F2WBLgLS4GCaEh5NpjPExjfx1WIeRBg2maKd/awRTlvmjZDti65dH5cTGDaW8byzNt/LjrWkeIHp
K98IAhbxAJ/0iSdTcKhaAkh3dInCns65I76vFFTCrMOlO5Wd4xd/IDXDfSBXS5AzsH2+38G1Utyn
G6mQka0CZg8ta/Q+WCMx1u+5bn85fX5+NECuz5mo0CQXPm3jWSaiinlJBVzwQrtyyExpdxzTfeTC
+B3gaiO78syf6r3SefcjPTWRdiYi3Td67SawY4KodTmnoqyiwBCJSIdMBAtFp1r/yy3GVDPQFxbn
MlQs2xto6c2sNjF60hDoWusbvR1A2/9669C+gJVIBMqpp08uhaqitREifNKehbVenUKR+6NsJhj9
9FHuFWzHLyZeasYZvPZLr5JT/oSb7NV8HbswtN66rdR6G297pZOffcWbJjoO0JIsD8O3OQyXO8E7
rKjy/BGzi6kpzYW92m34F6SWP0CRCvGurFVsSDZ2Xz43lvg2KUHfFngwDubQ2qbV3kjgmdKgO9a9
XPK613MeqEsB6+2nmIo8paRUELrUBBxDtJ9eEWPvm5ltZfemxYAMVFFUOwNBaxvIAdM/GnKnPGbw
TnAick85Wk8/PI0SqjNXa4jZ3dsV1g1G6/ahDQnk5vkVS942LylE0Cwng2glEZo+bHSxp3ldofco
WIbB/VEfgMVH9SKYr41LwcWil++TmoXrIaKeVW9rLTz1PgnG/IkdeCI18t5wHb7xJFHPt3/Hi17a
DPE79Z4xmeQcUlDOQ4pC/gbP5ZJiGiDQ6canDTZ5eX1oxSDqt4d/PmyG8ZC1QcVjwyJR71O+X3SI
djqM/Z8SAcRedro+hkFaLLJN/F4MtP9f6Qak4cDXKk3MH5zaYBu23FQEPBCRNDdoVm3H73SrjWRu
8F/byDpvQtb35HkM4NxPdOBldEwr34YxCgn84fVDdbF3i7CNH/+y7LE+rKfXYIl+XMOsct00PRFm
Y1PfeU/cLeCM4yI12d4A0kLakM0CTqwAYnUmKCam+AxIpkB/TTdrdAt/sCyNfpGtJQqSFkxxJ7BG
l+NcOdjxMT5m+n3a4DU/NtHRUVXr+MjGE+zHHF29W2+CXFOhJmrc/v0ViO7ToPGQc53olJfR3LEg
m2xRPccKlBeIQZiorzlzOsNZJ3ORamlmdXlhuX2EptyRgkS5YYt+MHItV1x+ZfzVMFW5gL4dH5/R
UOL5AjK/dQdlE32rXn561vGTfrnupPCuilDjUO4eV8+WcytzOtLlxu8e4N0gzyTI0g0lNwRFyZFd
hVfrILg1F3/AFm8kYcQRTWTOguI3Mh8zgZ9A1NnxztZK2LHm3WEtV6rLeE/ZZw5KdJIhhQtijH0r
c82+ma3++iJN0dufe0Qg/f4m5tUeaY4zMulhltXYR0o1HmlBAFyodGb8rqfylKxBSWDsLZeAL6Zp
xCdQhmTCKzJlSE4uzy6jMbQmEdoZbD93jw3FcSTsSfH72p1q/bbWRfof7BH3fkJPzTSzuQKptOvi
SubJSsG71Ga3tWUAJaPh9XA8RrQDQPGqyJnC0vHzNcH/yXiEJcKIOadHWYPibz2J8vTMx/v7uK58
LIb3F0TnpE2LJ0yH2EE+NE6c0b53GMSLPWnLNurL2Tykma/4t78yriwsPckEFg3k0x3S9+Rj2RWU
snJjC3DobZ3KW4C7slXLbqy5Pu04G6yXwwagzYrssm1nZWa2vNHe7xoluNGIbQc6tGlKCSsxGEfy
Jj7K6uG7iQB/F/Q1+7NkkaCnSJdVXFjJ1ScUSv3+ROKszOSP0VBzd4W3Uz0Vi2M4dJplyXu15KqH
eOmw+TAcMMqOJ55tsPQvSd/43U0Fp5S/34+F2uyS1UkWjuaXgBga/HKH0df1yKqY2jft2Hp6xb9n
3gKEDSK1E9drkqvtIJTHxNEqhnuKOE3P2QifDm0rJisHFITiwkikHC0kwJZGj3l4JWKOzKcoElS4
s94sZyTEWQu/uv0fhUiRv8d3CIvWNeYoTZR8tQYhN7631mYqjw7QkdoXDf7IEBKfUc4Mhoz8pTA2
MhGukpJE2N3SuijXQtICbZ3LSfu9bxiXIkt1Mw2CLIk3iMOLsQZh/BdmVoVnCLt9zqIEvEiiLiBx
d/dzyEyvRDQukZ0cpLMqda0iojO400xCrpjGgh+B5nACXAOH+BNnBPJy8vBvFwBkNoPoCqrRCWPW
LmWJaGtVkZT6ePiGukJYwoOOEpkx2Vo8lsC85coxoFkxXN0EFbXCiwh5wddJvT95kObe06oWkBqu
tdtzt3+mL28jPG9B8tIs0hO3QY0B4HHFnhYCJDi9NND/qvGdOpzUArqk2/6972y8rbaUp2/TTv9b
PhoCm49o645uB5kL0tAhoK2Sp5HQ4bPe//8M22u0h7gleH1Kbuv3lczHgUHIJEo+ev7kPzT5u/sR
wvcS9UYJQrFL3JH/f61SjQmDcMsRUADDOKgpAzciafwynxMG//TdmAnEA4MRX2kOEpsnVRS3j9Yw
XPN0skWnkIj3tq9MZSqEwzSweJEhzMK9vplVQeN8oXXXgMB0uEmqC+bupqw+/eTgSTV3nOniF2vD
9fF7QfmwL/GgOt5nCRbic6n77mar7HIHn9MjNwmOi2ak2DAMb6wN6moLNHD6N1EpDHG9ffW52dae
Nwt1oBXvCL/FcxlCzRMeWGpZfaoi8DgNVOV5e4t/lreLJ30m0ZY4V4Lt9kxZGmhF8R5yISTAo9Wg
B0K/Xw4iR8U1tfTton2NyjBBSfUE191VIItJuqNRhVkRWQzsf+Uw2duvDYdo8UXqpM16Vt/ujjCe
yg1T46LiGBEIwx6C1Y4/Fb/yxynDxDD+ubM/nY3M00b3HyKqm0/A0xXGqmHLE4V2M59m2FTYs0Vk
x5u+LhgDiDBGoS9tnfDNnEyx968+sKmx4YuqyoHLREEYz28/eZHqgxqLG4x/3zjuaBcx+V6TijfY
JlWMlbjnr8yZrTPMR9mGScIjdmABd+cLx5oJKGE3+jJNu+1Ub1QL7Oc98uxlepq49RFmq6fE+QMK
gQbKzORzywKjxBXIAv23UplWtg4HMrBHYMblquGJTUCr0zna6VLvAmx0TbTBs665MWnMBvnLMC/J
MprFkGpgJ+ODOFtakIIp0L6hlAVcFRZqS5FZfdC1p+Z2NFVHUN/54fwRHiZZvPBOINyNayr23hdF
BpPW8/3EdVJtaOwnffdpOfTZaCWIV4Pf4wNvO/9Q+X7zo5NGKBqMbxBEovxu+zLT87ns7wNiuGBv
u8qHxcqUSqbMBI+5DcpezwC6DdxOD/hoLRH+4XuaDkW5fXbJJ033aNyuYCUCVtpukSWe/F73FQ2b
axjF5KSXuX1vAVKwgO5nSp06P/QruiC1ftTbJdcX2wcIJZ/mfzsNYoFX8vQuCrQ4MyOyjtgunuIy
K/ABQm45Fo9WTH9GLi7d4CPA/AtrZecuKEaRgOaxnIaKArU+LL4U1i01JfqUbL9Aj9uivYOAMpNt
uwRc0Ex3UQDsVnrTa3YqJQQaBRC5tqjLiE79znt3TnFCFNzcDzRgxk93Js/hGLgjSQQ/VesV6CTy
4/ix2Ejw11cT+pI4xn/U5FK5I/bMnnjFgCqd8oJ1FHEz9ea57VGv3cp90X0UIaGc7EGYLed4P0vW
kVIfxCBq//k7S9+N8o+6CZ8xy1FInnaN4sQvMqexSoZeB4BHsFMG8qHoTxLAXCmiaSB6mbFJEg4A
av5Mzw5g/Bsd2wmYcaAwRryQxwQqqejfVHRlnHljla5WX94JyA58GcU11w0XGIRe2+l7W7CKCIrI
7ONrvw8KQXHuPans3Vc+1MvArrlSLAiX9Xe9x8ioWMGxFpFkKamwePo6aqbeqgzEfuIA1qyAQhtf
KEBd/fyIkLuI1Ebr3VCGsyvE5zlrCYVAtEEnjdCbGTUZev0S6ZWvzUKCATJxJzUbPRbf0GCWXqKX
uSVKCDMhheneNJJ1wct1KDDq0PnXxJI8wtu6+csPAEqxAEPDn2+Ew+57eGswNZ9GQ5chC/nnA91J
SYPHZQdp/PcN6+ueBA+4VTC6KCpQYMBZGcN3P1/XweNU+b2/tQ1q2E5Zkng0BJ9zvvAiDL/hnaS0
12OOUj6o2dyx3e4rtC+xYG7Cb4FqhG+a8xPssDXiwD3OC/+33sWO6X99LKYh3PxsZQc6yHoVeOLR
d/zudgQyk6fS9Ju5hU5oWfiI3FLI1Ch7S/fS/O2TGeViWXQCJmYMZ1Pv4YlUJMueqOjzztE/8dQD
VeU+4gT0Js3r75adp2CLEYV2xi7COPixdA8NW1SuAj5VajE8bQbAnEZdUHyV1zBn1d6EuhAKlLvG
gzJH7Gj2ONML7YqlxVBnqhGG+wx9pweNJiYnTCCGWhU3CmqbDr2ymSzxm973EGCYMWQlKHcHYC+4
5eFQduosOqPhjo2HHQEWr5EtP0tZoVkH8dcYPwuwNveKZEk24JWrEseCFsdnmINBUPKUqnZdAwOM
izBUmY5opIQ3t5pCn7fZn9QsdPKMncA4acSD8eiqYFH8eLrwQTT7fBG9BG5Yn1/x/QJtD/Eu8u9D
70iQvKMOOMZmj7SIiy2q2k7F54b0wHZElsr7OLfmpRxzxbDSIkbT7PpqImqhHf9brYeEwPU+beGT
H1k3AMJBFA1xaiMsS1Gzpc+g0x492QB7xUyWbYcJT7FepLfv/Lb69F2hk+VWIuH7jcQnFpby23wE
rgH5mM2PMRpdtYL4sTnj6XNeJfNVk/U5dYOZlGRCs3B9fFTXLQmi6b8wX0/+jlBsNecUaoSYXgl2
vzEef0FBBSVWOctVpbXAaLihirMkThexAvvW/0G9K5GLLhXUMiAB++/qWG1ocokMiRoVyj0FjFm5
U8ecxqrNJDn5EgCT+6StGvTSuBFbYw/FuYXMY8QDLv/XsIYhKr/aEekT90V4t1INdrXMiNvzK+pe
4Qvt8pK9U2VzXjFPIvIdp6n2SNfc4Or9uQI36nX6rYtXTm1J7FMewoxCDlfn0dvu2kqwwOvcmvfR
nUodYbO5BxqwxjANBcNbZuuzRSPLpp2Jgff3WwfhtjuiMYjnmt29tgJOSVWDjET5OEFPcsJuT8pg
CuaSLo7bpEtVgbLslK86+3BAiUQZzqPeAc+irrQcSxNVUaCtJFS52ijNiwsItpg+zP7bsXQw7171
NtNDqjJT+lqOgyN/OhBEw9c72EPd+0ykFNR9mjMxHhX60hxqfmLWwu4AlI/EmJ3RB2OhBn/CxWhw
MArgNkYK7VCp16EtC/hf24q6+w7VQtdhQKrTm2Oxqxz/Y30MwmL3laOj5zonxCl284R3xjakg8bu
EKKyHtqFKG0vLnpoSUwSleVziG8Tpo0VMeLkpkiDCyCdEV5AgV5A1L3n0mXJ4n4/QLHr0jdbto0E
F48mUYbHC8B68gLqhCZbDjFgtzPgrlTG2/fRqRMZLP3ReiXQQwM0x8f9cqjnvfbz3dJ8fze8sKXL
SWEtBBmGCZrKY+z0flAoCQtkFiAUo4meX8lX8/3P1M7Gh48R6di+FRChGpu4TsURW6oT7x56SCRe
rBE2+Nm+AmVMpEE7TlJQarbCNOjwFkG6mOP6n0FhMo2eE64Em7P60fXmctAPgNMk3D9TDSjc4Pym
nfOzIAvZp8HCljSw7QQptFMhm5SEvAu2wnTetyLWLfBh2kydhbd6WUL9W6o5BZNx96cZUiSEl19J
N0vPwUiimswEchPYTUf7LGjjfPndtDC8Pm5hu5DygayvjAjdv0jXI+m3mZKbuqwMM0GqF6hsBxzN
WEoSymCodJYcYoosczPfQLvNH8d8shcEW0SZ7sjppNoukv5SNgwT4QwZHoZgLn2ATXyIDSUspnPz
jLK61V1dUseGyLD5BjyDClKZUimTn+5/DjMSs7oq8UGgPGu5PTGuuI6wKTVfPSd/CN/0z7DJ1jKs
KUI9CqYu93AXDhsYEMch59VuOmh0S4exo1uddw8PoY3OjD/XCa6MIW2Yn7Sftcz4kXuT5ElDlIVl
AGylGcdsvYSdFP696rkPg9NR75RaCtifCmLpXf9carUMARe3gS3FS6FkxwjrChPrRfE0/6MxcIhQ
TVTGajMvbKQO7/EYikNZuZ9PIPqOA4rFiJ/62jE3oHdfXXaVgr/YhY7t2RHr2dhbssek/h+msaKq
XadhcifXxV8ZD+1qhKS7iyqugHboXyt00xhcHFp8vKyl+Wh2Ayic8E2Z1pIrepKaswSzSbu/fJxX
sREPcwfn1pvrkS/vQ7jUX454SNjT3vhD63wbbR7sXU5rUwKJuRG09IEI0eDmCkN9dJxWsy/hJ7Ak
ubBzY1MA4s3VfieAvu6nlIxfwue4PBbWhwCu9p1H7KD4ZgwKwvdyfMBZfE3VgDh5ynV1SmxQk1sT
vDt+dt7eO/APJXmMi+3woRDR5O2mNg0hWi2g20/A08NK6FCDv+qG4nsyWn/r7Plgg3yj66Ys9dka
sXckGz5o2uJxyExW6bvWT3mLHLPeJ+VPEFbdFtaiaBajfX1M9iD8uHvdENkcuuJbWiqMAxgIBXms
lkOEthpSPb2ZCgUTXWyf61rRv0VAYX7pXJAOXjBo0dGMQJ6QemoKGiJ/uWb4vWhrmudQa4oN5n0P
8larh4ux2gZTUCh5FGvgC4FEN4l0/+QqVdqkIHS4lTZgcJ1h5ZJsdXD6+ov06tTgP+NpHEwzcG6Q
eXiz/FrIFnG5qPfbCrC5LGgiZqWdc3sEuUGVcFYW0OBdKXC9XMPWe4Ut//+AJWFpNaYlB5IDkhKF
x4fZWnmB6QGJxA10G3I9TYT6l6jYC4Rwu4Up8pZTNIAWmd4T+x0wnLb/GLam1Bt5Yvr5nYgdc1kh
OMSscNtW4RmQxwqsVC/k0LyAl05P9iduU2CgD6ppMuGzZOpP+gfGMWiFmDnw5GJodCoE9yJ4xcNi
Cqb9Gp5V0UETmFqHU7wcXRncICsC6SlNrFrdwBvuYXfGLLgoOcLDssaq5WJJ1j9312QvOOLkOSkr
3XtLBy9TPNUXHCU9FLU/Ic6X6U1hrbVXAob3B6w+YsI12tbh6RzDegudHBRn33Jihgy7ZuSWIPB9
tGQteV/4HxJqS3ksXDKX77h25SUurYjBdHhsBFFiRILak8BPSnpfUPxfjEX51o6AuznR4On4osqN
V15W840/yaWHsLniOsc6luXaFBw55vJj3fi6zbZt2Id2vEKAdHlDkBxJr3xBTQeLncy6hvznENUq
x3eUVGBam0QTph4WngEC2b6IhAP5xJH7zUOS1/KhdfKSEeTaidYupYxwCquSgxPVenpNBHqJmmLG
CaVedNUHW+KBQgfCFyKECa26xi703vnQerQMy1bwcAQ1Of2K5SfI65Bzk0AzVem7TB/ccOAYjR92
Kxt87eJufPH+x+NDs+xTSvMS8ZaodPKktV1jsGiLh2+YoFpnjoVZoRhxdxsi8MMIhIqXl4ZG0iNn
ThWbwREUQI6Y/C/EvUzUOgc/bLycsAMbsmPqKGE/dSgUp3mMoyHmdTmzBnTtc/EzL/NUIaZ4TsY9
DvZBIhuDT8HURuBJmWdL39U2WAC22rmZhl8xvoaeCgZwuyB9BrmyhLR33MU5mOlLY5o+FeYuB3wk
A7j+KeJxlkFPcqBh80pjFjIPhhFua9b8ae73ajBaZPi8f0co2YW8uOtDALPJ8Vqprwocxh35TdOG
TFuvQ8ZFr4yEU/XCz+2t5pCVLhJa+t058HWv5bJQggGB4t9/mIt6D9ma6RWAJMhoZU1X5Uf79SRK
7WhYQjCxbGupRseiwelaqiSDF0jhweQAkSRsmeURvSId0VtuckioP+nyFQvEAxLZLIJfRZJtgaZ8
ewg5e33tZpvPInNIqlQqAVooVXSNGGPz/PH4hIKIt+sFtD7wYehqPWWrE713BM3hpJ/hL+Yiw20Y
3WbkUCKZWndQJ9yDQy8PNtZ+/sad5fW5llIIleA/mVWkoBn5qdRfKFZzOFLrDhYSJSzZSpGZygBX
+sF/OlQ8HJnypA0o3Uw+VZz33by+taWJ9gdQVj0BqRlHJTTiXLIU9k4iAMvBLjA8BwaKd9zQeSnx
0fN3LgKe0mjn4CgrUi5YsPK91h5E4v4GBETl1YHdx79VNLQLmY/pXzOlEaLtK3i9Fnudt/03P805
+kWkM7M7xy8njfp+ARc+HylVXgow4WrnvrSLXAO3w/25x0w/CHwFcXA3UuEPpW49D89M0a0StVSH
7xKdCqoFJ8OCIX2IdoM2ZZKYsm0md8/pO3W2P4PAM+28jlb5zZi2hA9oY8HokRnQlVp0xL6tzQ9j
WPeKBChQIFh3vbf6cMxSKMbJ7dnTb1hkIDBTcJy3PWZB8LLk96SelJuQcHdG1ptN9htljbXgdXqu
ANfz7Gms/77meyZSVBuhllEyMfH6liHcJ+edaYJYRX9W+A8V4WtbR13d2Dds/gBxEvPClNFl7SSk
LLlDo+YEyCwsV7zvT28WBUGNka1n9G8/dsglVAMETVlfENcXXD4limZzm07V+bENqI4kOvcATqSa
Kb4PTR8/8mh8lQZ6oZ80SS4T/dj5cpOCNvCRZmcpNFBlLc+j4Wf4Q9Kj2dV68E9lxw/TtX0MwtmI
QwrGgjOBgKWk13+xVKWgFcEVt6tcZDor5ybpdNolPpB33sPlTiYVDm8dbgO2JpfVhCRqJZhsWjyt
58uQSVxkBZOhTcILPBSOuHj+43NK6na3U2v6Z1xj0kbbduOxO+9bIOwHZDw7SRiOdv2p3pefldBs
DxxaVbrIysC1jwQfdQAGNuBtKg9pR04QE9mWa5Y9Q1zlBSX61Uprc6X9MOKBvGlN82mdtQHQrxt2
vq9szaO6H34PZhjGwS8Sj6W3TmTBzVnU3qW3NMX2wh0PPcSIxo9zNwlJH7pWbIBvHFCl6SQXz1sR
jYj6oBFCh88u4kSZy1FLsU/WslR6ex3/s+Ee9V3TUHHLHSuhb36BgPa7EXtgaPiTI5GGGvZRvNxs
TEpXH5P5wbUs9C409auGJW9weSXy7c96RqUukjTTIhI0QeGQt9bHT4A4OTkjT8LWU3f92nR7SwFp
Qod8YARSGNVmYujlCO0xE8OOQSekiy34PrnF08QjkYT80Pw6+HpNILz0XtmV3q3yKGyvNU2vZNxJ
IDG2W7LhXT+GXYz41IAMAYtzvXemqsEG3HJq/ZMRewWSZGLpAHvuPFG4X4cJhgPzjxIrz6PVvsBe
4zOHIBcJglcek68oMbz6VbRJlsoQl/RDzPyYx7eiB5bZfCDw8u9Uh+OKTt2rWpUrLMCQ1bneXf0G
3SH+XpKx2hFVyOX+QhdPixw+UjSPHbqKVADT3tyxseopjrC5PA3vkXiIk5uf3/TFq38ObY7pHB92
xFIn62V/jbF7YBjjGDKCcEKM5D0aINKTTGCjR0p+R5LtIsVO5FopyJ/a4kFenkVUtpJllmSSFVTm
0XocpC1RsKrkNae6sv5xZN85UjsMk8bR7xDmaUyaQ8Bftn6g1CmUCBAQ9EjIrhN/GaPgz+iWHptt
+hCRQu7ccwTdP3bbxHIdck7ALCAq/Vv8isknhpR+PbBs8hWm5Hj2CwPMRZL+0o+NefDaROWl6vV9
AQLEnaiI39y/anDKY4TlE2DC8HHB5mkveyPNLo0v66GIekmOUqewqlj9U8aUUscHgdNtyavBKh3Y
ImDM1qkuDFF6+pGvFyBpakWiWD8lp4+myn54jOUdg/RidVCmcTkLtzoimyiIOGq1cMZfBTpbNiCX
ER26Go3GwtbWsPZMFe6x183EFV3PM5ozf/htxB+Qo/7vQiDGeegoXArE5qGziV4Z9ojM5mWKLHCk
qQ14LukrNt75wyI6cBqDX6VoWcHq+bux4AM461jk3zaQ276Sp/gxBPt2PljfaLKTdI64YC7XYMXJ
fgHxFvqnmVsAFhuEnKU=
`protect end_protected
