`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RRaZQ66/gY1yn8Eg9tfIyYEVVuG9MAX7yp1LQHW0aRq8ZpzL75i+3jyHjXY8K2BxHBVI3EGaZks1
FSJbxh/p2w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LzmhgrMtDY2wQ1eWxeioEvqlOYynCwbFhXHxJ6EZm575LQOxV/7YDP6HHvJm8wBfagODCYLQIHPo
meDH8p7szW+UfwSEA3xTV3QCOd/EFqi35YhFxLamIHw8hFrznZcpF5WjdgkYZWd2ZQN2b/uT/xEk
EkLBtkPhrgr9G3d2mwY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HCjfYXZpsy4pRCieXgFxEqxznJ/8DKzir5C4vp/W4KR42hhyO+YGL6DHObxTwBHkNXAgbIdFUpRD
y1ehDZBUiD7Lcdhn2B3h7RBAIIBw0zgcZhC+sw+d1/5tXxdnKRXmBFTJl2sQItak8ELZFRw2INwL
roRq7m/1s5YRt5cGd+mjNFULKzW61nWkdJLlgG4qohP1+XxgQpKHtn6Rmnx4BGADxbWUKfVEc9kU
oST+MTUhxK76HZPcE03b/naRYysmqPn7B4dGeUJ2dEH5qzpmmC/hyHR+zCKR41lXbmCHMzZNkTwW
wY2YWIHQj0NJBz+CUH73lS1lBP6/tq9T1zR0mw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
r152pvG8vEC+eLv6PqkayJJPRGr/Glwbz+AjRYMBfEmCtKDUhE+VesIJWzICoJmDay/iTlU5iVd8
eTYaR/1Wymu/Qt00NJ6SnBeTurz9SMgiC8Fjklw7t2+S31CN04y5TzmYsGPJwM8UhtwSkwxA+JJ6
AA26OZyJ7Y+GgMWkyOY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A+fAciNlOclWyV3r1a4gGPGnWWqAH2O/F1soONnpAr5/RKoJa9DiuFuQWmFhMHAGXa2yUBBRssfZ
+KLSKDrzQ7OctM7D5Xmi9Nhm4lSdhUelo9dhfxjlKfvsHltDUAGN4onxJOgN0vPKSsLYh3fvk2cb
lwCNsl+Me70vblULgWb+6meHBp9lShxBkj0ertZUs43l5tyso+8H34wdld3IroZ6tu0mUx7jP69N
rOMhXd0cNGTw6RiyBfRRye+pUSbC22ejFF89JYarLXLELvUxOqLotjp0uvgb3vH1wnwoN6I0LrQ9
VC/xEZ7vM6Qfhjux/esEeRD0gclP9SnnJXCULw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12176)
`protect data_block
B46yJKlWHWEuEOALgZtdNlweAxkol60DzByq39DrS9uUhdbeb/M4YZ4uji6lKMl1WnUVTouR2Bf8
i+rb9CkRC46NH170qIp/RoJq77SWriWE0I2SH38Bmu9VGcchUdYRHxxGyJN9vNafAN4P2i2Rv3Kd
MXxU9WmZvNZYwdPWhUfBp66tSzOzz5yx0mb79ZCg0PqZ3xo0EmzFxBw7mLkba/NXRmNSQx40iKoR
g3EIBS51tAJ8TEUVGsqcUDQlxrWQFTxPgdhBVCPmEjfBWbFTVI7z/OQglPEp+z6NLEuyq2x0D+bN
TNpijR4yjrIJEAVZ0CGW/0WHWsT/r7hh46/bPV565Fxa2ZXq+dBwikVonYytPuHhOn9h/Q41qgvn
oyc4e4qWTsdwAYPq5NHL/YzzCJPsv40R1z+xFhIbcxBM64dZ8/0HnRT9wzIwrAyi6C+GkInRSXn4
81wPs1FuLZus+rigtgdD4e8V9+4jCpM5pTpMs+kpTr/i899BkeexcdpHSIq8kJkn2TPgwHirxb1X
f/kF2bD0m0h5bwh+7AA21sCtu54a6w+KP4Lt6pTO+G6MtuDSA2Nfg9zNkSxRafBIT4mcyQ5LrrNK
5haHxcIePc4YlMrK1IjIdBN63aXZniFN4tQUONwctiFdQ9KzHiXE7Elbw24aybUoZiKe51LA9xIJ
cgipCxqNQ011YIfG/1qtuLKh+srWarKdkeni1ivHskucu4boJ+ZPECTXrMpOYDMJ/EXMsfp7ZXFg
cSeYGsI4GojneIrhxMIehToYWlVWA7O9VAFfKv4xvpesabB6iQYJsHRmTMr21tWQP8EkHuWqcUTM
TcOE0CKsS/PLgr+IKC2WoYCgLM1Rhu/Wa1KDAFbPhAI6c1uvJPBa48fS3GOviPxPExmOZlVc4LrT
DbQ411JPG8xudk5JoMR3Cxb1ioPHuiHxH9KPcA4hMMR7FIzJp+MhanJ16ks6e3HMGUkKvqFKPCFO
4UCfyruQHJM4gF8cJE8DpQZJRcXGf2LoRpE65u5UUD6PwDSNdjAirIILXA2XgLdC78m5yg2YsqyJ
J7RdAR0zoY3li/vwwWClj8XuTsiEite2LE2krIspL8QXe9wUbg1qrC0uO5ydZPJdvPM8b5Xid65R
7rQ/ohV0h7njck9PfNzOP0hIq7xlS9o/UrY7jr6Tx2AdUQiGtMORQbmxedCUs1uKfuOl9+GR2+rq
zO/vr3Yz4efehj7CuxhFADSe2P7DatKtbVeUNZbRznB2Rk+HqJdMTWlHpDBnsLiYJgr23EhbYdKr
BOwlorQEBuDH2lc0DGIxjF6+VVrlr0/K6Ak4d+6c7LZueESF1iH3zA1fHs7Hlx52S4/wVCRoM9fN
vSPA/V/1DVoF4w0aE2jd1e3eAQwZECeYJ+b5ZAcd/zYLgsamewBhYx/NmaiI3pBePFnci9fqS4DG
+KM0wtDGuX/1ClAFDZOMOlQEVpPN5QUxjYTczFpH44V1fqTXMkpInt83ifmMevL66aUQUKI+Apo0
XwxGa0xIT47oCJujs46LA3DrUK4uuHo6LM3435gQ5OUJRfElI0PybngSmr0c+pri5TPP1JtS9wzg
M4RfXvs8IEq726bFe/iHN4rMAozXVhN/e2ka5l9yjLfhXVvIfgw85hKqe6oHY1xacxmmpKGRIzKf
8SeAvJQ1WUjw+fde5LRKLAD/YutAtR48N69WnrYd79aqBgQzTYIrUX46RclHRLDVLO1exEpeepl5
u2OvTY+r+SKxjwvleJW34TxIzDqHHWKJAk7c3aCXih8oysheZmKEhEpjSi2JI4Hn2Sh1yMzD6rIk
zQzliehs3v68EaOhO0KzU7bZF7Y+CNiR5D1BF5OB6VOedfnlptmyHc8B4LBVSzCz8fJVfogy/w+6
x6pzH2sxM14oZsWNFyI0Zy+XEWbZls7VpG4TexSYTSXO1sZOdTfp2NyLIsE09eUwOj7gOy09wltR
Z47CwyvEmi/A6qyTdRlGlaH4IC4fFbIkceKMGhnFprSDdwAG60ETWEKJfAuGoOT11CgQ6Tl0PTln
v5bltnEcF8ns/N6iZoGa4q2NffqmpCBCP71yQdvk3bIBdk8ypfSxnEC/au4JWBW4GMzavydfMvJy
LCJkaV6Jx+CAgm1sXk308sGqfkOFz12VY7sF/voJthg41iYLAn799Upzjje8sLW8jx8Rr64lMAHn
Z/Mu+vNkGtRntBYV4+mkDdfhwdJWYGLvcxpcGyzxdcMv3rtlERD4n1PExJ+OGmqY0FWO9zwqI1i3
t0QCt0cyuc9AAkfxyuX+6ulgQ7ARC4Ko2HPkH4269ffblvz5W5LyvJuSkLUHWq36tNQXYJoxtzZs
o5f5FHEBUueS5Mt+0DSFN0PZ3efgCa7lISzbGC1jb9aB8W9WddS2dXoB+rcwETfquUD9z7Fc8rBN
AG2KH0UHaApDNGjUmMQr2b8dCSKJA1BGxXLibyJ271dTMVd9hvjCtzK4qGPbnpxYw7vq/R3t1W8A
/Nm5tp4z/2ImUK8wgHyf2toYaNxGlLNz6nVzAP4cMKRq7QDf2HjcuU2XO21UKtJq6iRbBXzipt/+
MSk13S5Xcw9pv6tP+87B3hyxx2dUGdV4hzhSaZaVONVFXMkFH4xxpKuYA1C1B49quUHDmjqOcVAw
Xgkqlxj4FdRMiaTVbuZGmSsxcg+36kFwSNJpE+mayGbOuYTwnITbie7fYJ1an2K5xxoSR79EFNmk
klw5QTLa+uU1hyrA7MOdiRXRKkqCdyu1kypVwiUPshTlHW8ibTsnAJgZjO1OVlQY0QlvaRqJSN5q
VaNJex/I6Ql+IZff2TYO22CfMCD6vFScZtzcXQZJHwE8EHcaPEvpa8l8QfAkD8NTGNU1KiJNcHo5
Gz/g4XpI7EWzglL4bp0nymGK9/ixRF5+qjLEu3NDAXZF7E0MMjGLCoz9l7zlYjMW06lKMwNxGj4d
tdSiE2Flt5YN4/K6NXytH3dnclaFQRVrWNtkyqHlCojHIOQg138M8PksNFIXMB2e5mCrGzCAAwou
uZkLI4kbsmWde1RJIhauxD4wn58LiZ/ECdnsocFUWz3z5g1Tq/cE8ltZaV85g/nmy1yOv13FAnMR
lOKSQ0e9xgRMEbDphrS0n6dKVaQKHgJ92gmI60fRjf2DTXm3nH2g1ezjoqJTIWWteKRm8rrt0cUl
lg6+3VXrV/CEzTrCuEVt5cIQoT620ZfIFKBU8KSahjsmUVRZeNiO0eZcUue1DASBYyEBNlzl1F0S
bfKmI6z+GkY0ryyHzjtGejnXGW9SU3UrDjpwY2lqAsHkjTMyOkTA2aJqJxt7YRPiZzm/ZLa1hwCa
Q8sAwBXgMn2TJWX+bEx91siffj4D0lA6X9XTwy+sWN2f2pAfZlVb/ATHMTseKvLuD3KBQe/tDyY0
Bb2RIJvNc5Cv2UMZ5D/oy5sEN2PKtVlcBNIvQCkSDPu3x3LQpUIrGCNPo3TuWkKgT1z8TCet28Mu
LUdykcPFm/CgOeVsIXrwd9GvR+ZLtUx92cF2VJtQrXkgfP7fIRqOVqtkmMAeW0oIYdUSh0FV0fAH
lgpGsZrG5WFdGZpYMU1nDpeCLHNQAzjjsjojzLZz6HT8DA9elJwnqW06lYgY1pXostgVrD2kOVVg
41K3Wee6VZsZMkKv+Odm+t5zSOw20TADuTfqgjdiN/2HlxoAjMqsVAYeBWEapN2AZB2yDWrJHqfa
x0TxLFxLVMXv/irhjpmNj2/2jrQ6hOTbnHkybU7Z0xy25oX5Hx+usJQgRVc2OgHzRgaP2g0ZiPDg
UMA3YiaGvdnZ5s6hVv1X8cxZlMUJb8acfZgK7VkKaI+6YqraxpmboQQxX5dM/GtdDHh2WQuLQUOs
pkSRNecj6I93btNa/DezoARkrwRlWueJSZcBaT0xzHagUCZuiuhmhbe7JijCXgOBgJf7ToXcDM7G
+K2hlKA0Lg2g3YRgtmFYOcD12mBp7JKWJdJRIu48qMdlHaKlOKtmapeyh4fRFWF8D9IXi361ix25
iN0Wwng1GFDnsq2ZKeANZ3NMgX/xqdMyfs2RNHwydx+nk/Jj1bOYEVZq+ktRR855Un/LgYGP1ztD
ddY+4Zef/X21lG9DB+V3cxCcheymMjwwYaFvNtNWHuChvg8SdLff3B33dQLlQ3Bd8vUokN+cdDpX
bNqHm6dpnhWdMTFadaUkgbzKrWZAMWuC7P0bgx7bjwz4HRt3qqmomIiAPn8eIZ3QgJXAK9rqt1mj
T709iDmfGP64rI17DtIejz3wuo3xcq7lwnksfp8kKndS+EtA+kWwOF0osgnsbOmIAlxOUb27gvA4
4kkhOYoE1+SHd//vG+ntfl/IGwKWDcAbY69T1Fgj+NdaMnzo5zUI1qqxwZGYAvPLc/om9tjZi96r
IMAx7hOpEnrzuiaBVomsR3NPqSqDsiQBBnlYtggWB/1oLS5L5fZP/zb2CCk1tPlZEfD7iLcdWEYa
yFLlnZT2dz1bRYwcZI42atLS9RTkcFe+shsni1UYILCC1Wm1uH/odgD+ODEaxe7jzYJt2Q+4XwV2
lBiiB/0XNR/9KPOA5oRq6Mq3aFW4ErUsrSsH5phLpuC3r1WjJ1mcosofiD8QQ5djAMt6MywGrb/m
sMtbFSr8cNzJrrubHl4tp8qLBveVYWFLF6OM9R+EFpANnnQQ7vyi+2sLkVY+S6kx2Wd4+OOtmgg/
nXdk/z/cVAXnjpXcBojP/1a6ZGcpFdmmUuwnDAlKMDSJA81ESpSWI4y41NyOsZc44sgj8eNpaloC
Qc0HbZSj0H+huGreph8HifF+il0PU+zAj6e2DA+wMpYAib4sO3eMgzHdnRzHRoizaah/VSU1C31l
s9hmgHF85nhgpaUt8j0Xh8MBnkEG3epA6gsLUpsTe2CE08RGXE1D4nPP6UYqo7r4eVaeM8dkePnn
KfZZjWLldzi/mQBls5Z98hFiweN5cfayre07cd6xrDmiy6wAq7054JtukerUkELH0tnWcVXs1Qfc
ZDmmkIYgTQ6Op6zU/wPW45+aAsRAxfsA1q05Qn0kr9E4fEDKSUVGHLanw/Wx4dqhZxEgAGVdD6xZ
CV4ME5Ok/6/zvHwXa2x9G7VDnUG+71E3uVdDhFaBCD72M62bPCJH35Et4i9J/zolmlo3X5bDEFvO
+zMO2pc/nTiTP5rOnYDu01Dt2mejbMxpviktwRhbtqH0EMPJ0UbeF0P8TjMUN7CZV1sCnrxvyiOz
VbfLenCO7J7UHdjhdkWNR0VI1Bsrf9vr7zyht9IWWV2wfVpGZSVauq72GNBYNPYW8+sA3FpupP1A
2cyKRxpIw4A4minoxSL+auz3F8fgx9/Ode/FHDVAKqbhS4rAygsVAxOrwvVDsbFzVWBUzTME9sX4
278GFWw605A6GzEmmFgvRvDTNXySbotfTdRYaOwTZ7k8Xcs/mWaXGNbugDFXs9CBdcLzFjp/JNBy
J3loHyiX4/CzgPGRETtfls28fLPtLWR308L0wIFFpjuzPRvhiN5kYtTBL9v2uN+amuePDT3iKmDI
DeW7WyQTE8jtrbBPblyQapd8wsN8HNZp3bnc4CKrGr18zbGrbsHSUO+wJKvn5l2SaZKgy+HANHGC
UgJI6mkK6jxDlOb+yb5U+pMEsgk6HQrHfQ/xIVI29E3oAAVx/whIWATb9FWlKpU17VwgYQnA3EDq
hUrxtVmo7iHFDeBY/6KJXmqbJ1YT6t3pBoszO8Ary4tQpKz/Hb9AZvUI89OL9jx2sRaMrXuxT8Aa
XNziZc1nH5gznGJetaFaKpBhBY4b2vM8++NBSB5kt3bfbWT4q0PilquV1WMZueSxXAbz363R4mWj
wD/jm8kyza4xnHAxk0nzYC3brxDYv73BX107stZs67FfGTOHW52Njjyba1xhRNWoYUN1TOgUvm7f
DGb1JriEGqzietJUM56LYul5i5zenpFG8xI3q2ZqoTLWU9Joi7E8fG9IsDSyr71Sd1lDF+oV+55D
2R8P6KeerIlIgP3VBmS/Wux7FseiGWmZQ3CHXWmcVnJy+TwXHcL50klrbCEguTVbCJXNAf42ulHE
BsvJJZMCns+e79b5glKGbTeMCXA1/shm9+2OzmbWyq6Ys2iB9OjCxK1jg2sTCQLX1nhAevSUweow
FQAzfMGKsZ/tDyg8Km+4u3rCHKY7XB4BHeeCScaK/4uanmVqcCdc59KXFaorNaoLzjon5/mDUe6a
xsecrmbAnb8UWAoqq5CllTuzULc42yxRpUDXdCpRJpAB8uAzC5HSAOzG7T+EPmcMizJiFX2txTnr
/bKigg7cQAW3+Bqc8SgDBj6+xdos0a1iRtjZQifP5Le53H+vlFf+0AsD5bNhFg5CV9gU7K1qfrO6
76wFVz/U8h8ODVHE/riz2WlmMtB1wzs9NoGjCx1vCJFq/L85rFO0LcIBtVR535bknttkJYBz3eRO
27vYuNKFzP/Iqgpep9kum8CUawZFNPNIXM7FeVkSWBMeKZYN4Xva0snlOKTA3kxnQfFkC+Cq6soF
CXAkPRIqdkkna+hR7Up0BsBXQzPaqWz94KI/23+aG457iN3LMVIS967SgBGsN0sh6h9jZkfImyNB
80zGj+zCEShqbdIM7b1H2H0s98O15CaCuqIzTPpzvuGTxg54wc4R9Lf2G9rc7dwDKjzMVzAX2UQn
2f0Oy4cGewigZuSbBZpjMhOSjWFnQqOctAYjZVOC3s2/ALM06ygl50PrhRSwdJktMTD/iXh7BNKH
DU4GJ6gtu8Ysg1pJhgY+SpL0aeKzYv2uo87rj6ROq0jgulfZZ/3HxOZmcAp26F+F76jG971Rb+bS
nhF8rl25yGI/93/XDGTmRGN8zgRNOJTUCHAyOVnNzz24+CYkWQ/1qrziQHgNfcHFRPivFAsxK5zp
9qbbyR3FJHstx/T35KIeoRY0Gx0S0B6LO4ltRGGKvhr7/44QVbLCZrVjFXpf9U5ZhxX/cEr/jjpx
E7uCw8ij5TUaHZ2Q7KeYQMiwXIVaCrtv5Pl38nGG1F17DV3LjI+ITaWkeNcvFajVn4M6yIU05jGq
ycP04uHdEql8lRPB6oa4znwXTB9v63I3XYcyJus+WT7e+SqW0DdQ3IIvCFOnqyHnC1XZzUeu/M9s
mnO8cxRvQXU2R5lZK22rBZrGh2SvDc/JtqPmb4IjaH4Hd9/4o/wvFFiTTMupqAjZpmOoizHGzh46
cprysn9pb9GgR4FE455Z/bSNdL5VfDad5ZLhW/XXhzG2ao2fMvt9dcfoPeF+rx6nSaqmls/T52gh
NjKQ7qZixu9NvlWmHfwTHmKvY1hJoQ/QEGxc6OwJlDNM/FTUhmXxck0bVrwH/Y7jRmVx8W9n1VJu
0FElsXRriSQodCSi8sar+sdriElyinge3gkTrv42EBhx+18kYyf0FT+IwVNM+5rpuNFi602gV4oa
Me80c8FGV3G0AOFOFtpLygixEFlfD1CU/b6oyvJMuRLfw3AZ3i8LxX04aNgr1sd1o/V1fRoEMIkF
GfwigAx6mqcHgKcbVvrI68jF5DTmKovx3OM+Z6HYkcvzWLLKZ5yNxuLH8+ZxUgIyBge7+HBQYlc8
7bHhhYEADNItjffDlvG4jO1+arxsIMAsssN9t1zmjVvCMx07DJfjlBy3L4KE9XGqJ0TQtZaxoDZ6
r2BzRcomjf0KthZsbz+ex9IuAxAd0ovd3yvsjTJbG5zkZPR6rFJKRw5kPvc5eqKQsCTRefWCFC99
eeqfB9w6UkW1PO/oQqNWEbggibbmNlPVRGc3CIO+h+oMKIGJldGUakYesQozhs6PuNW1HFrWdTpM
gxL/Jr2rnsKv5lmb+DKXxenBuCTtRQy4jqrkJNI3t5LPCXS3BjvBStw5AYnBLYNFpVJngPQubyOc
xmaF4+UqB8QkngHHMgqoueGmHaRzAYKtcbM7REuzSHHdUH0VsmLW61w3AUbaLYZ4lgFmR/CMdR+3
/eh/jzSk6W+ZEOcyPssisqsn1u20vPAOQpWdb52n/tVPEbCT3AptQ3lU0J0Rgd4DE/2vRkH5Um4s
KaaqbGjisj2ODSrHJsdfjvtQckXLN2GwHBlskWULIgbY0ZkUrQD7qVR2M/QtUSTEqEq0dOS2uYAa
amt2k/uczIK80nPARVbpIatKrrpWY2k29P3jVEFmeNQvAh6s5cozrzt/9OKh1r2mwPnwM0ED6Myw
yRP12Yg7oWmyAza6zTrr4dCAfy4e1qfosKQzCbnPfdaxdmT2NI7bMIFlhSqy0oUlM7lEAC0HBYmQ
cv8R3J6tR9fawi9hBxNO7cpzdmoHAgig4a3fn3z8zKEPx8EOomArLgs8r40S21llwxX9cFUqbNXY
ley8PZtKZXuSX4JRVphfuXBoSMlgstB/+iNrfxTNFvijmuw3Efo8rp+HmKTyWbbcw+JEvovO3zSO
i/1iOmb0XiAR4pqGwrZ2fhAvAoi6BiseIkME/f1IZaAptlIXpKA8T+BEzVPV+CeKsIEirpT15DoK
VBEaXbjAhnHwVQW0/EwiXnVfsK1+i/4r+kEmQHOkWf1WmAUiS1fkVu+opQiXwbCG99tunOUh5VA0
5h9h9lDZZ5B6l3Lx68lrmHbtD3fMBb4+h6ErR5EIh2U98YPmFe16xhaQyqXljZ5GuJOKvv75wllV
7B76tgg4pAd8VXVQ+o/lLYL/CdlHZcIK9se13VFJQv+ZzX8gOGBmvTWs8CCxev+r1ik2kt3u7Xyk
0oAgFTs4B08g7P5Qf095sIWtnKtGqZSIz7/YuUspK7dkOfmteKi/pl0i/vqk17q8Y930xYWV+9dH
09iFnEoU+Wrl0VW+luugzilPEQVEPJonBvgfUi2I++Q81VQuIQ36rl/kpJZXSdDeWxyEQjCABDBD
PK7iltUsdIyOKuuFWT+T972JT8/jRvQsRyeCAks/gwytAar8+VECV8ls7W0nnw7sZ1JtxL1jLwnf
0k3jlmDZfdZmOq1lo+3wybdaxdMJFHz5UgxGPHOWdXnlv2Sopl27dbYENM4nJVxcg1x7n++KHezg
uD8iy4NGU6X3Ct828AP5Nrdo813owdNvc1NxNu9fXw8ZE03I+DrLLAeNI0QffjkyWb89qU/FRBmM
pebnyaxyPJiM2uNHjgs2VLJHaB32gK3XY/U+ZR5DJBcbx42FmYyo8kDWeUTw2W3b775JMvgsTvpg
/6GRFA7XGj1Rq9LA1s+Hfr53DbKLji4HEFsH0KVZ+zBgGdAc9k1xLK67qCBTAe33fNuhPhypNPr0
O8fTtdRnrnrpjeuki+JM0U5WbrfWBnzUONrBwUmdcNY4NdVaGxkVEN3/zniISRxC0CrTyRXyu3eM
fVGjhpovAPRHsvjjdD2kDt726gjkh8bikCI1Qq9xYotZN4sBVVbmzXvH0SqOFQHSrhdPfH+tcuIA
2P6p2SN4hWrY1RZLMewKlETPS6a9C+GD0IvBSN7VaphJ5tuBKLcvYYfXnTRhpG3yUL29IJ4/luXv
nQSpdgAzvZyvBSiDlkKEZfd0q6id/rFAGkG0v5iwxA2KbP31foIkuCXKhyEkPflfrZ0r5HjHpsaT
vaufEc+QY5yAIb3aLER7ZGL/C8PW9QpxDYLKwACT47zAwvJ61+31fxsvNz2jSUEd6fewinUGHWzM
qo1+fcNjMqG/+lJnhB/+blparqmQtKghAl6Pfwxz8USqqAopPzW2awo0WPdRm/Bno2G8s56d4RB9
lSQAlhbp9KNZQBgPPPZryxQcI4kGhGDmoNPgKBXOhjShMTAwB4uN0oI50kEfB9GwSGeD/UXwvu0T
lOteIu2n5nUqDsieuPJOLTieOel41zHTmeKzI+WavsxZvKjrO9tJALDiLh31DEJ3iiwPQhiB/aWF
/WsvSUl9bgaSSSqi1L4Yq1oJ/HxNnYL1KuMay2KQ3bfmiJSNf9L/MK70/0cyWXVNEIhqk+DTyLYC
4b0oUnK9WOjbrnotC9RrJGSRi7KubJ+cPNCIdImnG1f+WPOpoCiX/w64kDBz1gp4TGDxyEBtQ1m2
cfRJv4wPnlfTA3QCRfXBbvniACA/yaQOptwdb81uGuGPSm8P1azDHHNurhlKDdSxn+BIDWZAvFJv
eAJNsJRs5HoP+MhDcN/J8E+V9ZYAdUzrXPR2Y33zd0tjQl7LrL9kCAM4cBwnHpBkA3j9Cb2EllyX
OwZubrREthUYuAA5TPQfbgycc/SHMrqurrYB4gSx04Bi3bt3+BYyfoXu91IyBzCiQz5EtlasQRNv
8rxkid/dskjEt2v4BFX9V0bhPu5eHhDXb+GwEvu3REKn0+/tMphjjVncqBj6K0J/CAf6Yk0iCccm
U78NeD9aGAcnz9kacrqXy+kcxLdW7oKRX79RcxBzTJHdiWeeElBUjfclUxXiM+XIV9DyNmBa4NJz
+PWntSQPB0sWmUz0+I9yf+4CTOGrdi43GEZt9hIxJuizF8/CE7wPFbdhwjvsF4uXgxqw0nt5LBG7
e4PUMx9LSAZ13n4K9E5Ay4W2EhNffXKE19t9emdF6qnqchXebZV08FyYZN7Gd66bcdzZ/NE7DDKw
54t1R0Wv1s5aDP4ksjZiecMmqfMnth+v/9i/2pGl2N6zbVSjLuEeQZaE44+iuhjoW0gYWS1M5FSm
9/2hzIYmQHaUF84UUicv2sJKaSiF7ppnmhb5tLDU0aavx6O2rjv+BrfkrkAwmOxTo96wyAXrB+wk
DuTwI2FOLeqyTuqWqixCJY0m79JWvY3p7DFnUtT89ghYNePmAra9chBIdAC0SvYNTgKeVazqGVLM
Np6y30DTY0S/X/7W5kBJA8xNkTGBisvV6N3XGHQvVT3LsDpL0LqApQc1IfOONpNZ4ISAWLJmGZyy
Wxm9m6uIq4nkfLolSEQRo5DXrj8hkWEf9ODFbNhw2PSObtxZKJJVKm8xAEW4/ssqfb55Jaw4wRc8
jqmUhPGRnjJ/SLFTXXzFwRilPoHOJKvYGdfITX6HSPUkMgi29vCJHu8989oP4f+DWTMUv1KuWwWC
VqqL3z8eczd8qpzT+OiPCEt9sCoQv+vioKB9WJG9NmjueUFD3cfIaBw9gwmfvQ0ysUgeNevPku8M
ZA6nxuSDFT62d3AELIpPoKgBeMAcshtncCuLT16AXDHXh+F3CO+ONCEXaLrltT47rBHrtC5QFhUU
WbdHZmsNdJbfrfoouzOdT75R39cu00IdVQZoCiMxqXvd6brxJVYQn8Bpz0p0no54hxXPkR3e5Ckw
cgj4voq+remI2aVhXOjpxMp+TeK3AIXxmmh/YKL8X7GvFCFqx7vBtwx523KRTTOw88PINNgAno/K
9EtXnYyMRKdOlomTNdkNW1MKlqs0RJdD6kywulVlx5o3fhzw1mVd24FG/7gLgPftlpcHXVYM2riP
/12p94nZIc5bDT+LvKfKCnV9N1yKdvKmlj0WiN/8fc5O7SHJzUGJkXQ4nvHWWnYP3X/juqbp3iuB
5W5bzl5KejC8xoIKIEi7rScZAIC7ViYA5dYQgpzWfT1eI6wJydwsEs+tcCX41Za54eJUmC/bNUUN
9MrQE14JEqpsQTNUG1qdMEMt42sIl3A9IPVhUMhWvky4GX6Lqj3c6eKX15WkSPcOStzf9vSXG9hq
UTb7Rrv3d1WQQWFqt/b/yq7m4Elv76c3v4IxWrP/tGNhKBp6WM5Xx+pNxVWhzb0XzKFhUUHQZgEa
3dCAJ3Q8S+XCtQFxpvbWXxIcdcUdD/LXzti8JGPEXvSzoKiBGkOxO71hjh17OZLFea2Cehrm1dLE
Qatnn3cL/0QP4sBuFP9aYARJKYG31An7qijtGotA2KCdV0ng3lv8+xArDYwCCsZKkYt9V035p88q
wqjzPTgRszrM03X0v/9+UajPxqPb75DBoGRbipEOSwEsJiIEjznzMzo6E/ca1PQst/9uPdMdr4mD
OvKpupQWAewX1X6UI7h2lTdaXf6HRCgL1a5s+3IKcew0KVNeYrVZtzkOA/ewOV5brOMXjT7V3SFa
SsAul6QIVwp7so9dFMjb1PD9AHrpwTZMRYb9/kSDhfK07rx1TYhlVm+d6LZDRe49hxoNEt5nvGW+
wnwDI2vCZsWnUHQJzvSVRF7U1gjkRWE4Kg6bgkASitdQydLqYuHmSCbL9z4VA5YFDwFT5Qeaer8O
JhFcTvLdqjZxZJbj2NTkJRBIXtqq/SPWGgM9mfEQQfxti2C5TUHP2GSL5RwzOOLba0rzDigVP8sF
p4UHzAIj+abdeA0CRqvPiNxf86YynCzuwwdY+XNUo5s+js5fWSieEWiIodMBCCr/VnEEGVUooopZ
e8EioKImiX65mzhNoimDyYjHqdtRFAClcBpL24BeApNgvriKvTt+8OXFZROAU8bCGLozvOSLDg2X
R19kAtUSPfLpO4xpsJRD02NSKitYrT9N0V0Xuk55E5zWIuKZ7WVK0wifxB+1I/qddBYfy6huK7ri
9EPn9J9cejDMp+KsGl4LyEc1OrL+DeMESjo2yXa5hdhO3nKRtqYoXzgYsQAfHL8vuPMnWWWkaJ3i
fetbzJC6z9Q67/J2zfDsTWHg5XVM8vqeMS8E2hHIFIWGnyRhL3AdqW6w0Q6sgK9dRU/AhtjOpZzr
eRB2u6wZe/uOwgolwW6pztbbfBATpgyHd63t9MBVZgJg87sz4pNpcLKvmNn5JEqRv3sExzIZMyo9
bra5rWQYROVdH80EyYCVXFx2fFXCnSnThHsl6ayC57d2l7WDjeuTcYCHm6W7RK5g0ozyC3XUMAaq
gQhhwdz3fNecXW03iBbxcGlDdBaG4jF6W5d2XqiKXgFskhuz9jFwMpaz/bcMITklIMN0ETL0eUIm
kTtW62QVQkP7wdvCtLIk/t1EGxXvHx0oVcJ355gBZJ449z1EvBMHPdzW6VhoQeWT9MtkMRXQocrK
19G1isgX7y2N7MYdMKKAggLZ1ayxrwUC11JKl+9r7kipvPQatu5FPx7Fx9rRL28RCMp7pJPKLQB/
8je61x24eiNL7Cc+rW2+Pq6PW+h4fm7oWd32u60XBvGKh8wRlbIymlRYXcQD2m59GObCQ5PD+OLh
5O7JmcEymDdxR0It0CERZjW1tiuFq/r00RQWcAcvHV9d00w3fKWAOICUO+m07lUBAwX2upRY75WO
zZ+weiqV/sRQ2Dtn7i1L5IvfmXRI0jerdgqkJtUjEGbOYhdsNyEe7RgOyJqDb+9d7tzgyLK+9lJw
ukJDVRnK0x3izjIwjPw8MBRBOfIYyOGpb+bY3lsGvujcXTaqkwc2W1gczF4uEx0pvzUII+/wqQa7
Npejhd0Vg/BI35B2xpudiXA/XKJ92dcf6+7peHxEehIbJxuxVKWxz/WqYeAE+vRRRNKfofw8bP6e
JtBLOsQLWWmUROl8vKwMiqXd2SNcPqWcyQdD9/J6lv1OsOQMxf+N+Uo+yjtI+wsevH/ntSWueSOU
IBXgZ62h8w3SWDRiItUL+dpSAsarZU5PY4VdX2Khjtl0dDbHz6N0HXGTFyrUqGAQkCYCaUdObble
jd/COpbYrVId8/gZTeGh6Hyw6lP3ZSskOwHTf9NyAstz8UtlvgazYoPKAg+LpGBEewjzMHXNg0zi
TCJx0YgG4fbYFozwUKjT4kp3bjxMB4bQYBKZ9ZIP8WtH+UrUa7Zue+FpGUqwNBFMIi7caDAo9VQ3
Ui/oO+bjgGFCeJUYCuTqOMMEXcMaQnsUJ+C6lhcyxtUw+jClySLIfQ4zJepfbitJ/esHHYt72iNE
TQ1D1mI97tgFw8UUPnJncDKM+naX8O74BEdKFP6MUrlUlw63v1i3BB6b+L2zBWqANUZ+Wo2aUGDo
PgXm4CpyAWvSgyp5boFyvAT44L/yGITjNVRd05Ulc+1PYSGYi+djFsGeeZ6NDnDt9P353u/k3aB0
ex/AsJxBGMWun5iLG9u576yS1GnaomTynIPPJ+LiZAq/fPhdOMuOsaZF8j6B6/KKOFQEUCfclmDh
7g1QgSHmiVfTjYwmoe3RGoN5tAf4h3azKYce6gj6zXRjNMl9o+UAp4xe4EWryTcq8aRC4BB4BU5k
BNFY3ys+k/Pj+o7hJAcAWXoDz+x9JPxe6T/fZLFrry/O1EfjqRzA1ZNyid2/zreT8S3TNPO0TTyu
PVOb52z2uZ1BqzGu/dDEtaV1jDW/ioevuhHyy5EUvyIy6880I28WqndI09ucnkOzw9yMlJqBlW84
FkDColF6RhTPRRdYO2UacNNvd1ODFwW1SHgyyeRwLf0+M0efViA65H7yYFiKA09u3gqDCk6htSmG
i2kx5N44OT13wa6qRzpK8+7G7N0FQfUNbM/e6ghIUeJgdesqadSOg2fYpAScScrGJisJ8Uvz3vQj
ilXMeL74a0RKAM7sqhwgE3+rhWU5K/jJiv5MR2jk4XvRh5MMEY7XgsKY7DIgYyVsMZ0vs8fokhU3
p3XXpdH29rZKXsegCeVuA/EhI5xnZdoLoV9Gp7jzz2CaH9rglAyrpIlYZOUdQARDfu4DZ13zyCiq
CH+pQ+b0SZo8qeNeyNecnvFB5Q6g1HAR09z7SfL8nVlJzqozewpYF/OzyMKkp2paVgs9UlymaPWx
YDGNuYHCw6MtfZTx5ENT6aIsupvRonK8tYsedC/h0sPGrIG0zT0bLJXF6fDmKrgd3GcuUyVjjg3a
797dPgdwHq8ux//VtlDCxQmWk4BHEYzSIOUR1kU87Q0l/nYBZk6+qdiO5h+WCLRPDJdCHKtfK5GJ
XOU4mEPnB2gQrNeLFBw1Qe6UD8AVjEzkYBQcfz1+Clvm3Wa8FwWVnBIDY998kcIELorWnrDu86dY
dF4UuOmB/HzkP67x1dSUAdzCUL0RtrXmcwhfCq2LS3vknt6PJ+5uW9pOk7zbiKpgYXaNhybRBN4J
dK7C6nsJW8OmjkSg1WeB2lACwGlv+POlGUkUJUbzo06svAB1I4Oka27vM31lrj9Fo15RyElcRHvQ
3UpyXYs7Z37RxpgPtPWjhUe+yWEKVtZVyfUJaPn/wqN6NJqsRhOKGu9WU429ySA0zoLosYmXzYsV
bZaivDv2im7r8x6p1a9BK2ofK/1u7DG3F1CNjHTM7BDYDfLN7D2hAiySgU03lYhGygXsysXqnvY/
div+/AvxAlbeMPBMl37Lyovbcds3dReY748UvRjiSFJvIMFWBVeXb0d7lK7J60pkOruByuAQbCab
HN4V9Ud5EXIILpdGhMhzjjjSrGcOWKcoTCBZJUudw2TUfaCxfth3T7QMJJ1DKVPY6YyuF0Ggsbm7
YJTRGcrOjw8nWnE2CmDaZpwKLFW+7NPSNc0gmb8Pq4ks/ciWOB/irmoOjRmZO0Z4fAnYPJ4vF5Wz
FluiYlSoQNQGFLFKlDgcl4lzcJY5ainMURU/4h9i4xp4HqnLMWN07X7XGyaQjeD7h/+9RpeY3GD9
bcO9Sy137x3wxPQUouZXwPjVsRyQjdpt2GunVgBQZxnEgbmX4A1aBlSnDND814KW31cZez7WhiFL
bLqirlAnARDOqnyO17wpSkmM/vMwDZitP3bVaNfAgXhAe6EUJh68JhQEoIK73ypHc6GBdUh+PRdW
XpaC9GVrIJJyATHrU5Q5/ptqWLdB70blFGTVx4tuKWgS8kjigCM82lQeiF4tEt5kx1Fc3WRlF2eB
S+SPSCU2pmIxmtjiXvnHDeHEGWxBLWy02Ke9fLqlnemwopPfjxT4fUOkQPYZzBbpwGBpqemn1UmM
ks74uTw25TkqD9a3yEV7t54uzPmU/vGsET1fBiEKRWq5UfyJjEUnbuZLfx92u0JGgPppY7iXEn5X
L7LcYT4VGfsrjBMGrn7awz8uBFSrZ39ZA4RRK+5Oxb3wqFImITxEp4ZZ5F0spOQwFV1sjp9wgD4a
g65pgrRpNyCMYkEEXyvfl/pEszr/xjcLi+CSnWRF6lYfdAZbt0p70u1ZrsEFKBPosuCKoVRmAFFk
ME7SjtwbrbHh9jPJuFHgVA7HUqDoS6C+uAbfrZpEeOVWkCukq+Y5lmkHuFMMSI749ekLWlFPTMXj
cO49hsIVdM3do7nA6m2z4qtEzvXV0T4lCKLLenePohdfwIj5cWt77KxvvCKco3uTDDeFxngvrsia
cRQ0tkc3Yt1/psJMr2xkpNzwfb2PTAbTdLCi+nPzKzC0cItgydZufQ89MN5Dt/aRBynXOVppszI2
e7mbOGCC87sRKvnkCSjMYWcYAstI1LTZO/uyZ/l+33skoyg=
`protect end_protected
