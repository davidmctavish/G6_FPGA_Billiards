`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lvSE1wnTbUzcyFaEkCK/oaIwLhSg0I6H5NtAJDSx1lTgwyyckziPTGY5rLYavTcVFBRHCSV5wXpw
oInm6nX4CQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c46olHU3F8bCjhyybwcNX5+VAFexzs/MQFisGTAzMX/KyUASEQnIrxg8MhWz9kHjdnq6rKc37dVG
1ZjbIdn8SkMrZ6jO7IRmCdIwB2EJTzAsoK8YFSf+6vyLoMhBmoDwezZkm/1rHqzqGVbjJUUQF2G4
P62ohvDWyPWNNIgy8JA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kk1hNe76KGY+Tdlckns92+3icZXVsH8SqvU4x4kYPRWgztibTY8vqSlNrsqzBHJdsETPt8u0QfLK
rDuQWNGJrxqMHSKFIsyfEfs0bmfsNV+V/rvrW3PMMpW1qQmLdTz2AR1aqM9ak/yz11TVvd+gg1S9
8e43wm8aETQxbosNdhrNLl9/0F06bpoxxaqy9pAztWtvjybX0PbWTo7mpZOZXhquCHhDCOgAUoVa
iqF4CjXc5CNxWspFmUpLkXJoG4RQW+ZSYUNweVqwAL+zY/NPkwMGzKXDJoB7oFe8gr5J6WuQwXzJ
K4AytURqWSKZO1uQyvsgQcXrmvaVAFUnfFq0/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2meTUxRFJcrHQ0hBTBJTkVAXwoHUYJpgII5GQKJSLR9629yOWtHT1gVQQ+/1DiJqelxMhOcZUTQh
U57QePWpJ7XVAAehftRjhyRKZvvjOSXsylQSyb1EU5+M8QqtLhmpagSdkcuEV9aR6SlXtPWIwzSH
4izOxcUZHdfC9UgUzZY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lt1ufMLnNLe6MPpqKfqVCN/YfycsVOQhsMH0cw/qRDjacuyDA1nAr3hI5fo0QPXNktQ06ZB0rz0u
+2ScolNa5DnjA0UdgIGXLztxHTJ8oj+Me1AK1QclJZE9Fqj/ihlVWPX/SWC018RWnpzz+44QrVbR
6pYK2NFPTh+zRUOKCLlQSCa75ftb3OYecza1taUkBWsh2vJaK7Eo7Rco7jppMAvQKKHggXtDwbKk
/YzMfTJYfkOVud9zn1XPdRy+927MWTUJT4sKcU9WL+psbWvcWsIavw5oJ8LRjc2oHQ+z8fF8NEvV
PcXHGZfB8tkdxiwwYgEEQalcaKorac2nBssNUg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103072)
`protect data_block
r93pkmwQ4keiO3KnJmGKo/0rSJptVMC7qfHCooXUyGZnmpQMgubF2FBn5lUlH0BZeMcdeGCjkayB
PZEb93bs0+BwMMWipf8BewLvmEvcweXgge3ZEmci1Pc+J1ml1/ZB7k3vHUj/vWBP0IczAiQGzw5B
3Hgm700jtgNo5VA/SBjnOoPY8sYpipJbc+3COWXbw0yQ9c7LeEre7IzV5JczB5nWnO0a085E5/8P
RcVR4h8H7gT4JFRNH1/21QLg0YfLzunSohRovJAAAx0S0y7pVe8i63iFByrYgWfaKd1imju49dyS
Szf4aJ3Gfo6e1LBfCQLfWAf1AXDPw4g8SyNhm7dWlSXx0npQ9VEpZdM+qmKkYMpc5aw19flJmqKt
KVHUzszmr7SQirco9puQK8A/N3eQuHOKvOFpnpVhkgU3f9EI8HHsgAQs9z0kM0dXf4h/1SHe+VBG
3A57zaU2qr8V31ROWlBe5j9HUH2zQJ4sYLFuSu+ktUHzrnKUiNxgCVJHvus2cmGqRw7FiEhWym4l
kQlzXCNY+dS7UkdHlWhla4onchtd6WOaQgr9maTLmTSU/DJcWrfkIGDesREx5jMORFGD1gGxCOQD
+N4jm28aH1YSG9CgD7MxGci2LpSQuoVHZSU9k/V6oAwZ1ryY0YBA4o0qfOJ2ldmTjZ0WOYbmvaKE
MsAn35ee1kLORxoq3ZLevD22K6VfaHQseqgA6J77sfm/KlqwHc+3eM1o5eJJ47jAc9EAn3J72VQ7
vXMkpGCMfWtjbjwqhNTIy3BpbTSsLLmG3VK034egYqZy5XNjsySi3AFqLstQUCC8ZvnK4QgzdUf+
x7CTKWVpzhuKJP2qx64rIZX8LQllo2lWEWAXAPN5KpzqexuR+H5H1wJKuqHziv7ZD1qmzX/6Dhzq
HSHmOLTOrkyoylYUw+FtUJNWvIZd04DT7GK9yzkRBBs0qsTntt0TCCYy2BSfu/f1Bn85Z7Q9Etzs
J3XLTuNjJ33lb1+a2uOp9cDGY/A/+NmvajjxUbc1zqUlk1i9NcpZn01EC28Ec5A1r+2FmBNANdqY
foGuK3KE2nOahkc8/2xRE5X7uA0sn8z5blYq/8U7obhX8PZK1Z6JdlENB7jtXStwlN19wvKjE0Gm
f27ZltVUxklhTwfQYyGzJYB/mTq6LiHzPecA0eX/cF3UuvI5LK17DNAeZvn0XJbS8rVdWPRQdSSR
JYkIUrotxOITx3htZH9+fnoCOicJ9Dd3CYQzSOjI7PyTDGTDQ1KFcplNTgMKOiiTncRHW8hKzj6E
aEsCUqK+e+lxb2FnjWJJbs4aQkG4GQgQrTVZA9Lgr75JgYyaWcAnHnCjzQ6WwjNny1qmupHELPEM
yEshPEhUxVrerdh7pOu3k/D53H2MXTlDGZ20VqBVnnlmZxRfnL0AzI2Fvkd8ss1wi9UyxP/C/g8J
DxAnWKTPE/g/p4FGhsmOBa+rt2DAahp1E+SFU2EwQ+dCZoWzaMy5AhcT1UvTSOgWLbnp01l5JkKO
ET7NOQKvFSpaI9rXJrtdtV9UCfB64rG6Kg+lR3FAlX0TGoyubVEcFN/CDyed8hJz7xJnKm3fBhwL
Ao3LIt+AC/cC5dRgsXeo56OKVrSHlLlFYstOHq0atq7q/S5SrTUiu2WwXoRid1ZtEX35UMAuOE9X
Y9ZcphM14pGxJ1m3yfi3zxX02rw0i2AwrgWd7vMJRj2EBeMLgjbNboksiZ6VBtMqw+lz6623l/Xp
N4RxRvHiBgTsY3HBJMVz2jJPe3WEtt6qXrlnGkXOx/eKwX4iXu3cYTU5KDiOAyYEVX6LVyanDamL
ANF+RththJlPmBxFYBGIG64mHK9tTvREej8BanU1UWtGe23NR18l1G07nqJ0xoR2QD9gHn6uZQOO
nc3+8Q5diAmcKpqixUapo13820RbL3s7mAsKbdTyuc4RGDngOcaAH0BMdX3XkRbspDRznFN/M8Yg
YCgc3BX+xAs/WtVSjCG8ejo06w5PzmpqCa7+5BIBja0g8GX8TwZaC4Wr5ngpUhATpc56wLyzY3w5
NO6/zCDWkF61EkGmSmJWC4R38ks21MYUWz6XIuIALoIJz2Tv5uJN4HWFvUSbDYon3uMT6YoT1FYW
1uPK84HEC3YaOf3NZU9orhAEpdHFR5hLnVVuCq/2DMYxIihJNl1sI8o/TiRMkGljJfTTvdwI5qwy
KwS6EYfWND9jecMecesCPShKWX0Ch/AXLaMvOe9btJ4QnXU9V8kxbzzUHn7SgVjeEIB6F21RWhu0
+wiHolmT7hPmQNHva4iHjtwmRH2e9UGFLKIba8kjJtTb1BUCFxZjVdU99tst24eKOmnBqISD/grV
xl1EpuryRLB53eERr7+GYd1UKDkAIlYQnXlQT0h/TGvXeQNNm1aQpxm9yZ1aE3qTxn2+Oe2e74jS
syxbeS0vMQLPa0nmk49kiDKXhftTpabTefI7G1CRBf9uqCdBDILxeeI8MTdCHHe48DcmhbqbUgI2
Tn+LWyUUL4YYF1793xpOB5VbaBPDDvem+gVsUOnvMpHKKGHZ90E3To+/eGhMTNiwJlRfAlqeCkUF
9dvhVbxJUvQHQm/WHnmI8emHGYGPA95f7lQAcFAVXKKUY+S4x3W2HbmL0Eltbf4vXofsId++GRuG
b8I2CMOVMkm6nFnNagBqeHxl9gdPOHmbLfSSSnlQ7yBmfC9A1DRs250d3pI9QnBio/vIoocV2vQ9
kumCp28KsiLk5j/VZD+gcPAqmfZJdUVDFeK6Uuy8/HAXc43fiaQl8HIYgACSLXUR4qXmjUvZGsPV
tEasp2bY36tKMnEzWJOrvURtI/Q5gA92GAieE5/c+E/Zn1i6SKnC6NoGVqfBmZrzaHOMv2B2/2ov
9Cwmq2G5UsxG5O/17p1Wo0s63DUROIIKIqhlGVf/dRApU7VukRTAGkT8Cmz4FYxLP+HUhAxIvv6J
kAh2DzeySKi6OgHeCsOwWVISY0scMhhtjACCfZ0rHIOkt4P0c6jOgMJ1JTWtdN0GBLIOX6+/KRZ8
dPw30evv0tpNOCev3A/mB/g/lMxF+VNgw9WopvWDaCFTHrxPx0+QLWDkKsiCqKfPly5Vgi4pHgp2
d5u2/GtrlStOBjmeXLkxOFNM9+7UN8OdVwPLJuunNy7gPo336djDsQBf734A0xNLHada+gEIDED/
FMarmE8skp8FKQblnsuA9iyCOQjuP6KV8GW5n7oRgZXufiEhU5jlVWL9ynWqjOd5Ap41V4osXqXD
LwGO36jX4iNqxv110LkjES2jCFRYmIKUjkaQBeGkTLsRER83osEH16oVHq4M91Ug/uGOlGDg9q20
cwMJagwo+T1s2n0lz4A06NwroJVaUfF+Ztizl86XgValN0mNKTn3gNzsdXFzoeCchU+sEinq2XEb
i8MWeZnsgYHwLnIdv3VTwEChIKKhcnc5F9w997w1uDq5X4eWxdyd8yTcu9EY8yuwWGw3dlw+bcnJ
eqlCThH6Rlg+jeAJlCBsNGpnf11lJetZCwFd5lY88q5HCF58taqSqSEcnUPt75Dg9EA0VnPSdBX2
RAYNtz3Q+nUnSnpEvBJ0knMwd3xuVyYmdpSnjvKkYurpMFSqEMACt2KvlXfG4EZRiEr5tXfAPCGx
ruEQs8OiYv2jjphnbn9ULb2FhxegBoVFYfh4QdOXuOW57jPaUnvujJIMXORSgLiyPfSpZpyWjvdF
GchZyo+85wFmLPU7TAGzDVRU7uFOkBnHoq8B+hDXbGhTyW3nC45s+TY2TKFw1b89XvxrETx3phXw
CwZAIlG26AXaKc//kpGmbR0TM5NetQ5/rsvzkeewedADswVF5DLIOUEPTBZV9s4r0WxL+NKg2pmS
fqZDh/OnOouWf6SoM1wmZ5BMZ2XTENUbcO1s1DdhIZuFicjX2fkAGS3JsnLtFCcinoL9agswfrTZ
vEXNrFKR9DoPofPyarzN8tMWfZC28qTTkwr5o24PSCnsJ72GQrmHAUewX73KZaMWTxEOEv1TrX3R
gyymjedHMi105iFpgCBC/qJ9qk6s+w84hoiv6s/nLAQJCimV8U9nRYREL0vdOEYW+YMk5E6Y6x85
sjK4s3Ea52cMDnxAeQ9IStz7/M5t2qRULTwnWUFrqBwhPbINQP2VQsMoRzGskJ+kliGbiYnwGkAO
LYs1DUepHZpkJx0SZa3QycsXi8/YTvbWPXNFX7WBZGaV3B/0S4kJuhHMve1MQj23F/Gn8PzYK1oz
1wNTdTagqu1cLPGyG/aiBRdJUv/SByrxqGeyRQY9MWGHqDkCFfeJbO3+aLD0cFCUAMHXRV1ZRlsB
juDMNSZ48NdfCT551T04HMARRtBJfjGl742Aj0uab1Zjjmhg1NAMHLhrmtwqV4xiWklBWJSRJLhf
oNNP3VSJhZsC9cJq+00ADR6gM/ucSLNbz4o4x4FTltdAb37KiPnPaucqpYspURwvKW9IiyxP4Nlq
7Q7hQdmSgxMC0ngV5FkkrqY/Z27xKgY890c+eCAjx7cZWELeqU2gDi9HLDPKcs46NE1sKz5Cy7ln
o1gpthmoHqTDr9QsIjlnpub3z9BGhAvr0Ik0P4E7WDCfCtEOXz7vvz8hGpk5h96E5nlD0XHvLy69
PRmEqr4y4VnHXLguVn+vx4ocG3F+M8DTOx0JIn4QdmtibZF54Fq4pFw2zxAWdTD4FrYrBVPwh0wT
wr5LcNjr63lXS4/DBxf8PeqlGhc9uhArmY6Ing+XIiIN81OEJSY111ewtaJDnhrja3bQuva01BR3
/wx+BJ1a885VowVDiXf5IUPCzsssW4ES0wJSAB9p/Gd7rfrBWIqFPKRN5YJn24kNSXLHeIhKd3HW
6dfCSrWgbC0dxAqcUgkGiB29G8kQSKFjqxSCKKycxEFld5GdV/BMc5yvgMcvSObELi4LfDEpwMl+
quJCRwHnCUlagL4xjE/qbukgDLKt/g1Qvn1dh/XdDmxSgOOvypsbbiuq0U3N1vlJI99TZ8eOEk3G
MjG1v16+8t5f+mbh82Kud0yMJPEwkWsInvXQv2hFBXP7tbAp2FsATNNZZf8zxlbs1pnAxIP0WyL3
n2llnq+681SLlJobq4c2HBKCw1bukD+96J5I4/Tg4F2QS7FH5ZvOYy4hO7nVws5BCZZmV5CZgTlL
H20u1akV80/2m7L6mdtDVoBhkoub+SOWyZVRBNKSEKeqv8a7DLeEmwv4L4amePk3cy++AwiPJm4h
nFpOS+Undf+hgptWBauuUa/5q3USwpiT8FLdehbGrBnYG4p9mozFOuHXrarpOF0O+xxvhxgf/Btq
z+VhTi44N4QdFTaglH1majCFMn0eAdw4YJxuR2+0Te3YCl+as3ev3kFofzaFub0+iK7tNKUl1s/W
1Nig3TIFNepVow9LNFEdbTzKp8o/481WTh6THFxjq3QBNN4boqJEQI+t7Tap8nC9qT5o/Td7PkCI
1ZRrILLBaERMmF7hjaAOPuJXvmBFmXrE50YYvgsygcG2oZkkcyOlJo+sb6a1Z1lgdwr/9feKE4gu
9alaYUqxqt02G9zT1wZTjRcIcY13EDGV9t7oys68h45aVUhifTGD9Qmba3EglHtZmutzA+tUT61X
lNHhhfueZ0NJwa2CF9+pIDyytf+I0gFnubdhq/zRQFvyZNafh+qvOPItom1pk/jufK63tnwwcBhg
dyVb7waAaveIToQhsBEL+R36hL+iHHZboU2dfkZHN8RSybxeQPmh+xjyfbkcdTLSRKGJuh1iFP5l
UZ/xulsq7EdaoubyxWJLu8kv+SyM4T0zAmB9tJL/v7G+qE6cdlLrX6Kwha8+AHo0ja4W8IvyMAvl
mUX02kzcsyT+dxuLu5YUuDDqjSMueOqeyXeu/q4v1PYx0RqIwU2JzC5wdL7Kphq5jhokjGplu5gl
RuykIzocwARHJjpTloKPJ1kd7dJTY+NCbXKEP03+0+CS+F16Y2n58waLNtdQ5aEF+OocthdZfq9L
HfW2y+9dYytJxp1TytDkV1BNUzyv60c9861adJ0P1+eG0lxVUhzEK4ZmlmcFYppvnfnJvylOEfEJ
HhHrN9MGQ1Cb3Si5myf76R+lTgh/yas9neCgOL1r6hm4b0jYQTMQc6BfIwSIVZce8iU4ttmTagM6
i4bU5rGEeH/PjWvHg4J8ePAXmnrGXLjdgTLUX07ilh+24GyHBbaDj2hU8pX8/fB8rdiyjvrt+H1Z
JQ+7pJb1oDtM8RdLpAqBwUv8cPUVt88UC/3kF3vSkrPjjxyANajWXyC3KDPovl7GtDWNnPOx1v0+
stMvbdESp9MA23UFpksNXe4lcXZzKykDKgtYjJ4ubUSAIkiPFfimmn7PzBQjdwkaovwAngwfdQYd
Jer1dLHnn+v6Z85PT0qCyx18poZHiKWiQxkXoXFvTlKcw8OUqkLQHoSg67rh8ld7rbGPuoe3dsJr
kh8uLkXrxtQRgVdoNULGCPMnAnpDExNulL3O+VJf3fNNhPBj/7AhkjHlby0sW7TypNytzVnFUD5K
cjkbR3zaLCOXPQs8ZGmqjqr3IdePOvQL9w43IVqEOiQzxfmVRVQrL6DhLpfYVhI3gmHKGTsWIk8E
4H0upXQu8GuKY3XuZvmm55O5AfSHS73T2POoAjHO1+4kdYcpG/ybzVdZ2q4eHNVesxxOYD1HswcI
VZwECHqJESIVHZ8CivDELZ7DptaJjQdxm2r3xS+JNrd3yAB4CjEdltFDY5z33fIhOk3kQ8Y+uPw5
2JUsudX6lySVHClPMEXOFZdBVToC4gX2wpEp/+Y4dsHGCzOF+2Fy894wWvbdtZAtcgvYhxRrzpeo
yCtT9vqsTN0V/zNXeGy07CSVm4NDCtGa75V1KpiQyRQRmsss6ZgJsscfDesJNSNhhfmT2YlZW31p
pRKwE8Rxq9G31aBiEXlnx3YVbUKUrRJXyytxMG7d5cT3ytMHyawVcYkoX+Jg637voBYcg/DdWdRC
+231qH5UpWI/wEMKsxUDHCMR0yYzmm+YSVLeO2I2T3Kvaa6mkY8KgycSq3UictkYvSgjy+XAovxg
weX62CDHdfItdkin05uepsNbHwAPirqN/0XGAQcE7MbwH2PpWWEvXbH+NsEzeZadWCDD14FZ8BxQ
uXzyYRMnHh65I6+p9SKIdBn7ZR9BjPRcayjLdW3SSV1t3HOrj19HGlwt0eWPpHITG9R6shhkzEGX
/hD5AsTPwwmwPHmCvdmhyTZhGFHi1FZNFzWVS8tzRlfFNgbB8sdvk77H4mM3msZJpMi0EZNY8GVO
hEqB1mAvD/uPXa9PAJczASR4B6zuyyjJscELWSUG1nGinVG12TwxVj0oOx220MYqCwsxHIuttiQf
n3iSHeMW5J5g94tYNbHPKcmnn6jyxT1r+d8shB8UdaMgvL4/ZgxBaLvhNouOY20iIiR+aixzWCi6
vEVrqlO8VL9AToVT+hMBR0WyN7xlztWC44Yyp985HiguppZ6+IJSwJPd6bJRJrynjur/eIZOIRo0
s4BppfpNexKSxXz22RIYzWBqvTmJE4nLcj8Qe/4Y6x9UgZmkqMWO1OmMzSH+KtEDEdS819DhR0/b
sLXm88BYHFTJ9YO0y4W3CwOC7CUd56yY54xP4hdkO6FbY8kR/DaaQhCLwXGPaE7q3MHIXYplscvR
fzixpfcWeYZ+ktD7E9Vke7JqGffXa8yo6rQgVYsYWWLA2fUCO97Ex/EvsuSpC7SCFk6UXlmy3akf
BelVK36QDrPIvyJ8ZdNr4gDcLgOY7Zf7UpeAD4hkeIuc3hmcHijAsLTVwuDNVB8z17CbeLglQ6vH
b51fKOcl4T7MH2zTCr1jN0qzvP7FKSbOQk5ZJYiBGTKGC8oo9/h+eClYUf/23IdGGiuBnTpYGQtD
fzc0LAbAcL28tm6X82e2g+ejDtKX3eZZldWAxSLtUHAcankHRC/TnwjUXCj/JD6XXQHYu3P72LTM
MmZdNsrCMFERM+aa7O9KhGQH7/47nj7a8+qAK+uDK3s76n/RhDxY2lrdv9jM6Jv+nkR3MOHLx6E5
L4zxveE/xTkxuq/tsyPYlJcCLs0M7Pz1mhMLQRZWhs9awGrrk4vCjbVZdacUpSwg7zAhul8jZ+nc
4lMfAE8I3FwHLebXwzrM4xjyHKaoNioXF81M1UMDkqxxyORnvI4/oIRlU4IKfdNvxaYxM9FI2ub5
qr5s2JbZPzGsh4wWXQLeFzg8oH2ES9VT8FYs3f2PdBKpfUdhU8LvHbkgExKq/v7B2u61bTRPo1GS
rhsc4GNmHjkNQDY1cOU89+eTMKc9czufiJoQT05opufhpnQrlWZJhSEq+KZBuxfcpN59gg02/k3V
tzc8np3ncNsINvZIuFgEDHb1KEsk5fa36k2QMj9ZQGnSwJ9EifVlJDB+2csgYA02BMcW9Rs6OzdW
p6kZa43coiC2oJtx5EIk/K6TdkpsRHeFnNdTVQbUdz5CzgDmBbz2F3q4xv9PSdpEWLqtPmSHo47y
+KAVbxIyOcf+pwGgVy/2zod0n6rpYesJm/pxWD8+mdYhYYNC+0GzjJj9IkCeLOvuV3pUNoQ4lbh8
mDcRYyOS5kadUyT87e2vDg0OJGBIXTJwCn6DmjotDdCa+5WcbYJFaNhJmB203EWy9McqddUK8W0P
cACGmNKPyrBRb5ElS5eAU7EEOpreRoZCsuNYF5UPVHZIjf6whdpZ4snLsG3oUEuRK1YydasGhodA
WY82u/JMNCXpbVE4Dkqlr4bVUMXCXpMJTRYi02s4cWC1XGqgcjPFpr+ar+7HGasIR9mQqCZDs12b
xLw/HjBP+AhFjfYLW/z/hMKsIWTUTf3Bx295n8Vbi5+kgQsfmZgEbX+qWva9MwZFtxrm2I7rH0vW
RKq+rxUFgXmA6jgFeafvLcCocX5+roxffesWam/LSJx7BxtspLhQxJlp7BfDnbC6REIofFKUyd9j
0Pyzf02fd4S7hiIKqXwzY/axn4MlXGDfbjzUGb2ax196U08O9YsyQSjK2Uzv5lK0dIv+g2FSl37e
H4R/TUYlGVwbopq/NnLiEBSh5Vnx7RLL/mZcBq0NOTjTUpbDI7hC8EfnxlJIZXW4cPtvC3HFovBK
TSmDEDoXUGVSR1pSfTw4W8/nqYhKbB6GWSGwCSYbI0jP7XNrx9g07vOzPEKqTYPH+Syip4ixnmVK
EwiHvICGDPM4Z2dowo/3MAgEs+ug59xLhUS83lF3HN64PnGIgdwHoH/xJqI5/Q5BjpuxAZLyCwb+
yjUsgcewi6DkmEgAKuSTQsCKnqjbMo7S9Ld96/0aAXO+LCXnmikgaLK5jaOOY/JgP43HyW786Avp
lgjDwVwQOgdMb4GBoDtsj+Q+87XtugDfzX5fIfMaI2ctSEghzgd+8yWOklrDkm2yB2XcrQiade5B
PCnj/JIzKVqSYXcJrxh3j0jhT+YnIGVG+L4SUxHSohSchZ0QmyFx1/q9jv7m1lPQYsYrgyOx9LAd
dCjONH7kIM56i46/6prBVxKAvV+LPqMiu2CNQYERxIv5ts4aacrVKKKGxS8nF3TbFQxJ4+q8x0MQ
Y8V52zZ0QlovLJWyqLyvsjd+HZEPrNdHx8qMFnZbqaYKySyG67FhlvvkcOgvIXbqawqBuCsKhJ3Z
xZVJNSLp5gnOzCQt5iwauKnbC8a2qntKXDCbC0VDkHZ0aC420N10BhJx9+toM8ltGXX2btPDNMef
v3ohaSlLd0/hDceC5T8Lkve5WoUXmKJ7E3n8xJDBqS4cLpMCF7Vqk2N0GJt7buXphz5Y88nh7UqK
fh/jCR2lpxGeHN0csaY3bIEpLmvX2fT26aAE7dPiD6jLZTvM5XqbJNmgwoRZa6drzM1ADIOKtHOa
EJrFRQXx0I/FSPUgXlXhjicGfKR17ClSCcz2L39dKdtqkFywozfpOgX/56ZIzFwMMBowoKz6JVKN
tihD/OSmNOMKAYAnNMyMe0/tuH7QxTGWBajICuZJcFxFR84TgA50fPxuIrgjNrvrR9rAln/38VYJ
/7VdKeNVmi+BD0174c4dXZ03HqpUvssl6I0EAFs8S01GMsES4LVMkXt3UoZ68VxH/i+JW9GZmQHd
1YJiwEaeSRYlUTkYurzKhxrCP9zTf+8kjva0FyfH4lWhqAl33Ezh5w3FyG/jLcMjNULHDp+2ZJyd
qs87aMh9UdloA53HJcLZioBpg+EHA5UKmcLPuF0fsPQL3l1Ld3rmP9OMZVFrBXA/v8gnVE8VvMK7
TWN1AZxlzpJwpQHkiA3PZrF/eV2dTNbNoySHVbw/RFW/ksfiILGpEFVct5rpD5gXy4z0bfjohf0k
NQKgi8kgakTkeIitXz+IVYXTVRL8+nxul4EWIqWAo5H5JvKX8cja9V520JyUpTcrrStQ3ww+g5Kr
gExF1n64I0ss+UvY0qu7Nj5Hu+/O3ILT7sl1WUeK6qcz8hPHSMAtH/Cw1KxZx8qOVzgVP9XzxYQB
hZVC/8eME32HKFjNrZCUrRm8IwId18vqoD1jSluZMxZwDFAOYpfK8Ss0mbWbg1U2fZ/MsQLmnFav
meUSwdR2KUlGGFj0T0orxoHYLLWgkSNGzOQ4x2xYP6SinjW4l1BITdLij0jez6SQLSHhHNLS0HoD
WhHcO7CJI62YaDj4/mHBmUi09eTYmSznskjP0w6VNWAHeYB+YN/sfbi0b+2Fgncmoq/losm4r2TA
MEzI3j+FCdQLVenG971nF7wNxv6CsYEPbCT/L3tTHwDtENWIavAUmDKJQ/YQVzFiNxYZ3/s/pvR5
y5mpMMbY71QA4YTJu4XDrMfiDTxzlgWcdDCs63CYDxCGKyIkvzd0Uc6kVF+j33kP+EdMjUMo5W7b
svzADzRKn/ZXAL6GqPczLF1m51Dy13ylpwQW1QZMq68bvikZM/5ihx0RAcx9/hpYfmGR73pJwGZD
Jg+atm6CK5KaEXZiE0bRFbEELYGZzzy//8wmUEUY95G1KYk6leU4BOyyetdKjKgyF4zuYHZR8QK9
ibLuzJ0UsSO8IhfT8zpgi/LqVvT4xrUwF+fa74fER4GOpEF45Tk9ZIT4NJsQjmizKaqQQr+Zum8P
gdfG7jIuZj8Lj4xcuscNKdGkfFbdMeJszTDNleecldIfBichytympzb0eYARjauAF0Ih4GYhVI2s
lRmJMdBJvzVpctpgjBMhBfQibkxZZl+JDjmJ9wd5Pqv8+kQ5vZ3xA+gq0VV77h+J89Mj0vO9ZUww
u5rdUPJsspOj/VBunFj7OdQaYEBteeM3z0/VD9a1psuMe3fZyjVGRL/gFYQStiOTgLGekY1UoMUx
lvJ06UUHT/LcamlfS4IjePZn6sWLP7Hqv3Xn6mPyQ1xjsCj6tKNT9EmITzOUDPGDv6+BNgHV1nDU
Kj++Nkzm4QQHcCw5111tIzDv8uL6IjwJNeL8MmSVy7BIO60KMtw5qcq6sNFcfTX9GsDZcX5WdegN
mrzT0CraeCgV+fI9siIqqYvu6kGgD32Io2LBn4xE7Qc3DQw0nuSE91rqryX08VfyoZpyKQNQ5qZo
uVPSYzvoouUThjr3KiqRrXua564hpcvE06BHSWanLrDy4D1Iyki0wlBmC4+rLusODACbyXzQhN2e
JqYThaFst3DeSXmV+XZifdtRsHjVr0Y4NAVFdDQO5EwuuVlIKAnZe9Uc5a4vap5E8RyMhvcVCVnj
VxouVPTNpg2d3gVzRyRH5LRTk81nokgwlcumyo6ruT9gShidNq8CsCjgHK4XkMGmaNddSFKeap10
lyGypeqP9IyG8MHSMrwq/JpSjg1wKXnKPYSolBmCx4PumN12JcH2JDaEqWBDTo88tV+YqFHgJ24W
faz6Frs1E2aRXZhhOT3U4l74tD8sghm/0bF7KsRIBWCvqEKczcbk1hWaR1y7Hggv3Xpr8fF39/Di
YDiEE2sui4RN669CquIstQgCLtAeJGSsYDfPva/aclkUFyUwg1dbSRZ2xodBWef0dVhX/pIjlHmN
nE5X63uJfyCOwCswH0IYbHr0gyxC/ide+uQY9zD0Lyn+PuQvWwk+fcJKLmA8j8r+x+e6bD4JzimX
FVif0sVNM20xnOVAeatffZMypzAIvW2YYBY7T2xsxdEjARlGXSE8gUxSyxmKplpaiqO/Sej1mlLa
pmibGhUozy9WgYqVWhYpggI0I0yb2Db6n5L2BbSwHk6R6x3TS4kCtkK6yJZT9SBMdagPdAQptWSd
gENpyZs1ixNIVf0mpIujhdYCazRyrW9y7b3aaE1hen9sKy5T/I47vuq8N1KRklPl+GHhVYINultf
vGl/8V8tMzs/PRfeToZm6dVhiWfl3TRhd5cnl1D8ysRDYMi9hoZLWRVpO4hM/imK3JeHt9hVSWUC
uFOT5Hph4hWWZvmsQa3mjJ1uqzbMDgW7zV/pQDztUZunP/sftVZwysHQq5My3mYUAmXtffmeg9NU
YAOBIRdZ1UrPoRDyRoHQVDS9VSPYkN/i00Wubd/6CckuO/k8Ma278cqvLoWxrSpplttt9LtIMbKN
n5uFxSXldqsrA3e3nQo8Dxe1PA4S4RbCuNgz9ESzes9LNbXIBJxipZKEbp+HeJkGUtZ2Jtsg/UgJ
iG38hb/eTgCCM8yVFdPgqPctV7MTcJIdgQ4ui1JWnJYfhBkoyWgx7wj5auXeCM8HZkCx+KSagaFc
u/8ZYv/ljFc8EO0b5n3FQaqenLCPFZ9bbtfAnGluJGmJKZPQYB37KhEgeL8H1xPJpYJ5JBxIMHSa
XQiR771vNyjKxJluBtJEMNZFmW3xjpH/kXR/gfJ+akgG2cPy7UldtzvqzjWTkv+txJV+afu53OhT
ZLtOSmD/W4Xq+TnDpg6lD5VKQTsik6k+FVgNroHO6IEWrd+dH7vDvoV3HgaomdoRvgbKpBKsxnCq
/R2WcPRIi6rqAcF7X93508giBhvsyQ0TmlEGbrjG4I2z/vcjVVlc9eq0esP+nu4uMm75YZsziN/X
xjf2GkIwbcJuJ0v6AyPSrd8WwpWk9DyoscaOajbyZeV4KGv82HPK70CDlRYge0GZsvqmWc4H0jSi
8uUTc3vDBvnYJJTd3AY6hDfLvVQ2tkKvOlYcQp0EcKtoC3aaep7FByQSUzOntwQ/Xqqmi0U8YU6L
PFPtZgLZ9f+XLbiUcJ+FAJ6KKnM0HuTM02MkyJkMNBaYjZ7VGfqUhn1JL6AdHusWN0zm2px+F1pH
hfKDlbt/FaQQD1MxOFQXVX5isXkXggi3vVWsQV/kwijQ5IJsi9bDAOGmBZZi/gQcloQk9ijKQx2N
CdQsZFKWXkdQ3LUICfWFEmzW+JegOPqtT2CMQgHXZ7pyQJAus71hqyZ1TvKK6vsFIXZH3HDeo+Ba
LcT3NYLCTtJ2elEANdV4KRSdf6NG18grd5ze6vNdDa2qvSbUIDSEYU5AuQ0mFt42KtPcJ1+M+aR9
euZrD5cX9Cy1x3B9VG1ebQB8IX7L67OE3RHiZZb/sBuX0bcJ4PQxDHtmxNd9XvfGvRD/2AGxPNw/
aLNjLpQSV9eAllRg9LnC+u+p0eXNdB6qxxkGuATPPNmyEeOcVSEpqfxxxf/raB9njSu4O9wkjodD
VNU4NExhE1o2gzzw+PJrwGjz4DxZKGYoyEzkss/4MmQZpDHFfe3LKHIXzLDHostsRQnXvQmqf37r
kdBympBMdhunosnIm8a/Df3H3WtCCZfH5xzoFPodTET+pdN/O8ObB0qhhOoInZwBrfeEUSs8FY3C
7PfRvuaWK2EThMg3OvpHgqAFA9ufWNnwV6biArUvm8lPAMOhbQbPtOcSBeCTGGIL8u0LF543rALF
7XwccuradWU58zwY/hmnRFxBdua35yjHw9HiMsmVw8Z3ofEFRkDDWpBQdQAdqqRZOri9txU8DbjA
CHuKhZ8sZrVvhshqFbH15zqcq6GxU0j6b3kZJt9glrZN7e96j3ANM2J+K7FTBCsBliEIlACJJ5En
rVIrhXq3j8qDh/veUeuROY10VDMBY0SBnM1r1G18kMO74ucobAsoCky5g9xaEKnasEiI1nWIS7fk
Etyehaq05hvWHmX4oXrEAjTNu4tGpNn8VO94u8FGMKJsTtq0mFLNc9yuL/vc2LTRuikiHPOmlLt5
YEErMUYpW+jwHLiS3MEx2QyIvJqPc5dCA3n8iO1ckkGWcWb0nHk6KJVKkmI3hJOQknCMnPkiE1Te
J5WHo0BoB1qqwBnSseQkTndCKewOIYsFrqCpKVUXQokaZJmks7yAolYc8265M+/dna51fIs29N+/
KYkrMz676kqh/i6xgJycglrdPTBZ4rW2eZ1pjjrapd9gIxEDNgrSIy6ehd7jw24R/DhAvq0Dxpca
O72kt2BFeOy6RHmX8eDSPUGtiLd25fasvL48TV9KYRznGnqPYN7tyeeGowa/JG8LCqwyzlfBcG67
awxjc6fHecxaN22rXYpzLoA4KpY/zr4mlzIMUIJtKQpiUOCIt34d/XB0O3f4VyzEfhkpPaPlz+V1
R4OLN+IzN5DEoQgPbzVrC+50STy41wz+wG2fwnZFv+khBGmwFdk205CBjYEifKJC6/45uSdtzXFe
X3mviwuqZe8syeK4IMmixDmMZ211E7M1xdvd/ZK4VBOKqg61rWgQMz3LveHpksjl7SLr4FiQFYaN
3G+InvOdOPVb0VZ601vOSoffmw+hxAi3C4SmvOsJN0sR6fSZUYV0n2QMhAUjTDIeAjyA9Kre+AoW
F0WUaa6Z/POIClwe0cqZhYu4ceOigXPJJjjz8uPqWPVYfcvjk3vILott5z28YSi6XV2NbCJvgwjC
/4OEsdwisuu0MTs5cxqbE1rONmrWoRikooBskHn+uSNl9vkSGjiryifBDjYYpKDMoymCbkgvyQox
U+/NcM70lgECevEwhGfoX6Tf6B8FIBTNztfr+a8j/plfJHpqiHQpTGyGJMSZRtC6p2F5jFoNeuTx
S0zQYMIRZMOn5K43jwG4RRZCl+Gl706Anhc4Cwpegy6tMfJ/1jI3OcuJfWsgfRD3T+Ia+MeWD/+L
fs/zb/hrtQvKvUlEEszjqGhKnThL3JN68AeY1j29BTlro5hFgt7nqDPAHiLmWSmYDLWAqNa2ixde
vCl0WjWwlo6xyi78O7mjbWdN9f2GUFTs/4pfRzXiQSSaHgP+juhYeySI0v4JJU7BEZD2qoLidwR2
GIzaL3w/OcrR0ZFdNVamzfArvGCySNepoeEnmGmYzUYxRXrjZ0zv308fv1FAB12F0vsQeCBkTU0O
MIKjiUGEAf1mYWUdgjTYDq81FOOhz7hFeYXy3AGC6O9Ps2FFw19Nor9nNTv4E+BoVPcj7UL+CcIn
nufvVjMAf5vi4WJ3ulDtnMFTyFd99y3wiQwWhklGY6V8qJU8nDER3BBwv7jT8DW2z7t8BIISYzno
XlCKu2A03xE/WncWXNTSa4IvDoRCsRF05AEYpMKjvGYQf+/BlFjap37NXLwvHI6rmM2b6hR8jfLG
T4+Dje3oTWYGFGGeNxbu9eBD8siwc69LmLQ+W5tm2ntC6CiYG9yZvF8ovV5Cc+Mxn0vxNRycwMgb
7qm077OrHtuzUAYr+lD4YUmypGp4koBSDVgF8S4h00HI4Gz1Lc5qoMFMT94RibG7czoy/1AFeBLL
KQiPpjfFJFWobQQbUac65EK3zW59GkvhDcI3/LJcFgxufwJ21s3khSSLF1W0FvDKg0o1k807srxO
HiYcQpWIsZxt/+QfY330sTUWeTis0UVFwwOOvp3wpUKMJSyXG46WTkCGw28xKZdVVEJrH1sphs2V
x9Aq0WQlg+mhp7aatPedNrI3dVIWjbr2Cx6+LvGy2LRsQm8g6PBXMe4m34tqFBokCA59AVPhTbrR
TV9noHOVZzn+PzBTbqnqfc2zxkffsvYQueHQ9EMRvul1A4juOMaKOIjYIkTdZXBF3mn/dVqEc8VI
XGtX0p2AYsj9BJPiAT5AjCvwUOih/axfRVV/UmJ5LUWpwilQupdvUr6E0fKPJOTID3j+jQv3bBdV
40pVhwZ2VKnww8K8WjSNkWO6bGWYEicMLn+ZXyL+8hIaplKizeyIx/RwLxsUME+CiSpWduk5bKVe
YK3t6ihYTEn6NL6o4xuombVIiAXPbRcXDI0tlItGjpNFGyfcH8lWYbIfvqVm/mfoWOn7Iq0iCqJ1
a7jpc2Fjhsb4Xa6oJYv4Zlu60x7n91C1PwLprjeN7fPzcw8zGm16GmEvMJImWbWV2s6/vWLWvQ71
kS8kUhOESwQTExFKjy+qjZDjhgFvTIiR7XqZyUC8rWwGJyfH0F2BZqEHSjJhIrW7BbIUHHyovy/N
DVqSK6F54boCtbTSLBI/FDhrmf3YMuzhQKM6YUFqDra/pSvP7zCYQE6FkOB1wykfSj4BIP8ILacv
VFU9quRlMJ4aQ1hnRjBp6ECX2ihOwhtRtv5mWgRtDO2PdvDmQmJcCRjKDjLuKKOoJS+jC3x/MVO8
24yUhz/AQaeO5Uf8KwuZOG3yz9DTLA3/EanUY0nM9AY4sVlgxYceJtlJUcaJDtStpEonNyH8AC6B
dyXWPh1Udu4ZulYsmYnnaZVBRTySRc40QmM/t6fzCanLJkRYs1wb1veSdm7K5j8NoXuZzTX5SG1e
3E8sDYKwR1SBX7XWRg5B6ptlPx2ekdRpMtGzzRmd6A1QNRaO6YrAA8RmsKJjGvPYZ5vwB93zzHDp
PR6ydMViuzPOgHb8g+8bwpUx7qA4XYuY9iSJzWtKYsbNvi8tXCuz0K5+fx9YgToi+UTNKojHDmZ1
WkDYwe/GIZVidTnSmrtXhUvFXPrxm57Q2ubps+VGcKYIRR6wbfSq5cavAWcZ7mrdJKrR8W6Jlm1r
pkbDETIgMN1iTMQAV/nfqDKx7rsC/cFagWtYbAZ12zlPvJOD8JVKWsSIglFdiYTIJFdNQzDM24V5
shT+idCO0mXLUFmzTngjPc+VER5eUqPm5gDbtQUaMKV4TlyIIE9NS0wvR2mDTSnlGVipIl0AXKe8
i1sNl9DblAWAOM1XEWhGTiwNxxkBxp2HKaIQmMauUNI4MNmpCarMX7rePgE00E3pOKd838ldZP16
vl01EYxxoLgbmvfbMiRk+zrUnVkXJuRCoVLYvM47+Ul31kjT5u+L1BnIuTcQsKLEDweKX1L+5mBE
6T04arYW+FZ9+XG8bOQJHu0jQa15SySXvLj02ACuDHVgFwa9AT5+RGv7D7PVLwnQlj33AP/5YZNc
V3xhY1s1TG8gwvZOqmVZWzBIkRs+1wgrTrzE2fYS66Njhip5Ev65W5+gxRiGISMA65tZ3JlU3vIx
XA3V5rkq5vW0Had5UIIP3iWoJUbBQvdDG1Tzz93n0SZl5F/4ro/926i62R3w6aB3/ypmQWj13Dmn
1/Bb7UVBJQS8DgwyH/qp6OXPFFO8+ansaSJGis4vQp63mQgydrIYyr10FLsJvcDJS+lJu0ailsu5
MMsnBTTm944nB8uue7TzoNmWGx1kPU8spRKdegI/roM8WaL7Prumbhgj3XnMNaeweazxcsSCAVXf
Yv4y68fA4DwKj4Md/QRaAGc/CNW/ciN4SM2YpwUECvdoc1fWkw3M3uQss+/vEuKguYNVI6RnmGGG
1Lf4NINyZeB9siDsnWSBrA3S+WvxWE9eO+O3gUZHQyDPj8yuZNVQ1+IY6BT1+OX6eKDNfEt1DcCi
XD6vPJA5K+tqyBWxpJJdeEdA7O68N9OpWO1dJp2/KrLib8OjAisqh8+6ktH7ZgOOiob8rLaHMB14
EpUtHWWTsLAP/MX2zyFnsh5kchZtdmUmS4YbTNhrXkoIFOZ9GZYeKb1kxjAyvr1bH/DKIpbOdVD0
uH6i0DYI5UDcIeYvS1mFxyyztgKKjoewBjyg826tYwyCGqMRZfchgVcfDEC4vmVccmGCNPdCAcCr
XlwbIeOCkCXLRqPD4UaPTHmlf8UeWbRJzh6i2bIFwGBq5cJsiZAjW5s80mjTh5Sri2bNqGH6hI71
/bC6Ze2DYDYHD0mQdgBIkrGDejsvNjiSenCpfumpZt9YFDPROs7Q6dlyNXcldqFpgZ5txvziwgaq
PE++JYrrTmAbV09VyH+oLKKFEoGHBH0yOsirMV+TsKUKFwUdChbIVqAlQSiLfJ+JpwGSmMVkqSqp
yoS1CaWSuYkVAkQ3pfRUlY7CCD/7a/ldZyF/IsgxvxSWIMERVv2/syENMHl75WP4/1dsh6GxlNTK
ZhX6QycFWm+rTm4N3fKjUKI1uVaUlL0sHwx5KG9l0E9+27ADdDGwh1DMl01trcbJwBZ3eOO5r53+
4ABWW99nhDGQV/W2zWbX0WLyfh478kzHR+e89hxol4qvhiPwfpPXEGCC9JitS4wBzftB8utiVgG9
bASnK65BmLaa27WvLIoV6UNEijwnGLf2IGKzD3Idv64jhGHSqM/C/DQqz0hqG+2/H5MogKua3Sq1
HY5qbf1JwsTuUNjrijMI9r+5cAW5CESJ2/hZ0hLG+Wnhkf09dkgCZr6W2TMcQcW+eQ8ksnALsYAi
Zrl55rVYBq9zrBMTWg2thr1008NR8Xios1d2+7ddJFeR2yciLteag+TNssWmiUkkFkuFTIiz8rzM
drb06w4mGr+NvdJUoPJv5rCWD5NaVyH2aXlQ9TXRxxr38+rxipkq8FpceWESl+hkVGwK8PZe1JEN
aYl5gf1czGYhw1NFtndjeFZqPfFy5LqUtF4o+V5dp+hT2/E511iPQRTM+fv6CnMJSxfmSdbh9c6q
DJHFnbUXSE0/2b4YqZW4nAYbutlXc6xW9tLyTnP1plOwQK94ZCEAjr37HREu/LgUjyGGH8n/BWh5
tCdwKwhN/JF6Kmk0MDPy7ruD0vKiYL9W6zUzx09XMc3LA8kV4OF76doNdUKhYOzhiUkjWTk+kF8Y
ya9wne72tN1YZJyIhkpT1yQCES0RQvVh+xA65Ez53HGI7wjMAtKjyQ/DAp8sAt1JY79G3+QPb0yM
w4KRNqoE8mQujVCrTO4wNQNU3VCU9mq9+437eCV973Uy7CkCaoQx9oFLYzcorC6NEwcPebUlxD5w
ErPiJncnMOTCxV7xwezLoYYWpDbQGRSL2AjzV6VHhB/ASuqf3og72+1UjE3tmLvPEPYpiWexQFvK
pcVciy9BaYtwD5nsv64OKDnqy5rjjm9TdS2RY8uCsh0dGPOy1UH30brHvL3Z1cbBucWddgV2kEDD
7ywxFLpE64NLP+143wmasQ7BlqWdvnIf0CCRc3PllqZprukSIRDGFvBCnE7op8OuLpwfodpf7Vi7
0UZyzAPO33R+O6P3RwT3N9XVZORO+Vnvl7rj+41J+DRwKbMw2itT3phcII1cPLsJPd+9PTql+T82
x/87EJ/gzr+ezYUPTkf6gpULLQZaFO8Od9rxDx1evu0IXcdyvOKKJkMAI/qTY4L9/F1oVG12ZSQP
YgC4vmNOpjhVPKB5UiqOjNQnkTIwYCJGgYQn9ZoioEDIGHG8ybpJOdo/zUsQiefCanW//YZ1ZUDs
QhWAMUvli0GaXLhwBZbfGJloUv2xunefyLCt0r6WPn+nhgmVwIaHJaN19+FhIoLOBDmrnqaDdv3f
xW5mF1C5V0+75bB1z+nPjUKJEE1HCjJZdnfs+osoS+0entWgDG5XQecAzjX63QoWIVtG94r78RUK
XAMLbZOX0ldOlmnnCOu8YLP7c5+pJM/l4I0Rcz0xW7w5n4zIKpUcrb7NtIS4U2+lxEjnzljaFVoH
PfwHpZNnS75qcXTTO/rkVCxGeEPp0X0xmjosX5svNsmJIBJOS/y7z/1ma41HNnr63AwbvjT0HEh6
M0CZHK+nN81iocZJXwc9AbpyCJS8qMRrl8UWkRR82zaN/rc81iyjQmw2yNyvPV9foC3Bs1N/aRhD
/Z6fYl0ZRVdR+8re2Y9PjoB8JuHr7hSN3lbv6XLQ4t29jHj+ulMvg8SkyFy9Elzi/Zunf6llu7id
It/C+9W3TF+NXj3Nnfhum84AgcWrtN8FbHDDK89KT6kmTIzT7Clm0/0aICU2dCCdcKkDyFSpqLDa
yeOIJgfB8b7cmicoTrIeKdSzl19aYdFKqVIQmsrcn9UG1AjotpzGOYE/Kh11SCYJORPHpgcgpqVH
gV3hpuVOcJWyE84/rgnmFtgsEGp9OyUPE5yYxtJNpNBUhWn4NY1k3ZhSj8XRefcmezSNFOSqytyU
3ebrZhtsFjSa2TVkwURJlFiVyDCEB62sAVChpW5N2raU/0cttWPCvaNA+tQLtUK5RitX3Xkqv5TJ
+y2i6jaWWCK2Pmn0O8JmBeUqMcvFGEDEAPXOkwVuezXcuGl9FrE2mJqDibiTmcGB3GaapRjwqKDc
q5WY6moVZAU7BAUe6YmzinEDEIVz7lp/w8f1MWm87/H74QOQrnXpDviPKMjA65MN318l4zlFGcbc
pWqG5inretfepNO2Nd8sKEHYAbsF7g0x1YlbFORj3dWybdeA+h1nZQcsoDONTUwVB4xT7nurCBL5
j2f5yIQGwQf0ME4XvK4uQwCZImHbBHEihC5GJHDEMYufHgjbbZQpqqe2MhxzAzw+raohEhJuCuVP
u5VJwq6QthEFQADck3/ElwuDO6nraL/Hz0KoRGIWVQqkp6YVYVf3E6VLBARFxJk5rykAmkZ2Oo4w
nGHO6DNWBdj5n2wYol61ReFxCvcVMWJf/E7hzzgf9CycKixStgMJl/5NDotGXDUpO6nAyqSxRd0b
4t9RpfxDsSZ1862WKYPWRRQ0Uwk0TKdzUBN3fwdJtEVa60q72acWk/P1DXD0NYH+zTAxiIb2CLJD
1LK/XhIWYRp5iWs2CO3tWVRM3+Vjx0hlliRUGnEvwLH05uFY1v8dKW5uIKdShLAebZqYav8/buSU
nc9XBuCQcbebMzTzt5ojOXAixaXH+9JbB21S6v1nDKPX2/NSP84kQurgxXU3o9+AEQtE+qNGqg6F
o9if38gxQtXnswnSxf3hqLfUnmhdobhfyz4h5G7If8h4nXay99+xoZbTLlS97VmrBaXFdtM/ju2M
PGxL0szGKz57l+/Fhg1Gdisnp7QfNKREulsq36idJJx+mSayZ+l6OMU9qLn5wh/h8v+d59g+o9ZS
cJdz04TpDt0lg9lAF1rHu0H9/e/eq4gmib3+BA8+8dU070z5cHaInjNIKhJbXvAFl3oGNH7ZNjUz
5wj7x6lqf5/8WXtujxANV4gzNariUmq3Vx/OLwU7zffR120mzSvnDbN2EcoF3Oi+x/CzVsYMxy3J
64DgBZUtHQIZwHNJDwev/LAuftIRPyly5M17XD2aZkwmMaqugoPeICkNV4sQz4Zn2KEbP0XypvRQ
R/WRiFvKrzAzXyo7ZeQja2SFwe4FiW1u1uLKFgyYFwaIXVhOpZUFrGbobp1/dAWzROiuAFAv/nbz
IIASJ/+PGYSTvkJDlR3p4Ea79XKxdtB9DG9PfI/rMneSXxR38QHFYn8SEtLHmlSXeeNi89Ru8OsS
GKvr2gfOquwUcfTdh84JdytjRyMGpRjsw2cMTFp4kz/pKecyxmTM/Ai5E+fjq58znPJa0HltXMzP
f8jxypyOy49yRE3xfUd49hkHqNmuVW1Gx1gSBUdXzFAghjvhSbTQsR+95qMWhgjUMpFeeyv9WDu8
0Ao2YbDOtTKvX02UA4VHzL05LHuBCWEfucgl9UVelvbD8h+cwVAMQhDKIlVYFKzczxfxzTMZT4xt
Vhed2T/K11ByQjhrZ2LBheG6MXqgU+7epl9uGGmgCCYZ5ObNNBPuTwfzFt5V0++xzPPSrnpDwsRM
Nsow6ahZFjAhzXCBn/fIA0CsDU4RBC+ahDjZigFaFT84UVdzoGePFp//kceotgXgOdGBPp2XN9Fu
C8tD12ddZDkbg4Xv6m9s7jrNDz3P60W+ikIgLFmTDW/rAJ9BuYfcjFTbahjtQM4V9Bd2HbYjoWRl
xtEVhY5ZHeX1vCihvybYomRgkG77AyVTJ5zKClLZFD8IaGMAzNZEbUkMG93YMjjaNK5l7eX4WtBR
oV2frXJ8LQjKnjuR53gFNIYNvirYldPdfzr5/7vrWMV3+2fed3DOJbd/+U91z+HuCpYVD7tCc1On
20yGlQiw/Csk/N1T8oCh2XGiGaeNIWuF7JH3CQe6QQA8lXrNje/Q9jy/oMvA5s4/PVT8P3NkZ9ze
1NqpK+RnBvuSPqeM3DzoI5eJ0TugvNwDTzegRu+VOpPBhYiVR93jawGEN0z1yJFvIIdWGcGfa+B4
EWtMDAqlqvZjgK05Zb2lB3N3wstH3Uym5/AbCowZQgO/giGC6wiyVwdDp9WkMX8PVOifYWC2X6ap
3QZnMUvQWscAbKp4tuKgwZia0utY2xpSbTe26hqZ6i9yPPFovoYJlQRLSUq6T3CcEe6VevPQL+3F
KRBLXHsUvtxmkO0HclsyjgKNJCYtbzFyDM8YSp1kwl/N9Z8ScrTt3uzB+jB0nxkGPylLzxcXVFY+
NfnU9MXlPJ1U9GjZcA+Qr7YYWbJ4WGJqrYCKrBj+EpXl+QEnt57q4Qfazciz1pKqqiZyYqLMkWJc
1QVi+b7PkIw6ua/oOSAkCDNksBrhFx92njZoWW4lEDQZLMnngKCTSKgckOwQo32nhRZmeJPsuvgy
N5C+zscQo3zfKMTFE15wE3O1PHySjX0+bnzaK6YVyr3ic1VeFecatP1g+Y4U9dGEKiU/vvrzFyR+
maFNi4YjNGhkOY4y/OdrruYtilcxbRCq/r1uOblJey+ZO5+S+mHV0BdPqZSPlnTkKurElUs4/WfW
6py4REg1XbhLEyWu3+w3AFdrPgwo217wjR95HcUTVH6JU6r4QoE3l7J1dn9YHipDrjLXnYWNMVpT
ikpkygHDJ9XuG6e8HctHJHm+HEwH+nDLB0RqmtW4N4oFpWXKvtpMmh7h9BU4A+jiwiKWqmA2N41F
TzA6A4ShZka/I9NSeQoSGoqyzVMAYdM8ncwsSj/uss61GQzfmal3+hbMxKRLR1W1v74k5lQLBn6B
qg9hnJ0ilwuOHPh1+dLLNH2HJxVHYSmC67Xd53prHQ8eeQyE27Bvul6AQB4XceGWV6H7Hdcp1KAk
bHGIGONnyoPiUU2OCr1mECUtxxLHN3Uxtthgo/PfjncjpUqGfTxxUKiLtLsWWION19Mkf7tJScRd
tP9FcaM+AFhG/J1LAiPuEG57B8bSGByxenzlqzP9+ocB1dP8GzEzi+iJWig6vxYNxlH6tJUoSELt
rNYO21Q5cZMdyfHIEeKU9cBpFPWP3l2DvgRym8UKG9AF1oOeZfOTkyhlKzQ1l29Y9JeDShDLZC4y
I1Pxcsr7c3BZR/ukl0ou44qd8z+/fJXsCKQbgcnBjRhQMSpK2WtnnuvouD42D/rvrf1yYqT9PvRc
MMLSk35KyYncAAbFeuqMqRjLeQe1mR6hm4+nbQ+MgaWl5i2rD+nLRrVveEgd2tZ8pI6w6U3AcFPE
g1hEuZjBEzv5qYfUN2ZtPaluVDGYDLfJ35ZqaHdJKIXiW3bSsLX5V3FJzItXa9DsvwGJFfyjqf6x
/0w9yn8pzz688H/6D5GuFKaYAPjEzXso3vB/QMYXD9C4QloQKZw8+sX/cIo7jiArcscXw9i4//vy
9MH2ftFFlFXNqbLam5k5mqBhaCVoZOLEiMvtZFpTz30HyV0EXnlcVrg5PCGa0EvrYEuUHTjnBt0p
NUuZuDj1uLVJHe6301ILscu0vBjksH5t8W56HBwrdDVxoD8eQVpWwWtPjqU11N9vboC2GXuQaXvP
huDsWZUxViQn5xX0GU49njsB5ORTVhzC1vHm2wOt+L/4T6ZWixE6b6F+Ltx7CjCl8w4FjrdIOTmP
nsvdRjOAiuWSozWC2cxVHK615M7ivZSDNMFHZ/gaER1BoStf5SpCewI00bTFyPQCN9sPN353ekQy
5oKIn851XiS6qkZnHlOy7rfe4n3nKrsbyi9IHhgyRLANLwDkPrBh1IfLoaGYb4z31GPtrnjIbG7z
XSwcjALggZrKnKyJsdatKle4Rf8wStYIQDeIDRHWdidcYW3j8oy/6dFLXOrMXsg1QYLfzZBmVbda
XsUHcRkv0sAz84QLk4sTtWI6NRyMDTSH2U/J91ux+MM10GT+tBoXQ7IHjw7OOB76WQ6AcrHsusol
uYFDtasAAqbLwNuchWEQ4gvRIdOk3HzAXSRLvVTiptz8JOnTCc1namlyqC61LFCyuHcJwjjXS4Io
W8CWGmHsCb6ihjUY/xqfC+S2DkzhpNH/Zc6TAWBcmxXAtBQiYNE3BeiMPOFTN40WV41TvLi2V3mH
65CATJVaYSFloJFd3SDytFGuvMZ5//cpeAicAejQZQ+dLxXBaV+Z9qXmW/PAAz87CtSKe6MCIFaT
8J7u5iwr9cQESbD6UBg9TDd2dGwwqVKyuDrv2VnMQJ27Y6rwF5pH7cMm56YAYQ000D1GNRYWC45b
VTbbgadccD0MG6UoT11jEJ6QIx3cRRA4u2PlFxaQykuCHY8jKxRC1fcIlDP55tu3+CvNFRXRCJ3r
2r/81aCqEa8SocSIHDXqZPesUPA2wV0C0F/D03ptoyKVb0lt9GpuHe/fc3uBsKqF4YJDUmRamYRn
rbC11lUCKmYin+sl9RTtnGkrNOIVIkS4+7QPyBuu6+sJgWRypE6PK/5f1xoXfCebkYtffYlCxhVv
8dhOBSpw8jHNYHOq/ZjOnMuBOJ6cEeody2ESrAO4+JNwlCml3jtMhI6wAVFiyq5KZwxVnSuGnV8h
jSo5uqTaytcikCTSwz38mAAF57ha1BtXWqcKh6PjRB88QwzmC2C22mz8XYDWyBF2LqVkd9lP0bDR
Exlb4acvcAjo1LDH69LSXwWi0VhWYEwCbFtlKgDB27h7LJy6eBjCiNkqHzRmN8uRu/V+7TuOZ0Du
Sx7NCPwT/LT9dNcU8hwfdhAnPeeBEPwnQfhcirn0x9+zHPCqPG4h1LJfk+N9dnMUr4+e+ii7MG5P
HFHVrK85Tc8c1I5zs20Aq/0W0uBa30RZKhJxDQEeONFFTV3wnFjj1klfuZaoH7THT4ho9XLd+iva
64uXPbZ++n2FV3M+D3fKoCV8nbZD5WRKga3/lRwVmHIgNNuJ05iYGpcvBwuQ5EJ2l/5aUn+NbhOu
r+aVL24VAU0EdYfAI+/Bp7rjBJrKZvVDT/NYoxNzzSLn80aaAzD3bhNdG4auXmT2wd3DbOJFw2Mw
FcMJYN5fg5mfWTLA6mHFgrBH1lNhMQE83j3UMCgqUCK8mLiK93gMix6KPnKwczuj01rYmG7BEyd+
OsTq2I2Hy45eXA9Ecs8FKgPdqQQdkuYqn+oRkbCXt5KZgKZYNBCdNFvY6hdRCLKw699xoTHm3zS/
EBaJrDqpdZdi+K/WfL9xHQJZGdUg8jpAwL8VdNLHyhJFSpEgIE90Br6HrR48Q5Ext0FmsCSww/+e
+FFErrQMGfKSLPiYHinR+NFxW2WOFD1ksbLm2Gj5/W1KmSOb2N0gP2RyZ4KcyoahM1EEesMJPjqg
G2GrBlvhkd2LuEhMN+mpDF6OAya1RuCeE13tL6nBym0b1fLx9W6RRfZIANaX3b0Um9+muZ2NDGIc
5f4svUsH5jwxr2TpRtS4VWs8LMejwZgRzz8i8MmsMg0u9IyWhp+QwI+vOYqtl6Utx62etzj1wZBp
agkq0oJWoqmOLCEKnUZ5hcyq5cNPqyz61RIDTNS1A2KMmR+rdaJVY5kqqbNWmPPPQO7nRpkwE8I/
I2D1DPkfWpLylgepNTgko0oXG4wlR7XSo1i7HLpz4KMZqorAXUd/EO0GqpdEdzthvPtHxC3yEVvA
6d2GrVjVtNfbsHIDjg4ZY9iyoSiamySLoXDoSt/W5o5X/dR9Pnkeh1aRI2hzCg3/wrU7V5/Etlmv
k5UbtGNKZYiLXv9E/lZBlKREbRyohRNrU3v+6NCM6zApDUeeeYXub95nrE44xm1yKeE/KaCal9Re
Clb5e8so8yQGqASLTx9je4vh7yLu43FPbevVScjdQqUu13c6eBSWtIOjy9g2smd6jdFxcpZiibwW
jpAE7O0wNVwkq2jkKnijR8/Yz406Wc2d+VjPMfxHOFP/wkMKOT6ZeN9grbE0yrEZVJmnsh/57JNV
0VNqxZTrnfkDu39Ab/qZBUID3qqoAVAoGOAM/EuzjdiDsRVdbSr2FI9zRuxy+oLVyOvb6OO6QScv
p0kUKiyDYwranGL68YhTnDYZIjVuDTbkWlQHhAvHf+5jV4yPsZE6izyrFEy8azCT7Gp/4jHYfIdf
GPpexCRHcp27ikPSz5+cwr6CJKwBAg9siIIn4tbn+dE/Td1tOhXc/jd6KT1c/0SA0uPD2sNp8eYr
ho/hv8rMMaCjpFJYtTWP8hKk8gKvl8IVSzK1QEhDqIahGgGMPfC70szE9dlYDhds16PLK9pqJWav
TVScxWypOwpE2Q5OyFrJjinWedsD78478hF1YGUD/xN8gZRs8rlJBiBxympiEq+Yq27Sz+s4c2Lc
Lg1HVB421dvPpq61dE6IqB4H6KsMDL8e7GymXEwpKinPCt7vdZf1M4612nhyNwRTJTGNDfiNyozg
alhu+cHQUxKJ7d6gGt7IPTCDECEoslza+2BMhVXScd+BWD/bcXnePt6DFgCu6CBFH2aEkAVKlEmc
xlhWWzDwJ6BvJnYNuQEo6VZ1gRnknJbYUcxb9eoolv8vGiIT4vbZj2/OnVvEl8Vd7IwtxDa3lzJ3
mXxSBr1RA6ElU3laEdvtr4qzOzDvKGgnZ9dT9vaLxtzhq9HOIJ3/ETb3b+OOQ8Y95XLAYgISTPMk
wYnXTc7/K9ZBXI/mi0JEGyUHVuL46M9utBerZAxusDNd1hOFj4St1wdAJzUivGthl7XF6gtq5/Xg
Cty9tO3fF1tDv6d3KosEsMM4RsMbs+Lx9Cc3cIAG1ljYEXNuP6XxHLXPGK7EETElM/V0oUG/uWEV
PuyYEtAIzW5BoByODyfTO+l037lU/sUtUC9z1pzT7DtHMuxR+v/JQ1p6F65dKgg0UHegixv4ltO3
XkQGtX1KZ1QkPahaiiviak0wNUkxBXYMBPIJcSYI2YNO+go9rCL22EpdfBUxDRyq8WZeyvOQlfJ1
/ys0bAHDZZdtZ9+iNycEbMJagZkZuwGP6Ha9ZEubnQp7ogbPEHUdmbaBtqqrxiuhHBpJZV+WI6u6
oz4QFwe7HPIBsd/7EgZdBjNC1V2jYhb4XXn6nBE7u6H0AMl6Y8jjhimT8vVemJON4kgaRlYCHQgI
GcczdTUFBWyr4PH4O7QevCNASbS2W9O+QzsqCCwh8cD7UVnpEVsAR8N7t/pQtjxLNwa3rwiukpn2
w6lSS3y800psUQo/u5pUvwneVI14uQzmX+qcERg3HgGpc+AgwAssvp4NqOeKnLV3gY/YEQWCPFTd
0XP0z4xdAhPrhkdhV+RgCH+ylSEd6Nboc7FgDP8DDnucNDr5LyGujxmSWheDjL7JhB+DIa2TjpOA
o4ghEcouumK6dwQZJqfMXhfp7/SEj+vi7BZBT9xRvD7iDJWGB6wcAFYF7MeT5KgFCqqrXQrxMrNA
a1x5MwuQ/tbQUe0zzw/7FSHm2v8SgRxqq1j6UOIXrPiGrH7YyllLwFUkRvZd7IAZpA9fn+bPlaS2
c+3lt2BotjbB2gkriEbsF+lyGZzgw5AAP+RUzNYj4L4fSy2vbV7b1whA/AZKCTseLiA8LPrPuTT8
yc1AQgszpxyagi21IDOEgZt8JHGJ935agaOAjUlaDtVd0ErKGbCkNrtzeb4TtwIjX4h1EoXnaAti
gykyMrzY1f0kaWw1IWxpHTvFkB2Te+BV/Dq5+CqFXOs/w4nC7X08NecFxzEAuPvmhSUiItlgxBWk
8w+M4qcmHYBmDf4BqBTx9L46WAeUmqqUJt2xXJkxEmF94ur37xLgF+lcBpQeEDOFC2CUHRjZ00qO
507jN019NkyyV7S36Re85SaHH7g0uxTL5wFLRSI8f0We/i/9VxeJB8cfpTNadcKgx75WVQKEwXKD
i0KlRnsjIgIbTzJpLG/88vEwMBdgL4IbEGU0YoIsU8FhG4VfQWhmw6S/ec/Arqt2TE3sUo56jb5Q
UShtz5ISPz2OPvW+lx7FIe9cvIy5Ui0E3oYDAHuBG/FBoMUv9RnLVx6tGrLMvfy3KGv5Nqh8LGRK
Hm4rF9/Hy2cNjxRAeqvGG+B0cXcdHPVNPSCyo6IdkLdBQl4qrK43ePgkCN8IXBV123GJszIbAf3X
TmEgiIGYekoLeCcTTkRUeRYypDLjulpVtKX4V6Y/3zx8LnUAZGIXG8wMjKEvVwCAvCXPjctmzd+c
PAxEDySGy8w/oicH42iJihtMM8melodJoSL5JuSA2i76duSCGEBG3xfQlh+GCGWvG3/s523MzDv9
9PpwXPaIBXwCYxGUpM3t/o3l95ydFi0F9vbsAJmX8LoUk1+U9sfpciD/RlZxGLp1vblly+lyIcs5
8lMbBgfcQkxLf06DNa7jrYKg5RTAp9h8NHexFLTRfq8D6AcW/f2ejOKd7zvPrBPFWOaMoUAeeROS
NPmLEWKHwYNXYJLHxE1z5JQNNjyVTCsRBi6fPJa2dXpwLcTC2XkT2NTsuuUDur99v+DDdR8zREIt
poPsLWmIqaJhk3JwDwlxveVB3QYM3M1YIY4cPQLbi7YmgB4/yf+/LPlB8MGrGEdJ9HpC+3GQivL7
DD9Q6tMG28dUG5wK6Hq+Mg0kByL09OUAvnbQJCWGEnICc+28M+A9g6g7vXj40dUFoYaft4i/KJqC
TQmpL1NjO0r1ztccz/XZrLfZDS4n0Y028F0t8HQCcO98T2fQxUzPLYEPQ4LJpbSp9sF+wcA4fKIb
DIUl8ZPxO1rUqu6JV5ja6eUKbsjrpTqs+gLR+fKIqcEsXuPGi63cxDqLNY4zI9aGSE2imGaLB3DZ
P8zFpVuvVYX9mFKW+lRb2d8LgS4sIpFM5XnPKWlgT5K/1m9/nZX4JI30BKfYFQG7D9tWnotRgLRk
n1qCohNqFHNuVgqzDNb3C1f9c5jkNRLKpyeOA5h75w1QHtenCw/eo5HpJZjvibi0BYkriU9Cqf0i
UbUr2M+ag6b1BDhV111YFa/ixdlnp7OljMks6kL0xZWRbHCcRlePnu+PED1WhH18j+oxBCr5vB4P
NGRKvkfRFUVt/VwWjKSC77K3PmgeKsk9qMP24SdMEkMZ2HECdyIyTeaj5Iz5RnBL+MLKTkCkTXzO
pHnxGz7Tx8+UBuVwawKemr4L6wCKq3P8YsvOTvIIB4STQmQK6PUyd5VuBi8b58Dyk6qDD0XWIdUV
5fshI8KvIT0iZ5+t7Q/Sp9m1eZc6LnzyH+hYdEoAJzF6/tTiJoIrUssYcBzJDSiK031y7pPv7pto
m7EioNAueILKcyjB/OUEssBYEANnmXUH/Ny2iGDN2iNevCwG1a2tTA4Vtm7pQBBXAT7zd2LskiJT
S124oB01j6sPhy4bSoUUmSgpmTPemovdRTn7vK5fIoKIfgg6f3TfSXC7F0ez8Dy5xqbPCZXS/nra
Vu1nD6T9EkeknyWYkMH+WeZASimwEFIY9O5X8DsyFzTG3yPnRm5m7istUinlmeCaxcFMAH2niLCr
r1m0T1e5KV5ZiJMahH8pl4khXrikDIVD8UYiYIzn9+EKGGJCxyuHOvme2cI/4OG5zYys88eZTM2l
GrKkOhVDg+v+tDor/NgvYUxPVGVmU9ZPhJCFakxDuaicpckV3AgWnPYDZ2LkDWUNRAdMfknG3U4t
z5GFCpNy61nMgQcUEsqGIjxv5ziu0C4eJD1dAERCHJpybNzbIUQnDvtfJrswO+AYxEngQkC2+U5J
8/S6EUYWSeBIdF3r0pOCa+YbQr5UCRAXsCQgZgEBUkz76vCUCQnPN+DUuZAFhSQN1HUa8rt/15+G
Pqr1daVF1XFRD4ccfnctIhaYhNH1a0tYohN941jf7rMApfLw9pRumIskFyGEVQ5CRV9jyrwY41Qs
y2GpWr+xqgYqoiXmK4zV8QhcTl4KWYGz/Ape10m6DSAhKLMeSMCxfOOeGk1XuuIuyEG2BT18bU90
DxEfI3e/LcV8grxZAxeqe6ZxOGlaNvlqIA+nPDopOcrNmmHCfiVxCOc96tNHC732JKBXnot5MniC
Z/I5Cxk4QmAOOfRDMyb77l2nkUCExCx5hwwYQjFWcAxQNA+RPmUDv4FKi7wP7RUPuBdCU3mThxSQ
grcu/7dQUrfk5Y+mlYiRLrplNKlunsOO67TEhXhCro5CPCy/gJFvzQoDHFEiTsa2HTOw37Uzn2qV
cEdvg9A2WdoQKF7Mcn8QJwrLq4A/a/Uz1tjphCUnmHcXcdiqGmx2diQtPFr90kN8nlZU2EOYxM6b
OtJkga2UMkN9UyYIjbd35vP5h/rb9C+b1VKOmo5x0MJPXnsvl0AurF8NM2MUl4tni1q7tsF2xCGg
prv16l32MFTbhyHhNVl6+OIdP2Xfwh3+/IZ5hOA7DUpE0NdIGUIITMmGC1GDbgRt7P/B+7SNDMPX
ropER7uHqJAzfhcdOF3KUHPUnbuARKQvzFRjq+QtgHHAWbaw3HJrsS85C0216wxMhMTel+O8GGBF
j5ACsxKXCpfdW1WM3DnklmMltKoIK/1vT/lAizui/zYExBDR7Fr9FJSrmimq1H+8MqrJADqamB5s
KQHT/8OSGyKG8MxbNqO/1RGwKYXxXW9dvqe3+VcXxlqEnn2xE7QnocG7+qHx6XFaU89dhB8l6fXq
2nLedOjNI2OwiWAvo/UBKk4H4vtRJit7VrEyxDr+pdjUx4LLBXKOB36p4vse97FLysO2gtFhiJSu
0aekHYsXwLtvLimmLUUhx/ryLWGAJrwJsuH6FXkldj+KGtQodRAKMYqwNH6SedVZFFRr6dEAgEnv
x/ftEOGuW8sdEADCrxm/e03asCuQhgGdGKXKE5UtU56Xlf/VQJuxxY3ZMEc1D0Ts6HGwqpflA1KX
uTcFPYaBywSIjffCyJENxvq059jyEURxaXKrpEWE3tP0T8rUnizL5OLAo02iT7ho4KgyhL+apcrQ
QzkU7YMHqfHPsKTdcKlFeiHndvIZsI34lyvSWS5m54lpp1mesMn0qgclfWd2EYo/54tKpsS/IIRV
Wl5MwzBA795X+5qcfPG08aneBLldKSe64TV8WsuWpsO3nlSwp+0hJRKBhCI3HB52S1ErYbzAA0Oo
Oit52MlFYB+PhnwNYyJYkXUMacH8vh3mIuufhrjOsJYi5eBp0xlEY/LAXhbzbJZ8l3MOgZ1JLHTI
GTptd/Djktawt+Yb6GX9kPXeMNdBZ2sut+FIemy2cXhAFfWyqFxWOipv6xL223xh5pvitbZMuCfo
tZxFNQASAUVsK6Up1vOeEbKKGE5LBXMY/QxXDuVAewhuRDEa6a4rg5tt7vws9grU7bVbBVCMWfIX
XUiFbhTpUbhmo9JNKL50QCSv1PjpEVnbhjFwHO36NoxIDkXKeE9daiLdkpil7w0hnRMYl3mkj2CA
U0GciQYuWJ4jnbUljxz3IAq2IdOxfRX6K+mlESKdflhmPsIK2AyLE8bfTJ/DcVzgnt6x7uk9yUzi
JsjH3ddpJuHLvuvMxvyZB2uQeQWHl/8f1wRc+k2xpol+eDKOW1vN8f/vli5x2KRRofgJbBIcbpyt
mMYja2pjV3ImV6I+fVOs4IXVJ62WRvFU28kr23W1guaFni4xKt3suJSn/6JzM1iArH8eCp8AfldA
RJYLX0VYHW4o7d6LBqAH83HtlAVGDgbslJBTlcCqBNudU+xHchU5qJcCFXt1DWqVQUd+IiaswArs
1Sqlo1aRuPBY7MPSNGIOue8RcFZMqXYEKU0hRYhxcvdBjzZOTkTOqB/d7kdmB8m0pUscJ3BxaPuE
bHpEqsxt2CKMHSbQAS2xnWkwxtrW1nYZXhTew5SvIR9C4iBfQYYnqEmNa4LUfBshWvNv2gquaFZ8
Z4y3HDYy1RmRbEC05/zWu1FFSBY1m6tw097McC7M+j3feT5iRDFAK12RLD4rgLej2BgMqF5KTeuY
l5T05vMxiJfTZLyibOToLj17jQeDdBqFkVEkgSjKhpXTnSi7MrhU40zJ3vROAB97ngz3e05nBwWC
iLB52oRjmkC1DWImU+lID7SV3+jBLRwN1qeX8CHCbBg/l1U7DnYCNmVhoJajlJTgbbDGF4q6qjYo
UFe9nsXLV78YdWUe4IwWoQue2YScDkGtsemRnHvZMXgJbl+lvmdNoCa1415ZvjPvQ8dCDBt5DCCu
3ag+PqzuEV7vrkJ/i2VBPnFqXBQOd2r2leUGX7CEzzbMHmAHRwuZId/zPffwT8uAsN672jnUzwSq
LQamERc3aZeDNiATc1+HPOtf45UWQT64AkWOs1QU1L2Nw55KAfj92Ngl4apC9fIgZzJ2/mIjtLJL
Zb/75lg40RZzayv7QoLsLMGA/cKUeZc0kuUpXIHdUJzCZuIlWn9L2QFIUYP07geJKn1iHgrJlIip
65xDhYCK7CiC4OFCY8Epub9jQUeRNWr5L6DgHGpQFd20HtXyyutPK4zn2br0PvgZ6CkShWZDu2jN
tl2acBJ//Uyo6VFPgcnPeExoQHViqvG6+YzMjQmX9Qn3CMK9hSd/gtBTvaVU6l08MnRE+bDgg+yO
0TgMcoCcgOPb/at0fBwYtGmBfAjHpzbjaFyGL6RzsycRTHkL+fa74Y70A2xxZqU0cgb4LJyQAZdh
/748//97pi1Uc4UL29ZdhxtOTI16MfY4uECIj+jrzwKZmp+EAyegHaAe8r+d3MfH/hfXm6+6QEd2
zKqdQwZOgzcLAz3ViosAU8wqXpOXfdONTbVBKBZhowdYIMAT9tPC+5tXip0Kx6TUS8Ap8bnnFhM4
8kAadNTyQ761955rQGWHIqaaLNX7t7MabGqJyqA1gATnBxy3hFp4w7md7PCBFgRjsPDJWiy+jeoN
ZwCZsVGoVKGgjjozxFlwoxADxjKe/QpYsLtam1Fanoapd4y4bvZ2r1nXjjy14NqstAdOH/rkiIA9
r1cjamprqlC+u8n8QUTVdIKn5bYf1W4eYddczfC8WQS+2CJbu06XWNvSAI9GccQw+fsPS7ruBwcx
vScVd9qrbdFg3vkNWZaZomvCsMLTLevpRyuauKwXKDIIG4mU/BaLnkzxveP1bmHRO6VbVNckfIOO
yCS7XQjdaLtMlNT67YX+hpC9WRTkFuFjwxulDuPCMm++61WsxTHRB1q4E1wbqnCyka4dPWGtOzc3
1/Z3nlJuUmYjQNgT2e3EnIyU/b965j6yk3A1babj0KsveGAMiWg+3IjWTj02mw9RPFalEcbEN6TB
nTA2XbtLTEpuAAsiXTOVw9dKzR5iYZiNP1D4rhEDHs5KTBiUxLLe+6z5q9W3FPYXiy1IukiDkcvo
2PGQjQrWhPLwo8NNuC1fENrKZWTjeTL2sZ9va2dLKac62qGqW9rpFNwZUxGbcFySh9/gWKEAeInE
pQiW2PO8Zb8CPczt+C+OCMzURs4Cw0nE8+65QyVIcwoorYwpyNtsnt9Hb6Be+NuSyqzjPy1Zw4RN
bpEQdSGP0ERUvHhn8HUJd82Hi/khM0HFWqysRdc0sfNFb6Vtila6q00mbiHZxaBEu6PyUYn+K4j8
6oAGDiKKc2zT5CC4p/nOmetIjHhoOPUgqavORuGegsO8svNxN9FDJiMe9wdAIU2lvY67j9MWoFnC
IRjPscQR6icG2qv7/Ja8KPB5M8eNUBXCGmGVAenl/jwJtEr/aleGQtrUAfM5Io3pwFoHfPd2IXYW
cnT/i+XELVkq+Tp7gPJoPfDDbm0QmRIGasNPjeINa/nPw+wzFIi633NL+g+jEq6S5EcL8yz1FWDb
oGQijXdctc5QuZTslvYWV+8fMtjxTwjAN+cgP8qU5sHMzVrRz+VPgLK5bsHmAANXBP0WG5bdH6Ob
RjqvnYtI9XrLQlUzuJdm2xBasiI20n5cR4RxQvEXCUtvvtJT/y95JXjv5EZ9EBQc7BSP63cssDar
Mb+KZlFxBZlAEGPulEyS7oGVrOAonhJnu2UZEHKJvzhQsAq2sQ1WyUsmm+Y+7M9VaIsFOUBoRzEo
idk06nbwmwDgrQL/vyvUqMBOEK3/cpgHJaDnjRrpmknCNthtIwf5R+g3rL55SUidjwvDJg7HujtS
TWg34g+D6eH4S5SMtj2UOsnckzvFKBwKVGmb5O8LeoBu4p00usm60NZ3C28gPqmA5CpNSOnSsoJx
htW+fXLOuzXx87ugRAZ+W5eFPPzvuylBthDJBeC0bMJhXLjNzaO7wWcf3QZq5GP69vtF7mgJ75Xa
8GhxcZo8YDNBEMRSksQXJnCU8PwZYuWDp6rrYwxtjDBHYcUt/GRl45pty2m7CJN4lLExcIOXC615
i86+lpd2J5whHMfOMQbN4i4K7CUB0s1SuS4RscRbNbw2VgQs/8iZwYDDFAWp6Tex0mgVij8gsRlI
Ooy7ZNA7GHbZyA6SzsC/YFpGeQWJri3CbBe9HEKelBzHuV0L4G+SkESnEMlWTdabYaTB2FY7kmHv
9qd11iNQxzGt9LPQCjWwB0+fWT379VXlFFvi2nxhZFaXiBYX9Ebx+M2OY3BBKPrww795lmetUfbq
+W9HZJrIpwxdHbFRCc/JldfeN3E9khM2Cf0vQ7UO7lYJG8rc0QEbpMWUXSH1yvzg4+VdjXNrhQrA
auw+alinxjCfb16KZlOcsfwhx22CFZBabiIigbAWchpGQtyrR2cLiacakBejEL2Rx6eFdRZcOJ5S
TFdzD6p25PrlhNzysKjTf5X9gHLWtLdmi6twZRGqf8YwBe8Y9R0Nh9D5OB3n7w1eKHQFgF73tb3g
C9lOixLmQ+28J925c2qAOuzaDiVh3Ptzpsa8t5R7rHrPKF6ATXFyexOHwa9Vm2zqK0bat5tpC2Jk
168XerFXgTxpFTS/k+V0PqElLqCIzV0+q6vEP9/iAnq9U4+WoS5omTIs9GqlWCzEaSVBtQrc5b8p
Q3fAiavhEGsSpEp0hF8rO2IC+Z4hUL/RQhB+KUZDkHeopp2QW80XsHbC9Fos65GBdIdurTtwuL38
GUoNHToXZ+uSY6jqzDp8yEAhw/0EZFARujJaEcqqOLUq5/8OqnMarjW/fb8DEnNVpFyBEtgryOaE
EkZoQQQVbwo14lXhyQGVhrrwMqiO4C1ggAKX33QsHB8ad0BQ54dcaox7KGuOJUekE/5QN2Vj/XmR
NE65KH8hQdOh4ZpJGXzCJG0FNmXTmnsYeR163pqNMv/Nka124hRcqRZ+WvHqUw3GsaEYgeSwjEbP
IiRUxlUuM3EzOQ9TTKdCgWSUTuYHpkI/fcq+ppKPlW/LE3OAumM9/kWJSr8XNG7qAHc14PU2kf3V
iCPp13dKBIVe+E74lBrXURvtAKLP7oQ1UgI9pO1j/OXf+7lmMPi/LW94BHNVdOyUq+0EQv4G5IrT
NQTb7AyVJfXfZJ0C586u12w2P2s2Kj66sMkvgadZLx3btEhwMDOxqQp8L+nh77y2ECnJZP4pBruE
u3mbp30XKKiCjpq0b0s2XCBd6RRwmyxpAkVyBvDCEVa8BZeCcdrCIk6Y7lDxB9As19lVAc1ij2FJ
Ppi2tgWQ5z4PKqE8D2qUJRj2nUeGGw/uHmQq8oo1zeKuBB7m50zi/Koo7yv1j/JK/2P5YR7pGNof
0w8F8HvH0YOzM6WDMlPBokUGhg0+cQzKJkkRfsOHTPjn1RF0f9Lmg3a935B9v+OATY+WEEx98dT/
D8UpIuGpP4MXXnA7VgJLR611bSJIOKaMlt6tDVPzWsV0xmx3PRW7XBQKwpyBs4YCWrn/qBTiO4VE
IW97Ut4QrlDl0V6ULmpmvVkHCXliMFgZ6+SG1QSL3V42RkDeOE38g4JDHe6IuZb3vy6X2rXJ9EBv
X0BRhwKi379SMzgkiTb+zj0zScL8fjRz0oGL/4M30je3/VlS66zzWf/8als/gJ+xzsxbHTkwMmK8
7G+qiAuNsfIPJ8mn5UQl61oaMYEY7FeCL2KeL1C+01aDx8F1gcqGtdIbHyrLJTBDrtdV/h0vGQF6
t2JLT1stva3boixYK0r5m5pUqjGGmRMek/dVNvg7tXzhpeZHp4LArE53hZPV4aET8xhLfyCjm+RE
t01iIunWTDIitx13Ub+j2WBo2mF6yBYIohrHC3VQ9SLGwePJNjAPDDZ5TDU3Q724cMGf8hoS2+P9
rnEGGd3gvnha/3JILZHFLnHzdQyASk/1TBS8/z1KNGVKjuAzRBYPr0DUb+s/ZM2QebrVffoYOTNk
yVS0WJl8KbPfOq4tjYGDfsSAA1RlCkgDELQ+jzCB51j9Ff2W7D4kcMLonrs9RHMt7BUXw0xvI5ui
AlM/zApPVOYcxItkNqYRh7shYN96CdbBGKbeBL3bE9PFDBlWS+O4mxoVNXfC4bCErTD8odVQDma9
tbLowecUFy+FRo63Qrc3NtLastCGxQP0gR7gCTR5K/qQRVo0RzYN84sohXcA0ZYGjUj2v2hSnRp8
weJHisiZI7AsLS+BYtxWgxCnnY+WwbXSvLvn9aoPHBZ+tU2FWwj03q3d0Xj2zCrxoaYOTCwDK09y
8i1bk6UKFtz2VGkWf4zZx2gpdbS+sBDOT/0+vXFhWYCebZtxnhAFr/iiBmupoE0HiYTQHjH3kTJ8
GWa3Nnx10PQiBsGEcInGq1rVIoG/UOAv8KUsBLn4PoVXb46VCWGgJANN0FQ/blOKiiYEBYlQU19Z
EmyQx3yddDQIPYGXP6o+dNMb83+iHiIdN0t1zAKw5kyrWep7+/6fEV6Vvt4W0Hha4mBCk5qmWizh
jt4p6Nd7G7rwPMR/sYaMY5qK98hbWMTXT1TSiaG0BNh9qMW1lIA4ca0kSZUzlpRK19W2hdA/E+1W
RxGlFeoLn53jAkNIwyEjR+Sm9AkI1GuATx0dDUqUf7KxxTS5/oJIPnYHJVhtAaP7s6EVgvVw/Lxd
oIZ9LpJNKi7fioZq6v2BLJVmnE2cEqpM68DET6Kn6JhdlBNazanYKRM4MfaxLGYurHlLaigfKMkB
uE7te614p8k7rv5HXE0AAVBgKE07jJ/OGMFmPs9nLvAnSWc3P3rTgfs0KnmhEmzmfeKdh3Aii8GV
brhXVyAB+ki7Rd/waS2lzWH7wzFujFEcMMU+igfPojqj+YzMjCUCBXuW0MqJY8UQkqFLBsvC4mKw
tLA+TWD5zi8aiKGj5bs5JakKCKEiyMiTS03uul2hkpUNyk8z7tvrxdT8ShSs7BWHCXBuwyA0hXGd
yZ03/EABlSp48m5+e+yRBtDmHi9cOuSvG4AOv6/WZQCZb/uTW2MXJtI663YqF71DUByDqszv/XKW
OA9gT35/2dTbtIwCO3dRMfBRRYI5R571qb1h1A5YZ9vWgRR5MvxmQDgAMng+gyQr57FIhpF1sFHz
RzeVhnHqhMURAX2ArZYaYZnCYwIlqj/eyr3n53Bqz8CbdiPv+fKo6/2fYidN+WM6cfEXEHGIuE7J
+/wZ/YDvyJlZmmX24f8CF04drJeN7xbnhqeTOJNuQko/KOjZAzwh0b77z5OcSp9Jh36FV9Vx3mYT
2DCv9cvwFn9KXBMTkdEVauyT81ES3Pe+1vvzurK1BA+PlVnqezH6rPRKy8l/xnIFVkLKHR+Cwtw1
ENxfTPQMEcM8aGkuIidclwjlAwMSzbska6QSkAVTFoVO6F7z9XNJ4Z/RihdrS4q2vr7BEkEssXyY
mEx0BnFuOkcIlYM28C8UsW2lDl53SIsxXseDjMuaDao6B1n7ZMhVmDyo6sEB3OCFgCyfNVPhkZSe
NvtFL8IFU6XcmV3n00mSzISL/VVJJr1fhvXyETozj28jx5xr0cR5LCJ5B2PbDsBtLVQFuNyt8YMf
ojlMaXqSldnNcplY4jKL9YQ7ZWhM2ru/nbvbe0pnD/pgfKfa1qHtIJscPlSeJFWxVJj2Q0K8zxeI
p3ju9qfH7YtvOG3uG4W/6KU3fvNX9kN4X38o3blWN48nORW/+yTWXO2GCxRt0ypbKr/XwGxlCOod
+DPUYyqptFYCTedA4OxksA7WJP6YCOZpxGozcWCzPl4nVUvEN4hKPrFnuZnY/ERT+v3DaOsqLmw7
jvz8DeeOTIjZ7AZbhxNiixg21tyWa+8InQIaXFuVnJMpqWY/tQ4LUAwKdKz9bgT5Pkx8qaEDh3PD
wluAWIX+PJsg6ZZPr5whW9cARHajcDvzbQABluSP5V3SD8oe5uSJcU7JMKuw+Q923NwBG/h3WoiM
FXpa/JK9+YQpq8iERviALr442NZgu9RzTw9yz+PJEqqpJqkS1eEltJucTsfd9hI8BPXxbFsgZVvi
JSQAp7FaX2HAFLexoDEOHd802CKXkMmw27uCPo5KRi0QcyaiYPzhzO2snZm3Gnfu2mcdZThobxpn
rdI0UxGbDij3HtEA5kbLKLM7D6OqtOiyTqePc9lZxU80Jnm6oxsIhgSMVQREyzPSh0VUVp91wMoc
8591WckVdXeF7LPNygVPtptiInnZO9RjNuuvFaJyurmTm8g6zMkfTWsrzSFwRh2nLVk9176+r4b6
CpmaasLaGe6mTm60JW4WQYWxMJg6KGX/lVWHfDVSh+NnGFNCMhjHBLiRFZkx93Z0FPsr/qFrXxGt
Y+pbON6nolf3zfCcmffhm1KlBtejQra1mmY4+XraT+jdhYQK/Ajgc+tvVk8iIymBDPNJB/jgr7rP
JFI087/ms5Nc0QCiUBlrxmb9vBOuTgTxhyndP8k716iK5nkKBQU8dL6OSqxuXo9XT/Ey0dEcLDSG
fsmjrNLWqIV9ANT27goVv4mxaBbr8Tsl4jrJUnJEzNGCTWT/f7WwvdDHWROTFtgg/AUUw7XPed6o
IZMc9Cj3EcLTKJ6GE8P/1W6oMwo9LDOcquls/et7uhkQmRoJpksbbVXqwCyHpV0JGRw8I1UrE+js
qIiBE2F6xd7pHCQYIIlfzdBPVWc5XAcVJWZBmpFkogXsqY4lQ68T/JCYcySytzq73Qc1DNwpIgTb
gL1LyhtKyBscXayXp8hia8OAG5JdyYqp/TpII+2MWWgdDVwSiX8yV2NikzNANy1CiPsSNU01lstl
0xRGuARt+kuezVlqOm6J5FSJwVp5bT9GAN+bZFfMPUb+PTcUctnwSH7GjNOk7rvuOCEovMOi6uqw
MnKIAD2tBLHYkMBgdU4VQrpLU2ak6aGFwwushxlSM11InrIS63lO8zvtNLza2FfK4S1AaXpqOB2o
p0g75GGQcEshGAMXw5vnrBN37bIDVBgpac52h5QK37A/nvcHpQsqq7lWonD4YLRZ6MzPCEQDT2lO
oYUOTbp2ZWmJRNx1WbbfRp8Ae+7rimbiaHa0kpBLbraGmVs3Ki++R1RgruO83T8WJu8um/EGBGYW
fyfPa9XXtYBb+cBqymfece8vycet3SY+HsXYNJhC5D001rQJCBbUB1iplUEklnp8snujE4JMXsml
wCcaGKgnkZoqRg/cItshEQQyqxY+gnMiXeTSUNf/K5mbihe6w9KORXMwz0qEYqkskynY0dcFX7gt
qB4vXOD4GnDk9SM+uoQXg+kiU+LOl9O38++RJlJNkEE8TCLQ3nFsHW0il/wM8h1i6zPXWEa/idEh
aZwzUUzK9pMd2ujdmexpHXoYSITi/uD/kpo50HTybv+iJuHzK6urO59Q4hPiEuGKPOihr4Ch++ev
biHT/t4wxVenqH413p90en+4uN/Lm5WxKLzX+KJDRZ8MNQjhS6MQ+UfCRxkG6xx/dLmwyHpkpcVc
K2FuBGRrMx3iSTFBHG4my1hcPtIlsdBObyjeV2GwtXum1TDpGLMMgmm0Rn+lJhJL1pCk/YEeZQtv
QlmPcNKL2/o7u/1yEJGgCVurTXHxfbbXyX37NaOc7WlTLlJZOu0bbEfKUIo++aUf32xxhFHCRe6d
F8wzHwlCcdJoSseayyLlOKazuQnxpCDq7otdxDwvUS7wZuQgQOkKckwl3tgmI2SO422rtWMWkhir
nLZAGJE9EE40/f3k2a2A/+1F59y7wSYn9/EwykClLkqnL030LIVejfEeO+0vByTXSoA+pKlj+Rzh
lbMH8wpc7baElBDQPbdWGluZI3Mbi2DES66R9WzQ8kzrL2mVItdBFhmydT7BGMAQPK2B11AIg7x2
ThCquLsHOW4wEfiaRkByaMZZ+QdEHiIOC7oCHs86enoTq6aG6gCAGkTodE8bej6KDAsSF3NWgRDL
m29su3+zUPRMdURdSBv1cQ6N856AhbvoIIQkOfBrzbUl1WUPBS8C0APFAbInJjNDlkGtip/J8jV/
Hi3ovbFhwT8TUwfa53imkTbuQRHCFw1n6+54hT5K5lRUKiKAlKX29eLrLKxJRs7eLMedu/9/cj5N
QtjD6o50a7NYG/CfqNI+JdfNoLGfq2sb/+xgZthfGMGaTolD+goWfE3SL5pRxi9W8lr9etAGVqVV
Goj9z2UvKL24SSuLtnObBT98zDGczP9gyNRXyAwBHhRJ17Xxtl3nyoKx+3fZpuIMg5pfFqQK3Yq6
VyXH+XAF2iBgqOH9GOQbmBX9ONdOo0ZV+0ka6VR55tF13p+/nSiyrHogtyR48W/4u2SDubDUG6j+
VASViipEJiBWgMM4oXRkiLLOzgXvktKihiRMaQcWVrmZn+6jiiMhZpEDpBeM3P9o1CjoLZP5Jc36
OnamjjllLZi8YXKEASkFlxRYd7pnnJ2AXmGX9KNZnwlyh9+Dx58AcKH1RDbpSQwsP7tTLhdGSx0N
t00KxgwmmKDq4qzV9wEPCRgTsk6kYsuP31WJHhFaKnkkltTdGIAsKBhzczQcjVL50UuuFI8LieUV
xgEI1tdhcoVMs0rR4Q/ZMeiKqcY2cPMFItKZaPJX07lSHD6xEoWGNuHj/lxGcofs9jT45B1XnA7d
Lx2YFi/k6v91HQ8PfsiGMZiaS0JKZceB4huqeHANAWusko3tWE7Y3aggSEapjMSlAedEUB8Ir+8v
7HAIEzmHkUyjcN45Klv0//yfDVtF4R4LZjjMKn1NqxmD0H917l2dUgIhCjqk5uKc7o/Doc/QDQFm
UBNL+PrtUUWOfMAgxvGL2EoGmojIzTEcx9XXG+EOM8X1cJ7A9ICToRu69BzR7gNFHOUilvMfsANb
ICk0lwjfa9BSYOk7SOyGGi5L3ZseRajUImrksYOIlExTgW0nfiiF7gLtQys4467uNkXCTDZuYsPH
0OdLg80aAYYf8+GbF4/YSSDeUDjTzQN4uFpTGPBlw4M3k9nJ6hInc65UT2N2uDQzrl+bMGwWYHpu
KJGPpKfHH9Vx24Ir3VDLc5nrauEGIJUglPyho+9LKgqwpN3orF5IYBQJ9ZZ1rBpSWKtkvQIuQOOg
wP4b/RVU3m1R+HdFbUzBFaeMBnuzC8h8MpM0jHoRhou9tDOifye4vjf9y7XYr7elrucOXQESwY3o
5l/CON/DrruL6SmmA9oTaA8xcwmkCcpW56Z5UNs59vLnHDklA1OFLb1tJiJ8c0Ls3Iq6FqAGPup0
T7K5K52miuxnXsE2EEA2LBoNGDPybicECNspGWSZRuV9v+P4U9zJsAS4wQ1rKaRLna6fRnJS1Qox
SrqzIHJyOq3Qiho1TP3CTiWtpJHpOueDA/zVHgbeZFm3vY6PTrdvmmfVEI43g8sdUmY4Nzjs84qi
ZxUsYnwuXoSRRLigbuCk2GWR0eJTv5TatvQK7nKiQQKyD1hbP3NP23lqz6vDfQD4Ooz2Ghv1HD3t
zntasghDsqqKrn0r4kxeHvDBVj6EYN5I+eUJvaCR3yG/uvRml2t/waRFFiXduTj2ayaJpp7hxXKI
9q37F2eTu6F6pKogKjZq8CrQnjraJRsfwsv+3Cf6N7tu1c3v7l1RciwBXG2arXOLsxcZk/2p78Un
KXgCYtopmOiP9f6KrwcxDKVt1SaFUZvtnwe+HtTXpKclWTh1WXT+5B2amT0TGBKGgZaTpPG7P8mn
edgLqt3mAW2pybidfZ8F5/R68VM8OCrZjvv5+8lKaUNUXADfp411lbiSqM/74/uv8VmsSH3yS/76
llQ7dV5HTyyBQlOOTS4ZawdoWj0ylt7CMGc+VnD2czMXetuzht4wFhKqoKuI0vK30Z8MnLU+PvGj
oifuMCqr7JbU0tbo9Ty7nWWev5+yclDdcYvtOpOALrLTw8jGx6CQTSH0cfvt7farUVPYHRVa/TkZ
jjLg0vZSDWqD+0sXXUEq//oWaIWtjyD0Ghp2DSssICJM2uVDB3TKWFGK8vKTduZnUUNeDBrGmdZG
4fLq9sMEewu/2EEfkpCKLv0xrB9IZzXEO84gJLQZCKrMk2fyMDBZ0eapODZRkgV+xtjwNmOtBiDr
F2NagfpUMMHbieuYmSDxXf7pTZZ1qgnL/6DTxnyzuhrSGJBDestgAqADLciChADZXWNygpKogFTj
ZX7qqdoEnN3irqhuz7DD8U9KnWlz74jSYsVAUvSFjakJSyDzWJQdiYDAfqKq1zaA+CJYjG/akxFV
D0m/YNhvaeWOCZ2yVKNZqhMepTwIk/wck0C6lg4Kov5+0XRqs8+iCpRPiI7XPm5wiSpfWzbaMplH
QKpKvIfgNCxuXMzZgRVduuFQ7VCj6CsX67l8B+lWcTN+ihqnbrXFTWDGiagrunovDOYq7cn0eHuu
fAskKGNEgCSrUgr2EX0uxxDyRRSbMbaXlUUgx7aYZkPAQu8smbWabbyQz74k40wteLeWdl9GnlNf
tMcLTMLZJMfPu19xOpF+kvFRNZPRrKiKDiLpjsJ27aflQYFH6EsAW5HzuttuabGE/81b9Kiokbd5
VTJ17wi4OCIfa/Yl7gQyIWHF4m8RC4Mct/WA81KTJLznkxIdHPNAq8Qr43nNX9axmlYZ4EGiSa7k
z2opCbg7M4u2INYfuSmFmBI5eFv0divArDYmbJ8Do2tDkVNJSpQbF59+TRvchg5+cZeI6Bak4qVJ
Y7fSKivfNHvwtJA4kCJZnyQ9WB9pOoE5Vu3LBq/5/R0c8hPRGIMlDaGtOs6GIQoz/SVTDyykDo9x
rghkVhgptlrC3AcMBJ3n95ZUOotbzQWOKHM6yN7bdDZAGXSdDXVDuuDuJDjHiauxE8uyKRiFcOk6
3XnOwV9meZCpmOUrEoE/Hl4NhrFNcwC+41qFqjMG8n2cJ65GK/rLiUkAfO/ztJfpjLS34MpK+nTI
EPKyf41e/GmC3KzExH0j01nUXa5DgYs9Hcnketeu6Ly0BffUQf64zelQyUhfRMYNuRAURSS0hQNw
KV/dzi/cE3crM1YLDgwpsERHoSlfnRw8o2Ld+/YBaCRR7FvIOcKv3U9x0akwGe2kPVv5GFMM0tUm
1IsoH4t1KgRLo40GssdpxLp15RDabRoK/gNPfP7xg6sUVkxs0e0DlIrMxShNl8M/SwGjWn83t9+t
toM3qMXJ+T1J6SIa40BQknoRToplt7OOnsnLQYZEWiru+OV3eU4K7jzp+ScvIEBjssz8pItJlcU6
k0QKZgzYyp/8pfngyJM+C73gSmCKgS0X6vIGpkL0mp66mD+UY+cFxIT1TMEA6jRmIfX/onUz+ZRo
1qld0F1u7BaRIESQln3U/RDVAdUuJDMHYrm7EYEGkd0VQwaXbIy61AWTT9adY1cgkWOKTp4oltjz
iCp0cj5CN1VM0QH0PWafYBl2ErYwsJQPteQOufaI7kDVJqpg7G4WJwPIvfFmdP5gfUW7AxGFkw8e
vD1PTVjfBAQHbdZn8haFopdiZuthP/IzEgba2uVBnyTeFf2fZJao3wokxsQ0mMw6CnBCN9UjH6yH
taEQ3Fkv3ja1vTTNceB1uEw3ldXjCB1gkthnsOKyPq24ptoHQ8M0UgJ/IYxbqiLjo+fHxWKjsgF8
0AABxK3DNsMowxYfxDOU1SA+wukmVriNB8f6DgwSZpeiV6rivL8VxM8EjQoLVAUb3hpEQv/ANb+f
sB/kjnCpfbrKb+6jzf4EaalLOrIRwbdzXc/cR2jGTnUb1X+/uyFQE7bcYAN4GfW8PvJh7L1PkfLq
JPFqRzPdq9lKWmyHRJWyFuYKIxQCg/TYvWtLaQ2OCkYLM8a+J5P/50f30jluTgV9IFvb7VKiLT3Q
n7fXizvmKceqAw+bv9d7MiA5aSFmzABSQYm0Ti5jv1G5zs8nwnmc9PEm8gtVS5DQ/J382hp84yqr
rCc26lWU7Qd4Y3D1whMQR7BxSvqcQH7ZjTklT/IHcFOuJPLxMX52uu/gCc82Qn6ED+XBTX9tFnh7
aJ82t//NqMNkUSrmeKoy6VqtX2HrBvKi9of6i92KEZcxVwgbfU5wm9fltPsfHhT/l3A/SKawFnfH
Snxkbz/6Gt8FDfOGt5txSsRoBOn7s2ilvzm7JOCN/Hzuo97uPkYpExC7o0sC11nxsYjdIVC9atQb
SxqpRVkI1w2gcaUh/1nXNKR9fyjdlrMJp1ofH3Vo1PV83WQD9+eQuC7PTBo8zurRO3V3mD0trjAP
Lm0OmpYNm4ny9ONbIxPrOJDpGDDeFSyWSZkoJuOJ6Pg/Vc6ynPPNnusYYGW3C92jwRxOCqt0aFrt
5HoXG3HZNrhZiV6aWKTxhKd+cFr/jEf1eb5cdzWzyzlokL80oNMy/ZFur0WnxBP79QfKGEl3OY87
rNWzyioRZFlIKpnVpyeqFSrXfGOtafhuYN50olPupQcum+d0abghbIHX0ZJhFW4vgNf7DqB3xhcA
oI5rWsGH1Nl4l0V2AO6s2T1IKdTugQRNyn8xZZcHwJh7FT1THzY6cP3B8msmm50lv93DUStiQlQE
wjo7ZxXRsfimWRJASppdsPRW99/fscy5mPPzezc+9ELadKgOVUeUVODgvSnIqsIlS6zDg0EZ45qV
7PvisM3jAK8foH1QR9xw1p8pB7/SI96XSd/NXhxNDo+1j7LZmodzt9zmXLFCa56Jk34s9xN6dy7t
KJM7dXSOJTFb3SqGqy8SW8Inmm7YoIjY5ndhrdbOLkoa4AKtZShE4Fc1ZArfDzYzjV/Rwl8QZLjV
I/RNv/P1WVCrlsFkLnYMfI4qSl0oxko5fot1ahQ5z4CXEYE5/+IoGElr3+K3mN5v56sqVc1i/93i
rmJ+yxe9qLyKbYXSha9+rNVWF7AHTgvu3fXP61RTxnIPP4ElIFzz2fggWmCN5IKoCf6AXUaseI+f
4Ezi0jv68SrKDnnahq07l04RMJ50taV8wn/p9tVut+7QqBNX3zVJDvc7HW6Gj23l6yqBYsxw0xgp
SZ5YpxqH2e/UjzeomE3D9kLKn4szv6gT5RWbCLN4D8RW2+J50ZqwjHy9kCtT59cfUfKgfUrD4cmU
fh2ihhqORFlpVWtKDbArhumAAV6JERUJh8VyckDFQ/FQGFaPrtseQwC1siFD+OktvdEuFDVXSFzO
CLsWShmaXePz0hiuzo1EqWVPQ4Kjw/zZBUT2+k6aNtDz1b7DxnxooKyrm6Bno+h2Y9IV0n5fmcz9
S2citcXrzVfE3uvQRHJVFa7/pkk472grf7wrjVZ5H2hMlnA78YlCqrix4mv676RyWrIs2tVIG/6X
F9S0av9ngaafBkqUZm+ron0tlPPgRpl7Ubrm4uC3dgaI6KTmxD+i6+DHo64opqdCLANclsbXrxdt
/hc3QOWZ5eFElYsc9n+OrpqOty1DuGFrMCe6okaSfTa2Ud4WAwPW6B37InP9YsaY9XFsLnnCgs+C
Ecmes8FPRa4P9RFZ7l67QabWyY1seHgsA9jUn+TLims4M4l5nWMpelMxw0RiOF3/P1cZ3DmU5Ch+
USd4kzH1mqjf+DRkB2fcjh6bhhj4EnE83dKAYkYuVQAB2uMHlX4EGxmjuZry2GD4ISIk1c6jzaoi
mSjNYeFjfmq8VhOyLKsQAd1aoPZxSpBqPbFA3u7nWLsHzlJuuHgn/tYYrr41R0M9ZNnOlHKV9Hns
2+jQptj/BkK5kFtyJMFIymwlpEMxt/iwJeY+8stpbPy8LEAPY3sH4Lgq0WSLnTWNOxTbvn4+nkcu
BnrJvTUIb40FhPU+zhOYktnW9JMyCbzOIOvuxlY0sz8JNYjnBdLkz3cgqIHLOtp03XqxsdFkpSnV
PyJptu4vfReO4N+lAenP7u8IlosACsAqeOxV7TUl44Q0Q+sWSpCxtUi17G6rAG7gsx/+HP6n6jcB
VIqcTT7eOjcyB3saQYYEi0QVbAtasFUTc9hqjtMxrEL8bNLkAEjlTeCH3WjsajWSziax005aukjG
IwHwcG8BWMkqSknvq5w7keSEa7lSFzgByxcyDMU4GmrniUlumm8wYrSkffah8YSJXACwtyB+ETYT
rWRYt4P1Vj6MAMPxiSGtTJlURzsnYj/GGMIIFyWc1gvM7yHy1xD4XoWK6GkVIsTG9fc++4p/rKdg
2GgnnZR+uhyOnaL+5p0h8CLRweSxjjpUDe9/TkDb/OOjIz8dd1vXGuZ0BEDo9Wv9MxYfWu71e6YG
nqKwHd2U2pWeQwn4HoeU6yI7JdTpKdceprdRMTvhYI+XYXZ/yPbM/w0wT6e1EJW4kPNLomhttll0
DUQCKt6sFwMFNJ2CMViI3H0BrB8XsHWXVB0e6G3ohJEZ2DinGxZ3QrRuvOeMTW+Dg2+JIoiwv2yM
Q8evw4K8NOEl9QPaGteEXyEzG/5H4lye8TMNMvHoS2b5v/93F1a8b9NNxAMvzjKvebESVi0o6v11
TWhNUtLQgfSn9Nd3OqSf7qNM6wZiaJpe7LM2bDJ98z4GCUJAS7Tm/DDG95r1Nk/1IGf4GQ3lmiSU
c30Xz5i+V1I+aWSGeYtHLPeKVJWx3OjXax3bKuv+2wBBWy9QNeoIClI4JaPWBK4qP31x1LWRvhr8
hv8n6RrL3RoMN14OG8JsWYV+IT7RMs/rK3RpAKx+B9naW9li1XoLKJ4mlGb7NgKMqNGJ1m6r7F+m
ovpJCebDX4yvu5Bs616SxeDlK2wbd4eZyufYBxxlVqD9zx7IaGmeDIQkQ+qLNmY90DKusQb5Vosl
pX/gIdQ/+afKl0SJsX57VEC6Id/7iD5kcQE/pax7e9i5yom/6QD6AZQuLeCT5DlUOJP5PBPoyc9G
ueDM3vkQgGVsbmAQ57rqfDqMKSX7BvcFzU5n5a+rapCisLm8NtmPc0g1JwF3bd5wAccpr/t9MJRI
M0sZsmbQegtzoAk+ud6K6yse5EMr1qxFPHTPA5GZ2Fasg0SZsHQXMKAdAwo1Z0ond1YmXO5zVkDN
6o4+I9XPGATusop9g3FfkANrf8lVs/OHK2fG8s5iXdrPe/aCyjc4ZR3mrOdPnJuK7igoYckZh0Nq
Ia7Hccjpuwqs0Hbxl+GvQ4z77wh8indzMvBfim4YJZ6qbAAkC51t1bO4Z6keh93dfqjg9uXLkHVd
Pgfh1t1VbFMaIA75HQEDSFH2fDhF+1EMZM9QDcMj0ULI24aWCAhyQnAJeyW3vFTmD7FhzD+Lhzj4
tG4Gj1hwn1jQwuSfeli9NuzekvuKJLMWy1S67OY29XsKwRVTRvqbGaM+heJaITyZFZHbD5JGnz3U
kPdxeHqFmOD4EKfOUgnQlzMPQtYHMhQtXmgO/5Xo64W+Y3q0heCnvOgj92TwSV9rwgXCXFZXoAw6
r9VTfSgcMUPJdIQzOK1zp9Rh7Fz3VQMIo+BEIA8yhK4bZqKokXtQANwtmTQHjX2sINIw3lhQNZZ+
v/L6HZIuGUr075LoddCcFzQpD60hCCQ5Q1Mw4FzE9vo+UwtFy6wLUfimQtGRMGD+/rxFGr67QCI8
uvZHbZGmbiar8wqeU0zYRxlpa7zj0Hs9eJUmYE+GvEa2ceGhD+kcBXqyefomex7UdtxEtx2HC9cq
mGCurl+zXgO2b+pGnU8VO9f8alLPNiRNhe74V9k+BRR2U2Ak5nw/OW6N9xAZe7g9kuhXl4xPlkjq
YgXseggwgmPQkBAkiX18xRLHTNEg79gRlUHrpOBcQmFPscYHUCfu/xKFLJg8QubtrSTQlh7o3hcx
xd6KmkVgy2YEvfOBcygHidRvrAvQzke+JQPMk84rGV6vxpSOzmgtyYZWKS1TiDf0ARq+MoDbffuB
/mgb7FEILolkEO5pPPtNLZz8Xf897HenM2AataikHGNVlYOod5UaXxSH00otnFBSlOi/BWcDMsLj
L42DfYVxWbCGfe3i6oeyDa2aruFp6jlRPSkbuNj/TeoKvYY1AALKRhTx5Q7sUtLEfrAiF/Dsc3RX
m1s8f6Ik7BCC/6MqUEvFPb3WjL0bQqlarMq8Pj4tgREb9/oPmNY6rk6ZchmorgI9LkcOWzx59jE4
jBWAFDoDuOipK9XZYVajiBozdmzjUrq3kTMrj/H8zeND5x3Dpn1OdYr2t1qd9Enr6Awdw34hHxtv
3qAd35YypC2qxAdobEC5BlTbjQsqArXSWLKPD9suEiQ3iY56MGBOLKFIRrH2x39ZNTog+az0mPiN
mKkrT+9IbYPj6z6AWxJIFrkGblFy5wJEHm6wwb63OYCG8kzk5aRgUbM23FEf5eJV7xT4gqoMwYmW
lTIcWONL6bVnyuB3WosSfNBajsV5RQlA8BNAa5nRo2hcLjYIqmmGOGcEMP/oXCe4yIYY0vbcRERB
sF2FIb2c2x6QYtAQR9AW9VeieKuuzyBy+HpObPvibzygmjZru5Z99fEsI4s1J1hfkqlEdXQz2iwo
ZUrVlxH2ffNxS74snrX2zaGvFVY3Cj9//59B/DzqdTmFbCvj6t6xTgtKMlnZmrqxHZZGH+W8nYE0
uD4rx7MDOs0oN7jGROqJK+GIu7YdhFMaGn7g5cLFsJ8i0RyYrcg0tXBFo5qgqqKXkoKh0WAyYgVu
Kg2cTx2EbWzO2cOW2ZpCEFZ+f+3bCVeVt2bzmo2fnwiQA6IuDeKp93B3c/kkoiMhaWpWSv4GUlPT
l3N1W1ghxoKQvSkWUzB2rxPd0UAA7Y9+hKbx91nt1ZRPpyupvCT7IQYNEit1NziRdRkUt0kcc10O
Nx3l9C9hihuB8E1jIvaVlufj6C1577Vz9xRZALBBREsr4hjb9tVNbUFMLeqR3cWmvo4DngEt7cd+
blsfBKi88I1NPAiQDazUwhRGTeizKF2Ng2ulsgxXapfKR0XGcadeSgRu2YqbdTI92JggYWt+1TOy
5LB6RUy5Xh7WTbb0L90GoDEwwSCs/HZ8EKvLR/QHgNLZezsWRe6P1xYTB0HlKbcAKSni7hWjZXay
8LgUItDabhFEj6MchRN3TugDRi7ldPv4zdmqB8gsy8NGoVa0o4hFPhgZlZ5OJFVMdeeRMuCikFcZ
JejVkDNo+1sm7Pn7VlWgYdO03HOpcSZ/pQT/PFQ3rs1Q5ZJLwF9DROlq8RhL9UE0CwpYaWBgf1+f
OojHNLZFaWbEuzZJsMl2ZSM7RskxZVGowisgO4LyoSNfe8CdFp9mv/KaHL4Gw5i7YN8gQl20ZTIb
B2+bqKxkJnl6vJi9Y1icQiGHaEYnyR7Qebjq3eo1/CWC1Qx5nbpfVQn1E/Qdg7mumvzz2c3ZyArL
/SKJO4vAPc0oQUbtnIi+OIrobFkkdG1oEiWrzmE3gvp0hGLlecKEYN7zwXWtJM9qm+CWJE7/VnPn
UidehhLpw6k5mio9mXvKWSNjwXxVnkiMmuoX0TPhOWevN5MG0pjc21VQxebQKCIc6AmqiO7hdH8s
zPxY5Sh2al1DE9Dq0RSM3DQ/bSqH6L9RvQpy6p04o0nSBXlI3K4rhIoR4U7JC/pJayTsA3RzdYWM
IEeb2rr7Q9DyuzqVGpXl5/p1y4o+XOTfT8IN3VErscsbi5eXr7iv3Kh1D0iY5HqJLSNH8Qn3XxrY
Qh0T3H+0rKMQ4bVT9tpPkUS2vWPVAqXm55kNcEf//W+xIOQqNJbwRdOZ1F1I4GVFpiiIYmWO9xjg
9qpwhiJC8bfdjjA5vFF5hyOVBR/Cnjp0iPS3tumbmJCsuJqk4MYOzvvBqMkiuLfxa7RaQwPo7GNK
UFNsuKkfX9PLaHD66dSG/WWa3vqvmadbY28EZvzW9jXy+zxXkBeyh988rGrU/jde8xszyhsRjUqy
BLhK09yX49R7vaCee9h0tiW5fXpl/bT2YpZpjkqpTmJTkfEqPXWDkCGmQP52Z6y4oHcOEBZkXVI1
NQNY2OuvBRYUm5a/MLr5sVl0EryeiU3H80vkmYwGKkm18XNMrbqd5Hsy66+0NDrDXk+eGbHgIUMY
Yb9ywk4KDryuatf71CHk3fQwzBkUmHSSHLLD1rdaDUxXVTIQCAzRmY1jbrH+23N+OAMltXielXw5
5UdqMY1syboRpkfBMexqevpQd/ScDXnIfR0103JFBd9yGfQ2KsXalY1hUWReGoo+R3d4hZnOoFVz
2y+gh65tINZGueCPDeUZJ+qyqFm3Hrcpv4bT9QL3rX1D+oj5ja+/ZaaJbnvvL6UOdzEuDAcFCA04
GKUPeF0zalDj4l8ZcwFNdOLXvuhFkqjfh34a4D0N7BPWG3wco6wmPC4zE4yors9mWfUV0l+UJaQH
q0ukiakFUGfv8w4zaK3eEKpJhWFf8ZRlEYPznJuOs55ko1+tUq6fTjUalrDWeaiMd81kWrF4fAA2
M9fO/x24JVo+/j0TOUC3zzPw6t9mhUoTQsH81ozAdieuVvA1C+U9knJPmfOvlL+HosYtDYaGHrgB
OcBct0/Ln9G4GTcxxrVVBGxTs8K6G2WupPdI/LfllDOcJQMzOJj1eKI/w/5xPh9zmgSnu52u/RQh
K0G6pOY3AcfI4eIuAp7KSKUGSalwiEXly+fUtsOfpVw3AdOV4/XUTY+/URLy95yvGBZm+2RK7EYa
JoUqt4jDelsj4+eyjX/QYBaPxrFkRXqmTbb6KrH62EPKT2VDKwo+Ti8XKdXYa05DciCsuZ2+TGKW
LbA0HXnqaLGZW2YJFSX34n2vq1vliGxT/Fpz7j4bidXxHr4j4fOOgqZ5pzb8Q9UeFjOplzWficdf
Q6M71u5g+ul+zJbTBuicB8y0zS6GQhv2+pZiDfZfd1Y/RFbisu+0tVXQKGjju1QSiOeaMeYv/chD
P0gRhQX8r1WfGe+IykxcZ5ih0un0MzvdoDfQlDM2cqHg2NmCH3M3DSw+9DEFlnm3Y5Q7i/RmX2Q1
oqgNrJCkMitfsUHTRjPhakfUfHhsa+tNpAsxBz8d17UNWgKuC9Zi/0KEjkgB+WGT0qGxWdp1Lhxh
eR0/ZCsIYku4sdnOY1AwcAoRlgcw/eagdGKmzzIbWZfMBx+RGQf1z7/tcO9cfKDa6COdMWUwMLTC
+7JpsYaBw0JnYLDNiUUaP+jVmmwjY61cuPWjtQMWo3bqEqoZNZJyW14b34W8/vU4JAJq9ZhJxPKc
2tO26w6To5qMg467qTo3/OdzhFCe91Ubjjw3zcT8vOCIxXlG1pUuxrg6k8X/jVtyzynqSYm05eZO
V0257By1zPl0pBWRfRY81VYolIZGtvTY4HPhIO890rTxZUwHjmNIKU/fUS1+AmWUDi//ASwwlgad
OQ9S+/F8v/r82T2trG5d/DAQR1hdFnsaLq6oRTHIpM3EsrMZvIjzVZm/QBlSRU5BHDsRlruxT/Jn
5ak6LVLeiGgAPbo7jEcJbBAl6SOrqt1SYxB60IR73UAgB6rFQdHMs5XMhkjInp8GjKyjO789EMSE
gArt7UdHdhh3DhoU2en6qUv/HdDfuSPVgO0p8evxIMR+cMKZ99z6r1tdbaqmImmivYeKxgMgySXN
cxyx8V395Sdhf7kPZt0683C9UmvOvHuEc9NQMlzKySfFBcJCbY24bm8Zg+30+AIXIkKNfo/5aZX+
Y45O2Ym24P8fnmkHKPck2lK3laSbfaWuXU5rnXhBlkhFLCUYCmhbzTnwpaZ7oxyJtkLxkTlZ/SPM
O7wdWezlFAwvJw1jevDT2CT31GuSkXrhemmHE5X+Mo6MTKmaRt+w2j3AYvfBMLmGxB5xnGG4KX6n
ttXaGSuI9ZvQEk4RC7WhVLQU+CftSpN87hNZdVXN9FzCXogZBa6sw1iZFNSEvCM2jIdFs2vw6Cwk
R6orl3vMhix9J14UY4SPaBh+/CpXOjcJ+b9y8gLRKsQqzKdON7e/m/v1UQaOLwPeW3aoWg4nnWjl
wF5sbbMmMhmJgwmr37WIxe/971GQyPp2CSISu1hnLq70lF+uwS7P8VFhXv8MGm6fxduYFSPPQgt0
fr5blG0qH//098uCkHc/804ceUb/J69Ds+sPNkKU8oXZiO8Jx9bf37Est2utD7zns8pWYVJBht6P
Yhy32/srosARKTNtizVrSlH7XQFRphlI63V78bFfHj9GRLMIaZwU+w9a/WKWjZ4if8CVA5ZPiv3z
u/7XLyf795dj3YHktx9CJzg5Uf79rZZy+pd+CB071IcU/xOZl+iZ9EEHddspV1GD93WOHS78Ojjb
vRzSkLMBSvZwtbP0FV3oTziv1CIbU/XaRAo8hX/PFn8f5gpOMTVdbd8RBqCXGK8jGr6w5KnoZXcN
/M0xMVpNvK+9YKDYL75WmmCiXFLs4RQfnIIeeT8NV7ILrrrHr73WMgIpKlSvVGgfHoQaBkO45/qI
eK40Hmn0+/vyupCPKyH2AMH/TzZLyzQqrIwFbLBY6vp0C0chiRGztwkv7kvHwwUjvs5gOUjARvaK
xPvxAgvDnLr2fAqVQIesHfDU8okMIitR073laWZorNTaaqvXCqcDLPUJn3QrXHtqBO7Nbsw3xYV2
jM+cSuoBuzsV0MRuPjbw2w9StlP9tqDgB8sETr1fl3qMDvuU3KYVtfYRgRcVlp2U5ztXH/mm6bWd
dVg7/7wUR4RjvtoPUGKU+VV3J0ETKHDRh9u5d42cw7V1mV8UGeNSwsbbCRrw3lcAm+KKT8p07MO6
xnhF8/EsxjmNWf3Qxifwg5vY7faqpXHL4/vXupYRY6mrqDdCiXnCMXh7K3UQJ6NPXAowQ3dU/mxG
zp0YwMVY2F+sdliO38Ynt4cAnOrhhD2KcZEel0sUxhZJ509QSOq163MpNPo57TKBjkdcKZe7kA5q
asp6CTdCSRNOQVx4en2V6eqhXbDZ7xzPHqBeFCOOwCwVeAFKf+o2hScwczKeW76ra6uVWBlwLofR
95mfroRR8vNSENq3fEX49VLM9mtca6FVL3UwVvaD6Gz47yrC0s6oWyI4vhAVcBuqRkBFiaaf8sJP
9GRyQQR9KnCKMcI2Q6uinb5MsyB2i0MGrdO9+BVaGNRQ0MZZoS2uLvvI55PtWGNU4ZtaGV8KgRDb
2Elpb3s4fyQmVIPOkDm9lR3O6VDaKjCEOaZ3uN++8Vo6lcje5bX96NbOC2MDcNrTNlnk2Her/p9L
ZwelrbO/YVgLXO1wtx+fkFdIr70B/f7tXXHgCEUBcQVfQFeKe0foNcwfPpwBAEgG3jx8vVPoyUMF
Az0MTFmgQrB3BleDzk5jubmpiWlK6qvx0wl4EmsX76LQGB0YxetfqVqBnKUamMSfFR79OA5dl/aU
WM9kS8rM6sNA0X789IbnKwKzQVfXbsH2nDgxVgpsYjRkLJO9GDfs8JdW6pDTvDh732NVEPhrXazM
Ls7IpF+FpEq+cDIt2BBg7lqtOtG3A4OwcYwp/fD74AVHXpf+HHCcZxsI3bbSiksDxpViS5Vmln0Y
0weZuKUcu7ON/D2C1vyJJ+3U17ptujoCv9xX8Xm6nNT/ipmC67SvJwHcVhWj+cjKsEcjIvVBWVl1
czo2rqjt4bTMpWlnqVogFO9yP+Z0UW4NEeMhiXLlVZymRTcuYz0vu64Y8+rTjRudARc47qOPpUU1
2bNog2sdwtBCCzhOKYZcsnsNNAjWy+5AySyMZJyY92fM5Mmxao7f9S7Z0xuo+3piNPIOZuo3pDlF
rJ67YVmPPd8xcsFcXoeFEj4Pu2egHt56NotnVGQ1RPXzYUfQSMgqToiKUGpQDHeiObeHTvIagzcb
dlKyhAiFRzq+bfRcQtXIsn4wbmJ53YxsxBPdcupzhkh0mDIMGl8Y0FLtV1IK5sOm0wW2MDL04orF
nv/U9v+KltfllkNhbpxIAc99xM0xIGarr83ya7s67X5jzt95pTxmJGY4At6lhopB+XyiTOH2xzV9
Hqoieb9CN8L76fhwuaUb9sZvPLc45NJ1TAduylXamky7dezP0+KM8/PPCUwWwsqRM+HxnMAU9WPx
3FRN5DhGovpCBKOi0uEMSTBLfiSZRqE0FtLGgbOTFyncvovpmVEQpESgMYRhDNJ5sDbrHvB3FCiH
+OU2ugz6D/SkYQ2jc98SG8SVyMzLcNFd4/k7NHIlFqdn3r2e4XEQDHA6YJNQEtSZmP5KDZv4LWpx
kS6Jy94wkH1tWWm7QVTmUm4Kg/LUsgB6IJT+T7jVUSUHm9nvFxe2c8S2/oRG7OxqXS7cp7ItJHnj
IfVsCFKWTykgeNcjBtfqvzrl/YG8lk2L+qOrx9BX8H8jhFENoTHkTQdJbdLvsNf7bctUMd6+e5O7
9zplKLgPwj6JavE2hKrDv36H3pt1YSCaSVOeQDEXMFalkhjmZklOp1UAmz93p+Ed3Z4pJY6pQBEe
sXyc9BVTMDbicvMxieloRsiUDiMTKDLSWYqOV3K9RTLcLmL5yx51hBN9jATanL32RqLwmSXmkfzW
gdrfWsDVi0mfzhglbAUDa/jLi5TzC49Fv+0tra+GOu4X31iJbH4uaQibapp6gYeYfFBqZEelXEsQ
peeseAhqndvlASmLDOX5Vc3LlDKoe6o0yVP7pvjS1LVqmCHWQvphCywS6C9l7X5vSfsqOPt2lJFJ
Wclhz6Kt5gWqvib1phw017g9pv8s/mPXh4LnRlqWucoKU+f4ZanW5Nmjon92ULTYBVqbVqZXF/+y
1SxrLJaqG8n1hIKu/hZoRxVT5GVJXRRjykvATghZwRjDGsqPEjJf0244gWYs7kWdqnU4CfEy3fMt
ffSc8FTMfJGnjp6S2XvmYyRwEsDE24wwJYXUqS/ESCTNpkcUzo0soGwX/IsbilQzZETQJUBCq0O4
wDIZoo6Z7rBbr/963h/P2ejOAmy08dGKzXveYOifyX/5S5pSuXt3HwLrjCXZui1axW8UdLnHKpVq
SarTs8vok9x+64unSIonUZPdRJJYh3AHR2TXeb48rmRPw6QUAX/dKyhYkl1FmOnQGmjSmqiNIU9v
zvba8sNrM5ifYr6t5BLFdx2IzC49z7hyrwMNtT6gpc07F/vjfmdzz0WGu9hf9SwEAqAH7s2MlT7v
yyuXQY/+FZWhVBJkYqUSQSfV41+Fz1M7WfCUY6mpRsFMeYc8g/IMEbnqM8tOUGUJnkJnT+dU3tsn
WzCzkZGTJox7PZZtxoOzcK7pQogC3JFN4vSaA3fgvK/JqnLALnJCMs6FiRBldy1qBDy1APxFLdv/
bO9lWMhQRdzVCcap6BZqsRpHuByK6PEz6u0SV7bSZyVXjz57vzV5QJbhTiiNIcd4nlZZpdLiVIEJ
vC/Ajo/3LVEOKI+Xn/oMST5qsiixqMddKEy/FrAlbrU7LxwZElmZ7SMyrC5J6rV/3p4m/zKPgxmN
Wh+fsThVk4kIKIlg10RF2LBq+q/WHlinTetOnNPIPS1tUWG8pYCK4IiVcqDc07ZsHdlnVbY3gPj+
O6p706NTu4nk00tdEEZyl9CtoY3c3FuczNz4pr+aGV68wZO7wRxVd5+e35NTiDZRJoPeRtWl7Iw4
sDVc67V5p9jbhIr+r36DOdSsXHbpJsY8vtnDhJPpJKQoc8eWCJ7+xQJYQhzoyh1LfGgYEm9qYFyJ
mjKkOXSVJkpFTARrwHc5c+R0xjdw1qcCc595HyKjXbaM7tFMt1oSiezkchRGrGjvzk2av94ZQuHl
nrtpT2+8J5VtRxrj+ytWoBhhXQCEz+LaoK/a+r74+YIX4wOA3nNTgIA8JvrZr34wJF1OAyX4CD4R
povWiHupStvUn6z/EGTxKboMqVJczwwAzdufFsyyGb6PVBZda57O+i4MCMvNaYPQelYGqAYkXXeD
YgRMUdJK0LBm26/8c3u6xZ4dx9cb36/rqaOYGrWw4A9OuB5gGxSwhCZSymJCgPzVPja7vtnSJXdG
HF3ceqZClbLYIBEDckbyrAWvFiCObe9snyEDq89CCwfvY+KDZtd4LF9CqQiRGPus2eGgMtjAUZHA
esju3Xua184K8W0At4wDIg6gxJFVYj7y2AQUyH0hRc+ctGQYc6xMt2XPewkhFjV0YKEcDyuFhGT+
95mTrOT7tyPLXdF2LcvIb7H/4Y/IjllADk8fgGGECPtzJCHEe+MWe4WhDfuuFOwAUTgFvWGv08l0
LnUG7xxQPAQLBiEJC+wEh8+wbRn+NpLMviE7fZ8jJQHeoCLoCaWhbuHQ3gHCZmf7CCc+9yM+ggVv
aJCr7McC68uVyKpVdlK6ZeNQit5S6DrUdld3dfWc1hbaDwDjVS1lpo1e+fDf7qR9atGfYSj0h2HN
aatEgzQmNy9l7GmsbAl0wH6TjfOSP9AKWJ6qtTZQ9jEarQroR1hKYdeD0i9xFa1fpwGLTXi4Futv
DjcmK+lKvZBX846h2z+Td4oFx7jhqsk9hrmvR41IWAHOOijNfcEQel6WbibF5tq2FU8rbrEQW/L3
gIyKxscv2hoBQ+XtGlxjNMfEVtxdEZgwTbO6oVGgDpAPGzBzO0JAYVZQQlC9/woOtxCyj+EcoCxN
untZjQzN6tGdlVg6zxtKVrQmlkA3bcD/AkskLSxQTBnQKo61FKoEgcX7dpjd0R/RFCJI3gX03vBj
WLrfVCMiEzvn0qKN2Ix9CWzMPO2Mu0fPsJMR5LZsutzHGQgrYRgnmQCqcoq9+1BBdfA2FfJhazvL
GK7YTb8MH7hwAlSdArK3rS1hrhargtZjhG4E/C4NsfKO3bCIi5GSTNZ9+Jk+BgUjRWxYtAtIq8TC
CPw1EW/+hrznRy9KudxYtjkSKJS+PqFC9/LcSt5Hf9xjOZ94av1Isemtlr+r0hOGr7UlpAx27vkW
BKH5/v1gSS/py9F7w3vIjkofdd9CaaiA4ZZF9041yFIG7IJxFQQ2QE3G1StM3Pwl9853zAO4yBVm
IQK9X7VMu9CccFP168Wgivu+BBHeyGdMWcLlAr4BCJy8LK66Ilz6ZQs7klHyiF1xlD3NWEl3O1m7
m3LnANJmdTbtROCywVKnG9cVuIsDyoVdFrvJ3ePYuL78qP2cdtol05VZI9h9pBwRVjSRt2CejsgA
tJ39LnIn6IT4OHSL3d+u7AlChKOxdsWxT+KZypfeqoOkkcS2LCzSGtBTV6MJIkd8lfZU3HoNQEag
++bUuxSNT3GlP8e4d0McebTaMc4Xh5eGOFZXgAfYTnoNVEpX27LhbxtKYmdimb1Oj8hQomu79q4p
UnIK8yAHHak9uCIDlmCKzlIsdxEQERKYJHo6z35z2E2fOsv1asYv5WQftGxgTMmD865UAViXC4ko
K2Bi/yD9VvCdb0iBa9GaseOurN/GUVzxrZF/krsOxBKhCTp/0wrNpH3pXs36yaKldhc4oUT0NEW7
5LG9f3UoOpxvS+w9Y1p6dZj8IpE76I/PldKCejSHQN9Q/foVrKqQD57v3MEafLlKmk1WGHIZ4JS4
uag/sBlltD15CsKC+2fUu0xYtfO4K6zLQDNSSeQ+Ev/SFsg5EPeiDXyhQ6iwEzmw+Uh7U7PY9FIq
KTA6sfnFjkz7bkscfVNk9qj2HVFCl4/KMytTMjpl6ui0MenoI0747Kn0w3JvU5u+kW4yvIIdpE9H
89jgUXkRdjel108HCrClmGtdj+QeMRyQLHiS4h++wtMikqvd5FxGu7T2kInoYBqtB325/4RUuQl5
VDXJh+HmyMmKmlIK1T2Maw4icuvs0f2UbuTbMyyX5eeEDVSTaUbfljezAhcyZY+AnocZRZvDtbdn
SRkDFiRSdpspPdsMSPz10kxVCgWy302qXgxHFBa3mDLNYVroMfY0SBeuLN408bj8TDAj9b6dOsVz
bjbr+XcGAGVscktUE1NGi1y37h9c3ABNPruqq9xwYMxwDYrLWcvj76dV9gYnHmEhOxYlX+HWZpw4
jrg2Z9/IslGDJjb9tiEJY1ZHWe7bl2v5FMKY3cAaYWhZwtXODa3gPIS66H26CsIg15Ru+jM78pP1
tAsAVqX6vF/EEWQMT0uuu4Xj2QkM6LW/wSm6HeaHARskApCKcsfzrEfRrvDnUipMsBjDKQ3p1FhC
Eo+WEyBh3BrYwnyiR+7Apf6TXwiM6qtVrDOnGcjwdKMXx64wTNTSeZ+e6Jybk3+TMpGX0P8HGHuQ
CQe1rMwWFdEdgs1YK/idYjfmecZuCf+2AmZ2clI7T3IwxnAehOzYyKC2C65dyquEd89uITsWD8pw
mVGwuLj3M7IO4J+ABlVW8gILYuiBZhMLXlWgAjl5dsR+WwrLz36Yz25vcbVhflHV8i2m94BqErbp
u+lh3tFajbPxhoekSSYp3FTxXyBCOwB41eiadughs9oVD/pHWHkXG28IOVZdYGn3lsqGMKqjzRdp
I95C85JvZTjOMpaqkA3qegLZClXREedjE6ptH6NKnC0SBYaVPcRLE3I7pbNF7LRccsjsJlfO0F0K
fjs3BYZYUbQOJzFDRrZ+ub9Yg/vyfyF9h6I3dnbqtpINZdW0OyxfwwvtRELXcySuusocqefRg9dY
c01TBggo3sCXOa9HGWxtC8oUlHB9iYMEkxvwb1eqVnZ0MjuVJAtgoqgpTuYxgdfUF6ihdj2oivsA
QJIOdYVRUSk5fyqhM7uZVV4CyHoqw8aycPTxlJWfM81ErHEniC+uOLssvObWK+61YRGiHtY9DkYy
zuTx+Xr++l91yQJEDCxN5LMGJrfTZp/n+c5FOwbo+cFQf8H/+Z/wdKtNI/XkeamHNT1xVSmbcCxL
PbZMFHNH9QmXIRxhFacliFfWGO/xWd7NPEW8fkv/7uTDiedGreaQVlARgrQr7K1WzG9J/iS4O2iR
Etnr0l+GHPmeZTJ9E7ZfDvmwLkqt0zSIMhvhQCgdBtRnWiTW99U2bincDrHOmYNIliAQnGIkr1P+
OYVnhWro4Whmq81MFlnmwHyQy30Uk7G8grPt98xWXkGaeJV/U/xxdLlQxUfPoxVKArC/HGoefJKt
xHQ3DUueUFFiqvECpu+qOifwlFnBe3cFn2GFLCrTobWqPJO3YHHTSzelFBJtmtpJmzMa3qNnPk7T
d3oV6A8o+mOi+MiPEAdXPpR6G8uYq89Nlu8A8CTxb5qfCpVqfT/it+BvFZCqyH4XAUPMBfGQQZJM
VwEnfT997uTUMxozMe+50ylz+N+N2oaq8MF/P+waXfy91ybObWAdoOxCeUPD7X63FJrCpaloK/In
csJKkiy2rokBmdrbobRejrRjghMGGxi/JreowbnQzE7BwB1A5tYtQrr857fjd3WSuWPF80qScZMX
IPoH5AfQvShfC8Z1x6qyuVn5sw8woUZpH6NwQKtqCDUnVnSAZn0+1LoMnYBxCgp3KIrll6jqDrBH
shUggvTbaOaJj4lQVrg7Lul8lpQKV5kFM+2KQNr3hIqPQJrgd5f0n7ogffnxHrjM+mWl7iNta1Nh
RNPl2fVLp8pUHdv2ARlqVgFlqdGesW2sVvOgTrkgVyItlq7YWKgp2Rq8m9d5e+X1Xmg2DNim6EFc
GHmHz6bylA+KJqZuhIg0phFu6314quOEL4zpTu+7mWMNXvYJDTh/eXw0nZCtWVSZEO88No02nzzn
3JHG5EgnrVpyhLI3SgzxQnH51TjBGEabIGUi+e67Mj8ZxcJAZGkX9cU2Fsq/3iKib4ZQWp0UQQ9M
SDD0tTXzD2EXUPAojCiOXNSfoKqrpYRItN8MQzicLs2zpXV6V9rne0qLCAzT6YqNkltJ+Y6cpvoz
/oJWtnrNVPVeyAAj8fF4BMBDESTiEvMBglie7CrXySQ7ee6QZ9szO8Qf9/ll1KiSqawmKbYMdRbi
WgkxvREFQN8vyOZ2+iM6vDzBg63EnTY8ltPUsMLJVKMaBEHnAAI8fubyxk7Y/RaaLieT1eHMhYhk
njanP0zqsUkef94QaN3lnXu1dukScWJcSuL96RKJPVUxPgoS8KKCt3IPcw7BV1uDHFjjveRKP03t
GkhpQHsfa+ZpgYurbo/6GP2GzoYgwECp84SsL/5csYAh0LIuFeZaO41ZjpovlJ/WulBRkKjXhOxX
MTSsMraoB7YCl9fBjNU5nLkmQrG+x28w26YjCfwLWtULeUvGcj010pAaoe40XfVVJ8LsAO/adDdT
7hT73lZLhImehP0/mVO6lVFw57NDPx+C4zw/5UZQJp/W/v945g3LtHEEqAxRczqdISXRrc76WvrA
cyEbfYgf7ejVP+8mbJzMyOWcfEHPLWPWG4rilZyKaz3wYAtcbxjRTno8xJ4HBjtVcmpchnpko/FI
mfEA0ayj8QTxPuevSHCJOJebkPFAHoWp8SWbcf8jdPVai6SxHgz4SrFgvexxsfVW3Fcl0YH3Y080
Isonh3716HgKSxSf3GHjY4FssB/f3NWGrgPMH2bC7BhV9EapjHU8DRlqhvgJYYzFyjgTlnNq8Bes
49d+oen/BHp8FrEPQ1sIKZvI/1yF4MlHKpIGeoDIFsqUWDNV5pBS5ADaO6TYHR8QFpichQwdiEbT
IuS1NZ2qi4ul4lm760cUY168rr3VxRQUolIhRxxfJoWv9oia/tqY1DpkK6SkioXCyAWTlDCDIBkK
nrX5Ch/vj+nk5hhwgg068lA/MOa0u96d8fPlUeivv5UogC/VxW8FNkaUhwEIT/DZ9RRCQjbNmTAD
ADQ0Ie1MaOOVT/LV8BX4eh7kAZowL4kz6mCn8qhVHo+E+uujuear1MMdNtId4b7JLNuytLAm74u2
EpVAobnoINyBcj6n44mGZGiqU88owNxsXFWuWFeY4r0t5z/ov8g500N/HC4zMb+n82vVfi1KoKLr
VENUvDUqk4aJowwjm+t7jzqyx42aK0ASO5D/RXlDdUwzwa1ZOLf1rettLlTTarWsoWX3WN1iKfNi
WC/r0bcuNhllO924vPOc3+Pi7yvu+ld/kbNp7alEtTR2525Zyjf3/kiUQVGFbr0WuR7SCujdag9d
xGSuY0Hr1x+oSBInl78IgpYCFO8lsdAmePJRckp/66+JoC6P9UHDXMCpHsNL34CkjfG3jETurgzS
lUDQY5daS2SgRbAWSxbcJxzicHizj/IwvyIk7Q5/RBL8VnTV6/I4Cz+V/pASwNrCUm66tVmUSHzB
ZSl/BJi0rTdXuUswiHWpq4/yVmoIPGEunKExW+3TOUuxAhoB2inMK9lMEK6t1GLxmTOUqwUQLWLB
hq3c0KG7WAyHtJybKtr1L9iG0qSc+1GXApYnM81gaQ3c/XOmZYYw/YSpO7hP8O0hF+Cp+p2TD4fY
5AG2g2LDX2iUpKONF2Exw4+CEsbj17R6KcelBkZhzyd8KaTNLA40n5290wK8VNWdGw3fm0d4ucOf
3DBZbnibKMIGCFdeWHCxC8fzcmYGSwKK0fe6Ter8zJlaW5sXoXQRW8/DmsBTy75zAsM3pWG3IipV
6UtfhRdnsJNwuo3EPCVZuuL+mTRyy9eMVLfZLWVf6FZMQ5hTJwb/rJVpk/i6yMYgRHUb3sOQ+FlA
Ob3hX4vtzixmG29153HiSRGPDMj6ypP/9RYCvAdIAh0eTW3c6ejpzck0Hu5Kit3vxyC5hgYeqff7
q2BGtYSz3ez2Rqb0rLm4pNcvYuHaS7+0iSaso33BFbsRuL2lZ6O7jBDUkxuo3KCFxpRmImEzqgwQ
Bj5Xml1ul/1WMK7cG1j4NR4+3OU6VLpu73HTLn0pVBFr9mgm9Rvi0aHMkdfXyF5pQXsCmfi32K+D
bGnMB0AmS/f5rlD9q5gZc1Rk1cNnZjxkzYVc2cohDxt53lmFeoHXBXr9hmA5fg5pDzaCuzhDLyGI
hH1sH4eoOyjMtwNWemOpjBUEryUkLPSduQJEjVnOjzGCz0hDbc8x/+4ppe5hIUC7Rzqmzaf8HiBf
/iguRYq1pUtiUJR2ljOqt8e+inFObplQFJ7Wh7AGwO33abUxY+arcUxuPyJYgQMSKKYom1PAcxVF
GAm2LdWjGiDrMMtBReZVkm6m7JGC7X/lH0ABeCRVyi0t6X0vYfWqNBH/2ZlTYcHpWEjOwb1gChjR
a2/lbg8q05oEmHJyKOC909SYtxpO5p8yGTuvTnYNf9PPV0xYq+ayfhUNvikQQFIopBgwYZ5QJFyh
mKueD8V++tZ7eMze+1xAqxvPkL0D4GwJ2/7F0vh96R8NUjp005TplBSMbQZ/qGudgpuRE9OffZLN
030j2ziYvj4tj67o3iDXTyn42SM1B8ShQvwNPiUDKAPzM6Tbfvm0XWxPlse5qv2ByZmWPf21tERX
f6zXmWFRHUtBgkG0s2rFTxFTs3GSWXbptLCNpLVUKLQ+qFJ5x2+jIdsOcPgsnR//XrltBEjyX81f
iLhe12XVv9o7LWOQC8h7UYUUrzOmN1c2Urs1RuMZ1Xrt3YrspuXvY7NFC9+XACwU5aTSH1SSq8j/
lm3762wEk2vu8J5pIQHCCnqFHZImVnyy9jVo3TDuFiyBUsgDaANWC8vjwbB171SmqsRPdkPCqn7M
2ELLCW2Ydu5c9DZqxOWJZ0xIwKZX8zA99+cBC5hYzjSwTDQePovU2uey7sxSR/z7LFIw9kRy3SP2
TfB1/x20U1UGPQJU6BQbkHnT/drjTrS+vvOisCDJtPpJYuDpsazzmTEN6g74MYkZgIMn5ZFSM07g
g89ICcw8vXeWwELLtsEz+KW9bkbxR1sHFfiZgGEhoBJaqAtahR7FtQBgkt4eeVPOcY2uyTJwLYr8
6P1DBHfJqbTXj0IKi0DcuOu61mJjPhtocg8DM4meHb/u4mIz+sGGq2lAOSc4GIbP6e+sYXWXELY2
Pv/Xh9eal6pjjeI26sK5q0MbhzscJGL2fJKSqaVQ8hBbSyOUWeFhuD+bGXak2Bg13w2DE52oUm6h
CRRwNOlbAqHAcu1QlhcXSin7I1mJw9GKhX5rv6dza3u6IcPDJV+1NWto1/7SDpHmu6ijFu7shjap
orev3w4qXsWi1hUCbnAeLsQzlEeAHGxElic6Z7o5TgNrRANG3jXTrX9cLfUFxJpiOHiAlOOGHnS/
N7Zr64IDDciCUFvQyyUXJAkdLRYCclDmKkfj/ImVB2j8deFFHvQBc7PoUVYmQNm98G7L31XOHwau
Bvr7IifAGUucvyqrjncqroeT4oBF8Yn/a2+dGTHlcToFbs8WnbSm8NIWbcjU/MLP2Alaz5OBOl4P
8mtuoSm4Bgsl6OUtFq/vAOs0F03DljVWqB25Zx2Wj2ov50DfF7mO7bNmj0Vqh7PL6zLS9xLrkdvB
pkkzYemDNWEFfQPQp45XftWCoOsTVmpNV3u71LQavFKo0ALI8wOvkPaHfgWt9soeuDk/+2L4cz4O
fd5gjmm1sCf58BVObzzV3/6KooJzonEItDApvLu/q4XT1gE1m1KTGg9mDCxLgTz+PL4pIzreL1+t
5ebsVZ47qzhd+QrXnkNHOSJI5Ts3GCKcAFucsE6dKsvpcOeuPXZo1ZLn1gru95boun3XqIKg4u9B
fgfO+cof/fI5ngIVy5h+8n92fDQOoQ8/C4RNdvmKKCJmln7mQXQWVNp1E6AMYfB/8x2hWHu3nKDl
Yxx6DOvm3LTy0b+XZmBlvL+w8bn+5Uy1NYa6vy5u2XNp/b9/JZUYcz0hb99TCT1F3kx3ESBvP8qH
Z/OMpDKcGLBGN04AtNCgov3E7H6VtJ3Mqd1mMFtpzfyb1pBDXXI3Kx121z408gUxOA2bBYpTwOSW
NKBKGcqfCLQWKD/97oOU6ji/oT6e/UWPeHIzv7LZVo/3zowIzxJGfoXbOeSpGozolT7+jHU2b44L
8pLwswd8F5AMESmIkFaun2PLVCDXcxv088XQLDnEWfKFpxURWHFkCMHKY/rj1iN4ljYvxMudrF3G
x2YXue4pFtRosEKi/C47nZb6axzuP7HKHR8V0phYYInwJewnb/L33VvZwDv2TbqnTQI42cbOrQpK
yXxE0uwcdBlPrD+uvIe4ylJv8Jlj85KiwphVlriZdXTYE7jj91CitaAkRYIv+Ku79nNxSAUwQFxg
qzmG0zMYoCBTtqWGpQGMjWutd2hLpaWV1WHK+AwLw/7uvWvldmX6kU8Yx0LtR4hcjSgnU9/4kP2+
u2pFoduJvLYM8VBaoaqb1OiWTX7BOMznqVPNFAiWCXIIYD3qt5A/iq7Wy9pILi24ge7zIQJ1ovGd
SMkZuAmxxm9tRleAWxPNZeRQVayUkRMCY4+u6Pj+UdvUULuOTB0raq5RjDTR4bbbUS5wTmoBCqcK
WjV4AmBa/QvVhxuS7XfxLS1KwDA19IiDAHp2+e5G8R1ofuWasgJv2mzFS7W11Pjlnu7n2Jn2pmf7
XsyWlv157FZRhQCnlaVeyo6bf3ILggn0LjaR7n/uWDr/WEQIHf6rvLOefoM3q20hcsvfAfDSjr4c
D7wsSAcsCVGMy3Ocli8qAYSBrvxrXSkfOB2e/oYxqM2MlJs/0pusIerF9dh12tVnN+68+LN7ZePA
XtWTdHdCLrq+LcbfaeLaxb1xvCX8A2I+J4u/DKQm2k6tQyMTo/2svSYsVComo6WZPHBEGHY2TEHi
cSLkAAp3pHuL9Jby/luzniXq8MOR6lUU3RckWEH/T7vF0sxS2KNKzhYq2CIDEbVUGikM/uSwxOVW
UmqgLG11attHn0h/Ac++w/L54v0twqml5xnb9Jcya4i2gEGbktGnKn2vulpqG1ePpuB0iv+t8Psj
uez8noFeiKxWa4CTYetWdIvMsqYz4lfhMUw5p6uCNSF3ml7n3G0C6Jj2b+qi9ug8jEX2rvz6y183
Bv5HagHMnVPEzVjHumim9VDKJ4PTqLfcenfo30uICBXZtHU9/oXPEQ/1+/m9kk2RwDv8UckJQUCY
Szs6HGl0G9OemsOuBNT1dkBLiHy0MAXyITUtSsWLyPKV5O4YKp69M0OngSChlXsOR891EmLldW4T
rhVU0Wuk/3NpTKTnohp12wBkt+gPDWiwr7Bk6u4iFHt8q+xBjfuB94mWL0fVR3FHBVas2hcQX3Ti
YYlgjUbDAAs9AsW3yawU3uRNpruVId/IIzPNp0qfm+hBckQKGOe7D0PYZ6f6+V/2RjoL9dXVPrRT
FFWSYVmPtc+yiK1hfEbyvpSrNE9DAw1ZQiQ97OoQbS81Oyet5SO/37wmHDC/VgI9+OPGUKl/VuSj
H97dxjevHpvE/hOk/cw99lyQ9/q+twyHR+E73LvZ774pLJoLHRvJMvEGqb18QMbVSmk061FahlUa
l2CuI3DFNF2xRSKDxvq/HBFfawG7p9z93d15HpNrAl8M9v7bWROHzbbPdC/ug4DA/eiiUQyQSPhl
0LD2SJMvT9uJPMIwuXyEKe3ZqRRL3B3d24SU44dI01cYHUxWRFDprohn0netTkxpDU0A/dGBerwO
2pnumwvdfssCAwU7lmKpTbkU/mM+a4262q8babmZBHqiX/yySGDy99uwS/MBeKoxdcPtotAesU7z
4ytJcBAtXl/yUzhIZ54iTx0QkJXotu2oMsdHEwb2h/UZYTNALj1d21rWXWZQt+yBUFVDdwt/W0Cq
q1ZGjLeD2/ITdZdXIJ/nvope1eohuFvfQgEBUmkG3UDYeMR+S2pSgQQ9q9Q4GBF8YdVy5WuBXlXe
kN6nJneI+J3Nh72Dghud57TC+zcn8CR0iiiqMUQl1AxdbBKQiR2qpYWqruGymbIyw2W2kjP7Sxzj
b6MtZ/3OkLcEk8p2rUd5W6/0gHTV0lcoyclojkAbpzwHRZ1Ic/4+W+HWZOJOnJ8YBtsCElxu7OBE
WD1u5fRkfFX1hB5MkAjcOKCh5+ohtksduidAuycEgihjuQVo/YmcJLtklGkz9htSuH4KTO3VRqbC
1mNaXB1TvGp/phdN4/fGZRA0zVg/OFe2gc651niUPBaaKza/DRKPypVfevdI2UEXqlAw0bLpE3pk
m2LGlDr+yFxjHBlXA4tkKjn9Vk1OTlr1dHeW7L3hxaGYNue16D975I9WUFUqfYR07uQlCEtNC4R9
vNHPIxhcM5krfUXP4lx5B2rsOd4NsTkM39AFkNj+2w+cwRb7iku9I4BSrJsAqOk8eGAR+CdO6sR/
a5pjVbXYtTORDBRH2v+bhcwNVU5UC9EcRVFCWPJ0v/D3tI4VtpI8qUQaGnkq4Sj2IGXfckPaaor/
Sr25eQ+TZAZRKlUoM8a28jjQFAOV1b/ielZYmyCI/2iQD8J/lXFgQm1QpOCpALFDm8VMbQyCz2CD
uoJEDLKb3qiDE4W1WOgNcBEoUyeMnM0u2ZHdP8VNI+e/FmNk78Qi36su5ZbvZltYENqhtLfQWYW8
QS55y+6NkpbTK+DpHtRUNBNPf5Vy+RnAdRc8WDHBF+9GCnJF7MjcE3EoYyM8yAZ94wAMXIJx07oG
D0oaTqg2WVZa6EUlqvO02MMD9luOY7Bkh9zmDIFYuxPRS/ocF/e26RxJPwu+kZtcehww6sfOIGNf
zU3hixWS55qUcdNNtT+qX/W52TXBkvspU9RIWoXgBZi2zfUnU7zJurQiSXvO0VIl/3Lr1kUuNnz9
frK1JDsW4SR7HQh9CRCFlMVg18+7GsbgjLRXO48m6Euji+qV1K6RzoKqeSdk/9MBaTw2NhP8N36i
SJF8HJ2SBUJClCxwq+jSkaORXypKXz/qizYtPap/bBbAa8mU69HTZ9YKkn9BqsXcixDeiKLBUu0w
Eh/57nejJvVeD3hmh4dvv+Rrr65HThFtNZtybr4DHjjp9dvLQ41N+qd7Gs21Tk7rXsl4vBUxW5bQ
mGBqrRElvWoREU8VDJht4B/kFY0YgP7RWqzKjcubjl/Lgz5xDPcAgA6TTHxdxyNqSmIt6yctkZSD
7kgZsHc1/a2rUiaDMSOVTjmZaF+6RjjP8tFlmj4fQrkDQ2BAtvuRmMe7y7ZSwe7qAb/Fs1sl7/Eh
+mWVQtVwmZgCLG45vVlBG9ltfQh2xWbaHYlwAnQJMpCmTKQLfdSLgLDGBfAVgA5Ez6B2+7Y71BKW
RLXJCwZPOGVMs+xFfyhgk5NuHMOauCd0vwHxdBwmB6clP5CeAFFVPFxjCHAm5FQiDZePECRjZVJ9
DdwrG34WJbC5bBXlfDZDkU6Aq1D/oG5jRjOUvdIaRW4/IlUo9CTe3E9/+0AN2EaS5poR95WuJIag
Mnzt6EjYStY2qGlq2ay96JY831UCE2+UCIP/yeVblTKLk31grlfWE5qq/mVwcXaMNfOVkTpF0nYk
DK6WD7t6fNIV3W9Kf4+hFKC+cAz9UNSjxqmsv7PERZHEWSw3HvSeehW0kE8IismWlTPXVFJ4HH7v
Q0+l0BLcC3h0JZ2VVGA9EEikOdCmBkD8InDEJs0LP8BHoAKoJgjVj280udghl3VP7yV+7ZZvBfnP
jM7TFWt09eyWYeDH2al/QEFuFLlvb+W3phs11AaelSf35T/yVKe9rbVBen8JftKe/XG5SxjCApF3
TrYZIsxpRU/1ecMgmk8yz1sL0QCJm8u/Q8LNn5ax8kDnVV57Iw7kZTR+ed0YzeosG0TiWOw3uNuV
yVl/GBVh4GiQwdrtyw2wQC7o/n0OZEuVFlB8ucb/XKqnHliSi18ZXKMTF7fxceZAMyglkA09AHMh
LumTvdJLfna5MNFSgBFaIL83otDmXn8RsXHuYyn7u4j7o+pv47CbjHjNhBkFaCm/QGiTVAF6m0cs
EdDGHK2zCr4UWzPeZx60ba/bXiZKMz68li23nKdJlO+BnpvCsXdAelxZ+PBwWs5gbbgX2yOYFdC6
wvR8Dz/wbd4oHCl50ABdJkNP+Smi/FxPwhJX+Fwwlg5/QJ5CpaOP4C7cxQEuA/0EteheOYXitTOv
xfQlEelmnLbPhGvKaXXdYZvaQw6XtZk7bmJ3QF8wdcTuq1tKHCawIwRBZGOzcR3ck4ksUYjDOImb
rMRa18zaHPoGyzhuMBqaVWlI1urd6FgQi23haQZO/Gy6YWO0kmREiNkahIPT/M7fC8LE3ugRb/6s
dyu9rRATnFhZckEN6/nOLyWsNGBi9NGlrE/hRVles++o3QoWtepjlu1DpO8KDbcexumBjuw6e0xr
JyVf48LfSXIqc6/LMHYLT6SggVQimDKwx37bvmbgcC0tRG1OvNMlvchTzvUTJH9f7nfbQxuhQuQt
fxsk/FcO9HL7oDrOjeGcIrsK0yIraNL1yjOL1PClDXX+5RzagYSm10RUucTb5DCxn1Q0JHvKnxLm
FIXLOHwM/uN/YdJrH0SlvY/aPUBT+lXdy5yKng3GlLRaEftemOU2dUOyhJxFy6+GWySSBru0yynq
212iYEjorQuj7WMtyZlYG8NdilbcBJVW1teCq8H9OKbtX3mMdxNSj1YAQ/YR+vCc6N4Q9gaBmFCb
6zTKLa7AUqrKf3bUQWJOY1UtSN98rRMB430wIOLWveE6TzT5KkfzG5g2JzBLdRtssirSRvAxZtiT
JDZV2+fisTfJULR3O19ZL7LH+0sHI54/903k291Cozsss5cfq98FI42f1KOEzXjh1i4DjoT67ZFE
GnE2i/B6tGRHr0tZ4gj9DGry0ojV7x0O9xB0rmNEEd8DH3vkEjGRsoSsUNsaIY6VGlkR6vrJoIK3
QF44iDnIE9e+vSpdMpzuiphVVy/x5QxYm/Y0+9HYQcwUysaF4BUxx7b+fbuW+DH5Y7YKj1TImk5s
qLqsNMP7D1WCfwwmkbsb3iOGu6X+tvZGb3KrvtwRJkkxoNZbM4emKvfmZ0rY6s27urXJE2LPn5br
N2bK5m8Qs2XesQ9KAeW8ZnlgSFhuQtjoLzog2DnJcT3QJ4BoFRjkAOBEbAQZ6jUNf6QWOjmWFxrq
PJEX/lGHDbylClkw2Fw+QgRYcR0wdT5Pzh8OHNV5A82Ch9NPzEKHwOI/0/jNwFv1LZ4LA9PDrtd2
TPpAm2j5VTS8O4rtsNzKjdY4Xdoyi35OuJlJouh/TAeXDbZfY/wjXqETnC1jS5TArFVpZYnnFKJ2
rW+ZXulKT0OHfcjZ1GVIMPOjdgRhCZlWQxee3MovW0IMyXGtisGvv2gQwczGkPXBIcIwQ8yCcdQ7
JDJ+jMNQyMNzStEtJ4K2mRYLDg/1Q/n/mDU8XJNkp3jJzRFIugrJQHK3PEwTzWk5aanVDoD51ymf
cDMpS8YGhxzoQ1g8SDEdAgQxWCUO9PucA3QRfMdFuNGTAOOVv7vyOXzbUuEWHMIg152MT5T3bXYF
95aDFpGka3LySL4+mxuKnbnfipE5b2rovEAN99Aa9rzxbm2tpwN9JJZd26MmtqWFUHyVbkFki2RJ
EBsfkNZfmaIpt+LBDyghDv7kjt4uvcoR5MGwWIt/jhCXG5nDYCsYa5cn16FHJPhAGi7ZZbNW7H0/
IEhEaxpTWadNzlEL20YPkQT61B0zH29Uz5szCTh+bhgvowRjU7qwuLNqH+uO5yVZFCs8dWGxYIzg
wcUT7p7pxBBbPrmukSSwKYEPZ/AyqvidZ1iTxVruptm3mHAzhwq27/IsA4eTxfzhD9JpDD563df4
WoMzz3ckjpvn22KorwCI1RcOvHWAELT08GWZv2oncOV95q8875CqN0QNiUiun4u+j2K1QI4xpkwN
7iXUCRgFvug5/QzmyKfr1JnfpxprQwJ5uBsB+Zw5UnlcD4HrJUanObjm18V0CmunOaAdIIyl0n9C
OGQOpvP/Wzz5pw4qqP3SxVSZVhbjmTQ0VHfuuDi39pRke2O8YG2PKUAObEJZC1aYUScpTlhzXBbL
j56qLNtfsvH8eYiDbGK0+TPCRnXIDwgxfJQcRYUjyDYFVYFWbnOsPMWchg2PEoJzULGInig06785
ihSH33R8zFmOgnraHD4cnjdy73QCxn8jHB+ESrYhUEsU0oqUP4u7uBBlp0jlDbgjFDyopPB+uIsA
8EN5Z2u8hFquZu2vzMpjoT3Jisq1FZtZUFZ7MXQN1eeH+AFfKd00aTD/MLQOPFlRQRr50E5U4lsb
r3IujvYbskHFf3Qwpr+krKtlzAbsf3tLQKN//EYmp9wWEyqUESZtcR2G76sELCNoT5cNa8BPyHBw
GzbwaVSp8dQrSN5hiIX4o6fv3iChaHD7cQdWUnwyZJDWsMqnpmnb12OuBwxqDXIA2iodXpD2MFU7
FhtNm3ItiF4xHeKJGoRDEEJbJUcU0hhGD3w83jsxpnrhkyPohYmYXw0ECka42oMckpULym4QfaLi
dVVpHo8p6ikEzAk09CikEfHUNoPhx+f2Lg3YNv0HtomD8Uuc26pgqJQ3V7wkUr3KtPUSQsTUrf36
18u/S2oP0vAkx4lTLixaBjqP8mR7zlaGpvQvj1ufcKJD4oXGyT94y8Z+lcimI4j1L9fZu09PQ26b
Ikvq0CoaIeLnZ9nLhEN2eCkkyX9W8l/YrVBYouRdjZEbQyqo2ILej2MJTyXD1J/pX9Fp5o6w0La7
93xHZ7ln5hSNNtb3uZzRQjAhGL8Sxz48XIpj727wrb2qSzEKx4frjqDOvuIi7UGNfcDKAAh+wnLl
S7UZSVZNvkBWqamLgpy2ZxIcxb2Q+KRcVqZ59tLTPuyJMOs1Wy/HXEL7BjoTb+QlgkhgvgK/c5PS
tRVoZsV87zsw6Lp0K1nvKyCKQE22NvwFQ2jOnT1etHiZB0KUc9fDxfJllrUd1l1JlNQ2vV5DFvN3
WRebGB9djlPVkrZmOlTKHFyCatJ2jxOCw56/l0NNDtzQhXRlf9XV5x+Hq3PrgTQ04zHZPifUwcEQ
4HUM7wx9iegJScml6k//f7kaKToaZUU47ON7FwUbzs8TCEfTwRDNe6/eKpYC8t6CULMA457HQcKg
aQy8S3Kn1mhZ52ND1PA4XuolSLJEo+b6uSwHcbqCtjMRxWwdMSczDW/kf9J61Xq/EsOf8KLklYKS
cnK30nkFOlmZ6QJBaUtAfhG9bzVQZzpGI1mzLhwiLrqhdehr22WfWbch96CvHth35ehEYx3DIUek
K6YaF6URuOuU2Q0YeF52VaP94cV5q5yV+Mcvf6RwSO5K6pfLuWa8hBD0BmChnTDn+LrdEcjTAaF9
LudjnAxqAVxymXP7TkHWiqOebL+/H0iJeHxCOlwO4c95LaFHQZhzwV40bNzd9zNc2D8+l9hBJGZF
KheOtrO1+z6Za+qw+6vEXEt+oD8l2MdGUnST71olUKBOwx9BJoZcwbVSgxdk06LLgZe1ZkZUzQJO
og/uFut6aXOurgdZ0gEQ3WhzAMf11Kxa2yi3MV30/i4Uu8Sr902djt+PuHo3hw/Xn45Ksep/ceaW
tqAQHjuggW6ViyLN0Gu2Vy8hwEYlwYoJ+9r+L39OiX5cEt94hwQkeJtukwczgO95US0vTAkiUGE4
8EMtwCL7ZibXsw+Wajh9nULnesRLAQWbyLTBoInFsn7l/1CVjic6rBMD2cIL4YFQGVEz72SHrEEE
5sD1TmZmvo0nDzc76GaWACtRtgzx8qYVf6IO66/O61Afwtre58ST7/HRvnNQ9GJnh41ZOBnMlijh
iCVncH1OeAdd461NDlKD/DBwrfBsYZtMT5gPGB5ZT59ZqmOxabrNv2wHD3/fgWrzhYbQ1fe8B1eE
v5cwyxCOEqLtKXXabenT5Cbkk6GiawAgsqWQ3VsgyPLPu1HpFIgQhsOganQ3ZfYUowBRp8Wq6jZp
mShlcki0xk+Q22TuCdfgXklwDfZO/fqn85M3ZddXR/bkb9vcivK75upOYhnfBKJNCNGkPq8vn1bn
FtoDQ8kPS749pkmNztKSg+lw3QzPZrmNovQvXfLwtreHV8QLJsDhbhvSwtUV/KMDlyg+EiELtxsl
RWxQ8TRhNUdsj1Hc/BhwQlCvfKEbAWFQPsdbjGTa/UE4JCGFT1G16rRCt/jOyniSPG7Nfzxm6LdW
dSoGKs+fNQOhIY8IYWXO3s2Xui+XjnbU/1xPhKBXMqdQP61l8dJcpbOnxiH3f68PijbwO2vUzTem
IOeAoBVrumaaBWqb4QDcshNHlacpuz0H2B2UeKqnuXdrOLKdJ9/4gZdLNrLrW0ChlOEmx5cNUFZ4
5PxhWlwOM0MHkBVZRDXgaZhA5wvu1UvRPXo95zyO/6ll7VxLd3xN4aKQ9sJ1v4VcC7VlLsymQRph
b2Z+fPZ8pEC+y+wP6ETd/Uel8uJZpC4Jwq/7rCD5DSCsh4OwFNAXo57YcodBVtsGOlTX6/zMCMHl
nP0czasiS+LrvuBv4ydUUonPUdfB4j0sNMrCt+wpNY7R7keYJYcrHf8u07FaBGi/Bg8cUXmPxF+V
YI12c1x1u3Igv4l1jMk3Yade9Z/xlHfjTJcOvwJh/P7q00ntuDxtNUzX5T22vA9F711/X9UF3zRR
rf9cx2CvOWc8ScHETObsK2RFhIj+MNxQ11qCd/PUCqgKtW2ok/2Y20aE5Q9JG1urK8hM1sQIQqSS
BJieYj5e0bxwFcEbIthsMAD2pjcwhCg0yYz1N3vzZ7z2eZ1PzsVMuQVgB1hz/xp0C0MFXdx0Nq2G
6BNZSAS4biLAd7sESOWVPejCq3P+7ClJ0hwUYT45dYlCimCPSOLFFovvGtGE0bUK74EV68Iiam5j
O+c0qwiPvxpvwxy+YfuSZxkhgAW5RDgS7KHQZz5chI97wvO5Ox/sP6gTVqc1IbQCul2r8hAUeTpY
/vqpIv8vrjD79y+hwKksMe5E8oM3laNmHjr0c8PlbEOzVmmzzoealEIlN+FfvMjuXO34wzKnEHCg
NPXXyPCp2Fv5ceoUankJYtcDytgBMqkJDuvWYjKlZymwPV+NNM+NSatlBIRGTRzZm1p3PUprKqrc
JtXDVeqjBdYq/PX7Qv5KB2ufpUOXtpZDvGRsgEnO8BBg6ma8rXUi8GPgBs3qKWEzJj7Er67Xdhiu
SCthPWVg16lNE4ORtZAd37CzvPErDsi35Ik9dL9bypRj+N8iT4IkPmZ4XHIoNPqeXpUXTP7tkFg4
/RnGkbBdH95B+PGFiEm3j72AcmDFAIL7/yW4eNH2hVwqPOEX20scbtkGcv7iI4cBhSfI+gBcRi5N
E9NODIU4mJt4hltFlQFzokfBPg0oPL5GqwLGkMqoNeANvElXY2c0V4OHwROLCKz81pc1OSaDA/iI
PStSvoMklRo1jGEGWen7iEpiCQklhENgH0aFaJ1FdrIcOyGe6rwkymlqvFe6A9jpN2OUOgdKXSxr
jSpn6iZrBDaqQc4TPeMMma/1amSzacEEbbxoUfI4H+DtZRe56KiPdrwLtYhyFBovOroNUJ4nBNa5
CwqGtI2z21keYWEYz7PuMM79ZXfYOn/OFkvOhHczF1HbsOso4WxFNxx+J6in1LaDak/ISl/oM2ck
HasxeeXZ369MrTHT7seEB6zftAkgJmRpkYsAWEdy+USXN8gx1HdpCURjaXqc946amigwLpE4Sslh
vFcMFPn57VJXi8xDQM4R62YlFJfyvW7STCSspI8CCd86G1k592JDm/HqohoKj0k7GJjWOFe2BxzZ
OgysWTdAHqIweCOHIbrA+498xqppyOh5pa6deuOx8ZPLh+RRypcZaFxmkRy4fPNOC18eL4lyPKlU
ilEnVJSWHLSwE8ufzGIJ0ZQDBXurL31b19+HQ3MeVR5jJIL3FJadcDQX+6ZXGbltR+qN7BzkGQlI
MUQ8q5yjZl9am3OWzRe036YuOvpbMjgh6X5IkUWE96zUMvxls0DylWsoEcHzXuQvQzRtmaXLo2Lc
dsIqWy0S2y03BMIm3+/bLCbtznhaEfQ0F/opCrzgakVudbV1YNbAX5gXnTd8QHJjLRNlCkk1DAjR
t2QN5kMXeC294+S0oxluL11KbaLY7D6JPa6viOqueL1Mb5pYSoJjNO1G9YAQ0nWGVGl7wLes+2If
CjEbXtPdK+Nx1/K6+YNxEmoQ8/nwS6PKZwlvbzsd61ZOH17WNGi+7AAwQNwlIc+P8I0cq/VtEgek
XE+/hRIUZPqE2sXC74sSCfACO6L2KWPuJzemg44mHnw9bwF3NkofTQcXkAAnxKxsSueSPwtfZ96g
GLIFkoEoRYCgbXbhEqXWrVRUfHE6CVNW+Lh7uX9KMPMP+4eaeOSA8L9v4GqjnfXqTf5DPsJstzBH
wqOG90oURc22s9PBp0iRvRCdJLJdUOxEiUgQbFKyfor6Mz7cX1TAn80+0vIIHNuyB7XXN254gCoa
lSX1R8aeY44bsZwXBEQ+9s9SNd48zUoIjlaQujoSMHroDIMxYZ05M/S3tuFymBh4Hoi7lLpI/CT+
vMp5geiLeqWrZw8ptO6louME6kGEWf4yIzQvzIYPwh3F3YukVnFja5HfeQFbm2dlHAC0EO9eL+uG
YFr+KlWlpVY0+kOEY582mGgtGPy7xkT7/MpsXJ9UR6rhZQ4IeWRaor5IkU2rvpwlBpPisIgkNcPZ
QCw3YhJqK/KrIfKUmLkGlZFQVCpHArhfaCUZtGOYLpFlXvRhrtnQYZG/UIbBvHvaPekK7VA8t3Aj
AUOXPzl2CwrUdi+1rLdHZA8jf9Gm7ADRaI69+6YOS+YvzpWZ96TOQ9qsFJNI9H/QW73uR65dgQ1R
IRIXSLVj5TwP5M/cClExyt7WJaiq5WWKnfD8HpmfCdAMI97FFu17eDeLl6jFPwAx+W5iBZNPUt8d
qEJczuJyJCWle4WjJdQuV6h+iijwA36uIyi8YksOHx7KdD0ywDP25jCrLUpgKrdHG0zBciFxHoWi
3t/wCQaPHKMVyZOdZUejpzyS7/Wvt+IjOdAR1jy52ciWzWLgcj/Du2QWQk9dWFAUQkWYnyEMZQcS
hy9Yk9yYGJ8yD7VuFoLcI3ltrxarFbxtWEhzxQAP/p0B9/s7nb6Xc/LPFuAX77yr+I4VnRMSJtcb
Bx3jiSOMzRnig2Mv4M5ZPU5XsrhzE940hvJDJQgO50u+M4Z1xr8CAFjndx2YT3bVlIiBtXS/aCbp
aTyC+uVbLIkKAJdrG0YhepSeq5klXCHtsc4MPp9/zvPyHuauGQzeOmZ3s697txND6YeYdPV/EeVv
64jsliOq97Dnt76utNyqCTbyJRTzDL4HDU+SZwBkE34T9R93UqEKRIDi9Id7bdjNmP2CASfIZtmg
ghR3QROUs5zrUXgGIZrSNG1RGR5wPf86WGfCWusdP32PdBfwZvCR/dRGXmLUpwsI0lwZgA0OJZe6
6NR+R9hQMjO3NEJA4b7yzT5RDG7ttJljiqk6wCGkpv/WpIIoZ/RfFwfIj5xa5j343VuwH9dbDsTv
C/SHake6VrWxe4GMPLCRVFmrpdc8MpVK1XWggDHMp8To3t0Clti3yKwJBJXytWVYxP9T597hTdCX
h5lf9lIVb1pRs6pLbYl1XHVpj7ptMF09ShZxnSEvNyVQp6J7EX1nbKKfO58+uUI+IuN7py1yrakY
1rCysqsX2nNQW5/jhl5+GXQ38ruOnjRLF55WtC6i4d6lRUMWG8Vns4meuyZq24yQ+hPPL5zoplay
GtEw7KE3krygt1ZStkPJHKOvm5tR8ljJwmyx/IYhV7/3/eS8V0pBMF/y6VWm5aMjTY2gaHTbXG5A
JF0GKfaeYdDtW2Gq38sgNVyE5cnE8hjpYLWjkyon+8R52+OEikPjaggzFER92oWcgNKDXrvuGIez
xzb79UjudTGxtGqM9dvBgk22FISmGlRTX27cNcVfbZrDDqOI2GYySTjAa3exSm3WAtkiaxh/+y5u
iBaFfmBo0q462uUlEMfFdnUS2cGiDlygBoF/KqeR8rpF67jMEYEi8wsUt+zoc3F6ecr0eESJkrHt
FYDRvlTua847yNpsMNaVZP4N/D6FKBfTuR6y10aLt2Mr8tvkBazS6+l4dHRiEd+hUuo81Pk9G9YY
/OwROXI54Kd5PmAZ+NkCVY9Cjp2mOOuCXG7UqZWvs1SA8wqzfRGf5QqJdje+cnLE1myLCZhP2ajw
NgGOAJ/12x+Bs4YW0UP2lup5rcBKRqEMg46r5TeMO4/WLQV6J2sl5g9GXpU68Rb4spOdNMOjBhBO
hedwlvvHjq3RojXtIAd4afqDPNBiOTeCjoHQWxC9mirJf3VcStbf/xL4W03x+mhPfzrqEbdTziur
ix3J0g5ef0HPhUNuIG3bo+kjrByFKj8nMWSZfdrtWtZhpMeHiu+WTENz+dtCRYR5uverFnUzWMRE
LLIlXG8jw1I/Ep8UgNm3g6whu0W1s0qlk8CwV41dWrVsTcK1h9x5xC5GxFitFGu+wWzJm/fb6ZFB
AfzEswCAnv70PHGQbbdKvTqev2fOIFsrp/1Hb9FsPt+PFvDtDE0SQTREvcWdQGu0c1Sy8cBNSqzx
LmfUSfEYC+pWzR5etY/P36oE9QIOTk1u2X4jrRaDCWeliMQSbLk2gFRzchwXanWHUlsxbH3C9Zke
MqX4RCmstF6AV9V3Gh02+i/OxGmI5RoYD2mpltEN+szpSQv2WrhiKgIZspRMtUzGrJUpahueGQjo
ROlYZib7YWfsYzOSh6yvOwfUPbe22Th99qZeNu1LW96qUTOunt02T/RBHsB6zBSqsMGMvc12zopu
Lrf6NwTfHG0WdGrOBd/BSK7ZIce7PN6KfiOafRXxpoJyUYDW/v08VN4iCxVABfzx3FFHfpdnpq/1
WLVOrfalAHh6t2dtVe3c3pTgG0mnnQmoaCq1AW8LSou81iTv15SN9hcWzjUYOPb0sZAAweGCacci
ryezV7ywbA3GfrMofn590S4sxSHOqSfjBZ1lQYt5GOrlLoXDwolCyUE0GqKhmPoQMXilsbXpz+jK
537BZdv4oUu9p6Y24T4vJilQq2e0VIz5rSyNwVM9j0bCfOPYbuPSkJW2cBy/8wSHsUgibelrShPZ
ItVEC6iWypCSmvXtBxgHKFg+KovB0BDH+18Yz3rILG2GnirXEO2zhNFAOUIYB6pu4OgN/lwaE/0a
yF7KBAaBoSuMETEuapMdxqJ4kBZUxd4j7Oz54R09aGkQDp7WvriE4bQ0uKmT/EElmFzzVdAsJcOe
6PCgvNRi6hsEJiySiCm8+w9EobagC7+G6NI68xjrTfXakyPmK2bzX7sfM6k55S25Ddwijq5gnRZH
6qrK5n+KJD0caeX+60WIc0f5UOOz48uHBHlMNSUGfuE6AqZYzlWftIJHtcVkh5G9oiKgN9JTMuAp
hII0Jq619fVUjTnN6mZGuk070PknxmZrRD19A+WO4G/yDoRnYBno4fweLyq/hpNcNYRBjAbIVIOd
sQTksmzbetHpv2PLwc2v1o5WWJ54dijJ/3IOt4Z7SiX8aKyWItK6MQ3YagfeSfb5Tk2V7fWCBJTV
iRhzG1CpVtWXM0OXxGC+L54XnBjIuDicynvfObZ5wjWQ/O5YqLztvsdw/AX9cL/rREq6kaUdvPu5
zBh4Uzvj8IFvjYpqT4tQFX63qRZ7+8Ep7XhWDNF9oKCvx2JIjvjYoNVAUEJW8Ge/GHwiQUznXPTI
D5kiXaI8EB9ujXyy8JwYcis6vpFmeVecd51OCnUUsUthEMAGrDwE3QJi4eegpCDjl+ykDuY6Gb4d
mG3c3m6oo3y94lIhtFNDZpJYOJPL7XgpYhvmyQSiiMT6uz75uwigjcono5x41/8uASj7xU5J4ure
kcp3w6EOnQMI6LcjMjPdvpTC+TWJtwAvHp2pBlxT2PznnvV2dtKeZdP1fs91e9ecRjyM1ZQh79R+
V3aqwIKfTBJOETcW9Nr1j//mbBgdMjZGmfIf+xFZeLu+G+9GbtpKP0Iy+m0LVHjxl3A4fTTZC0H+
iaHSGotTIUwXdwVom1RjSOuSyyIFwwEr35Sy2qolZMkcEZ9infr7ldEn/DMIHDjKIc5Dljq/A/UC
9RJHqJ8S7zgW4DHrbEURWbt8AzPpzWSfOnFVPdRh+P4ybpit1igTSL7lnnRE75K0VAK8aYeYz7L3
/PCmPv67G6Vdtx84S/Pojt1go2d6jSZcIRV1Y2Wi8uvFleYaDusyAvwfCVNePuJ3nNHYwt7veVrP
qKTtMa1NpTMmNRCQzI3HVY2j+Br49NW5r0x1YHmX89sqe924bOR7kN952spruPlsgRJ5wstpDJ2a
05UTgiov4Ygk6zWDKpUoYLGv4BbPVw8M6SJ6o+qgciI8TD5ib1rdrfIo1DxU8X8qEVW5NrpyAAPO
COGbxjk1Ht2DgVSgk8/2DpS5In6E2oAeI0r3qN/au3/TwPOlkvKXdjunDHqXBRgC65vpsKGlwev9
4RhQi6LvRn2BSL1Ss3Rchkl0WLBbRahYxWg0kvddNVNmaPS2VXqak917XaLOw469ZF+RGIP0W68L
N7usftWkVlR1RlRvcjAegvy2ryKrSLK7pJCsGT4DNkYsB3OkMcSp4Nzf8CjKSqqSlos1LbaySdyd
9kpXLv7/Wi7GuMQRu01RXVofMPw9A3XRtzUvM65iAKOJkn0/LF3+Zd48IJoKST1cseHMTwuFrbbM
nEm7HshG7mJ+tHkrTAQTbf5OpPZVPF6/th0kuDQQQuBbd4Br252Svafch1DXSzX+z97rS9DQ1NWM
t+S0Lgl3VB0hqxWYhDHCay3IUiya+tSxflpAdNxhdVkGLIpUy5UPwcaHabOkFrVobIBFIF0caVrc
zla79T3MzOEs+w3Eod926Y4KsPUX5CxwPxIO7SrT02Gzp/BJMOwIWIq2ypBaUKW6vLI3SxJJwnCK
DXyA9D78FH08ld7cAsL8foyqvjOCiTmYKdhd0BRZEOBHjrFKUnJdlccfcqOlJEfLTqxEuY4zFeMe
nuS7/1bFvbbMKmCM7w+1ftOw6/+XKlE4xkJg9ZJk03Z/v0bnk0PPXBJtk5ksytXt9m/vOCEmTAix
cRnsTqQK4a+U2XgUQjt3tVgdRs6VnnWjyBJGbHouYz0fL5ROgsnD8GSFhzYRchloU4D0+EZffVh5
DdoX4AeIRp7Hj36/PV/sGuireUuaghrwwiTy2ImZ6rTvifoFK3TfjV2CbNfhen3UZ+1z9XoSUUS3
RfIsjeah9MPpZlf+ytBgQHc3Xaz8Bf+JB2LHmU1aX35Mkdou0NGOFIS6Xxut8DNt2zji7Gb/kQkY
Vb60tCJR8raYEcpXiEIu1Ae0rp1F3yljaunzZV+v8erQewq4aa/j3ZhbIa8uipxt1DL1Tg4YYKCX
p8h+Pfby6vTh2JAU2eV/wq0/mnVDOZ1uuVcMCV42kkJPQ8NATT0jYleHFCHFV58SW3yHAl98MeiW
E+2qDiLFa59FfAmcRPHnxchOKz1PcTOh+2rP0UQfGFjmMKRL0dh/myWZO0R6vuCDMqa7lMzXsNl4
Bbra2Ef/hp0I6CNzQt4d5EBa+0jmAclEXbxpKNbTQIyB/SUet7A2u4dYBP3jUVrbutZ40wGZ8xVU
Vz0vhP5y1Xz5nQrKmDVxA5lRcGWIAVJZXUw2JpCw9SE3EghkwEa5Pqsy68gkreMPMD++uhoSuO7k
InDZpYOWOiYKYGeMkQx1VJz4ubAFP9358osv2/2w9urJqor5mS6veAQJcvdaW0Y8zXUSlXAcelN+
9gzMBwzizC5E1argOF3bJKYab02i1UuyMotNB2hpkKjuBdk1nvX6qwyyjGCL4FA4kxRoHDx7ySgl
y0VKASyKDXdTJpwp6rfTjhXQB7qezaU1PQ8rqbEmEzkZ+42mVElpVP99IDfWp1NCK8/N+iuVOwFt
GAEUeuvFzSCq8Spq/F2Nangy0rYt7DzTiT2kJT5/LuCSLEPCmK5kR6ZL9NYKCmmMT7KZ4Q3GGTC3
Swyspb+C4FTMVP7gykWww692NLQ8s81r+1Iu7305u8WQ3uXauyT8eHcavGnYw01gKeqWItUliYcU
NDRr3Pjln43X/H2FeHXOpjDXUAlM2aVpsSGhTsXM2b1rxXbhQdWL9hsi1QbTGHpKc+uyydxMZpb+
Y+9nmrINro/OstC3QEE1OlSoOoLEfdVwEt0uvckv0XWFcvqilHVjgUIJiM5v3jlPfbo8tUM0qat4
z8u2Vabrnp9l/1juBM7Bof61dz1ETi8SMUjmsTeFt04pbO/5jrllKFQwiDVOdjj2opkdn28HXN8n
qIvv7WHajj+ogSYxagQuRal9TU2ykPGzbZmnTKnEb1oU4nG9N5E9vJsPcMU/7MeEhvOkzA2Lj6M6
gJnyjkvWk0SOuUHvcoShcxMRqMXCBiiC14v+TpwPxA9H0JfUDY7ceqhGNgTc3A6gpsFN0SZQFpH8
iYuM/bzppux8WAI2nfQemYhM+igLDqzA+Z86+0VsPj+YPnmi0483J32GpqBg0q3h9vJq+F6+39AI
FmzUt7ph7QhYJWsSovMWE1wLYJ49wf9ETMlyl1PtdMAbramjaUTi5kzDaqkHBHRPWFBzIGR2OahP
cThgYpuKk5PRyb+9cU0tEnvMXoANMtKt1cM2w/eKZGy+GrL9yX+AfaxUOW7Gij1BkJOwKlCQCqEl
4YabhkHOJzXIArA+zIkFkBDbZI6rwoiUg62OrnRBFb/ysO8tWwDZr/mkQ0lDY2QRRHZYvFpO6SnJ
V1m/a+OM7TR95vAv8QIPIiXbIU9xUGozQuQvOkwO3Hr+78wuKX/1No7UI66acCIHn+WaSlQp2v6K
Snuo3JZ7PSwoWoEmpXO4DcndvdlYdWS5zWkW/sOqVaFegI6Xpsf2YWAVYk9V8DW7YmuOSCkNCnFm
MTPFbZGMLI31yaiwvnHn4F+4aS8G+KqwGLqwYxEJ/625Gr930kIN/b0aORAoEjtnf2bZjio9sS8/
ehrg9RbUgadMljQj+F8KiXQb8lXWl9eUOQLraCbmA9LMpLTOdUzWLDWcDc8Zyk68pxNl7+PxPjqo
ovDYRuo8bS5VTAuMUvInjNiIaAmXAGMNbrPuPXrllmq+HsZnp9lD3AtkPdLqxmKTZMhA+9Wuu7il
tGnD/ESzNy2PJ6h0l758Rt/2nQdF64dwiR0MleBJe8BlIx+/O3KwV75SXcGera9bUf9AnpemkFIx
uMcLAD30OI9Eg659ilgiHsG9hCbRXw1koZgqwd/ovJ7V4UKp6VZ3epeC6bftLWiy/Ie2Aw930e5Z
6iLJjV0eXCbX0PEuxeIvs3nG8AdfE6Fu8PSjll4c8168mWN6jzA5i6JXVNLYCVjM+kNqF2X9NV/F
siDaHFraGR7+Bk+wJm7pFKD+QhqDtDgFtp8/QlKUNXLFCGttvnsfm1l8DWqT5Wn9Dz7DHS+T2oZ5
oMFldNw/ez3909urJDjTgL2YgZ6N2PpRuomGRW9efXa9mY5SwBKMtOr/lSOEtEDxX6PnJ4zJWxOa
2pFk7kPimeQLQCU9lrIPpRw8wzktVh4Vwi6GjMymdHT/g1TsupxtJzRC2+aaAL+7yLSNUFJyKBb1
R0AQ52aHzh31wt5hhyPWfjznLNwF7OfvefxT95gqHCyfb3BL2N1gqbDueg+5K6qsfbAtFPb68tpc
Xr+5APUQ6JDyUa04TJzZOhH2KiT6iAeOnhRNwjT1ZJq2wWF50RLK2J+fnvA2IbRfGuxwC15aBOst
aUrEOInVtSydyI/TzRO/t3Hv1xAWuFLvmmFCmtyfSRaRZRoR3nEaFwaUIJTZPlk2kutuYMGvigjk
W7tsOuNVYQSaPE/C8rSuH/Gd3O/ZcdKSlOMETNyzHJvIZZEy/0RxuTyYK1ELd6eQtsyjT4etn+OM
4wG5FaB231/Sx78OLpEVQsw4RBuMIuyycqysXXGRliT/RCCGw43UP5PLZcpUOodYapE+8nsi4diJ
PZ1SXXnUHLamdHrvlntnDck+/GleOdTVZX/gYyVCe2MUWdEODFlPie6IfBqApTK549v0QjVizUoJ
+RKopqgKJMDZqQmIunRE27vJaPIATYGew3q5kXlCUEw2neoG1V/tnZ/Y7RXtbhyLBAUa8y1u+7Ee
fftaLMqho/02q2YS1mumuyMLpMTfCrLgQxqOfSzWJTLg8c8gwk6swY6FMDwWSpvIL+Sa1stOhDtq
Kql8NSGx1eE6k5IkOUrh8Qc9heqt7hp62izQYxIJW4Fo77+wZc2mYn3IXoxLeSf0gx4doNpVty5W
v3FbM8/kVSkFgI47oGJY1eChRlplZgFGaMR/aTIidsRxthq+9Dci2u2aEZxccQsKXzMWav7Cdi1L
2BlayGdrhBYiPs5eKuHAMxr/Knam3RZgqPROuS+3qtxpLaOumokWkn3BXXaa7ds23vswGOwJoWGe
tJ3PJgBYF8Ts42qjCuDNiXwtS86my3gTb5uaDwNDX3uwWSxUaPNSBPSQMK+aJmvZjiUTxzFrs/QN
zFkPRtcqdtDRPrc0HGEDHxUhHU859Qb76l4JHvXY5YJWpuq887LNQrdufWdYaZMMHttpQyqB9w+H
6owkXb9lVNyDa0yOsj6mEnfcdqHg5QC7PMgVnUDBZImF8Jf7HEYP8NTHwnqkzlnpUKwsNmTLGkmj
du7GQ5RqsfM9sv6PbTIj00zTedAbSDvs3fIWaModc06TXjkEi9eLHNqy0hYibTnrKyEzZORftGtX
hxlgH6BexpV0SIyDxiz8ywhdTriIkmAcw+A6MIazblUguqv/nqkaJdOW1wBlSKG4J4aWAHqhUupB
A6/bAzsKZznVR3e2iv0oyqf4ZdJ1AnLx4uNaZ1bO9YzYwtBsqt7PK8K6dXaOUPrAwV2eXgfFnRFe
ulXxANjEeUCHBpKH27gYW9+mnc0KUzWzIRWM4Fz156IHOqgQkbSvD3bVrSjmKvGyAsoRn57iO6JE
Aoa/zfSJhF9Hs/JuUYz3vSLn/AAAC0qNuHy1q5Py4gih7eBvTek+C+GhkeKsBrocWlbjJAGSLgjk
xkQKAVJYcSP8lYw1rNRhk05+uH5FcYyeX/yab7ZRFPK7EEbQ1xGIOOsPDkwNeqBxeSupT2bNhO02
NUFhkrUQWqIhdFFFGQLR34v7MJZBKpvPDmYH0Y7XM9Qtgqt2ijTrcpx+uAm23s1oSZxSMW5hCNJo
TiDeLMhPhWXh1zArf+PhJwS9nWz0L/DK4xsf1LVbKnxqTW6YyOX98q1dWOesmpSFJX98sBuoYsWS
Qan6VjYciKoxIoPe3t0rLJ2rN4Ud15hmpeEymhygFXfqu6W2dRVhjCQgnleF1WujZWTFOBIN1Q7L
KSGh+/8txUYz2oSDY113BFT2PzaeG3g5jyV/G9JRvWnUv3albR2Ufu+dCvGVTeliPIJ4cOpccc6R
1KmanqP31m7puPm+rl0iNLqQ6ruXwrG/Hq5Vn476hVC7c52frYEgUnL+ZKhe/AiyFnN9YHcwkaW+
Wbvrd6K4BZ4tlnKPEP6XGivbAjUdjDbgziwXtHJsrio2qN5NJIsewOYwpUNJwewdGtnH8hGPTIBr
ytJM6drf8y1SXprLUhwQ+jQbHy8lEDbZo+dPDb11Ge+1JR9m2W6xh2WB3eJ+0grE85cxRqLfCX4O
cPlH5P6QBy8zLt4O+rrw+Mxghv4EnpTiACQkbYVEKa3NXylDKfqYig9dFwepzXaL8kktQlWrPErC
wDMqE5Rxnubm83U+yRpBmHYCoue5wzExrUHR9NJsD5sw4wxKHhdVhRoZLLdJbID3MoZq4Ijz23n2
D0Xvp4DZ7zaP8FOKgfzx/ees4qhddzuPUlfH4GtAQWNCXxdHinY4rKesng5+KZ5ZX55kZNjlt4U/
ty0PkuvFEnccHcP94PN/f7XfklvD8tYeKRL1+A3xmflK3Dc8D022+xBgXmbGakK9Tj7H2v+uf07n
agF2ukMhUWlYaQ8M0SxEVyWMHn1NxDM/ckD5MA1E/MsMeB8xnhkhydJSoEI7xtHQoEzjMDM/NgEQ
WE4niXgn9JrepDUyYJ/V+rZ+kQTzp6KIPSR+ICO2LyNKRPgdZlaRHxDE953RfXHFrHajVlChpV7E
RtlAvpbZfg+7VhSZp78lN5ujNts2CCGBg+R6GPy4N359ePVDouGzqKPqTdFOtP77NPrSWsB6OsnI
dW6zODN60VAJXqfM+DNB6zd7cIlg7M7fU7mrsfnhZlpY5mQK0vF1V6dCJnYO1BjCrzVMTB/pp1m1
uEkiMyZssKGyEo2u6B8M28S30fUQGPjfUhdBmp/A2BHQGLeYCOxFpQolppgapfBiKtr9xUP6BTuC
95WpaIChSG0sFVvrRghrLAPRh6T11kJekGysyUkOf735/lcnx8Nh3sU/XBpoNMnaWAwUyOjjePvT
ppWn+n/l+pxa7+nSZiCymb8XzD8UUruMqxYjOQuOYQ9qRzhNDHdyGlMPinfMBqhRyRFRYGmxrzLE
znXhDT0WgdQEgwJY9aLW8x7ESN4zAG4BUjFXTtnmVcefFONmyEfnTl7RJXI9EA4DIBI5PG+EcH+t
iPRSqvy6stcceYmNV1O1/GGaXeuxylB9YUshHLh/4QQaF2IkydMsIazc7+RCUUTmdIH6/Mix3Sfh
TjAf2Im/V05NLU3w/7+S3It+YeXBP1AC0mbaVed83qpmsQRd2RQpyMQ7MNYWt1NHozHMLn0sRj4B
8WWPtLVeRtGnwYtwUueP/BsQWpMCIiudKvsLnek8rwBxmql2dL7hOzhEFRco/YbUwIoLPw+/hkbu
Lrmkkp03PP2H6xO/e2GF1w2oWdgIhL3ONCNKnqaA0HCjRiQ+hxPEcXLu4YeGKfYb85UixRLkU/ga
HSNEjUhQAb4WMcPfaJRrCn/5litB4dwf5FSJg7FvsWTnptiiwALd263pRIw0332Fn9Ce8llgkQqc
Pms2l8ivgGTXRyP5hVwEQ7Zj78taQgUF1bg9NQrrUAOasZIaSgI1VOY+NUhrAoDaWHrAWNENN56S
JlW77PnovZ6ymDYEpzmiSpbX+96lZTN/MxDCv4vVs3jPl+tHGeMZlqtkt2tCidSFm/KtN1xG7Xyg
PqrIJ8wYIgsRZemCrkL3oougNX8VvVaag6UCNR4T1sKicumzdnikiKOSY2ReQMQC7rKubRDAxvTA
9neVwiLxgiEPLhf2HrfxXz0z/Gla/A6q61a8m8HJAbSuXpJEjH+ziBYkFIPIszb8TsWMPgHpgNHA
ajYbgd19tb44lflgPkKaTXR3ym+HpM4kds8xozgQF3YQ2X68/mqkK/cC1FZUm2kTA/0XNFLfdSaz
ON0PulrBEu1d+y4xDgpC8RgjKMh2zOXD859m2YNY92avykd+FOxw+asKazgQ3j8zs3EEEd76G8ud
fTmcFppX9nYXXX+wiEpNZvysdjIgBapMIMPNHH1ssYNSiSz05z+BCDevLod46IMxWsWg+Bx5CJn+
5r4+fIeDV16QaZb2wXjXkYnzA8L8dprfc4E0XqdSWRF2obUvA7Fa627J9BP8qY2lXeK5w8GArW7O
Es+JQRVA/icflMikn2A5n4sAUn2OblElOAKVooA7Nf7yJCZ7DKi8JtjHfQsMJdUKML0f4iGKnivd
KPi5VJS/C0882v5pgzGwsFIUoRE0M/DEhoQcYGHo9q3Zk/4GGMeJUcGn+GXpPI1qDOg9/RtLodMV
dEj/XlK+mgW7dDWfpKVJS4/41I/B+OMmRVSd8RCQoEy1NV50wh/Ymn8cP5vXuPd0NmaXSKsAq8aX
6tRLZGC+ynTm/rN9fn8o7KvuiUhHiZk63EOJxaT7XyhlmyLTdpAZTGhHazmaWlHyNpTng+SDWqYy
zT7554kbu2l703pPNQBBdimhBWM3GkvKN5bnEDJGzaQpEAs0LY5SElkvBlVWNBSkIx/GcpVLoP+x
kbZDyY5+YtYjUyP27STqatXzEyiMYAIYT+2BXVOhnJeHXw5Vzz0+mz2/pDx6VbLJkAs6p1VhFySg
Z9hypPRb+NZRuDFMAwT+PT7NDjshh+U5WTN0OTKCfUdwrpmPJFXLIqIWean6q7MlSO1/KR+Tu61R
CioAskKxEdi3lUN9lZyiAPADUhPMuU7+h0UoS5z8VkA2lg5lOjU0wipYsTDzaWpmbqeKjxgFScFG
qq7LZAayWx57Ctcvzsoi8Bl/oXZ8JSgnZy+1WNRKUjWBcOALWQuPTYXyqwIKko7aeH5HGyPjaCbf
mi7S9KfPLTWu4GpkOlVGvx8aK2BTMggJZssbs+jyrp0wCN7MsLradkOcQX8M3yZtJyxTUzxqV1im
NqJZ55frULfcu9A6VI/CcuteCowb1nppgil4DamH9dc71XEbI2q+m7MsIa05phn+PR6fDpZztVes
Ap46xDXAfGmwLFIkdjaONnLpJHqVGzq45+cpjKJWz13agV72gWy46vcJYerC7tGJJJCKwJCY6E9n
FpEUASM7YIz06ZFuwsYXamodc5Ptr2qXRfG5Mw9HJ4rtXoWl6vvmqnAxaUnrZuvLoEeCvspmQBbE
DpPPgxnMvjd403FpCT3gMIT+qp9+DDJROtlybPVi6UrrdPmHCsYjkj+MxjeCvZ85GRIFlK3N2Mzd
0/5nGhxn38XADsdTM39uZuBdFdSPhuyAzVKwf5ZUftYYMaYrk5kJnDxCBP0+LszQck0i9jqTYzmp
ZMFrwDyb4etY9gp4QKOQXqDTI/wx0FjceBokrVdOwV1C6lL5DmlwnPx+YobqVJz8HNW3pH0sGjez
cPQ5zsQEOjLIKMtz59685pdN/Tc8WfNvEV+byFaZjAW6Gwq9HQsyUkp448+0WrU8aM5s9carfhcv
i0f5K9DeUHq7rELlXlVjYrw54VQ0X0dQH5ECTNgHEqjp4b46gXjT3f1CSRmF6AtGXX+W8xxIbaa5
7D7b6pX4P0YcJCXXjh7PlYh+XDF04WP72G/8g3w9DX6FA1jwoBpa+wJyUHZ+Ty3jYiJnUgchGocr
Ec2Rd/BJANLTXAdPqKC0R/HDs/cLA+Oowbb7iBiw534kb/AkNZ2hAHzVoJ0j5xYRSilkSBfvOJWP
WHG56XlMWss6KniUY4E00OvwrcsHgihu+Q601jW/PqjuiFTyn7Ve+avdZgNRdaMYZQhKlG0YSXlu
nTy28m/aJQgggIk5xhNuhLDCmcPkEEAaF2BtFlX2GF5CqP/uj6bXx33eFBm4hw1OVwiZP6ZzBzrZ
D/aVbpZt3DnReV+ofOo2jTaUrS9MPv1650TgG8f4miPV9qLNi5BtE/mDMT4+vafG0y62cxsQ1ASJ
9q3PLhsyaFoCqpEsHYfFy/OS6oJwE4QKWIV1EOFe740SpUgmQrM7mrny1VsIQw7HdjCh34113E9u
pTnB2eRVZIxrJRh8RCcoXZ6tYYZtlDu5BaYuZVExf/l+EfW9FGeYrvVXjTx+xXZveeO0Cq6MeDO5
/yn/sCLL3dUiA4InXNSKdSqr9b/vknOy/9RZWHIvIHYlpljRK6LBeNk0GHloFfzTgvUSj55gjfLG
iiqs/r6AhLM0L4Sle7HZu17wYzRCI9IbUhcHLnWQn+CxaMxpvAQ2dVRIBKDo3aKzpLACaOU/6ICX
FgcEUe6LOBaQ2QZ1rnf8zN/6nvqCUuz60JYZB3h7LQSF7mIZX/OrBy3qn5MDMTQhivSfyN8eoqCk
LVf21Lr1giVKzjl7Qhs5vVsoOJUhLz5gp5YxGki7d0YisjizEaSgDFoti5aQ8rHat2F71fvDoTM1
7P9oBxlOf8JAvYB9+2kSLYvse8kexwW+HPDkkv6BZlJxPJ4OUTs6e0x7zcEoJ9XnYEXVqClDmz+m
Kx5wp/DWR1RRggCUI0f6Iq550Ikd4VkBOXQSqRCpOWRG2umQAWAdW5czkDI4DXBH7cgy/fZzsnu+
2SRStgondeSMlg/kFeNwV8K0+MIuaru6Go4DeXk7xwl6/fOUUYWKGZz1ILXFzMhdKG/AD/WTXe4O
rNDK2dgYVwZ1+/kS3kPquwv3E+QxYINCPasPR+e0Ckw2MHbPA9FK3UHCz4zQcuJm+w1hrAva/Yy+
qNkWJmHvcyJqypieNlEDnCapDV4KQ2UE5zJunCuVcFWAqfx24ZkpDzsC2k656/OqhOYJ5vUk7spd
TFiKnZD99D0TUhen1q+C5fze16H38ISnoMarqzBqQCY5OBYjX42fcyBThLehMpU+sVKpmmgQSy07
RCI39rHqL/qDfYpBC11L7d0aoTTfX/WhsneYUy0r7CD69YMFupPHnFf+y9+Nf8KZ1VYvVSG9UqHc
H6X1omTCO9xRc+MVTV8Eddo6JU3G5uAWCOrclEWDG4Bnp92gHl9Gf0mdocbxdIrWdhLskTkSVOSP
9nIBN2VqEnKStMXBlByWPyzL76oLJwMFMmOSXSwTDUYI4IW16+X9OqPd4v0F0acl64BEOZI+8IGw
VJBaXyJA4oEWCS3CTkg1oxp2o4IxwhKa1p266Xzf1fYEj0K94jtptSJ2YqIokF1nnofj1kkMZqkq
6SBRS+EwNtmK5nbahz2U2oHWKCerOxR1c9zZl8OkZAivoEALx6TX7YHjTcuqmmyiR+T4Oi8ec3W8
qodTdbVKhDReV2mkJ4r/RNblc6Y1Yg2PRrYm9FGysRCeclJ4rBq7uzaXh9oeMQh0sQ3JyfTpUvoL
OzBgfeoBj2uKnb4JC4X1UqC01LBLFORd6Ey/7MKRas9zNkO/80aTLBDdDKtmOrhvRBndFHNCHKON
GkQdKo4AZKcKErrKFIUwbuuWjcym0epWZe1b/LlyBo9sNCSoKoFJ3CvfdR9gdO0jsH9/rBz9EqyF
rBlfgfu5YbYJhu8NwUrWjWho/NQLV3nJ4BmXcMxqXarXFvBUqa/hIu78CgQDkpveGoG9OUJDvtGo
FdYxYQqhgNQko5j+hEuQ2NiSjPamTlsAxv96Kcs1UfH1wnp8ANHwRkwEzaWVGdwUhQfYVSTUv7sh
pN/cxEh1JcNBbqUFPYfm6bcE7WaCT6w6qE/9KwXHCt1vuVJ9GJuSOEhu2bD0Mcd1rrhxD8ylBl1m
Jzb8rG4FCj6P0ZjVWNgg49oCz97Z9YFIcZOsclHAi08qL5CNBKQp06XXp5IzBXitKydCoddq/m32
Qgj20ztDll1ii2dzetaJ/0R8Od574eU19b7PbdRjQrKSVg5UBMYBOQnZbOaiIc3+TFbXGh7qcLGB
KPWYdebtz50V2IE8MoUGIF17KPhrq/Aks/dUnhTP1Nvkk1+YS5vt/BCdRA/JOk2hY/omZ5Q9Lf48
xqdawqp6OaMU4PIyFmVoMQHH9UlHjXeu+8LLnJuGCcQppWmC7u1jVwrseN5hfh4GsgFFAuQSD5UW
CQ3RZFO81uTnAStMFM+Myj0sWmd3ga6mKVbcwGGE7flMVZ1E/DSggBkP0qVGr6yL8fsawLR9PoQR
QlAglNrUaZvuGuaAd324U7VVduidwxVO3/r9QlLCk0k2hniN0mB6SvVkra0J3g6ivM+4dx5xVXsl
hX4e6QUcXZnOe9eb+FbCuhEY6x0tg3LUO69MVumL8IXn+ZJUbCPs5Afd9Ea3cF1uBO9AsbgRHyy2
LDcRgrnUc3h0uS+U5cEXEAIaWHP4iyWh15DhSJIvSXSENLGPL8cfip2hxEyLdQPrSJu39vo5Qf8t
YW9Z9b0zcCJSx+TA99OOU1HGN4fOCZ1G7XACQtkwKdma1h9DrEA6Sqr1AmSAmgEADHmPdc94vE5w
9F5PE9lH7ZVpKDEruiZ+VwIBYmhYHnUV/hCc8EUtM5lBiIa1J2B6pSIsd0IMxs/iN+Ey13mtnCR5
XnKldc6AifRpu177aXlFgDYWJ1SQXmt5cmNqb/G4Vyv7wto9QwG4aEn3sMNmtv++mWvaN0mzEAON
hFQ6Qmpth3/JgxHfK4vzeVxbkvGojG8gruuAO5uXBVHM0zEtZjpFDiYKghox0PjJ3Rf1nSFbEIj2
AqmVvxT5/ZqMKUfs3IC/rrR5aKjzKE7Zeq4P0laO4hk8SZVgH0vfPpJSdu6aq0QjsECiAjIesmoo
wMRtMbjnhSAAxnCG/8CJHDsNDewTd56GdfojAr0fp+VGCpfh5qpvsiPBVgFhxCQo3bQ4ARD3vSBv
wuDZs44nuVtEYQw313dO1usQpBImtCZ5bbXfXgwG/bRxRXXLku+bgfwN20SuAXLTRSr7jogNUE+C
mzEJzQfpVp7oJcHatzPQWPbRZIg14c94qHYX0EsphxY0QpdLWZZqRNWdc0rBFxFMZEavJ4lEUFUY
yldiLgm94cGA/k0LQ40iJaiyhpdwr45ktFQSsSUlbQnaxK5KQDOEqRU6TLqyV4/Bgi3/PB/Phx6v
IrUUmqXExV4nkYRgQnQQFlJRbqiDpE6rlRRBunT/+11qaaLwFupE38qv58E97cBDP9vwScf27NIw
Ulhp8Qg2HY/sdgdqfif5ogqUhwZa6XhRiLlEBQsV1eRmYs2FVMOe0FGgpoiSknYcOvZGLRzbnA7s
R/z7aTfbqB+0PORkcDszdhWxfOO2WdETO8LeED9s1GLoRAiLF8IYsO55bAHX4Gi266YoI3jjb9v+
wDiPhjxuPM/UE0fRBpCXzkdkS3gpLwajQNJ3GCiMPwGJwd8aU3Rnz6mvQe1Kc6DRq32KzGKydbW7
0jta0pwdeWRzPHfq2DIlgCamkc/jg+0c+wkAribukJKCT/sXaYqds999G58xQMH+VxhCrnyM4POH
vLIsp5IOK5eixUk0kt9cv8mbaujrRkRaAhmqq7zfhzgowRnIDyxlOinCku4Ahp9K0LbbD7/XX7MN
RMoXbY+fZTnsCeP8/v6qy9NORC8GV0bygxTRz7R5RqptZYFgaUnEsLDZGRDlfWSGUveNIBHDnBja
m6tX4jb0p+fD9sbATEMB8KCtKMkojgwgEdVgeJqRy+Vh2EVS3QCO0pKAqm1ecmwjdGeEZUdYs5Cg
DZxWKYovuTjzK15wYZdk+pg4EHKbFtrXv3f7PgV3eCA1X+zhch7WY53aRemqO1wTqUE1VCwP1/Yi
C3eVBmu2Wfu2msdII4w4tRMIzBLxcaD7nbLvI4D9lJa1PB99TzqKfj7pBQKWk5q0tBwscBDgegdD
YKWXqzYzNyKjAjxCyX8zxWlSgh4WMzWQQXI40TnB+7VomQPxs6ohOPTOwPHs2OVrOogQxiw4wfx1
oy0H2KBAk5BGTWXCpgW8/GP6AkoU4ZsQ/ijPKooy9FpAk7ZZ6VOkGxzlrji+rVO2WaNCafQD2AbK
uOvfw+qY8iYpBKQpnctInp53AyoTJUWPOOjA5LC22VYmiONZodJ9CwFpuxXbKApUc1xw4QwJ+fM6
vMQNahFEDOe7126AkZDgo7zH6ruG+iV22OH6sBf1DCT1en3QLuAhWcnoVtwu7Ny7Yuv3CrHDkfs2
P+BceDcBJr5vWWqQM3VlKMyS/Pgv6R6CBhdEClubV2tDYKyDub4t8sA0WoLoiBwAfgAmuqMGb6b7
j53xTm2mwOXebp7UxGsRHtif/znEJVDMtlVkCL+SvAKeZe3qialDZvjOVc/YybbQXGS99V2kAHtJ
gbQz3ZXMNLsCdKOxcMrV0Sty3sygJEJbCSgiu/Vce/hO38gxUdIZkPslvGk+xi4kz7R1rURsYaWs
ZrPTa/Slu712HqpBPHVFBjUdOwjQC8/X6Fz2eAi+VYuvb+4gOxE8jMK5T3f0SC3/w1+3E4/GIH+a
mn8laZx+fUkGk/AgbKE6t13xscjAQbm/KBmUDBxVN+YJHTiduiCXhGRqriYRAp4xMF9VWPdbGGN9
bsO/fMUbOMqnQo5m0cK/O1HsVpq2Cj/L7ewm63UmGVde7Sds04gfZjr1lWUKo9cZUWfs3K6AMjY8
UoS1U0VMaf/Ri+j47nBMbfFPRKjT11F9iM8o+RHBVXizaGFYjJqcVLw57UN7jYG8qHOIuaVWtcrs
Gf7i/0bUP5/JiIgO5wndeSNNWOBV6/yQT4XyfQyloa1fJceNA7x0rDT/ehLS2avUNRdihToMTGrR
Pb9VL3QkSzfdXFJMzVackbokI0BU2LVOgjN4+rj4WDPr4ZfvfpgOdIUDj4WeW3YvL3SB2HBydJSq
zV4JVa2SRwOsp7ys+jcrDoRzrXEBdnVusw+SXAJ1JkKSVSzhtZaT6NXnC5WbQQdhJiTiobBJTegT
0eJA1W5w5eunGXKd+ETw3kuUoEKSlU+NokfWCFbSb9eUORKUnxZCoaNZuwpT0n9rTLUG/5d8bKt3
TmfI51sv2ACgRx4kBoCJykFI6+oBT1s6NyuIq8Slpk1gUo0dvI3hDrIfC9ho84a2gPYOlGCLQF00
UmaIGE1L3wpMKo/7j3Px8AUXvViRy12/BmFSsi0zOkKsNUh35cWDnxZrdFwl3INk+xqg5hF9ymrW
z1nLC4sfnI0xJc3yEPSz/LabQioenmnOlRe3++5TjuM+lYoiQ4U0VK5MerHciEOjZdKDKGR2kU7f
gWp1Lge3aI3RDbJus0Aqha+KVrahnINf3x9DtOSs4hl9xkXdjUnr8oo47NCYnTtnxq9KLu1OL6F0
uLi+q9uzZ5zlyJx8zOiK0wfj5PnDgfMxOhxfVSEJANEsEMF/kJ9gFXtJ4IZIZvkmHcD1GyxqKFZ8
fcFbN7aTbifQURgA/b77jp3F+ImSLCafkItL1p+L6JRpeFpRiiojwi53pYC7NakW1pAK+KndhL4r
bii+6jUQGvIiZ0DYqI0UkvthsvoRCYVX3NJXFA1hX1f7/xE67K+xhuV6mghe5g6OcE/YvfYe4/Fg
+hsyS+RNxn8p+1IV6bnlW6sxUjAeLP92DBse7F7a0ssDgx+UmG8anf8GuuDs2yJ1tC+kD9vfEpZG
bJZfyZAgwflv6qyKgn0KsJKx4FWBk3Y5ul+xtaRJqABIpWtLK2vznuPlJLU0dFKOwlVqGLXNesrR
wubM6mylOxgX7/fv2HYdQSxSmGxUrI8G54MqJDSJScWs/ruz8djZ67czNbwPOjVg/JTLHzqMp3kg
4WhAPBVDS/l43BSE1ghncZ2Xh2tJTY95WGx7OEs4dwiFy4F9dWIWiRPYcG5yHtPJmM0TatBjFDaS
YvykkXu2nV1JM5nqK/HJ/8+z5EUbxTj4T6CeYNbSuHnXK5iqhZcB9TOUl8atDuGYPQnDABILVHRO
22Cy1Efxilb8GorRTpN3HigTosFeppRmiCcpmh1LGxmQi9M0pI7Il6I41RltyyVuEQs12b7devgu
FEd29TO8Oa9MS9EI8z6Ic+SdOLmVXgkI4tEW07iPlz4MV79M4ajnsabbWyf2EyH6qHkMWV84GnaF
EvXLm/3PSPTqQg+KD4E4zH7/AUaU4e/KQMfnJS1ebTl+5sJx4SvDxof+xBEnPC4x5+I44ZJoh8dL
9h3y5zuk9QNpdt45x2pubKXdD3+cM85MIXNOBdUm0j9V1tu8GkOwdPUaOwew3p6C2rqTxQ5PisSr
PjmJqk2tS3b+9s1/wWnkgjEghatMfmbq2Ss3og4D8BTXyF0EVfcIIQ2a4ptoMKh3dc+9zH7PzJwC
v31Rmzh3oNnO1EurBToBt9/g/4JdczHLzcotoRFq6m6UpZEHChfouOkhqxMd776LYFct94pNSbj3
SqFV3fbYQC3zYxMNaur3XEjCrIcaIsk3SdPwT7tx3/CqzrzcZ8JsOuI91Y66qhU/zKlDpgktba5e
L6xH+I0k0QSE2S5vRWUEMgs0SEL30bfAAnEL4Ga6eQ/UrEon/RUr7Ea7q3vrcxe2VRnQkZvky6d+
8ALLhgt0SramTwv55kxqBOR7kRCpwB7MePfSKZQOGFqcB1jtH1znPoJu0REanXVlSxzeBeyY5EOx
vCw46VlETeKNP1JrFxWhRKxBl2Ps0hcBlsQraA9yku2Z03Ks0wZViHnBne011jIQLdRiAgyf4XXB
w/WCkbALAjeUKreIsWD15UTZoPppI9IRcM8CoYe1Z8RvNfUPgC13dUKEG0COHeKgaWE7Lu0CP63D
tKzfso3kHwEGi4pszghwZKKLRH2je/Pl44TJw5JnReZdBagBlBMKyYJGA4uVLNYTYDKn9G0GjpKX
6U8QOmkH/a754lLixpmDkAwNGQqGlp0jvlnNvEu44Lit5fyU6wy8uVS9DWDfXcKYDTE4D2K88HZp
XslO73D0DQKqIVs/8w9c0qDhMx7QMBx/sXgxLU5R4WY8R2X4hi7LOgy4vecozCIB5kFWSrWfqAva
pOJE4nf3bjK24CT0gvQM7esgVjOy/utW3mBgExO172aCiRcTdS1h40ZeklBzq4cghFsIEGAti+bI
sIhL123WyTLISbkdoR6PnrODTTM7d1x+W4pq6Fd8j2eIUTBQJgUEGjePbRAH56p1/zzFHfgsW0HB
8PGfWkr7jHa25SWM8w9IaB0Blzu1sLm9LCWOdmgn+Bc7wRNfJwgRu0VwF5xt1SLuqlKxb8jh5OOY
wHlPpAk+xHno0c2r6KsiaVBeczb0Ww0uSPuRsNO9d1fcY65yx+vaZbVWmMBeuya2xnLh2/fCwQ/t
5jo13B+ATaHj7Pexvmz7CvWESXTJY7pR6IMryOviMczGEUkjEDXmh8HYMUXuDcY4odW68VYJQLLZ
nfq4QHAXL+NaDFfkleUp3HKt2lN3Q8OPHOA1zc9kdwEljRgf+JG1Ux5/JGr/p7LvjGf/43TGNnWs
cwugj3EfLF8vCQllXRmKatiaqmYvXKRJ9Z/CGiOQ1yGTqoq/meu6SX64ZkxBaaYsbr15fdVoqJ4Q
DMgYD7kg4gX2fe0gIozHnrDDYAY5VE3CeI+UhNUefn/9t65sAZnB8bSYnTy8Urn7h9KyNoGT7dvm
1GnLkpT1TTG4eE/FCz/8PgYpWQhEyBFwMfgwMFiO9dshcaqMRjVSrpDH82Q3Jje4gkt8X3MZ6/P0
sxqxVQ6UhJv+4U9zrD+91zLwfBR4j7pIGcqFVr1hBl9bjdL14JgeiDplNlHUESRnTDwhfCPD0Lxg
MHHH2GtinwBBH+kF4j2kVMQIAsV4aTDzH54ZBUJZAAA7mam+K9LNsfuDBnPVDzVxbaxuZ50aVhVc
U0TbvLVoUNHM+oe6ohTDem5vY1HMKo9AJRmRhBHSsB7EQKRyqTlBXB5VijIGAGkCDdEaQ9j6S7wb
f9dUKCuE9lYAjsKRNcUPiHRn/R5PDquHJqOckIZT7xWODPrZqd3PLyFYldB1lGOHQh1UonQ7uLnB
VbDF8K9IcqYsd6jv1j4LZLLSR6zbVP0K4oTTWcjfgo/Gmy41Z6I9bZhk6lZ8CvYOWS4Jc804qluF
umh0aF/WfbFp8ZIPFEHQS28Y/JJq96wt1aNGVTCKzmGeTZauJBRRHNGUJ0Moy4GOIOpQfMs9MgSE
AcrE7xzbzswqz4MsDQ5txtH0+ta+t0emPwwoeqHAsfEUiWvC3oSAyBlID02nahCs5zASW2Coj5Jq
BFsgiOExGibNAOyO1z0TCPHPrNFFDGCre8hHtyXPWko2CPjfl/ZFZ3n0GyKw6dO2nJF3Q7D5ykyn
xSonqNzlWus4BaNg4tQUDCcezj4frq4/Vf3oc5TSRcv9CW8L4YxSOkq3gghm5HFKl/PcnCFtas/8
jBBTTKEyDAmyBDMpQrc9ZNTeETwPdTfV3AhN5SS7EdOwWUUvTZVC/c4SrKuffREA1f/SLcWyPyHo
6RQ1tZlB37RsHeTWsdBAljQ+rFLIcPVcU8DHuPXC1PeNEfDQeSP6TOySjIW/pfub1o2K8kTH9TcD
D+mpMjJqgh/i2JcVuk3wGBeAAFJzWI7UJMVilEK1I7P3tz9DcwiV80GD/RXLtXGXzziZe1c5mzyk
42kw5Q1ghBxVjCIgjTIcI4Ru98cD+45RRUxGuEkIewqAx02MuxZC8D5FP2/NLZK/UJIitNHGw1Q4
wo5yOC3kyl3Cw2nkhDMLnIBGQgOmp/ZX/k5LJV2XYTxMLp1pcKMyqPVOOqd7PcJDE4nU6GajNwBl
5njD4ITvG1ThSllbCSWeppry76QKgxgKI6pjvtcxcg62eWpVoQCpdWBVegAVfwTelKdQ5jQiFvSw
d0bRl7x4ImDmjKZPm2AOPvj2Ghy3TdjAwM1jab4Xbu+OKZk2bAnqbmv14xCYY7cHbqEfR3bpdVsy
+eQSDXuewDXHwgsYUIVRRWG1mIK2FY4nQFiJDZTRfO7F88dj6nsunSrLl7PJhjYHX734bOaq+2P7
KuTAXwKAH10J4G/CC2fEKSq6IDDpp0DOj55zQVVsvKNCdhaCaH3r8DsLFJtSxB4ZJGFPJWgsru+S
KpPgSbed/vURZNM5Q/G0M6UM3zwkmaduACOedjUsss+BQTl9qv1JYEpnch2zQ4xUa9HwZb+uW6fE
4vij8HAKGYmv0OAug7SzVlmGXjNdtW4EKVSfDk9+ViVbR1FKvBdVViLZs/CxvuKxTdJ9zpDee3Ju
mNmEIJRE8qCAm1pK5bXIHHv7FW3hpxyP6QksAV/yeZCk3goJdmDKRuGMFVhlV57TdZ9NwDE37csJ
Mp8ozjppJS4M6xACfDhVn8n72LnnCEznnFseTMWnjIm3B17bnb4zEqj3ZIHe0g8lAcCllndedVXf
SsqRxZ8tAr+4zPkn4Mvkp+O2WC9/SrtwhvziO13aLwu4Pa5KUGgctV92EwTTuzWqLR6zvQT8XXxz
k2Bi3Axuv++waLGp/RxS6grEbq2nuw3aXwOsIeN0xPXSrhjvvuv3t/hpxIZ/UkfW7NTHc7HbxaOI
bYz9STB0JnEWC5qOkrEpImcEotp0X44mZcqU6xCxTWSZFTUF27S3LRa3t/ir3/DY92442emd6lXy
px8//Uim7u6cLERvxc6cg7FDJKRm4lSx7g6t3ZRnCom+WvrCo2y4ulpswsvl4TxPV8EFG844hFCp
Tzzgy9uDc6SQLNZG9rht2bIgHBwK5CEnzvqdPNsncItJS1nfBhj1hQzNOe4gq+lqj05/sWrDAdzW
QX41ScOTmIk7VE4mFqbFdWHCtXKmelQ1HsoE2mK4BkkS7SzZhaXEsq8wWN8Tb+2dHiOVDCFq1KeD
FToC1j4xlb92M5nER4U/XquvQbRqxUd3FIk7qEeSmZ6D2gHVvxvR3r4nyfK/hNQWPCk3RYtT90fw
aZcOBC7xivz1QrVupffxlvBRGlkML+ONYy4PLp5qGb15+lKNez230whjRnPnKCiiNbjY6TC9oLZ/
5t1buhukovV1i5dxzRKLNQmg62iEXp3Am1R5oLNMG2VVh2jXKymodcKjEJoaorpmcEx32iBo46rG
ZpnrvAlNHMPYlSbxhJA41B3YBhUTE6nQ938oicTuCpW/YdAQ9Tz4bdF2EE4h0euDlFEJksg1cEjL
YvlhfXyEXD+tQiq+qZL2/OMiT1Y0574yxFcaHW5Dq3x7RnblsSAeCL/GYKB/abyeXswUPlrweN23
fwDWRFdzJCLC/JLinpfg8X46SOPqkCCdwZknCDiMHv5TCtweEare3CjNVievRSF1gooWG3WkuqZD
RBuZ5hTU92LGqC/HAplUWWZuWxED71XB3UMBEzCL7VAyByXJguXe2LKEQN61H41ce/prMd9jW/G3
RR2RoXOp6F8w6hFwRH/d42uhHmApzyTI9B+GTncHvNP7jE0d/rUTjVzz6GxQvaY6jb+zKYI9V/3V
jhxiv7Ucy6JRH0rhPn+l9jpoHCuGhPxm/J91LYIo3cx9wskwa9RK0DTX8uPRIqfaXvzreun4NpGb
hRVVNL0IOquhNZacORYWRaZItSXhUc6lTi4+UxmWp/gJmLtoOtv0oBpbvfSdC6VjF35yGks6GBwl
LQDHBGJrIv7/JvQHiCce7lBr9NhtRIuYHVU8yUqaESPlAa/rbwQ8/4XO7pr++kEeB1ygq2o5MkFQ
7+jvw2yySWJg4Oylo1SIzairUPL6ET8nSSwWTp25xZQmjJ9JG/qN+FNR0VBWNFizJlNRumCnEC2b
sD28WypyOB7Sk1s/5Y6x3GVAfcqIuhBJSUS1RaXbi8IfskenO95rEyfRrJX8a5UXAmM44PgaduFU
CNRnpwDB3lWdxYC0G7NYvMRqGmjEuIQRwvG5kOAnqrNTMVy96cEm9fjynNMu5wlMuEg5nPYf6rSV
lC3RBbwozrWIStD0UiixdTXOOa3SGuk1QttI1APYu3pf4qIaNI636wBK6YZGvVOuqD1n22gCPCUb
9LoUR/1JbWYoJKveTkIKLUE+ue4qAPfPfrcwYNRX48kL00JiFUYnPyNdPZh+IIWSqk7Qu7jYa17G
woQwaECrYRNPFtf+DSs5wr+l1IcIqvuXPh+/OVKdESNQSdbEBVimdh0g/aWqJw2uOghwmvfLtXBi
hsVIW+w39TRc3QUrWHSxrmzOq5TnjqUUYx/LT4WgxYc3Oznq+L2iT7D+BxnGehnfKnqfXBtVhcne
dXz3wW9kqXGkKy5YAV9IlNfN04OSpmpvEV+qhP8TZHOyQ8D5z7Es+7SwGLSdJmRMVSHqb5zLxJCJ
9pMNv+vbyF8I+dZwbERBuoXW1xSlcrzRhHLHUq77Pxm08qHfmyaCK+yltxX8D7GW3EpC5wGbFYMh
BO+SV44gWL9gQBZwzMjoHvhNeAy5LFt8SGr6Nh2+nLT5k//3krqjradbzlCuTLadnDXko+8gBFCA
ja/GmXwOMcNQce+4B64d8I77Ia7WLkawwJasKIZq0BHFNOf/esYsRVBnNOkImIiAXkE8wXDH2rFW
FPNvrrmuWZIujr3xVuvTl5HSuLitdwXCXFrvD/bu684eD6z8aHeRBPiAjzphVUvnkDCrjXQURMxb
grnmNGKVlaOUzR1hH+7u8/IOy9f639dQeid/ASbVXeM7xH4IM2j2iCD4beYfs9gUkXmh7i8mQYfa
5OZwZ/Ll1Q+vzdzVRPF/u4gKU3kCVsHD32GJEtdVZVXKDwiEZFxBpDCFxwRAg6ROlUYKg7MXg52t
PoU1nOnZ4Od/p/U4FOkVNkAnIxUofurG9ga7BmwKXUZe4s/XsdWI2WRVV+ujzpLiNTiYFnPi1YRx
p53H8VuakvlcG70YBqH61RkQ1wJgIMmr2I/TNDOCMLxWGwdE/2xofWCZ4We+zg7yNOyaWPi1fqVn
bue/1aZqFXbfI5xTlECSvWfz/dB3TVDf+v4allMf8BKqx0XW2YUqtbTvklPRpzuYnToYFfimKKuV
LHn771G5ZtCFbWolae0J2U0esYVctvuMa93dA1LUYPVgFqD+3+qbpzXAunSm/tkS4rclFR6+E3EO
XmypHl5S3Xtw+AQo5V+ZkKF9jAro5ybOmNCdTikXi18kNYZCHDxpb38CgF+PM0u5oQl3VZipnTcN
7xB4KEm2I1Q7/GBLnJHyx9//gaYbMDEg2crpsTa+cV1LderZN1dvYXdQnrNiD4SnVwof1UquJoKg
rDTlQBHRze9tITkaLH8gcmrY2zDi9LhRXwVtQ6fjGzF4m9CGdpkoITINJO1RSkKf6yrr8Va4J2FZ
0zkfNSOR4CEz6z3R/DDeVFnaqQ3FxeA1j9GfteVYBSaYB4JxSipGA5MSsgAzZrjP7qz0xLy0fOva
0czxeLWXPzn0GPvgqy0l2GHkFA3fXZSDrpOqtxVcKqyijlQvri2vh5L0aLvbru3OMX/Yxg06Gt6w
EpyK6iIofRsnZO1F89xj8BG8V0cbNi47c+Kl/avyDkKw319lLhKHeBP7B5pZBzcxYKMEQIOjrBv0
u1Rsxb1f0QgwHRjQrdXh6iu8OMSLtp4NyMq+RWMWE7zW3RjxaIc5Nx2QqS6kzsQueYwHv3r62tJi
zZfgC7d77FeKdxPkKLpIK597K0EiwkDbv38q+DjFundYNSr0coIrIFO2+6RmlTJX6chnLZmBZA/W
oHiBHYjU77IR+obA0+XcE8zDlpQjH/ZamuoSnrOlKfceaWMvk6zJVGsNK1UUZUuGeRAppOWkqzXO
2gAF/gG4ggByn1DtDlxmFzsWtM0eWRTZmMRi5KtE4gwkgm75EmzzFGzsy6JYBBJufv79jgeW7OQQ
dT3AihWWoRzApPotLJ412Br6oAJWUZob3CTIB0Fc7K2LWqpuu8egTpiQMy9+VFr4rf+dA5MYIi3z
Qvmdjt3a7D50YmAwvohrBTnTA5TJYuK/uin3VtEL1loKTTwOjdZyhqIJA9RJCRuSgfenAYaun6sT
bbzJkXBoLaplbCIKvrbaI7tfayjmHaFeCEbrxsaUF4t/Hciy7JxlQAtsXZ+itD35ZDN3psvas9of
rs1gsP46gMUjqe3qjKj5Gh4UhybxtSd+oBbXiCQWGHTKkNkIX9q9e+Z4eVSt4CElc2Jsrrxu3bqR
lRV4ruq1fC7+cR+VHvg/15/9qtFRYgnKGjvU55XK6MqwSyjkZNhJ1Er95rGiaMn9+yHKwoZC3e97
M/nHuHlzNOn+CTF8OwbVYRaBbKoF119GsTZRFTV4hTqP5fuQVDeOlDr5OUkqNcMjeo8qfIS/a7R2
6puhx3xGDVlYPzHpmMc7sc4KH9y6jtE5XPFt9bCi8gKBdYdkd6DfSPx+6w7V4IufOIFuM3+JaPzK
64zPHYkrOrWb0XnLta/+8dzvs5zFxt/GUrSqcnv3TDl4RZBvRXeAzQIcDLEcsnAvdh19zBO1XRB7
F/O/NvTvE8bZqAq7eIL2hzFDV1Yh+kK6pUQGANxnzdmHOp+q3w1rmPbh69jKI9GsoVCdoFBh7nrV
osLgAMZbr2BR+l764UyhsgnwcV8Db/CvWNW56e1TX319KInQaItDSJacrfB5isfpLpoEoDYff5/f
7WEVRGZzzWPrHx9tQg3uskJEbOAtIFo7EfqfWPu1cDTi1RbJk6Nj20zDjH3ujlHMIuZHTgO7Kml5
7LB1Dmo4lh7wkr1HQuURPaPmvlIX9xoNDHqsboinNKvRLu8bbEHumivwDrjKPLIVjJigm1pho8gT
AgEuzS/2GQtsr6lMKnHJvmZHekFxfdoHGUV/kWHOMOeVGcsbXPW9/0mGqNCr/7Z5d0Ti+HgoT5fW
LVfu/JXmHXnd1xOB8+otRDQQwboqJlVVVgyFV2TUt34694eGmfUZ4LxKJGehUEMus4z8Nb8mIzU8
xbARioG5rkoRbcfo+9Dwc8qcUceZiJBOn06+gkXjeXRh/Ewq2b4rwTlunFNpt1qT3usC2qkcUpuF
EuTZCu+8aNkEbB4wKNpFoY7I80VozpMLj+1gBCQVJYyCiGO1kIbOj2lBpR0WP9NHFkp4cusKRgRV
joAdK1ZqCP2l3aNt7Kr8mDTuvqQXCbhrad/dh0wK8Nsayibly7N4NG06QJdvpZiXq0suFrzaDY4U
mzuawEEeHrRsTblR/i0zRLU8CcWexCW0OYtsfaXORcSUhax/EP1wWmB2wW/l7w/8pIIbhewVo2T0
yhi5Z2kU5tQ8DT2rB6FFE0vXLtBv0gyZHFHrnsfgrbQKEVlV2TGudTZY+ftBM4s/p2fD57Y+q2Rf
ryqPwzOWS+/2sxL+B8MEtW7NtWue97ZEp3RnbgmGqvpzyad5VBPZVUZw/4etlW8Eve8GElHajT/T
a0MW3HrPp9ZPdY5kEcm/ZvPZ1EGRZRSaFFkLQbiOPTdTW/HpUDVw439KwYub/ivBZSpqLHqeJqzb
eEo2OZmaTseMKikK1yr1Zp1P9qPKOPPpY1jszvOH1tQSt3KM3igzic41E5ooQuixZJYjzImrIjtg
ZlMURGEfcEsTmw+4dcZ6as7022cxOsRhWNBUdT+G6X3eYRMgbmPvBwve2B9fdMH4kor5cOYnJngo
DVRlETQhmDPX0PWZRO0A030OgRmeF4yepNSpEUTmuSXr/C2Ny/67WS40DH3aqXk2NuK7/cs33uC9
10ulTRuTzoEmTV4xdJUwaAcfyEpjmEqDWkmIHe6iLdQvZ7ERjWQCywOmCxpeXpsKXF382EI6AIzV
MrlNLTBTOZfUKxZkPsfGWheRPD0/WkVyrBNnUKXicRMtG1RV8K0UZOVtxGO3LDeSTbxsvjomHteA
k5iJ79N0iZGDGdtL6EbP2LSJDIOfwh75QX32aimdHe1cE0MVVBjVrHYP4v4PerNT101leszAtnR8
hZJH5lbxHGhVB96euBqpd00/R/Wqs/gvTNVdFDHTMujO2lwgUZjqXtUcP50eTm/xzIpKXeAvxP0+
Ob43YzDBpqy1NVFWWAlm7o8E+/ul9DLNXWDzPRJhYSDrM74F83vg5/Dtmt1LapTAIWSpO6AkdRHa
L521Ek6C6VljWbxa5moHtVQ4mic/Jp5Ccc15Nk99cJMDFab8OJjXkg/SzSZN/6MXjv5Z6NgNC07X
teSZg+BNvaCa57zQ8klTRuHf2Y7SAZuFNuTnwYjbKVCIq4d1OmCewVx+OVg197v1K8x0gvSXMIt1
TDTqYdiqiv7kXn7S+ltvoBgUL/+hHKmdRIBgcQFPEpqZcuzO4seJoyKCfqyl1s6T7AIvRce3ykFA
TKJRi3NP+1bCjorpfc50RLoEaCSzf1Ciqv90Zft1gYcGg6WDiKbEnbe0azD8DtvGg39BQ5JFgX4G
JkopQSDvdePTNe0BAxaO22dGOMX1ZvRjPBNV7RM2LqRsQkL9xMBkXMy6UUMDJ1y93X8++1aSUWmf
h1h5K5e4b0q74zzrlDZ0+8OlPtH9F8xIUseb9vqsBSVEpY7THnYcxCRLXECyc4o5uYgsvfd1kaLv
Q+dedFtkCoD5509u2UI5akP2uzAXQrLd1ohi//GSTvKAMZVjOEGN+mktIaEuvooAo5coQe6eOXRa
f+ByKZysTFsxeMMFNCj6afvY8h1maYBJBna5ZT4K6dsFGaEtX3maZrjTpdufv0J5Z3vuB2jLvpNm
e9a6VORWsQLplJCmDt4GRh+vdDfMTJuB2E1ypdWMkVrfF0SKajh1HMH6EGZgKhqNnyf5VS6kmoeh
7GgZvvt1tvPE8V+P4WxdUkT1YPk3Clwf7uyHh9xTRwBxjNKmU6ETRUznWsaJ0cc8tsZgiBbXfINE
3PKE8yp7Sz4srTLeBuxZ0vHTv2B8Q775BoDVRaFY5af7WlNrZtAfiHAFivURCsq+rMWEdRw4CAY5
neGPp2Nd6k+jr69BxF4pmnwrrtuZ4Oz1HpNOCwA0E9/5/OceOg9Z5n0wx7TK6plC6pHjjwgiXbvh
nVHA2wFX1CN93LxKGjVVn36wXkEAMh/TET1boRp8y1Y0ojtY8wY6H8PeJyM9B5NmabzDEiuOZZ8l
LJV5Cf8FpErcR/LmIWAGSfl8McTlpnnkKzVl+n0Jp1680Wv8XLtIYLx+NdejWCAi3IjQb9tYJ3Rm
FzhC/4RrdswxA0bxJUerZkBDNyQyzQbwVWpa55dMoZwQ3NeQ7T/tjMKWeJ8SKn+xQFu/ZmQK4rh/
wG6BALZU1R3q/76OuGtsBIbkHV5zIZndF+rAOYMuZotnKcISHhSW+yDXN/4OsV24eoXUucQLT5zK
gDto9FB5cDzE1p8X8hb7ZH1bjsVokrM7XlLo9WbBOxqAtn1eKZQMEIjoC8NTHVdZrrA8P9+oVhpH
trGyg3NCQA/YAyBF9Voi5hhoWAkAijdq8B82BItE5So9i56WbwkVeu0nds/nvrQ7hYt2OSkUddm3
5Mujh6qviQzD49W4RDp18fiiqtuZMrLGgu2ePsRA83EdXZrBULmjM8bt0sd+RXNUKOMBa85VU5rO
IpVzNH3EtEJ3yvKjfBRkdJpFaweyxPdzataWXo9rQnqMdHcUxBn+WptfhL6UsNVeP9qAcXkBMR5w
dixbcUpCpClIUITt64swYmZsP/hXKDCrc6mIv1UqfXYDLqqxPmV/gvnwe1bARLCianppDKpAZbJH
BvOiuACHRnHSr92bJwWkYy5BtKSbmpd/jBPBjpeFZC3OOdZfiTd02xgv+x8afZQNwqGQG3CDmEJi
Tc6hwzUVMx4P3QWB13cBKcnk5qPISC0TeRaAwPa4QArZQE9YXxHMEefPVxkUJlDS3Ex/G2NXV5S9
L0FmcsRpsnou2q3u1FDWaNjHC3Qi88VHSuCjmQtU/ZvUjbdq2I2Cg8XncbOcuSsgecVs5aL0Jtvd
FtP/d6fxkal2daqIaO3aBGqRfxwCkDtaJeryX0Trp28ExH7xxj3+zQIH60dyLA7CivSlHYnYIm2l
51qNBUBHNoDyT3zp155LtroqR2XhEAR/CuxFHg932yTaxT9eov9WwmQuAa0MYiPGzMMQlXlLx6kA
MOK9iwE4N1CG2xEFfj1tbUZTJ+2OSHOLGhAh1tkmGiiZe4XnBoHdWO2c9n6IdWta8my+2pocyCKX
xC8BX4CdaZ2m4txKD/c8F2mJEHAVRVclPAw8VkXoJihKQeRiCrVl8aWMUhWxP4Zj9nhvusuH6O6d
2jzsVWZcIQC3o1jZ99XurWX3JxoejcM7FxAKqxv/d5dvCttVZEEU5qHQ36q56GKlzIH626U3l1yk
IZ/TCqXxta7VyaEPR4JPoC8lJNhBf1T5NSj6RlkhkAaKYLGSEdHwun+8HF5bv8o1DwKjuXm74WGt
bbVv+WRYmAeryEUS/N+sojBdLWa5adxeflT1N31YlGQoo0L/BLH7He+fjiB4h2UYJrejvssPf6ac
m7z2XkpADTZ/tgvA9/otbWaXOI1H+OjYumS/8k4MqURulG87YLd41XOzPrY4d1Xeg34bJBhMcNMU
XeXFMFqdAIFynaxnbA5j+sFeZgCgO0Y8AL2ZMpMQ6sHeICrVhxEnX7ICHMMF+nkJOb/IC+wRmb9/
dU0FYfPWETg4uSyxJ5CQ8RZnLNBvzED/P76klispaHhOKR3Uq8Yn8vfUfIvJTFeR1nECFlxgQN70
Uw9rdju1EwcILQzpY18Cd2Nlfe2F4hWcj7Vgr+S3dAZrgZucW4CfrbogRLyxflwifffBv7RApXUi
oTYFTAQdJP2JuPVLn5ec7Xd6wkg1wi+opMwXdDyBxz0416vmBcEOQfWJ+qQUplg4qtERQZPpeirz
TIJbloP6Zc0+PBGBzy4xsVctx0ROqwDGpL4VcbSnSBohyqmYLOeU6y51a7LLQ+DQghOQxccIVF9G
sHxAdjZD89JPNPYEdvp1ctBXlmoBbrHdxQpACiPCEk82+Q7Sub+InjJKeS4hIkWQ9p6n5/N5yAi+
n7HrHzC91kPoFTIajcfwMJTb078h4nJGavlwp2Iv1xvHu1kXGy4/mnSiRGtcEVxmO78UlS3PKt0J
sZf67YquALL7JpyK65tLrHHaGE8avppWiLy7wfmDDWKYtPJFDsW7nyjwlrFV6UA60eYTemcjt/YP
PESj3LjhBLSE9a/01aecMZMpZ2Z7SYog7v3fqUh+etINFBBLGo3EgIJGvEoZNsqeBo8cie3N9u/q
KfjpPrsE4EVZSdYCJLjvPEkNWY5JD1CN42v230pmFOioaxAYY4yL1sTSL6auL2oypuyDv6gjSlbe
K/u1RPdMJD7LavJeSmKcKjEO26FJ5ioZQRo/jRqlYIEIELcx1XKk0mh+jkwaVzN5/HSfFfXp4QBJ
SEXRh83ywV1LGpZZYXCugJ5KpmPDDjC16PrYXjkcZmiNJ3mvFw0hAaajiORxE2nQjHAEv5RqJ9wG
yZs6IEg89cO7vKqFZuE44ZlcCvtyTZ7MFqLxVfDcuD9exPp5XkPJh+RNIkHcA/a2PpYW5utkl53D
VXHAjqJpE8fy/7zQR6cDTY9GKzOw7XmqR3rQb41FsrdTjr9dtN2QkX+0wCg+E5wWzuYFXimku4YU
VkjSscygeES8mkH1HSxxUUQS8/3tsd5TgH8I9C2b7VqKTCOcrng6a8lEz5tExdDNO4LGVCtbf7zt
9cEyRpZuzp1NWr6dWAeR4v4HRm4y0JHlzlh/5FDuv/EZIkzE1lHZIWZkeOAiRsywr3K35h81NCoi
jYsb9SNmK/OXzXWnRANpyTSDiDwezrhj0v800htn60uncK+/isQvZZ8DFBQbvPaVRWZTG4syvhA2
mpDyFzZAXwnwfYRuewQzcT+P43lwqRUkOWIszEfe77cJhM0f/jAQPJyqkL1EguigzED67EE73Gbk
R2XhX4XXjNAFX1w4Dx67QarSYoHH39OhjBHuu2fyRxQL3cwvCfITECfJm4krMqepokgOgmqKQbyJ
ERwdiF4YBOlbcxMngf2kbvEHsu0DwmDFyOjMDjPz+0RiFtGp3SEOIm5Y63dLLVdEBv4z8ICPPfUz
A+TXU91tYoKtRLgijYKDS9l0aP01k0vZVXcOmh2YcQtvZezNqVKf5RfaCW/YShdBKMuZBIm2xyJj
Zu4zAnezehvZLILqry0HGrQ+YjC9O4pAmfwiljtAM0pEkuN7/isqUwPmy3CqQOujn8OJwxC49W+U
yyAkt2//6+NRDRUMmSf8TugrvqI07Ov0+hhaQtUp5xnIrh69u8xLoC4TIaToVhg+syXQ7CjzmOaZ
sYdfmQDOHFhRa7PczTeHTtHJL/Gh4ivAJWejg0Aoi6nme/nGeZc2k8lKcooRBo3OocwGrnlWonDV
+Fk15UT/ol23qzUYJlpA5AYE2SDLdfbjqGdFT7NvXhe+dSSmTAiIuXQF12fLRLNoOiDPatYEsAWF
udne151r0hiNznE4+kTFO1rDu8xNVLTus0E5gWMdVZwWvFOve7d01/gob+RPUl3Yf/SUlFd+cINh
Ad24Z6nD+AfyTSMFJc/y4X2LvsxkLWa/htGLCxGFz++PJp3XRyRso3xhfQkLarju49Vz6lsa7lvs
LOEOR6O90fM9dg1Z1DKC+STn1bYnW+NDYNNaYCKHM82jsOdqBDeMgoxT/GQ2rhgCFcUaElbvQ7Nh
g9XxqLZvQNfJBN/zdJDRoFCORFpeGKwKkk+juZ7lATkcnOC+89XEZqz0AUdE6oj/IPgSePPeOVnm
SuuggfjSijgBdEeW4Q+6J+wN0npu1BDq9P1bBCzpvYGecsF+aZ6+353aW/prZnHYfyDyZ5xcX/WX
aId7r2VbssnqSVt2LLMhd9CGQFv0d6eBfmkVMZyeGkq2nXtxsM//wLdGHJS4P8UQZkJ1xGU93LsD
FddG6D/QWxZ+h1FQFp473fAgI9to7XFM2j+JMgJX3WzJeozXm2CUbxz10c1hwNGBASGgo47DieCA
AucrT613YjZlHN1/XIimqMYafBSxZZfthfLEj+qFHII1zUARLx9K76+wuL0t6S90Ha8JPylJmLdX
kTPXkV0fs6v69EEK3n8LNS8ohOl7dj0aXWElkWyjsRDxLzWp+XHov0+G9YaB3glsUFuARthNUnec
GbQbQ4nxn2kgHP5EKMv5YPsk+tZ+FxuyMwip1WpJMx1km5GzD6dNS8x+XhIha4j2ZdELiK5xPOpE
56S/o1zzcUmNSNrSdwlZs6aa/zYyhxNFw/liWA4tCu5Kw4z1TVR2KZHsySWiFK5qabrI9paJrabJ
JtEdmnYt9BRzv8XU1m4oIeHaTjP8i8ghsMVFiMYn1xF/dDWemOFR/myL0YlU7ZWvj9LBn340H62h
nIFy9zoDt+4+NIg6fdG9EjVpf/1Arxow2GIMB5CUKr4FSyWd7K1G2ommXUVvt8ylkh9yCBFWKzKY
+PVNTO/M3A4is7JVEsvqhUWDqwyKSyT8ITX8/5Ue5wuX1DYUijVrcCinVzZ5dF9cAB2Hok1OETkm
5EVgLzot3d0Vj5hmX3RgNKkOBOB7u87V5igd1ikcx9DUurz8nLEfsBSsqc3hXH9GggnQc2nenmGS
T3GxWNFIXKO8mKDJtOb08qOTMYBCqMb6cDQpYbpE9Z2l4DJX3x+vOdiqNWfNpKHZg/SqraIStnvg
HP6hR8tR0BqeCdLS8d6wtyQfUEjDlNXi/So5I+KTtmSAFLztDnv2SQ0Y+iNfQ1bbLxioZ7mY0T2e
NXZk+n1L9YjwZSr2XyjjRTU3KsbdZQ0i0yeRqFf6fOv1P6yZMA/oFAMK2UZFlnZDkzRjRCGoJdKA
Fiz7lud1D3j7m762gisfna+zb+YiyVsLQ6fTG0uUoLpQz4pAqgPVju6xt02GVNkI7Uk5yhkIgnsT
GpcG/0q6nQNgfh0EFGbzkgB8Y7yTyIesUJJxB25xjzEgNcxI1LkN4rbg39vI3DJ8Ys6aRY0glmlX
RnomCCB4q8IBAh9vD4SJcXty6ufJhuSgn0pwytstJ6m1JYhbS1j1IaEpGx5EQde28VWkwGpowdkt
Gej5Hl0s+C7AStP1MfEfByJQNysxynSIB5uNxBNSFzyvyadU80bwHQtAzuMo49OmZtk7wC0u0noV
0muvKw9ENcWdzYpQXuxKCHpJhabAk1e5WLIonB38qmmr1A3vcLGFPoe/5nyYtx+2Ttambf2DviJN
UshcYXvto8rnJ3BrTEakoQW74VF+oqhzcHI+wvkGmESHMlgmzeonhr27+MqR0cehIGGzFd5V3IJj
EGtNDfeHpha3MxUJ+jjH1THsX7GS/y9H42SwpU10U5DZbbkMzXXv4aJiNWuVQBh4icIhk3TQ5Jdj
S6mMOUrC6IgYJsBXga+HxYl2JG3TdiWn5MEMvF+tCUgNja0fxTKvVxf2JYD/mYwXmntrO0oDIp3B
puTWO4n0Ei7r/+cGRVJd1iV0SgLHtD8264OsIdI/qVh27CFxOLObAgMpPy6TkmFs0LviUnIddoe6
3yxbSHLEde/NTT91rGNasbsp5qbcLGwH7CzBLr+ZfmvrgeHLQ4A2Tfl1t++SKmpaqopglZVGalSz
yUdwQ43Fp4wItbrtc2cyFAgE6HM7suOzOIq2k5YKa29muW6p/V/TuGt/NjVnxZt52XjdmLzLe3fp
eotNp9WdHva5jKJdG8Kqf9xaLB6xogxvIrvDDA+fmGdUevSWyKF2BgJ3RfJcIG127Fz1iSTpCv/J
3xkx2U5aQzDpE0zlLQyO1dwB7SGn0O7i0g2HAxpFZd9Ee19AgWqerG0Kf6jaZIFjHRw7oDLb2D0q
NqQ/GlWq/p1dLygVOm1+/rp56Ir/mk1DybceUvCBGbcQ8SLmxlECFQZG/5K11JY0DYUmKhOgYWu+
IAm7qZQB88aKKDg9D58WE8cErw5W//m/sIW9MXbOQNH5SHQE4EsUE5THyR1eXlusT7WnGDIsQGuz
mY9RQ6po2LBOlAelYBfmx0TbM/dZjTFbxbcCDjm6kqN4MqFl+kMrudQmt4dTrUXbd0HblSWHLu8/
xnD0H4DQMla5QWJ9YSC45lb/LHn9ZBXuRKaUXyJTQ3GAAn1A2ur8TTkTttW9ks1vfbEJufiep5ro
Y7CCuXTfqwAmEvYOX447RjkGJlWup1ooXyJ1DFRXWFnpgc6+0ADN9Tk8XBU1+RsF14KixiZGthZB
xk2fMtjRuXmjWEMG6ZTajn+EFOEIF2E/yh7fAqFKLmdXh8TAKS2K9oIFKFbK7FtsGAmYmkFPya48
DCWxCHz5UtDuznvBp9c0WL91Q0+SH/7odF5SBhkwwXOokVt+mqVP5/1dFJunFKH8pPHyT7LU+ZBS
J6MTb92E/xAsrztI5bSauVq1/jcFdXZEvCFsK0vfD7Rj/6Ow9aL8OqDg6IDI8Ay/qu5BnFh8c/8E
vlu9y7JqKSbjzwrVGT+40HB6t7mODmDChS08A8a3/OvVh0oxbh5QlaYHXPBh8PPE7v7vlcunQsBc
iC8OYTLk/MojxLI6oZVh/e5dVXFo84hRuzyy7FzAfcGM0B4DQBduR8Sr4FmU+Jz2VvHNlqo7us0x
N/JAuf95biJ7xE5HyJrqRjkYtG47JIRRLYZJG1EgZ2w4dvl6nFvadXoemx4GRCPprAZJKnVPrsL1
DTJECnacSFOIZrfakq9IXEYKT/x/0xpFYm/Mqs/cIdDjaERQMtbIho9sT5oUR+RB9TTieZ3YYfPK
k8csP2p4W8TTAPlc4Z4+DtKmjUHW4ABZT+87XKRSGkUVBTBQh9PPkGU08JtC+PiO15GTPG1eAXHI
X0P8e5AGGwnt8rujj7VlhM8PPr54V16lNTMw1dXbdCaxEvSFgu2TyrQ0i4NAu+wZzCp/LNf+3GrN
gSlJHaq6TFE3e26Lbzho4mo0FVdJvlztVKlkltEjM9nEfYJKVJScQOMgjZfW7Wk7cm54fKMDeuZH
xhSJdqh+WqWZ9hbR0r52HTwrbzDkDxovGJGgkXb0gpo1gzSJ+ivnHf4RVXRSfXiLVhWleWEDlsx3
oo7IIEhQzD1dp/KqNlUsWjmTtojm6aoCdI1VsWnO0vzI28W2Qi5KdUwNDE14tD9Hf0NCOUz/8wzj
TbaT4gte9bI40ezk5v+zX5eAzFUgAj6X2sp0Va20cf4sJa+f32BWJ7/tmOOxkX9VsS4I3uKr10Wy
n1vmiNQrSlmsqxxyoewg7a8pPWfAjwVm+iZ0PrFwYZneDtJc8cmctog2y3EYrF9v9NFH3BEkk/8a
+Uow40yXGOEzOzDowjpagpvZLJ16sxO0kVDAexsCpzjpHwGQiUHZyvP/im01pemsr37VHg91XCqj
oj4aEFdt8dtnHlv4K01JFTVkXqGXutYeY48S6exoHFdSxp1wO8Res2CJ2WGtDNlwJtB9AhuWjCau
oPjp1crfjvYQteZNKHttS5HBkjvsMoEsPL7b2BrBxlmzaxEqz6HRhUwefrOcC2y/+TRxMeGX4fQf
jhB4rgxNRI8KS9vkFUTgnUo263HsrxnhmSqRVzZzhYNuPgAiNEbu/00z8hSXXJJkG5Oyfvh7yaMw
La9f5I+iG/DL+Ge0TugXjRulbzuoZj13lHOq3hgLhKl3711x1oelk/Vd89a4k95qLv/Pv1qPq4GC
SEYauTDc/Nb42zxAYIzWGsn5LwY4MpsN41wTGV2LaOEeBwQZnejfuDOuFrel54wM5L6vR26foAfa
alSeD5oYyHjDtxx+JvTB9fB3LbBa6Al/hzNn3XYghuPv75sg03BZwuNlLd6HsnpGteqUjLjV52if
WuKsQGQ+Rw6hwYjk7Vnx5ix5Z0F89lGd0qA3kWDnl9jcyebeAH5TGyjheiZe2WzxuUtvkLW7PNvy
5oCEn6hANqjn75A6W4QnHr354nZItvRiXpu8Ora4n/o+ECJZX0V8kTT22kstUV6dSJZWOr0DiBdX
6eJ29UeUxmT9bZ49c2EFkZE8CfRqro/q+wggJtMgZys2hDfWiTPZa0IzGUa4PHJ44JRMQMTwSZny
mdiqXFeJxVBe4WK/U6Gf8QAeKd08p9NtzUO6RDeX55+jcF/zlXPQ4KH9a9jK8dPBWF6m8qMjTAFq
QE+YISEMsjtLJonafmhyk7vINUfgbBLsLTRGs89Qxru9Jx9PwU1ipYsJL4ZXjTGhqSlRoT6uW9PL
overmqfDORF9T4Mve/aeS9M1O6Z5NyxllP+meHNIAYrhUMKTMiybUDcA0qUfosne60FBu6YafQ7p
yL5dPhGb0Ri7F8M88l6musIYDfDvEq+dZ5WIVeF3U7hxrJiIicECRK97+gpfyDC1c7u9rkFIlq9D
25kdKubo6SfrV2AwIcoQEwIb99biacuGmMTA/nlQqM7L0pHOdgweWPh5WfG+dUbLrknZL6fUlKyS
fCR1DurrhV2oWo3MtlG7+M1WYok+YLt/KpNdZ5UWcdZ7pdyzCv6hpb5Oy6mPaJ0c8VVySRya1SS7
C1/FtWnQCbZd5nwi097GdJF0tSqPpBX61D01gJAILr6yOAwsCevYe2j8jVXUHAKej+zFXK8JhT90
+vq3rLIaABviyLiF5kEbBb5ETE6EOrJ85QkIN9O0bpNgrTN9uNS2WrEmHzExVpgHhnpaOmwooZB0
fNjypLtiyziFb9ITPWIMKGIY5viXHgZvEbQDyHvDyAIEVoBPCcMwG3UK4Ob9tvObVmOEQGthpYCL
PYe7eLPG1yu97SRd2IeBARoCITONO1MXLjDX7sVuwuvMwseys440W5ahQ4a5vwX2nbg8hPnhBBWa
wj6ixJ9TmSDneboFdulpZcfUwiudXQvwz4XTLYPlpr5Mrd57wcE4qzkJi265IFu/0KN19DOdVe2O
XC/5n4WnJIMgQCLclKWZnTVnELTMIwNXVf6ZWl7b8zIJKPmJIw37SZ19YiP5onRFGV8RMSKu9bIr
1OnE/b2IUvj1hznQB3NybB0AEAL+/eqljzWqqhAVhomk3Yp2Ry09J0PyB6SXRtQE/Mpk12U+NvjZ
ATHYtLNZhDkYAWIyrrfIm3npuzvLhIwb625FLlzaf1WoFHvqtyreHD9ADSsh0YGxUk1OxrnsFrSH
66fgQOqp/69vEzcBEZpHLEk1bqWua8/8ryf3+gU4mstIHKQBt4zhLKkqOcthpFMxw+66EtTvHCab
K2MmtWQ/dBDuxJN6p301JvU36Z4Jv+EKlDVEOLIT6goVW6iuB18uf/DI8ArM3KahmrCwTrXUuP7x
huJCuZJ7kYFLYYe0sbXyJ+nrXDRCwjraBzAkHoi4rvU8y/lwACBod8Ar1y7nHapp0LND2s2UjR7D
BFe9NVELjmVh7PptMpynzbD1I4x9ld22CzHrLs7YjfQKmE0gMTd95Yy44S9HBCfbV1Q+b8aZf4vv
xjPsGKY0OFtprJ/Ah8Iw3J2cykv3Wwm0PQwJylvdD5MTyuvHG3SwptI/6gpOO/vs56pOin9KsQHL
JSy5wKDpBvNohW9oXmDxefxuAUfmVzl6g378pEae30A7tCXCaXqvVJ7KmnllV3KC/bgtGt4mOaoD
Y8w1/BTdMpzm14vdZtx6CwTCKeqoZnvkmmQPT28y90/LDcJQl3pveTzXl4utO5U+uuqvREp7a+nV
ftV8H40pfLbMUjCrL5v+isGBATrAtqcmSDQHVfg2RUn6P78sN+nD5X+ZojG1EmTFluKWdwUq8gJ/
kmU7QvRP8K6s0yBa8bkMULCuepXi5q4zbsKxn9t0VQ1FID2MtKYDTBWFfx4PHqC9Ap60vcH2mrni
codCKyLIID6zTGz4L7ayQm7d+Zt/xGaktmRlFn6Ve8rFj6HKRGJJ0Rh9jLe8FejgUbgQLjvHocfc
xPNIhobZwR3MMf/MFEtQwGZGQevaMHOvNSjJMhE5hdcEiIdKFGquJwo2J/1dNVLvu0G0ToukrKbo
mB7Tp7f77TCHcAIRy57xF+xff6S1SBWBW1BKBN+TrJjrKQJnPwkIzydBenMU6Dghc4LFDOJcTbmX
Ges3ec4uGEPygTs3QXn+XuOOk3HjNgJdWuIxEX6rPdbOukjYF7R3pSgMpOgssRU/lMEZrI7GN+AQ
FZgFjCM055TZpWe/tfQBrspTXbnse8aYpr6BgL4b1KxdNZcvQgVPM9qXAX33nC5pcW6NQwxxNubd
4klITS6FlvbKp9REqRIhjsHum8hKfT2RswCqgoN5hiYZC28pY257qeZ6kQn7v0RX9tsIEX1GaC+e
I4i3YRyVzZg0K6mz/fWpvUUM3GPo3QIHyR/upSL91kCIpxQeujQnbuUXj4p5NExblYG62CrWQIH+
Re5BwlM58Puas6vvgMdppX29NzekFKsi+BTu0uXmD5VUYatyrnXj4HJJs/jWs0SiRoHJRrzPpi4c
CeKbr+KeCPeUmA1Ut/UGhcAKFFN+1dxvrgd5+RELjEAwnUvFSm28hdYnf2j8ULkAEHdRroZRAxwh
UXBrhVZAuJNQWpCNbDMlvy19IY1ERa9T9KnahPBaidwL2JkkqtnywF5ErKliAbQfj/sLvfm7ufLT
vX3fsJv2EyGFsr+FKdULAA48jBg4QHnw2OMYHHH1RFtdyjgqXwdTMs1vpxI09US+vHDx+3ZSAi8J
sAZFXsv5RTAmCXexh4b/t6w+E3A+nmt1h6jzSdCluCCd6m+1PiRPPwExPJof45U6GSTXzMqIN1aL
JGiHIZlNt/OA4MfqxVCrIXd9iDQwvupeoqz+CjA2HRZG9vffeiBytfZLheLlEW2qVWlYMXNmB1aM
RLuQO3rQqnXKpqiSEEMKKm0yjy+VvACHmPntO8PUYJHz6BRObkLRKdohVvesP/vkjezPTrAf6RFF
5KTwhJ0MAT3NCY7h8RmIn+W4dD0t7F2MibGXIMfoIqdioGHvcMupE+KNJ1T2vDHxicdpJ+0KUNsR
fpHCADXSlwsp5/Cu2XQhH58xxvMkAmfMKQWHdWWqtlAuxLzDZo3SueoiJr9scj0r5v5VArK+mHIo
uTlotiGOm5zil5IFRCuWpsyPzpjI6n/ECbaa2WJVIwFTQpZ+YZ979d9wx1Lfi3MUjjZCxjt4HgZr
bT4cFQ68GwxZ8luQbGrrVDy4Q10VkytEnaagdDTT/KubBJdy/DQvjItqeGIs24EOxExXnIGOs37g
TjySgHc39sbxE23l9tZLxc84coRFYIIJydfObEMZ3OwdBN7m5EKaYWsmRwJdms6fmgGrwEVzWjzK
k38DPrVBByKkCiWpbWCdC9UEkg2yH26espqjIZnJn+8cGvb/R3mXPWDE8Mqs9g1xgZWRVGF8r7eT
Q3egrvw0VyoT/UScIrWWHtzcbGMaMYkgSIPCJ0j9iukEz4J1W+clNOC+9FiLe4WmexbG3KcyC1E+
IysmoeEg2/xrxA6astd7liEciPk/3nSjQKpaTfupPTEssLnovOpOLsgT1lXmXp+D4uPI7sAhjTZK
L9uBWLrsxqSxMw13b5QxXEigVpuil2ZRQeeBxPCRRBnpczBFC7B0ZGgx42uWFQuFrkZ6xVMfHb4q
67c7Km4PJNddLIpJBCEpd088ZouUb9WLtKAqJltFykd8YnFndEt7Kl9KopWuekz59XqeivVLm7on
rNW9jFqWZyLiRO8XPglQ0AMsPkruUvgjG8KpbsrRMuOm501rX0nkFzPqhYlV0mDHJNJFqHi+wzKr
/Re0kO3Dnf6STU8yVLoZAT6QJxlwc4EcyCJvzGA6h9Z8PHyclA0YzZ8DV+jh16jxRSfJLmpqRPvH
oSo7C03/JIvEc016wNkJOtlXqRGkAZeXxPJEMVz7yKCHaeMYCA5TfpNMbQ17amx4PGlNWYFA1BMe
aVBbQRIMA7mbIA+REQYynSHYruuA4lOxaBrAtUysfmRoQyxpsCBBTUOzzKf2Z9ZRShtWbSff94pi
+4jZn8QAOHux8GmdS/fXZfUruYCTHlKDLSoT5kAVLZv+jZHG3AVjgbQmOYbmwA2O1FjFKWCN1Djq
32aZETuF1LZWJhZiLRZVlaxBopOImsWfD77w7mZkMUxe1zQJVM+Ld3NrSCl0CpGOdMBs9P69umBp
KF4dBKv+96I8WfM4/CL8Mpa+igCA2aUjUk5lZW5owTWvzlDxDZlWCrU1uAa9tRgP8YhCKcmxAsSw
eYywWexG/li9BNou7oOsdnMu1Wsr7V5/JFqXTj7Zcw9MkJf62U2tnkfF1BUQmv13FPO03bAhVcTC
yiFZT2I+FOZsmeVXLfS/qcb5Z+M0Y1bmnsfkL+mVWvtpKOMymstDaOF7AcCE2xECVu2eoQPIHzeO
RXNtjrQ923MhNb/4iEc6dZG5CERTd5FIrXsHSq+qDpGLIxeZWAdmW0fK5zG/aD3+LKXvJCHEcexJ
V+AXmQKCgsfmnf2Ox7hr1WWu9mQcuP5KBQjmjXt7hdfpy2RPa8t9b4GLnVQmaSzcSlbmOTecWc5U
DEMKknOxv24NvDP42q5XOa/ziZ5GrmQ38e7xdbgpcH33bPcX8+3893kP4PvtPRSvHZt0BxCgzZHK
HPNJWlgOU+yFJcWr0+v6ZuYrm1bHkGfQmRiKT+5tnvVpyi4qWfLA43+CQ2z3YMNAatFWSQ4LyGRR
6sbUVE5E4g8MiQ1qCmEVJ05ZwyRE28F9ugUkG5F0BlsgSNa1khPN95t5Not4MrO930uP/XNzkwjD
2yIWvksI7jk8/5DMjLlabP8kMA3Wblxiycu3UWkWD864Pc1lgQjXQhwMTz8AUfR9XRVupXMTFv9D
WSYwfDFnRqgae+RRToibFCY7tCZA8CM0cFHDpIgwl5U3PANlbjCexnzn1T9Sk/1z+MTp9kPyCGdY
eJ9haw1MvGSwOaneptHlRgw8UyANakn/H/5KD87im+9KICPpY8AP/2EFfY9D4tpabdSCU55WrveH
msH32M4zR8PsferaQbAk3F3YDh9nP5mP5VoTk47z1itCb0w/gdigll5uRJGwJvJE7JGIlmnw7iXd
KKvv6oxR37B546X0K8AiN91uFtz39l8jCRg7FtkMxEyyjwjNNwT0a4MUpzYL1FIQhuyFQHAeOgUd
PahWMXDdEnLKHf9UiDI7ZX8pDm2jMiXd6Cz6B5iYXuS4D/Ij2xsUnemdBY3NL9ydHeoT/vTR1LNk
jBrOZLJDg+O89szxlRRUJlVAlu+cXNbC5fsw0USGSaSgzuSenuRubPuFoiIO1dungVGWeuM8dSi8
k6WSkp4GNKNgkelzECtso/0/hONsOf03xjAdvZtMMDfoQj3erfD6OTIfzmEn6LOZzNchOslF3myC
k/9bySaG5NWBbvRb+KhLlyJ8fCvAi6Yu78WS9AuK/YEdK+H0OoaEWMayUfkTdF1l7jMlxntG+O2O
khetX0APCqBrt9zXrRJJpa4SMaBWW9ad0xZ0TyGx8FysLNy0VPy1iGbWOm0E1cEtjoIjqaNwA6iz
Fk8NviY5QJ2OxwRkd2HCXTjLGp5DHC5gpx+4f4NZlaouZ3f02Xo4+7T3R8IQeFjw2C1MCyLU3ixc
fZ00JfeHZDbNjp5LNg0FL5Cc1BOYBNQIbPCF4Nqcf58p59E5UB+cPM8nDXcmkI3FKgdcTTyG7riC
SFxvh0fEr7pGdk/BGI75LQBd6iVxux8FWOMetYE0I/qAJY88QqxP/jCJSF2JlIBoi3Op3OmCNR4O
4/vfr9v8AHxPcIgImFitIuT2A3pHEeV0WqmBJ+AXBx6UjN2mbHg90mssGSaSu1r1Z/A+Q1HSUkSU
D+VVzTM6VmJKcjwSwGhuUqoKoeqifRtnmUwlnMoxiDJ8UomfPZBKj+lr5TvlXzBzMfkB7Hi+xZIf
DejBI8tezudvTKzm6GHPIQYdzeferretgxKwMB8QsZDAsAxFv3cSGthZZOZ9ibPt5neZxm0C4E4N
PHNVQZhPx94rEJuFp8rSJjufSixmGZyBK6JWnCSAM8zIUTagwE8fcoOD557vru1MP/2iW9Xa1UnM
QV+jXSZQtfEdV9+wlIhAUAA0NEgRcq+wh8+abDXZTvQWX2viEm6TixMQPvdt62MKhtOuHPnREf9n
jWdpdrA29LVSMs8YUkDtxVUMra85xUYdHH+ruOZN9UEB3u65BAEebSVIN7vOSlvi5+07S+i1Byh5
fOyKJDXcUuuXCvZgGEYjK/s0+UH5LEHg0uxYB+H5FTi520BMtvH/sQbtPsPboDTwohMNQuL7ffsu
gIWVLwWivKmTqqYXsO4L4Mw/Fo1aBLv3Z7TGNt32x7eZjyMPXlSX1k2I6BlWN6It9/j9WsLChAJ3
avjTHzBd+4nF1eikk8/ARnOXkAyd7/tLTCUkOWrB3sEHDCQl23J7L7z3iKb4F7sVF5mffUR4/sX/
ylmtLTs+4xDvWX6eDgJ2MQBCzwdX3FA+jG1xEMvAzSGMhR1mlMNaQvwK5koJm+9HqS/Mp690ZfOg
9cT0qN0ukcdAPvPcdoFQwXnqBbRSmy6IXAkdSPmuITCuh5s1RByOpX+zISz5oPtQNyVz57H4XW78
QxnA+g6wWrc3KC++VyojLwyrFgHGM0PukF8KtY6ws3UqH4ZPCljQQNSCAhefzXtjLq8eWGNGqYs0
HKl94dN6J5be54eta32DHSC75+PJt9evAnYZ4Drzciys6pNcgL6/Dcl+jpwEEWzXqr2hghLLfR5y
gxRi5q+xopyzVCy4sQDPH6UNgZL7gIAURTgab0pwZ1CchZDqpU4Q/nI+JyEH7tt4DCfiziaAXDXV
XTTeYD0n+FqVl+PVd001xojO/12mCcCmyI13LrpNZawDdlA1pYHgwMjM5V+4h4y00Bs6zX9bbXrJ
JXzjVqaytrRLz5f3OTyE2jwgCP87j84CuJ7AYXbwV+bUFbb+2N5V2nqy9yUaivkMjtvd2XWZ/l0R
Y/PcPixhNKfsDu+Je4tCahm16btdmCcKZl6fqvIgsjc5aFIxXTELOn1S5818kpng8YUBALya17Xu
jBJtTDD8VWpy5gQE9lyjOa0RCL5BtYrDcHbpGL1BTgSxcRLkS5fZFPpHvB8NP1CqyhyC2LjSJlBK
Md4brywZ8TIB2vXH6YChEAEnKw4KiQg78pCZEMkHQxxtLlLOYZUDpe5YdcV6XcwB1fozdkgfmbmQ
5ly3HENNJO6UX8sO3PM6TDR2a0GLtksLcal/rCAA2BrFQ1nQSM5hw+tUlSCnu1A1rLLuRSCe5/c0
IFS4mCH0Fc6Fc4zitH9JU8UEjj2h4P8fE5RleJWD3JXzh2dFIt2JcIXsZ3T8SwphTdrkYQOY36Sb
8UXVWCEZqslYG2IOZy0NYkV6XqCgTj1vRI/dTJuj1qlhNv4i+zT6mfDjtfik2OZ8p92WuGFlyL6s
Gw1nQT6AWN6ACK4A8kMYLzBfkX8waCn4A+MWWMm3EBJW9xmuLfuBOVGwWeEZzbSbGa1gdtgrcgHS
snt8VMPM8QZwmU5Ew9fitb3VHtgAq3Xavg+h28N74/JqhfCJJyclR2NtMdi44j2kRp74doAkFYqO
D0K4sTkrVEJYh/mlSm4AHm9C12h2iy3jBXGT7mItuhM3JNo8v4G/2ZeE2oOrcFypHFh05ElszPJa
wQsNIHYuw71sLeNJznbUhAI9IryjVb61OfLNHQvRbUbu900DYIrcEH0sBAjA/GmvgEAL1bwSv28M
nHvuOXfqEGNfkH+Dqrkb0T7geRnlXomluwyNqCo+wU4HuDdGU8umF5e4dBRVDcdtwUy2D8DXREbW
jV6+Kj0XNpI9koxG3e+kJt8KReG/ibsf+bM8PspUVFdMIJ20LkiIoGbrNUspyYhKr3PIyoxzW2m2
mP5oiDgM7Rv8/F7G/QYpIUIp1yLQd8plWaEnuRDVzDpLr+Osyj7AzV6FH2kWDLnUPVSp5FVufWXr
rJpA2SZLDxs/kX/MZpvCwRuJ7hDemWUHEUwd9f4D010fIPddfV1HDYzIfB7KEcmMuwb2UywTc0mI
HXIbd+S/Y8Nulf+gmDPUdLvGHe0dZ1v5Grx7/rNtwcDy/GL4gLqPR1p3dijMsEaASgmUjOIFs9F2
SbI2/mtOn9w7tchRpszPCl2Gs+dbrAMUYEVFSjGq6sy5DB+4mEmKza1ULuI8/jsk9EfIZpCq1oBB
6XwXuYbChpEh2L0cyg/fOAF/ZXriiWeA9gf90tOidV3xqeLHQmcPZh4LBEEYX8Oy6zVF4V/5qLKv
rJ7dgDzElc4KztCANbIJpd/14QgpVOBuae0FACaR+MkbvuZezyHN5ITS09ndYkY/pa9lRYoOXt1q
pNZEvBKk54PuUYGGrpmuEc9eMIAPlOy2RVYDeLBwPyO/Xc2oQklKNqQaLggJDafeWVtGAKKcHGXn
bXuwgqUfayY6T0h/Z6qvgnsvio5TpEcdKCrgCSV40JFJ0nkmm/ekbnsrN/QfB7nx2m+lO+Ds8nDz
pUbEux0EITJrceET3dVvnCpemKeCjw0DL8qaOdw/vtPaufouiKQJiI4KqwPoe8o5klRuuH3hkym+
94t0ARVEvwbcB86jOAUcbEU9yMTurM61jxZkLqB0Ws/bOxDKtPiHBCbCXsFO9SCKgqGkkJtl+yFu
l+yc9GwecfluTEQ7PtOn/1DmhGyrJNzvKq0Zv4asd4swcJy//GdQ0RvFX1ZSH3smd35cMrb5lBt9
515G8d6PSZjU1FUmXJAEwwN38PTk72KTf3ObSZken5wDzAVJiQ4kPCPFcQQnEqmu11xFIDhdrWtd
40tEQIFYics7blmkpYwvLa+Hbuwj6I6EAjgALA4STI2K1rL7eExTmIQRBtmY7oX+2o1wXaF+FEOp
GjyottFcKK0CwEBB3vfM33hbi46Ets8RMxOsdfg8duUaLQUiTT4xzmzNs2L9V7CtRxL8PvswEzv4
AwHYIet0VXIVLAlVoCxrF2UCUHplKJEC1n9xyTt+wkj7QvJ960QeHqtGVE1/JOV/q1a2fS9Qx6NY
oaeb76+Oo/jIfan4PZVMeFzLtXSjV5WX7BkoGTJYQxBFJNLmrNZhr0Xx64qy+8mRJoXVk5+ac2K1
4ggoI6XqQvCuQvtb60IS0r1ahEsefBGAGxuKsgT0efzQ96oY41DQeDjB57FUlU+9fHY2DXz9z7Ft
1TfbcLaea7ZmLfw/sYCv2yggBGJ5hCsiqm4hLsvuvWEHwlsphJRhMwyLUbAI3PBajm3+Ro0Gs9SF
HJXvEiZ5w67xJUe6HE9tzCAqqOBO7UD+U1a0qgzh9NWFhp81HFHpPEzl4NxyPrZkSV1MLBIzUusi
16yerIDnY7Vx0mJ7rIPYnwd/xtZOGAsCFIS3tLybexqPoQ6tqDNfkL3HlNYHkYz8Mc/jKqrjcKfq
oH9fVTElA4G0Hzvtd3BbGjuL7f6oDadb9jGVu+5ysifI4zjGupNiprTw9T2kNJOff1EQ1cy5d8YK
lH/HikGiI4ljA5iMnByUG9Z396vH/CHViRBn8+KGgsBspJBTQY319HQju3PPSsmcOh8f9IL2V3FX
ZKR/V8L6Ac+YMjD1hMKC4DCeRXSUCHLwMqwf8lJRQJwvaFYQuWKijCxWlI1eunjBfDuA8MkY49U4
QVNp3Art0984IQmBUXmAs9sNbu0d5e9iOkXU797kABRY+Cu6wBnERnxKOZXOFr5kVg9DG3rYboDa
5OTvElghgDkV+I+LQXX4G9zL4rVOl+W4KwIuAoR9+B5Xr7YMpNKKg5hZmf6Z7bTZahWAdZNwTPZX
kr37SGzHSpmqFkVbeG1tAlPh4GwababypiZ45Rc4hoXi6IQMGop8WmPyDd6qOLyIdJPr8oaQo/GY
vF6F5q0/Ak2i9aSS/Gig0Sx/edGC+T5cp0XfQ9M64P0x8UUZXyOEvIAtAQS02t3bUqB+MqtKYQOu
XWX91HyTqE+pGjKxL11D5sL3Tfe+hxWv0sHU13L/gU/WB2NMLeSSFE6jvNkdWLhkkd2fx6n4DM44
FcpSBqP9xXOPjM1j5MYwWxryeieH7fzOuJTjrXVLNWTGnrpdTGmGJsh1TfQaxQizFvjZw1kzRePn
TBczcDM/DX8Xr8uN2K95EuTC5ms+8lf/OQrzoOx/TROBvHadhFUa74Jh/gr80VlXs1GFLWhHl3tw
hZW1u8Rzgy4LV8cjL/5K9LPTuk4SNq79SeHIT4z7zV7kCw/uL0rhDInP7AC8GKXbqMJo+6wTInk0
ALVrnSekkmwVtkhA0gQ7O3vMxa5RERmk4Jj9Uk4adRp1YCLmKDPeesPtLGDZL5YASLruO6d041S4
LTa+kSNZd3cH8U40taSwyyYDs0+R8PV9Tz8ozKqos2S2puMYHA/2V+aKb+BrUf76BRM3Ww/9PSbJ
w6dshhaaTHIEVBQUQiHR6OzVzpQG3UMkzAwGgBycfrYnxkUfZgK8AxvDk0foebsaTy/U9Avab+ls
mHLxw7SRdzLixxxauL/4LNisrv9UNM4pxZ+yoDW/opkVdJCcnLYfYdaSnDfY0xH400JOZLkXhcDr
MW1wujHSx3vnzk8rjq5c2UUolT3kI58JBtiHxmXvmy8w69DH+dpnOJ9e70iNkmHhGeGooPuhnl5Q
MBsx8cIciL379a9gvRJ/w56tMnPg9whxVaIihoPiW2Nk5Mlf3gwnvihpfIykQVL0YpQMvl9XsPWq
U7IU2NgJh4UE6Vt8W8WxeTMEiezw4zpodb/aN6LNms5LEQkqzJStBXAj/VJx1kMgoFR+Byvgphmo
yNTF3SFKkOAlKGet3KFR3zPDyzoMKgB6MxO+4bmm9Ukp/LeLywTs2Yzx8ubZEH0p3h0VVTrUuIua
RjPqI9ljCfm/1nZNDBhirgGHE879/t80Q51gWwZufOoXuVlplwfZ6zg5i2pv22bjzt6/cIW82cmv
ISZSJnT/AKnHPJHMEAOwF64etL6Funb0nSQWHbGw2DiRyJGnh1C8TkW9tt7ZCL+DbDSJDNAN07iH
5C+mykCRFANrt3Mpv9w51XvfthwvJ4x8RX2JfLBMscdnmIiFdnkXT0SLfIdlQW+1CbYYgMVPye1K
4thIFJQOQmEaPZ3KwAl/oI3Ii8FPbosbg21d6z+SJL2TmZuYVeOAm3RysLOYuC4vt7mAZ81er41o
7glli7dxAR88XNw2QWVMsK1qqxabWRxHcL/pD1nrRwxXh3Bt3SdTmogKnO3MusEWo5iXBK2gTH4i
137Cz22/9k2sPDjbkPXmv8DjSnSfucBfV5fIFPdXYsFJdM9H10Z+vshCUY9GyQPehMp1BSnWKoV0
Yosqp8XloLq54GDro0ep37tlJShjYt4n5QWZJAGHFbAhDGCPFEtwxUHnt5fqmGiwKI2STL2M8Vio
HfXr8XIb37YlzPlq0CQoS6FIjcxMBGTjkYUzt5W+rEq0ZOTZH3BoHgGZD654Tgb9rvbJD+1tB8At
VWJfs3L2mQuE+fdsi3CWKnKPz9qqqG+lkGpAyyruR7VWJax3uZER7VL6g2+nfI9B6VOvKbyEQIUr
q+ERpGzQ61PLMcEWAD7f9VjtphRKvviPjSk2ZNjx3iFjsrgYGtsln27IFx/7aevDYyBypSxP4wb5
FKXldBsDdZ1cA9JDyB4TxBK1bIBZ8fPKG+atin0PzNrT55r2jWarGCpawWE9yLvpVxquV2XQLMLl
WTBv2o4zKCRYAbNtdxoow1/UE84g3xTAzAAGYa/QR0BmXwP692chZ2LIuEMy4kyVkro3uzY+O6ZX
G+qSPSnbnGEDe+n1fKg41HysiNFF5vZU33AoBTHMAB3oVaAuW40TLp6Hhia3lNubjg1yfgW1Rdc1
f4Hgj5DTZ++LvjSFA2iuwu20tZ9FhcGLXYZK2eTPUFguIsMc7+UzO7GjGvoqQFbB5B7UYP5CVRfR
si8fKTY3j3dqfNKLuOu7UZuHpkwT6jTqkNLWiO2e0U5Iq0b+8pwwv219yHIkFSofFwpmoOIo9KNM
xEWnYT/7B+iKShW1bl5fJyiuNCF2UFPoOCZL0U2WsJnznstO1AmK3xH+h1vEku3F9r8HfxuX+iWT
Z75lVJHSWSTLfiXmm+n6/3bZXzgO8Jq5urY9xolyMGPJa9DgTREPClpFcj41oeEUeonidvG+hKnS
ciujF94gJVJ51yNl+EpJtMuiFg/ZEcm8TdMDb/yDDa12tQIEd1guK3Onshs5WzoICFZmT2J/aMJn
EM2Yjt8Q4ll7/BwcOwkuHyBHAi1zXapU0qTY3f5fVPJFX9+D3D7YoLhEkkQy6Vws2SfDAgcA5dhE
tI83SQP8IZs+ppl7i9YnNZWEo11cS1SaGjOya4mX1wnIljXZ9bS8l8p5HrPB5wtH3Dn0uJClvU/E
7YdiX13uEr9QLnemCOwlY0yIEGbcSOn3WFSpciXmuIb/c9LMYELylPYozchitWRh9sEYFlOax+oU
btaATcBGNwuURf5sLE/VS2gmdtuj+46YodvQpYLYH/8StsACJoGzqKZo8VoX2Vz3J8yFHgULmj/S
GJGaGjrfAkwgtsoH7S3CK2CB+uAxhsWAc5YoER4h4XeXS0Kqi2vm1g73wCp/hW+wugb/vS4FWOin
qaM2HPpI8Wj9wAcGHgpORsuq9GV2yf6Feq4u8hjKCHg9OHTL21VUanyxykyF2adnWtRNvciqXwgg
gSYM4Q3VzgcAsF4+7GNggdtV8zoemsKJOLJ7giSSRlr5DT/ves2qXK3vLfARp4XGBxRbLrZkXUYy
dP7PcqQ+4cU1q3/y3zw0Vp9078Xq+mFqrbSUkuA1HjQHhwcEMc7cB9VnutRTnAzAtJCL72bKienp
GN2IDplNRKehLrw4k92Wd7rUe/o3YNIk5UYX63T0+8Yeli2rpGML9nmukr7cU3dn36gy7XLqHojC
t7GNp07CtBNRl425YJSJCp0ynCrFPB2EBvSEI1wdcl6Tc7L2JwXvgp/lKPhkpwEOwMZuUG1JIWU8
9TRXhTU3eMPrkori4+vGbILdU9GWJ+r6Ex8rcLdkiDr8KZqME6Wqfr0DWjareFoG2+pGOJo1Qife
2xCZ+3arJx31HNRbmvWDMvEuJ2+YU12Cp7n97VOrwXSkxDZVMFuawD5ezzYX93Uxy3+CFCN+cDN+
3vA3HpfL4eFn7sRff07hNto+aX5vB1RmdRbMS+8K9znnS6sC/0/4J9/IJm3B72qa1T4mXbrZRVZe
l7WK9yese5TJFC93Wqc7jFcwvoO9RY+p7czWSQ1S38ZpBoFBErNV2+iLJsK5V4dR8D1qKEBO8z7W
JeTNYqt5Ih3HiEabUu6YW8WssvulMECarasP57sSF6zDznt55/hfRjw81x8OBBi9e2o30Sy3aF+O
/1GzrKvBDneTrZLUBuLuCuDBaGtLV/67lVhpxl1h2FTxdkaIIiKsQn7WeWKWUW9Qb+Y6wbT2pZEo
RT1SyvjjZjcKs4qstFFU1uV5uRJUWCIxcKM8R9pKXjyY5SGcxTYNyQqbjUvfqsuu5mm9e3xBALCn
gPVeIRxu/rwqEE1yt+FXAr8JWrDwMObwswx42Kz5CtNKgjNyiEaNFLEe9/qeUpgeIfoe5Kp58T21
OKdiwP0Npwy5JNpghj1NWY4IMDr8qP74T/d10P0hbjPYacsKCJEfil4ue5syStioCzE6Tu3V+HKT
L6sa3RBDEunx6I1mIOAcyqsLi0ZRgoR8GMRc5MlkMhmtDS9Nr/g3vJWgEcJ6D68+/x6NLhS8K1kf
R+qZMmSmT0Oo7Z8aqQtXw6yRw6WgYhDbnWFANuitxl54JWypVOj2/eQ4KGQGX2d3GAUvyYk2UMHG
3TZrR8thLQ8TfD1Mn9Ag8vxpoOh9bHnJNHLSSE3RCiHpk+QDtH/ISA2ePeZUbCoEDnfbCipJHaSB
dfXxKO9gC47cnT8SqFO/qx+Gl5CJAIgrM7Cfaq0bJ+9CuXXojcVR3rr8mjZMSkPEfJKKECQ1lXxy
kcpK6H94QzrLTEoJkYXZLqmkJt7f4jQrWHV1e+dRpVrNu4C7KMoY84rIxWuORJ8ivrb6zI5HqnxW
s4/7RJML91FYgt4v6t6hWtjW4lvilSElASjPz+LV7wEMff/MUm0aAiM02UryffB326qRTu6dK9Y4
yyeJRP0FLKugU/8FoZnVLTUg/qTgiiBQd//xkKKloCIPBZgcjIBCCGZ5K25M+jOyt0qgTHfLMdMX
7BSbH8O77CjwaJK0G4AOdhzphhCMMkhuyL2K9NRSC0yZFeYjuQI2GxL8S9rO2oTNfsmbOxAoxyYz
YEbaPTsowT9Ax4KivET0FCMLK83oXxy8GIhzTpzZ5BeM4UW3WQgaKbbYcbOk8vu9OhJLhQpwPGgn
BtQXIP86oeXsAHbForxEDP35T1MVukIYWeQxWbP+UEo9Jcy4PBGggh4fwqvEY6Zrt4czGoutAx6i
XlMJJATY+xHtLSPMe/3xHXWaoFWTlVxOeuy6n6W5BZJA6u2Qe85r0gVhGU1VCk9q6Ua3UzcbmXP7
Zkxb9tfI/him8TLbviR0aTHnCa2sofk+vNMIUx4Dj4ksaPkjJngOdHlo+Z/iN539b0MH+Mpr4uvU
WsUbQaq8xEJLnlBpSx3+4snWkbJfxXPdQD8eeREpj7lHMfmhk/kokDKGBk4CQAUWfSwz67IaXkbE
BIoX8dp2RAh/xDwxAt76hYXk6MR11DlAa40P9nBp1SH9BSh24j4yMz0+67+tiMY3lGf+FSOs438D
ElUHvAE3PQwl9c5OCBcYzvHCpqtMgTEhB5xyNpWSDPQwOxw56HOgV7muOVs0nWoMFwIeQy2pVas8
HssUa8SczY6j+yO84tsanRCi/tNuP6nButIXLJ2EBbiyHtsBjSp86wlg4k0rXsHfli7XDGF51Ab8
zYUHNKiI4WJl6RmWpakDuiBMDNzUJ2QuQF72hqWPnIP7C3U4mmovi0LTDPtxVZrscFKaQtd7Bbxo
J1XPmzsKTJ1g4LXRvacjZrDZLOJ8JbYg27LJoiVrL+4M6V6rDAFbzprdKEtqFkCNm5SxzSTzbM98
NTsrn36MhnBcJSJ4CJ8LQkiC/tJLzw+zV4n38z/krY8EOdkakgJhYzBsz5Q0unPmnjUiyd8XtmL4
dM1KGa0hP3bw/ETNCGwCeCECqp89zq8dlLxF8WagUAcNfRG7Iv4axQ0R5AINtIbPbth8A6w/tegZ
jdBZ2aS/w57WxsKA0l3C+7RSpYe62lJC5u9GE9AWYw4e7UlQI138D7JqCRYKuF3N03h78N5IvM0B
dm42iuvpBy3HKmYKgSINvyxTxkseRCicLQB2hWbAUgdJuqSoScKNXrBTFDOukchHrGpl2h9Khv/J
COApjDFTIKqRl9XUdZU6S42Pdb7Xkqjmtw+RTMHnRkWumvF+2ac7r2c81QMQGJHcQ+eYxr/tLu5N
0mfPlbR9FraSMWe7MvH6CqIS9YZC+bV9tegEas4/kZyhw0edLEpg7nF02h2e8wItRFqM266WfL12
C01PsrykeYuw0FRInoWKYP4JCr3U+yS4qWsgBqRkirOTA9Yx6AakIVQl/F1ZF7u0xz+Sals/TuCy
RIENV6KgRZHqOlJOTGDHq2kwx2agI+CwnwogQf2qj75gggvK9pho0rYjUMTA+gmeFkXboZkr2gOs
cjrxM8R013unBoQ6Za9tscAD0BfpiKy/bQuU05i/PMxTdt/ZxY/GYnox9dNZkEu+PW8tzPAVHSEU
XPOi/3hGrXEDQzepHvivq+4oPrutpH15eMy9yMR6usTMUtw/La77pWkt/xEyKKrCbIVcSdQfHWrS
97ofx20gLaoj5Co5hIef/HvA3FAkTxt7OBmbHJjAaeHNMTR66/D6UW+wUSv4sUVwb20Z3Yz5BaKH
9XtCD1RPVir8Yqc8+LRgwx/McY3/dWYqJGCD2sKBz65/PaTXwoN2TcEl2Cj0o1nOuvO5B+AYF4xl
Y3jSoUx3X4Z0vuk6V38yWRmr6oOq+QKQWY7GLjM0y4Rv42MPhghNPFfnvFW+uvUq1sTr6xbuhuqd
B9FVG/ViqkcRluzJw80tP/v2M0SsOoAmkZyRcvRxwBrDO6ubr4vGdsNEm4QS139jT970Dj6b0B3H
JyjFIjaJ2Kum5snUCt+tZSBkTRbBuend5WlwT7mOJHvptBrv35g481KqAqMK1NQaQI9nIJof4KGs
klrhV6v9cLsUs5GFs7xLJa49HYwsTcf5zxK+iZua1vtvnZR34pOWNRkF4YgH1sEuo1152BePaACi
zY0tXOFn55MCG6eYqgVnx3OHKmYC+7JF5idEIl0PfLs8Zyu90BZkyig4Q0LGrW0F7tjHVu8Seots
D7CVRmj6QojwpE7em7Ys2hS+YTXpkOdFfS22Snd+cRl8Se9SgTtVbipu9JyemoPxaiGuIP3zmXdm
2V/eNSEmyTCTiFWeh78XkD6xzPsqbk7AkaprbPWAGjGO4McYTzQRtLiyI2f20NOsTwexfSeLqLkg
N/zjXL4tYjRUOU/TXpSuSi0ZO+7/WFcTZSU5fiUw0maojM7RgAHeFcxvzIkNMf6b6TFGgS7EZF+A
k1HgTsPP6IVncsxZ1H2ObfxYYd+4nqCuNarIxUqDP37UM3+c5XvTGN2Fjpm36bwW8rfhsLxWWmDx
AF7g8365GFq+cvaYc6u4LcfMwdFgW/jLV9b3iiVO9NT8ue2uCutj21BMscIdHLT0fYXXFO6qOOhM
pls6eubW+dCxcYMOmkKWvRnl8GpyrTvDoHrkji/QkscM9G+JKg7K8B444XAhDMz53kH4ej7dXwpX
mGHGXQJtEu/Vt30eGODxij9grtuWmni5qngrFcBP9IFdlJA5Bc99Q1aiemMS8QnB/FKn23MVrEt/
n1ydFraWYMB9YnlubMExrzome8JQBg3e1Xs/gIZNrIjT62vN41EeermgenO6/eQf7ktqby7yO6jE
UmnIbw5UCqPwEP9Upw85CL/ZuzIhgT234r9CY18U+klnUdzuARjUnPYli0rRgUberfM8YCpZCMB4
9o304QHZWBafpxtewzqQ49WMgpJxQRPD8/jcxH5nbQ31VEiQ2w/1+1goSQ0Ww+nWcQyxUup2H4Ln
DD/mYJ4vvAjAJ5vwk1//NqyRn0hlb9m2SErUui1/HdFSgQ9mb3WC42GJAddTPB9aqJhv2wPFuQgn
CFGRfrOfJ1AVEf3daA9SDvSj9runhmwUQy3aXC+yd46W3ouCkyx4DRc8qDbvfe1RnXD3m5pK3AKd
jdjLaEaBApDWMX5zF4Dx2EaEWdtxqjg868DHcYbQDV3TC+zSDtOVBTbgvLUcV5bT+/TkfRr5j/Mu
dXUh3lLoO2Xb8xSyP9bb/Rw44yXXxpIBeCZrVkHig8yxvowu/3Nehk2zaWhdEtbowBMvbkF8MSKl
JWMiutTDoKvAlfbLvQEwU4/a53hI8kJJMh07GWzmLKjuHP1G5nrTFj1VQKIu7IwVLtAfnsgW0yvw
hbUT/ydLGYNHOpk5Gu3MZKlGjE8i9pI0kxB36QpeBGQrSWUGCsZ7NWOePrfqXbdEh3LsGjkqKbN8
cFPT7aNFk+LGsLq+Gz7UGhTyBpfhyFQpqBu/KwInAcDtnjspBEvWv3T8G4B16Q0NzgzsA8frezFg
/vLbrhaEWlIfyNQdgyime8sUr/Au5ICPeG3Q8rlQ0awrqmNnxve1RzkX4vBlZ7D9NuD0NGemj7xu
Q/6LDzTpNWiIQMLG/woh9nQE5UyGHO/3dcO+MMqxh9R9PHZtm3XEZNgqDlUWMTFbLNSaS5wa6uVh
w+7Cxu6Cn1oSA4mB5Aj1qMPLGvBBaeqojKiv+lCn3chrp/M1XJcP1ijpUtq3igmhMIZ3jRYvyRAZ
xUH95Lcm0xhv0X1CKso8BYXI2okDjPkAgWS8TcTHVdvqHaMssIFiaN4ydv+NI45kdz4BT7b/swLn
7bS9CU6IniEW+4/613q39G8Li1OE5Zb4xokQRKeK/7UiYecqBMgzbl2z2sNqS6Ytd0pXlRxINqrq
xusPWo02dJVZum1/4MgEeqD4W6Jl0RRbAR+3f9KruvmGPqbuLsuAICROI1hrYjF5Zs1OGkLcMz8y
RJl1J9ba7tdtiTAhONe75xqSWXYlELmjOdW/+p9BqaADbjZIixfINUrYEx1BORoL7FTXTtLHy/dY
qG8+284y4TTF5eK4Aip4KHgit6feQw5w41jVYQ/afTkBoC+eCMF3AZ9u5qFAYpl0lyRts8iakX7P
yaFH++CJd8f81iwr518ajsHMnxRNSmIXc7LdSLxLckRC9fz+m17H87vzyKvtvUBwt0ds6XdBY7fL
eToXuz39jXO+osfU5ulwVuFUf7kkORcsd0U/qZzBu5OcJCethkIImnpoFpWAwWR2185YEzijfuWE
SMbYpVTSK9RAKmVMLLGU4pt/Y+hzpb60atzQ/Zuz++nlenN9HVfXMUOf/5JGN9hkkWUbjh3Vqvdh
iDRzhQA1zL9UeNCK2IDD9wgP804JmHI+vEDMB1U+s9UWT2wKr3rbtRY7RFMYO2Pqd/Q0+SH3rvNm
QDd+9yAExkVnDyzoLf2rvr4MBQwWqXVa8JuYC/padwIqdRKlUcthVTYnkV80pALwTfLoNTUEFH/H
N2CL4Eaz1qsNi6fAIskRvyBH19s73RBzD94EkZjdIslpigQ+lOgrUv2JtV6rg3QygnjsKTmiIW0w
fhcP3LDZomaRs+4cPd2Ne2/DBegrzAj2pwsyGnC6pauMW+ZDcIVjLhshplPxYORTK+FzcHoUFFBk
el2ElP5tS3z63eyIdS0zCMiMt2lU3X/dN55kmsSlFqdgPHLFoMJLNjSJFMHWwPX0hL9iVejokDGf
YHNndHQ6ED/tD5aHnzyUpq5Kc9RXU/yEFMErouz0RAfudhx0nFbZM/b/4ti14K9h14qDoaE/ZaRP
Ovyu8KThKDExMOJJ/I+X4cE2984YRP8L7BfHopylxrLivIdUHhTQPHyaZF3weoreOmccs2m7cGXw
6ui9IdO1OhD8CMez2fjGqp7/1ODx1eIrpfjSpAZw0scti5+TET2XXNdcAo8sWH4MKuwaZhochPL/
4LhGglmkhvDJzMphaxFPk+gbtQH1imB/CHXwesHg6t+YUqGSig2/w8ua9MFBSyRvuzNsBbuz/7eF
fb2G5VQPUMJn74XcpRT1N+5J62+ncNQlu2bWDOu4IByWEQlDBk9ChTI4rVsqXtgvsz5T264EaZZy
D4wIpAucb9B/rXi7OSPeSQ1jKpNva4R50Qx6NJEzLG2jvV5+g8lonWKhuiVRYca66Ks/UsBJoqdm
VnAPZsuH9OujpChCNC/ZHC8Y2V0g2jbFYrIk34Zd3SuKayeeghzzAAtPJ37Ll59pM3rEodsm6AM2
0AcFn70eEJ9jaGADDtMP8gFUoGwGm3t9YfXvswx5FelOHcBWzNO89v2R3ZH/wsBLPXaFl4k/mdf5
psVy82ufiAosLUFZmpJ4IHGWNy1IVbvIMayZj/DE2ZFXMLctMF7VBzonu4eklzWVhHR9hIpU3M0Q
iHkGCVNmd7I9zGJtVVGOqryeB4UUZOxQy/ZoZ4SE2s31OyQOZEwhbzv4qZdBAMZRRf+eUXunDXON
Jyl0C5+G4x5vjemes6o3MYsIj1k0S35JqrTpIwLteGIERw+aYhaBUpZe2SDUNhTe0MITtLxHeifW
lBsbZtoqJo8Goy7ybSE37MHKdtlefmn/D422yfTRHKg6dXR6kyg9uPun9h2mQYe+zbL1VGlgHQnz
RX+I2VR5Wctjkztj6bBm27hvLsVljldTF4eepjRbusr4LGY0a6RppAxMYHENBy13NYDzNWNdgdJb
mrxhxqeqAF8RhmoNU85fjk1pxP4Z1b95rzea208l+vewTLaRTglNh4RKUAnj5xPuOEYnXGaijqlG
GtXtnW6B2is0fFVqVH81skI0brtzGFKbp9d1WqRLSIMlOKLw4WIVG1VyzHrsPZenKa3pdlL7J0Yn
qjQqW8MxqhjShf5TKjJaC+19z60lcOk1qs+RQOwS/7EUSjHo4Yv9ZribH615xz4GyPxuYM6PDgG1
2YykK4DmBX0DL7FC5Co/uw626vbn7o0U6ZQEXns5nE5TY9Xn8zNLopdhDLb84fRWwpytJnpbnV8h
fauXdjWQM8oInvWwCJGzKcu+Gz6CTsgpQjd1xGxSkdFNdfVxkCh5EZtT1EE0Mc+ztuS6pnzOeAPK
SM8ME1xKumsHJBD7W94hcrJxp1lUUlgK3s/uMrQffuMIK83+2gTA5t9D8iHqmuyliP6lj+gC0x2l
O0YHf/zpOcYoGlwAy1fT4qdXsNvsnwxeNiGES4M314lk5wPs+SaxO29L66KBaey1TidrIu7aXqyB
eGX8jf0mtgLZ8elgbmSTRrQlo1RrzXoz6KHwLPSrF/6iwhm55jq7E7e+MBlu8c9bgdABrP2JcxkK
uAyY3suF+qO4Euss9HbnR4bCFHQOhvoc5npIAx/cpYiX0sBOskDWS1xt08bY9tYSF/r/lnTByjc9
qK9SJ2WzyrxSI4+htgU/WKYoKpJUGo2PSEXCkZPxGd9l6rptcERR+2nxXrszby1tuqHrIJmO+tPx
lJqD559EdG3kTSe4AI47Tafj/09qvx9SN+hUOoAiY8kArieh4NUX1yFaVHSyF66tNk6oOG8pNkM/
6Nrf6XNY71iUBp4j1ARXIHiFz8H/byRaHZ8HCtavyZiQhLduFVfU/uNdLQ8e4IyVQj+lyfF+n3kB
PWop8i4yxKf01hFRCDZq8x4N5kVp4iZtwcgd+eCaDuZNADvpDVvp9ap9BrrLGM7gLDtYmAW9hwxZ
T4Vh//HbBbSO4v8SPiPf2TAG++rUlveZd7U6XgbtxraIFN7R5Iccss8mTRwwfOFxa0BxYDjVWUcS
IovfgO3b4YAe8XAUTjaHUT7aFLFFFpjE+YzV8QHKvOTzDbg12Hp8Wge6iufcfIA1YzGp4US0a1h5
FAif4VS0hm4dR4gO/zVSWmOIQuYP39rnG6A5a2LiRmW8GgkEOdj6I6x/74nxgCMHE4wpsGbUkSSG
oLCNbxuhpkXCMjAUAb8ls+j5F+ta8ax/XOYVNgRA+cZitScnSGcg+rSMSr0L61YTDdWqT2nSBDpj
IWoZLqGP4S3IzNZngBsF/ssTKW6SO+1U38CPbp3qi0WMJ6pVD3fT9bVYlZ1zV8f0Ax52upqScTTQ
I6Foo0ZPV2D1NuQ4N32tI/Oz/5kCBn4m9oAfdzJ+NKUQLnRVUvrr0PtB3HX0kmo2MVEJ7xaq5+jF
HxNYk5gVoiWemNuqHZZRjKQJ30pdHBLAe6PMKeZxYSZKvcdNeeUTIfVN7We5Km7I8SmouEFu/YQs
IU8tgx0jhKnLX9hCxhKcIxxhzNexU0P0Rm3lTt46JHcHPK4ExH44EIaehM3QS0jgjvj0f8Kwqax2
fDf5XvbJ8NW/Wq4+slu6AIHL/IvionLFBbjVJbFPEY2Nf7UhIeHEG7timLbk5ReyeMHvga5noJdp
38buvDuCNojgmt8Gs1QDbJ9mWQ4s/MXhZn4LP40KJvLAYZbUIbPotiHogKlBuBAZ8gdkq1h80HC5
xlw4dWV+p/9Wv2oCITHEtRcQwNJgQkGPzhLuk1VtiSw6MYtcJTat985o1OrpsxGDPC1F6xwETbit
HMOjH1hhc+qc0hK0yKxu8ekBV7my03PpS4dXTXr9m1Vil3yqM1lOVf+JIUfOOih1leNbZjO7U4di
yJM1bdPX1mmK5LroASCHOmBEJMK5Fza0QpITl++FPNMMCG4bt7+EiSvV7KK+Q1ZcXrfxQgYJ5twj
hLqSGltNzeLcTM3d8424TRvFh3g24qIEB2FHFZyUOm/kM05LV0mf5VARGFKWu2ee92pnQ5G/AlFY
VLi5/M/+XMHsxpf3JGbfMsEGeBH1wju5RvMXamqn4fHqD7HxBJEAyzZ1I92hPvqJGdOvYapdwq74
lk32f78sQLhbltD6XcS6OshM3MVtRues3SY4uw/7f6a3xI0TWG8z2fm6ja2nTMlLybfYH0xupfYA
AnOa7FTrWbSqOPB6cs8katjrpV7qHhjL/zp/7jD9MHrHRkVUDp0DCbhCY0h8HFjP7GBlOaD7JCCi
KmaY/jd3MWPGSRvYXxQoMnrlvzuXUvpSq/+NuVluqRY95zm4zKsNWZZxDC05l/o+7EMwTuvAsMG9
UNw5bQ2xWLAo8kgn1iAcm1bMqemh+4LB3Bf4cmIilHCh06X4P1Ifnm7Pt3jH7ymAL/65x0zzU/TA
JC4j/EFN4IjhX2xhO+A/xPFl3uuJuDJ9EkOCaxG3q8mPrrf/gkudnCOTlUPcJGu48hNQhYxSAzQb
NuvysCJ1YUdfM0Q6/LxVN7fxIvX4h6IMfyzV6IdFgOqkZXYab+7XKHYVEl3apm7O77Pwq3gNMy4D
EpC+FCuqBhfr6p4qeEy6YHNalWOCjyxwpWsNJMZlsP0YwdQHZTPYJ1aWwGML+SuUoTdBu5FzJcp0
Tm6i4aA7fgiUQWmZTgJlD/dMMhU45nCvgHzJrwO2dkp516QCOcAYAyQSxHBfz4p7qzl0iVZWLPnK
ZncWZoIMUC7sdrM8Ne4pqUvlBIZ04Y+O317VYPCL7y7EmROtraLYu2FgiHEsddGGuDR6XVVIujF+
ZdjQ3sV+uRdZBm+b+8efBUWUr0AKJQsKcjKxJVOaEbguVss9TPtXHsjp88qgUv94ay0QzKkcoIZq
qlH+YrFXQcKE/Htb1p/Q+SBl3ci1CV9lnufJVZYTkUbL8YOJx2SxHGJEh7zy5kuyXlvE8TrrDmaz
L/+ubvFhNIutyT4Tu09Otk1vu0gDkfgwAw5vaN3KeDNlovmfTvYqUO4DRS0lEuQS28oFLgjiLR66
t74aNPTSG8FANerhJo00zlSMlHqE0Cj6AK6TVJnOGXzxHFKJFwLN2jBFmfftQLEzobQT1ocS52/V
NsWHrcHEvG8KfnwrDrT/voAqTPRjo569Zjch2Ow+1vG588KcVfpGNOCMJXY5giTJS5V58pIah7Ky
XABKyClISlwm7fOiuFqnImakV/GH4/B/6oBc21KJvsOxqq6cOyFublJwZ1QjviXC7rEgKmr+RjUA
C2zzWw1RNw4L5RVf93+Bj+dXM+FhNNC57QuFmmcfsX94lRe2ad/F6ILmDS2BNyip++Td+7Os5b4I
MnjoqAC6T+YNP+ukWOqitfl9EDPvYslULSbLrOEEyyb4Vrtg9VPlYpXmNY1OPN+7Y+nxTgD1/82L
lTqWLb5Tc6lY06QFvWqsCNjzKjnG/hVh0gFwtFXAYP0hLmqLITA1jU2NQVTKdWzDPeiGJt/ekcJc
gYHGwfztwWzk01+w1ZARV0+xuv25g60UVghf+a/E2ax62qO6opMLd73q/auco/96I3l1w/nOgblk
VsgljnRnUObgpN+x0bwhVPh4wK4a//WKYvnhNHFe6kkUw8dQ/0b8IGJ5JC0QHEdhQphk5FicU4LU
L/Ucm6fWe9TR+Cu5vRaCErJDofuQQhYdyiGJlAVZrrd2/CkZkg+jyiGbq5DeczlNm6/oku+7upi5
GWV65ivPq1OTptJkc0t9TJbSYO4LUwrgL32q0o3+lZaPR3LwSIlmlQ8f4IDKyzuSVYDCj1ErEG6Q
lt4dv3njJtFxQrc/b/jvq00tjHyHurRG1wDQcDAeDZeOJXacYj2d5IgcEDXjpsQrH//UejG8Ojvs
SR3wMuNcr3LDGsPBCUoutmO+tgGKR6oVNW49SyEHKmXs5CjTC8YDWutKAQkUMbUpkrwpOF6N8+B+
rp+j34sUJtDogDu49BQmfSVhWanvVXHy9XrmiTlY/opm7ylSVqGB+/KCkL4ykq9abyIYKgRTKmyd
C/9FwXLrFQ0dSNhxNlKViFu+lf8c8x0snO9RESRxkquDVipBY4bZ48+OcUXWPJcUl81z1fGAEUkm
vphvDOhE9oS5iLs1GEDeWJnSpZAgWVR7QxkDzw5/5XBIpZ4OWcb3JuogGz0rh6OsobO6jFNViZSe
vOJ/j4Oyx1OMZaWCrF016AH6r83tu62FyCiz7y4/N4W0R1RCELMJYsB5SLk6iVJzy25LKbF+sry9
HjV57q0u9BvK3eC9msPYQQdU9hwaAQ293dYhI7Y9lpeBpNwDnOOHN37y6Njc+753kEbOdyMng43v
5OzqvRj6Fa77fQ0tAzlWBjfZ5I+lRcCVyMmh2iYIoH99jC62ZbeK3eSMKQupvJxvmxzAOCPhItSH
3lix25MTsaXCXEwNVMLiY4/dGjIqv1mDU42tizhFP0HA/PHmpfjR699dogKdv+4eYPWyYEz8yUzM
kCw632+YR5mdlWsJrrRHHZKmMl9nikHko2BmOHjCUIiH8YUBBxxhyvaYtiwGwenl8R/NHc1K9Bze
9kepFEMHtnYQwsqEgRqOqMrVF6p8egCTgWHk3L6GQTgmH0FQ24Ulk9+8j4w9t9V5p5pizirN9dhc
Ybg1OwqHV5S4JBvsgrDchlTo+pCrGURO28EdeyK4eSc456uGqrsnlHojOnuJA8xO7RtTFVA3xEqn
RYkWXy37g6Ar3c+84v119y1JDfxsA51si2VNuhzAfYy0qEtxghX2f85nqnVu2SJ/nmAt6cVYF/RA
moZiyPd/sb7yYI3o43XPS6aGom20R5Kwhn9Kb+U8zkWPIRO+Hkgjq28aJ/KhhsT7+Z3Rx3p9mqyX
K+s1aETS5x3NQG5ulj/Sd8H2RScP+6Z7nzwXXmcFLNsUPtQkeg71fjovL7LnoqK7kP6YiSJwoYmC
oPvjx1Ot+fHcrCf7eT4/F5SBJDceRUK/3MYqetiPpCiRLTCCUeNgI8eUmuE897/nOyPdI5vE20VZ
K0MhHFYiBmuza8OBfovqLF1e6id+1YGTgOeDbmsPrPtOTDcf+5LVmJpVH4bG90iE59/MniixgNhB
vrn00+iC4dQQYDfbPSJMe8qHW3g+UzpeyaWDiDojsQW/6I4DVxMhioGEdGdYtWYaIbYgyePNKYV/
hdZGKE/d1kJoAY1csuzJ37nBtmuVr77Upi5lfnAowMK878Kh+y2jafZ7BrQXtQN4jkBarpA20Ir+
ZTx2J6ajiC23K0yhwnt7rzdr5Bnz0QCWXV9JVXSoMoOJ7Mrot1WBhmF4wRBNFMkaeFtNJoe3oNKH
iL/6tJ1IVPotQSKtSWsUDgARZSr3G4CJvAL4hsLthYOgh7CTCxzXHzwiQUuZccDepR6qnDBooTzG
+Iaz+zkn6utTCHOnrCsAz6DIMb3iFc+ihPYCFR9dS72jFulWJ0Mb4PdfoCJvxaNmyv+ej80FtuJV
O9wM5Orb6XqalXfOv4n3DmaxV2BVNbDw3AmxVzEA1kG5KQXdBcoygwY2Es8EHfrQ/x3R0nmEPHq7
E/L7L1o6ndPdOj1/3Rg6xtccBgRde4SZnUrRcS0gDQM6WSJRCJ+4O7aS8PTk2eyOmTF5iTe1LoMP
M1Xc/OGk5wkJWxnpKJ4BjwFQ9439NAarOGLC2FBMXdkUa4skjG9iCNMKXV/SGNkC5IGAFUr+9xWi
63d5hzdMHNf2VMPbq0H7vCOAdV8QiMgrg9sZyI5QPaxqI0qPhQbWusv6od6ZRFiBp05yYmK7YO4J
3jUwz+sunxCO96jXbf9wfXzUOluFHaMUpgB/qVRGJjx+utY2vYepH3qtaTtoI0imgJNNPx+IHEqe
hCgsBeBDkLsTuPF3fgLhl1s44LftYxzQjTSCBMyNa3WYEGhc0Ot9RjJCdTFM1GKr6DU9VunncMXC
SFtL+fKeYpxAvpyw6Bmy6Wl2PQSSRVjGESZGE+EYZFMvqCH8x6kTeNTV0FxjEZ6nX5RlkRdNuYfG
6L3VuomsYRzNZvmy5xMLpIg4YaZI1spoldwtRjqP0IzEVkqX1er8DDCv7etz12jjwMd6tC40PysD
s0w89XG8CMo1vcFcF9sGacGRs32DclX/ds4EsLAoepA9YExzL76nVhbiVGOl3sPn6tRtKhg6gM+Y
QuD26SuKsNcfJzUSk+VnZngLZIkzvLQsg2D7zlcZfD5qcEyUZ57VU3YjPXOTHKJHwthvegQphWQa
0jDwmahPYh3u984NcuSn0nEuxUIrI2zcFbZpCrVq1gHvhpwA0Ew/DDizUf7vWVfs70hp1PBgKltK
riuayNXlelkw9Q5tioTdAMHE7LZ55ZaBMzVnDwuXY+WLnbUoblQYeag2pSqNOzWeHL3CVrYMzvE6
K9Oos8ivZvbDxn7vfN8X69eqtw7slLpyDp9bebmSX6Sfwsk2kXAP6NuEk2mEeOb1OcmhTdYej+Ip
5CQ1brMVBKZmHMXwlR55IdmB647Ihy3+zRens/0dLgil1VoYrNRyagGFv8IepHcFlJ5g7x5v1DJ8
HDXNmWNCVarKkcGOed+JCwEKpd1ARWG+Wh32+OPYuxAQJ76vupfmenFS6BQk98yiE+KZokSDBZqv
tMywyC2VRX5pjtzcmUi/G1Fb1Uu/00OLsDCaFXVnVUSSR5E7Di5mQ4ih7n4NvmsGp5+VFkYKfvuD
7EWqAuVjT0/0G0gu7or88EqjcZqus9eorempBVrYm05Ab1cDqyAkAdzznt/v+FV5QhmZecEoCiSV
V2Imf/iz8nCneJIdkrtjiV85dSFH/RLeGtbFZ8aRuvQRAikxqmwDmiOnWfvHNbfbjg0HHR2a/5MQ
jdvGhsDqZizj+eEcvFRBQg==
`protect end_protected
