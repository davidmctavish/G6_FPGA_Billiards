`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AsrkS0Oo1H5S4ca0WhL4sTCo6Iv+T77FY/zlahr3vQbJgNLmLx51eRjFxoSkT44D737wvzoEStsR
yTRz+NHXlQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nEowrhM/X6423w6lmghX3tdt/hTLBQ3oIcQsCh7KSyPZ4IlZTVBNpv58SgAeLWAZkTIalAevTk78
Dtwt//AUYgJtD1CvoX2hh0tX2734LvpfsaR4hT5rAsyZ31L16MTE6Qg/dImZH922qdkKXc5MKZIP
VhV5ZGFAhN1L+DqJeVY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JX4dppZdQz5EDzEUdUpLYu4Vqk9DKRlA1YNF5uf+In9tkmRJcmobaKCQYsnAvCJaZmZMyAjJ+Gxw
9c3IOlGKOIFFg+mn3ZaTxV+JVfjy9ktq/d+39Fvc+4oTcNjBI2zFZ1iMTSnhdTL/kIaJmNOdsmFL
bV9Fg5q3VSRzzOTh4g/A1y4l8gfudyvdTFz1pULQ+oZtDajTp0nnEz9Ql5/uD86iIDYYvXpgYoDC
xzlG2hEzxIoGmyN6SYaq6sORn1nyUZNIro1cyP4ZHWrvDhAad7YqPYmHv2dbPxcgc5q24C4pyPOC
kF9f471dwtOS4OcdylOiukQcyxnsF67lfGDVLw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IopJx2bszK61eMePaOlsdG42WSEfLtFDrJV0ZWPVn16UaqAb45ocxeZu23MeVv7bHbKgj+EPT2D2
ViH8PS26rlLSwHEV1nyaCRLO4Si7DPGZD2XJfWINmWboLiAnvL+uV1K1k5WN/aMRwAJzNfr+i7VE
ULwej0zaL6Jlw4xC4gQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ORnUBoE9MEOeZ26I89s5ve29AZF/JAAupa7d6Q3ppaE+7HbMvaXGv4BV+mo6eDEByDhUKnrEmU2k
1HQ0uH1U95azzaM6KnEzxB/c/L8YfYSfs8Elyj5hy9K7JC/OqG5KpLy87AT6cH+PeCxxVwJMLNmd
9hJNaKOCXIELhV4E86ykfgLgsDPlh4tKDZEAdR+y/jX4OCFXESrk/tkYadxden315uj493BeXCLG
TSiyy1rsQGI7AkD2cxlE/ooinResaIJ0OoKYTAPwcAExEaRp7W2mOOMyOhr+IuCohIdEIpCQ9sp1
pkdT/juW7XQQoZ1g74VYD0g75A9wkUminK5cuA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18288)
`protect data_block
aS6qHccrZu8NMj0K6xicXHcfoKAIxQi8EH4cyRKm0ZO/1Zglt3Qeg5KimK7njmNA5yxpDn0A7AGr
RlfXo0E1kXAMpi3Iqk8763YHHx+6Rey6Sc1nD663KFrhEQk6yT9ctzk9DAvNyEM2o07Hht7nAX18
+9/47ibbLbnfkaA6sdR9K6MEXuP1lbx2IdgW+lzwAUFIQw4HsfHt4VXOd4O5xqMtJbDT6SYppDvJ
66N7OfW0hMF5UGmw6fCSwH94VySoFlQCmP0jDv054EH+GJ5p9p+7VBBo9LrGE3/KjqqzIYkd8oL1
lpSPLq5PqHXBTe8yPGYck4KetXIDhNAqQuV2nc4mLv88t4CEmy0PiR3yeDrnb9xAvK2E5AV6E+Br
vb91JquM479pSD8MHmIP522AyL5S9h4IZ5gvDkaa7YUZNL231MJTaLtUY3rPaj907eiN6JfKOMkc
5xE+4aG2XjuQbQSVmCLMCXSg9zQVdZa1SCVt2wl4Dtbkq3hHZ/3Lzgl8gvfAHx+OYjpsxoJICWCF
Nm5H0jT6VlT7wKwK5qvlR2lxDV1JbxqQVyINVN8+1khWq5mw7SQNrxuQwaS/8yP7lc/XbRCfiXVQ
efUY5eKTg2PJj8cWYx8ED193uM/7fWv8+kQDAIhfaYDQC809QvugqYDddlh1UcTB1NJp74WPsEC2
J2ACp3bVgxBDPBxJ34n8xMxUwfuCwv959mBlaXEhQG9QTP0ZjtnRZmiSSB+wIjd2x7iHInweC/QR
t2y/ibewEo/rQC9cIdPXFwo6W/N94RzRJN6GRyqPu+mE/XAu71YIXZzW1C1SwXv9uo2QmVzxwwRu
tuT0x7gwybKkPern2mm+qe6kHEfJST615IVJdoAd9pqdi/VN01rTH5SkRdHDnuv8/G6QNCQD2TKw
3Mt6CuQTWe7o1qgFzGjsnPrchyjPdvqn0MCPkjv9N0H48ViokEqefkbcChQZdVnq+oGnPE6+JzhR
VLZMEKLaMl9LiaRC5h2K2DLsED/6F0u+ROtmSf/ksgsGujxaNKk1btsorCDg9DJ7i2vsbo27Aaln
phkM8GS0WUGlpDcoE/JQFHiIJ2UGfoiGrGDzV3oun77QApK928bJqzsmoTCLiu0fJbJ8JyLUsd8M
1pyv0XQjoAJ9YpqxiEwOIufrRIKf0yX0xUAmiMveGw2Hf1o3PGHn39q8+C9SxWPAtUgeUotvmJPa
vbryKJHhW2+5KADQ+Ng3/hOCFAY8v00iBXRdS/5mQ/fNqhZvkXl7c8NLK83Lph0ghGT/dPGmeqrC
yP3mdb3EnEN8O+H3HBzbf58W0t6e8GSBnkQ8/HgrRIZnBQ+AV1/M39xKbsq470Q9GEr9CQHL6zl/
CbgMbLOuvzY0qA++A+niQhdtZWJ9RbNY0gyupeh/MkjU4cTm5Wez2DD7smzoX6M7Vynmg115C5l5
Oa7QyiPjOtH9OJBaEt3nh3t6PwDYOukBtWYYqzaZElp43scRaaNsc0BVese/rn221Zhl9RtWVtju
pc0YNjP61VT9K8mp0BtQwRS7mOGAR6uQixNkWYRxH/i0s0Yf0ipcn2CwQnkHEXMbGikXBGiUFYnS
VQzMv+h+zVJVcReRQfRcLfScBhVSPf3V2GcbC/Omh8T4UzYxppJOm7z/eYr6YUwm5ik5Xvg73Nl2
Ehqac58DoLkCgMOm0EqVNgJktMr4B1A5DYT0ie7wfUXon2duBQrj0WOqEb6TMfmWbwkJcD/5I06I
d3zYtejcLmf6D6MDbMu1+oMu64RRmOGhJHYpHyrtiIcTTnHHhS4QDjULm8UVgWE0iC+OjfQdULHB
F6a57cG8/mwwTlXnj7ZKob70Voe/gB2tz641cQfabHsipXyEWJkPcYD1F1foo7LAeBcYpA340YRB
LwR/LYz1E3p48ZHJrTVqLSjacPU/BYsv7xAuD/2Cr9Q811pe5wNEDb+nn51ubB91WpGJuU6K2tj3
E90MVfzfwrHTSUg/5dS/En2YjapHZnATVHJ6i5oiTz/WuMiwWMN6TYb+MCDHD+g3jXyHPYSO6s41
3nB5medT9Py3tWudUGDl+YzWsRp3IO/kl1fNBxzHpbqKoEymoYDZKyb5cLNUT4IePpduPpsWE3vT
x1Si/QoLnkWv83u3pmwqrnhD+QStNEY7b4n1ILV3c/0pXpM7UOc8D+bMcZO69ygYL88VmbyNYSXf
4m7fwLHq0a4z8+53KDH6L584JFnBqh3P9P90K+hMwLbiw2jJbbQrqf7aKAWntO3TBIkAmcA3dSlU
DGgUMCLIh8arwpZmVXCELRR0ks5I9d/3gGvg63g+V/1SjYp6zrPD7g3DJ0pltHwlp0NCroXDLIMG
euSEgoejAQ8wa9LtBAnPQIIBiQQfVJGxc+Wg/ddCJNi0e8cZyU/73JTiSA/B3UJ5NGAfXBakZ0Uh
mtPMTOlXYsW4hXe4ARO45id9UteTu2vx8YsZiu53eCFgCTASC1rb1FyJtqbP8ELFgBj3BiklT00d
q4uqQ+Gbn6cpRbPqq6vR/wOA6yMNpCqdGsZ+zJdk63tWLwvMxVqZ41JaJuq85ui+iVr3trBiwQcz
NbJBJc7PMF1Bwe2HvLoMleb3A43GSPTwKoIy4M1eVho3Zbt7yIe+ZxjPuIAiLvBFngND+otW0HM9
6G7wooR93B+0lHQgX1lKHDwkdS0o4QoRyO7bmIMhzYWtLtFPl6bXV6c6yWblHDjU9F2XEyfS7jtU
pYTeMZoWKKkhsk0jtSG08VboNmA2oFwSOQW00QjQidLD1aRoZ2Sq6NoVFi9rGapvgl/TEA5SetFN
lNIJbnQwBXkIbo+XmJlMG2IY724+UW7W+0xJXV5MY9oyOZQQp1pZCF7kl4IMbZTgFtA69VraGCGq
Mt9J3W7yY3S7H8U1ELiEXqYYGnhYzJzpUgs9zFfKhNZ3D/FPKiOO5sdqStEgxpatjaodS/musApm
bq+xds9RYOYhTnztaF50lySy1yrE1+i9aLsqx3ypf4UX/Wv1mDVbtPue4ZHGb1dh+FzrLJMKNbFg
jv2OtKjwMyGb9MsYmyoJ0GFZS6Cm554PnZZ/JnuXW9TERnALoqM6PJ5DMB8ZDp/Zsfbe51MQ+fQs
wr0t3+u6GAu4GhBwBBpsUGhOs/ZIJ6aIofls6brE0SEAS2Hf281OnIty0549kDBTcH9kzvOi3oc+
0pTJdqdDvLL8usuhHEtWFO9rhDu2O/CBbUDD0Fk+An139Ql0ffX2Cjt688g9MRMNeSnN1qJrs7WF
uAX0v4MIhJrzNiMd7fH+uqJqEPOlzp6M0ZdYM4bAHflq3WkJTlEceHfpAQ4FEvIWFJ6HDs6VfcyT
SGj01kuEh2l7VxDgZWXlhMWP/7HKioDDqr2C/2bB2kKt8ri3Hg3TTnElKpi1vQGGENxzjn8ZG4Ad
Kn9ks3ElKRsbIFNOrRbXEy6A1ZRnzaeiS1m7uUYhgIjYcnPgeJ87sqSWiqSNuTT4CU+7gi3nqZ4L
7y1n4yhXhj2Ci943YXhuPN8jn2xItcf7zAfHTzB9zl5bNSh1aIK1f1z/FxkiuYPDcgmNeRsSP3Xy
IiRsO9t8ikaRZCHTno4CZdiue9EAmXBtsl65wFugmNtn6ISl4em3WfVWTE8npKzMp36dsADAm9i/
E8xKNrLN9xgQa68S040dD2tHtI/uTGh7F03MkG4Zi2hGhOqxMI28dDPx/eWRzSWGpljrzQp3skmk
A9Dhh/P7allMVbxaUe4UbwFwa/LGUaT8rQCdjXNELfEeKenL477Oh/MkmzJWm0t3nOPDzkhjuoh9
UVxKSPAW6rzgu0OUuuKKqXnq7S1i0wR8zos4nThlopmIaRWEIQbvp0hlkjVaUMsCskHer+AHFEtY
a9vqU+CvyEC5+TTkvvi6bsMSWMeH8qTaLIjIVLJYlzg94UVoyzpViit7IX5Da349otx+IJYPxb/P
dxqo7Laa2beIxxphqLvIRZrwuXKyB68mLe73NIhe+MWwUKcYxWO3Z3Ojmv4BFbFfpsno/TSuz7bT
XmyYvkq1Nh77wLAnX7H38ySgOEZegpevzv+ZB2f7eC+MYLibcQ4v6O+/xFfbR3x2JYIhahd7oCZK
kyXrNBwDIeaDejaxFrKFU2uIse978q0yEHQkqUkwfbN5A9SfH5UWJkdUJwvburGMuHPRllKTt6Ph
GrM9/W1J+Hxl6JF6r5eODiVFSIDtUkpvf9pK6N+xMdErlHAbrwvB60w9YpzNGjv0KTZljjvjS3/s
2bZrm0L7IozxWJg0lxbYXIbszO4/LMGjh4kWvLO07cn6lN+B3SHMdJ5lANxdG2jmKlNbRwXPJP6n
tlPrx/b8IF1Tg83OHDHpyy2rNFAXuSZCL2ucADUvcjc5yeXiV2WVr5masEHTk7IHZCjbKQ33ZOtS
JX93xDk6BiLoQbcpBRnAJdYDWCa0guWLWe+9ZUKHE85oWd5oIl0l0Brngzgvh+D7R3gGcmyWEhI/
86WE2Uh+NliujUW/d2oJpCeCf9WlLqtaP4wv5+b5O9nhbx4mj3m8g3xPctSca9BGcuHFjMDA4ZSI
yjq9+qPXVFymz1vET2VmNtcW+nZNkDrN/Y2XJme3aGqURmCnsclDh2wcvIWTdBwmKEWcF5mIDMij
glhknXIn6JGQ6kBmA7dGLgu6u77RdnhLgW41gO6USIkl3IbEYvRHflft7oW6EkDzzESSAXESNn1Q
S9nJKww16Q1Sg2e/FdrPgR3ov7TCeWfsoEVSmQttL1IRWpOQOtWQD/Kk9l5ZeUDJKoP3U+fgJTQR
VXq2kGixMmXsrlwhS3ipQXO2XfG3mhdrp9X1Q5EmEy71TMlVv22ZLFr5i+JVw+TVSFeNYNnBVqWa
rpLS2jkvreOXtz6X6tDKIGbYM1leEfL9mIXiQn8hlX8nE9thUldWk9zHW99eGdhfPAj4ump0Q68l
0SuVanbvwXRb+qjxD0hRuxs82APVxkMXIp1ol/Jxhu8oDy/sRhYlL9Yb5DPmz/nPgS5lA6HZ3zj6
A9/9Vc8IMihIGCoIan2Qb+a/wK7ZXTOtFD1QmV63qj9uCsYEvLV+QDS4AhJ0cO6I0rNI9zTbAAc8
PIgDiAqI1vlUuRLUg6WvDHqjrADt6tgjMyeESBmtcjz4W+Y6TFLOlsI73Alcj+j6MhwRXwIFMKfI
67YokPFfWt26NB/xUkhQld4TUnt1f6DpVKkyUFlk/LQxLW4i/acAzB0C5USDKnyLEyliATH/JeFd
8dF3aRBVLRKj7sZibVkDPgKsgw8IqoAynpaWY4Rp64ipInKBKMovoWcG3BZ8PRQrpovxYvLjKBLY
74nUPi9JZ7B9Oda//+mya7x9qOuJ8roFuKcIyKf3mLblVZvJqX8lBk+njhMd4JseR/QHGnHtSvyH
tZNrvj7tMaFNNFvWVpyQVWRzzh9hnxDeKUuRMiogz8bGZzMgE2wIyS3848vzyS6aNQiRQJqcb2iV
Xm95AcJQyQS45lCJOz+HQFtzYZkO4lDGiMkpTQ0FqpInqORTpp7KV4SpIPAUOWghLDsRBSS21tqi
+6QGkrX6vgA6Y3FDGA9X8OSqhP2CYyboPJb5p1VbBGKkQ1UGgGrk9Wki1UA+Ra1Pm9Z+ovdE8ZhN
cOsedcHNXplhkLaoGt6Uk90w4j0bzpwd0VlGarkPr0Zk0YQqM/GYjWHuzPwBL8k3AggbJQXUvqfK
vNwAi2L5bDhwYUJiz1D8+sZ4XJaaz626BAQbiO5Le3Tc23pK3OS86+MXJCvdIGdrN2fc2x31523g
sOalcdAM6ErYvu4ZYcmLJvau10mvBHV8T4TFfzJrfSUIkyqxnpdqqOzXFRjbQuPOrY2PG+2Ws4Ll
jbiA8BOO+pHR9irToxP7fIQGZ3aaLBTX9IslJazoIp8C8jafBfrlln/xQANRpoFff00JQE/Y+ztM
KE7N+M9YTW9xtuA+4fRDg1cbWHkICx1Hj5f9sRScq8yYSRlEa4IOQECj5Cdd5P+ePDvEkvfNptqw
u7OmLoXkUt2CZFAMGFdBTd/c4djzGxRK0Bzc0JPnkt+YR+EyD/XQB6dcmPAMltfdlBZt35YFA/nl
GAjw5TCq1mInPCmN4DC/ULfvWcvmlZWCLR94jFTsBMJT0yOvhlzlTnRogXvZ69g7Vu8H4S/trldb
b53K56hYPfsZZfhqicSGVFHwaQem6O/B5ZAFjSTTjBotKQlmKMQ3DGTNWtgbYmfY/nj8OjLo50to
RM/0qAryhoLGGPRTzIbb/8/uJPOBYKuvQpnmWKpEumDgMWMoQ6vcFuD9rYrO3xkmLZr+QJSXEA2G
2YjxoGU4gnjlyWsqdChJ5pwzLgmIZtTNJyg5OP7JiTNseAckZCU3tX6iBSTln0XSg/Ug+I3qDqCx
OoJVgVGZe5DRpO+tkbVeVSrV3nmAKwtOcG1jZm9WgUdyb8eCmq1AvB9eTfS4/pugMEEH7xBDmMN0
HjT5prsVoODzOeYH5TBRlj2JIbGvOntuzhtrFPSq9wJ8e+bTKQItuy9E6M77e2FsNh115jqTxGdN
kVqtqxXqPFByy1UPEs8f7t5PqPX7jDNYjvXudPgIzLhbbFxUHfUFZtWYbSc6rG0t65ks+kp47gPb
h09xG7JahAkyeSJL7BGI633bmPKyQF/9B0f5SNvQUFWk9JUa75guetHSlhQTBpXcGVrvNAt7/33c
pIqY7ktkgZgj13wU6sWD9Xa4rdBZaLMCoop2wtDy1JnxB0VqIVhUtbkt/2IbkX+bVuxdh6paVWmJ
ODmViym7g8//1duRFquBBPFOI3Xr0Xsy9zwm52R8xccHlvaLULfHZWBvgqoVujgMhP7mmJsAG4AP
eljwqaznDRTtYj5tJBC0ju9q2SdhV2rILb3gG4ZTu7aRyl9e+glhOOUjKxEvlO3VEWKpn+Eperxz
jcRx6WjnJcQcyqwITymZ+aH0quyu9Nk5uOpGj4aKp2ZqbRO1fcBMEliRfqdY4XTcaAHWVxdlpOa3
HAhd6yOZk0GqViE79G1QwpbowhtYt1bW0+rXHUCIjprzKQjN+54wHAbggrXwvdviQhbWOnNx7odt
V9HqiHgBMEpWws6Hd55gotgWGtur4G74aEnNridSjCFL0yVTwzq7lbeKcNOqNP4tkfgVxPDpq9gl
ZJcoDcyWtTIBWwXLPAG5TmXyEdLszbTMTE7HdAhiphDnfZ6FRw+DQARzgS/YGP/+3To8pnvF8GJU
khAPSPioFBNfEKXjMNZ9dKJdmCaBwRazFUYsvwJU3vWZrSb+6bLlUMZjujFU8/Y+eMKAEheZjdk4
jkTy/46QFokq6oDWed8Hd49B3zNJQrFJxYz9xglKxUPv9lnVgXoHH4/ZHLNdoKbgD9Kxnaj3dOze
03PvqMoIEkzOjzeFsYKeJhIXa/7fGBWRrvaV9eS8oMeUOq62co28qJeMzrwCU3J/QPLL92ZFBijk
ubmGG6YweuYBu/NeAVAPqGh6pOAkd1CbJ4+ClqeDcrTKfXDctN1whqNQVlTxgYGDyjjseUR7hVTE
vTQMywIp5O3zq5R6q+ucEr6UTbHy9474uNp2eIZxUGWxC9M7HUgpxsEOiLik/Haf699YgvstOiCU
MGbVOhp+7uC+n8F6DPd+eonTON6yP+AGY9PhfxLwRdpOeaTC3PFcu5Sd940stihWhnsvYVfxP3rY
zivfmqLOJzx8sHYOeW8FGsgnaTweq64yH+7nCMuJUUh81DPVJkDMozpdaLHyZr/VeuOHr6lF2TeB
hUjz5yDUMP9uF8J8StJqOaY7PHUwKDXASpT+SwqDOMj1a86jy/p6Ce2AKcsttEOJAj3Zocp2KnAn
XHtE1N5mz4byfYMI84l4bHPto+2ClUiBt9Ooc6PkItThpQBaICuB355HzCxvchtVgQKAzuNsFI1m
oqBMtc9egIfF2UUKJyAPhQkG0SeYDA4PVrcv09E0iZYpSMgc90+wJngrEL0tadxQL7wMUd5zuLGF
ZWPW5oy6fv932EqVA5WkH/aFxara0UugnkTKvkFfttIxeC0Aooukx6DyXoJx48jqyAmMng/V4384
ECp9Rb8xSvHhZRNieFB97QTmDWAVrGlxwoW1ziZtKTBQ2sBTMMU6mibRlS1pZPxqS1Mew0ubixtx
FC7Qq+9deAMv9bso2GZtuwYLpTMWMum6R0KlEKfg8t0oGxfH+6KUxcfcurcPDoJz2eTjLlEARgc1
g4MktpNZ3FqYNHTxbxqF6Cf0gaZiiQtjslSyHOiv5OTj6jBJXbi3ypCZIpCtmYpT0CPaFyziB8YO
U+euzGiJeeeBPOOa0Ly8YAn9C/6pJogM3xIvRagh706apCt5VBx7BfwY31qutUFY1NbFjV90DrD8
MjawIG8xuueqFB+Umu+XEGDuCQVQqy5JDl1YuXIglnCL9tt2BvF40cg/45JpiIfm08n+4+kxdZ3T
KW0ZN6ygQesCxJ274v44+TLzQLWvk/vQI+U+R10CdAm7YhObnIeyTKWv57W4X5YdYUyNf6AC2cve
BdMsyw7l5YrdMurLUrYVnX8FwlR0bYiR4PoGpxdlhDTsYmb1/YcSs8nK30X0XCbkFK/XayfLRR+6
w8/88gpxKs2lhvGGosYqU2aIfMNRV3w1D0pnZ08JIixQdYMxoEr/gaHJtrDm3EKf2Fc2kwic/btT
MkayUW7zlvX5Uy6Cu+jp2x5eLVOAQ8frLaJsl3CdaCDXj7ZI/8LVMVv8ePSCHSYYJnnjDfQ4pZyt
jtbraTC0TXvbu/hPBPEM0hiPBQwlfM27M7ctsDZhSz5sxb3H2xppHhtjyYa8rRP2UvL/dmZ9vFGp
gsL//8Wcdrn2kIZ1WwTiyynYaR/BOKcRte4QxChXGcT+hJ0BKbBVYkO7/6Vmt/9bPDPPXHF58ryn
SF/0H9TRTBwQuyOljJUjFlJcnP31whNHYMRfzZO9KBm0ZVCGFcIPMXqaQ+EPcVh7qPr/t5BdkeTl
vJVlGEKNIhDEmc+QUL7I3cPkzntI+oIswdTaFUU+TWhtqzDpbMYG6DJvAU/GV0Rrn7SnKIs2jOLT
sqJ+FfR47zjO6Q2sPWu8BAMJK5VUOkTGvTW0TzX6GiKawVhpaLRkD5RhmTbH3SRVBEArvJsmTGfk
VTW/H3P1JkyJ38eYoG9syCbPRxN0NFpx4g9QSsw5+UXYXYxOrGL7cGUvU7uNT3l2ArKlEKuFQNJ5
VbvzNzdflEP6bAc62vWNAGNghTmV1YHdHjxrS/f5xk0pKCe//cJbMHK1XlnVxbj/X6CB8a7Ku/He
xvuiohJ3qM1nnBz9HVQAVuwfx6JKpZ/vGOXlRDpIF3P2JYb6bXxJuw4y2EW/JcMuG878/Cp+uBSN
GvGYyBZgro+rtZLDTn30CFP2kp7+duoFw+PunnFKHUQqWH5XODJcBu0ZpacZ2i++RytKSWjhu2oy
fjPTo00ctO4LiPnhXdwK+g/G525hfc4ou4XlmyHdNesHjkgqfHQYMvwCqXNFrmEFTIMlRQnvb2Vt
9Tu29hb85l+j6Eehy2pwRyprJnkEAiA1Cm8m6Z85JlGJkoRBmsdsdeUqdJDVvUHKOoNJlktEuhpP
7Zs7UGcDTetS06/stBRENF5RM/q7F6TBm1Csue9MbHn8ZyMWdc++CWRZfL6FYtBC//yJL2o9TQC1
spLoXoY7neE0nurZwJjr6Ym+mU1KqW/MDeRiHqr8xLD8N759WfOMc4kFupOlkkR+/ozXqpephBeG
ukqY6gVouC7NoUgVx36Kj4C7wLn0N4tyYPpDFeap20yvOFPnaNssTrz3dx/fw8FEu1HEK9NyNMmi
HU64VJEI3Bs1S5c3P/5baO0V3l43dCtZK4NuOq8tgWcNeulDAKlswEiBR+h6XnsUL5UuxWDTc5Ab
ZAh+FLlLwpVNYkDEKlW6sIfwvdMWRpCE/vkti+Gdr+PDBzOpm0gMNyjO7uy84l4AWwdjUknb+gNa
arCu2r3S/Xd/8QpjKEaDSvtBkMa/pv3ePzjzh8QbfY9gW23S1O18CBAyWOGxJAA1aWczXjr7vU3t
kJBUdoALsjrT/fHTsDTYilooWlil5m5a8N7AZkSB5aXTA+Fv7/2Nz+s289a7hYpvbrup+NtGbfX4
jYy2MqrTo/rrG7xjQF/8k+r00eB78bVFiyoANR1UO0TkrxhlEQg7b56tOzTTk4oIoA0VaFFZQl60
t68ZwG1c9+MTBNNb2NXebfJwQYJon/FKgm45tCl+F/2opiMICrWrA3/P3gZOX/NsF2tkiMiLT12A
J8z17aV1j8sr+HZKYJhf4y8pGmdq9s+UYFBQr5s7PPwAEWhnKg0PvhKos5H3CVkVV59+TLkG7U4r
8O6Dh7AIvno4FMVMGD98hu70JCjsZsUVw6Sg4xcYa7qOFZvM/kvquVRY8OOMwO1fnCyRPL1nVzXf
3HVnG2Y26KW4IZlS3C5d9LTkEBkzgm0RWdanJ7P/9GgCM5fpPkg52gUPagUrDEvrXpmE2nGutYOr
2ka9jX4Fi5+llQ/um7yFE5uO7s35fxIhvN2B1QgKtYmxhKqpeRrC6jiqa1KRha5fKQ2XtlVeTUbN
cCVNdx3KwgZaWv5IjZVgtI9NdTS+YXrBvqGHS0yOH5Wl41XO0A5RogloyK5Yd9T4YR3f3qLWJEIj
5znlrs89ZTj4Hn1ISZlfutDByIQUsKezqLtzcR/o9mJWp3mMGjQIp4PRsBteIxwu4+1Fyx2uHVoF
IM5G1tf8yNUlGgESA2P/2dU5qHyavAxjpp2YPffr2aAhIN5Qb289dL0JiiDRMDhznDd8n5RPdHkp
5EvzioWTgTVEzniCNiI8fWHhrRZCi96ouuhTo7jC1sf31Hc6gL8QiXZxz/K6G4yupPItqznbp0wF
GqR5arKwjUKB7hys3w/+01C9OU0BLaUyCu4cKoH75lZ6dVzo5holgQk+QMO2ljLUb+X58yWRlRev
2vaOglGJ+5UzQJDMOpW5IvBWL+rELYW7k8wN5TgNMIMjGtWAV661pnZQKZdNFrUsKOzIbx6AHqAl
n2yzordK4sZhw5ehbfCzg+5+OeQx8ZTgX+cmeasUix+YdAB4odlTojs0QHOn9fKcNU7msHWDv8cV
HhgsEbETvLtxJ641njwDgjTp5jD0HCcOYscz0ZBxipZbbudOV0PZT1izIpR0KbPRe4WLtx3F1Dmj
nUppG5wRz/oUeD8FvaPXNj7boo7Gp9W8KwloqixkEeCXwqgCDNMHVDHVe6WLRegiBBiaH9yMTNPu
5aOidoMgNyDCIzSmoX13lBfThgIvOmQn4aXVqhwhYt2/AIeZDMq1GJXd1oSkduHVY8KC5DThLxxP
AAKgcf1wSgCIYkEh0sp8h8kM4sDbvMECjwO6k6khmyOcNzDWLtwH9HF+0xH/n70MlIqKiOqL1ymd
vQVS19gWsUcy54mHW8srR1Mt0jQsCGMqAO80virZhZdZVp2+MO1KKtSP0NkcY/GIDYr9usucdj6Q
wsxUahx5rw6oYuEWpN3RuXm9Cea9iJUcnfB9Q89t1F1whMvhxnzUaAcxIYWcbew4D9yS/lpgvtit
A5ujq7OdhFED9Z0jjAK2iEk8FT0nfUN4bJ5snuz4GG4ET9ue0S+m8mee6RoNZ6WrKRmkmYzJQMXg
k2TF4YZy0QpYWLUEOcZ4jZku6KS7dgT2or7m2aYN20ywCrdPk7pQmBLGNIUFB4ZWEuXMEIKwabpj
bITlOZyXEsPKn2R7165K0SYNSULbsURGWPXENihDbxz7EbN33BVaPzTimqILBNnVdz8ch+aw8hnb
riJ12cyhL7v2HDH2mZH+Ge6JzIHBuBTRnsdNY04Pt5VMES2UB3hs1oa0A8MgD6XBh5OYwy5nnUBR
Qf7p6vXluELlClRKa3bSnLUse8BvUgNoji4oHaCu6Ptrz8zUowrCun7MLSqOXYj45v6M0yIgdT/X
mupRgiR98tCgkhpkOhIanVisrZCuVf/OnyyB99bZX01Svi882agC1QwOBw4Vw0tCSjIHNMDIZUDe
jhuviCFBoRAfeDlQV3L03QrtNfhQUSqgfgsC5NO1XwxZg+zEt1lviL5rBsyW82YR6oVnt1zS3w4c
bHpCNLmW8pvJWOYQYhL51goOG2HgpnXtW1Cyo7WEMCk/2hmo0ldaVK3gHxKiiv5lqnqB7z1qD8fB
VN40EDbTltJyqNTrk4rNFT0V5ydbpiYQOjCoMt3rryyPW9Nmpmwe8WaQoR0x246ISYDGESpGQtOL
QubVkBn1lmzwZqX+O4YgINp+bACY0MpfCYlpWUhbVpd5jDdmcb95UZDoJYhJ0R3XSYVnXoP8EvGy
B+nJulMRPzTRU/+Tak4TN8OHlv8fqmWc+NIjVFV0TbuFWJyEF8y2/hkeYrNeLoEk9tYtWCGu/ZII
JvZxMfAG4AVDjuInlgn94CrSgpWAgMSwlzyBnaYT3WweJSiBsTGYYuWAVYVl5bPl3eom8j5aY5As
AdSa0vS1fczmpVCjPXqZBnwYEOYuxkHdpn7I9cTQ7M85FQ5gwSIEpR+2J7HIpnWW7lqUgEki57yY
qVALqmb8Turo+kDU+P7ArpPQQzG2zdX4ieDJhVNcy0q10GZXSi/4lWgC/hA9Ull+cCE3R3UlOLIs
8yyJOMmAauQ6oj0VJPc16UnZLFpxI28wiLqpf/SJyzZQgO60VZ24HQoxLgosCS8cUKVkRBiWmX82
jr2EcEJlvUGY3TFc9HPUIGRMdO1wHgTxc+/OM1Jxy8/9pk5hibNBT5lQ042fpyw94NhORdBZZJcE
9Cpk22mfLP0T+AAwH8PXpAI6Ya2XaJ9kF3WKfnDaMiYMqZQFQJyHcM2D0d1ih8hNpue18uVXqh3t
UlIM0+4U2ocfvPRpYNsiMexnFBK8zqvnc8fs1bSjmekIfWotReubE4wEBIEyfrAKU+ElQj8Vk0d6
KIUXqmixiXE+IpJydaItvqjuvcqVAO4b4Lv5RhXHrrWMNewKpDeh8xu01IZlZbwMIsUhumOrF2hd
+Mta1y0jjP2IqxgLXDehmoCOITDDKyipyEFkeKpTrVYn6DAjaa06vC2ozAtsk1xoM62DfL4zEQ/g
pAcF7YroUIOL2WOaHixeBfxMeAxaG4+UthQOs7IlSVvb4cX9XSd13ifDJqApBJwQhYVt40XaLmsW
EQjiQcy13X/dULoclZbcfqnQZyWqICRq6xEqTGSQExqlDw54SC/+9VeCHPRI4ziTl01TN/CDhzed
hVxJEy78TCxG2FA4t804C88YXB4R8WO8srYOGsIYPbpUg7VtIgzJscEm/aDES4wsxas6JRMhk3Fc
PdGs3USZYwCLcD8Rcoub8G33fa9Ho7/kfym4RHDMDlbLaTGiSfi0FPDMEllcGpHtVigh0SHlzTiy
ck2EbmjSCptVCocPiTZSt57Jt2bIpr35cVe9fVf019GytFmXR14Nap7EksAYc3G4WpMNRNtPdAdm
2Y1yjHBdgbENbvQBZN/3N7HApYyaM6zvmhZXco1GxnuXOX/fV0JoioSGB4+8LZHwh5Qi32tyg9Cb
hNUpnZg0zpJhe9Y+iGoQ4/Yl2iO2GDJW7RXtpZFz49HbpuH3QFSM2wLddEIWXLUKzQbwlk+dqWIH
V62Q/+FrELRUmTG8U2Dg6rpU1q3MItUiKL8ONgKtfWpKkvIwPC5QjZZd7hRDzVaFsVEpA0vkgn9Q
hAQXoIGv0vXoHnthvo7Kn7eUfb9lIApV6E6/iCM94WJTelwBTS5sLuupxlodyw8rDytQdONQ3Blp
DtEj6QrIOc7BYniMRuKLE1H5Jxf2JkK2xX7VzhlWhDz9kyrGl9rAAOdUFYKUxe/hyNH2lwAM4YtO
8aweZ2JPtc/KAIS0kFwmPWCtGvAG8pwQfACf7lPGAsvPPvrzLB8v9icNfZsHEmSLHPwD/NoNas2C
N/GSwQkHbeUQH1NQtpQXSeuCzIzu2QqtgIzT3IKLWiqLXssl5dnj6RIUn2Er3f3znuZ4hAw6qxoV
1EIEKGyN8JgMHJXgH9sYcZu+3DuCpx4U+Oe2L2nY8VYDQYgq9ov1VPcp5+y0g5j1WVrccjyor39+
/iqhlIN+YISu0p8u/xHZC3eEbEwk6+X+keE3eYkQmzFBKxk4LOYf6hhgQ68iqAeGALJgts2yBzcS
PUx4rRQcR+qUrTY4TH81pLtiNB8TPmI42aLuueLCNgVPAsHxSPDOg8ErjEyc6Mfen4y59Mf191P4
J3aKO+jl+nNGHZKevslorj63QWJYPZsERYqbRoU8M5xKsR2OO0MS9IZX+wUlx9nIllD5qbjt6BXF
PU+R1bpg6ybOwmM7oNMEOVVU6pnOEHBXNqfBFz8tm+6aclF1vnCT0FleJBH1bUP8qojGBIngBJNn
D+wmPCJweDFTwne9OXjRzE/EUXSTRoT6/hd70eGgzPTR1iUvWZWpLFODcgt6+HkxV2nioW30ltOt
rrLpAAJPxhg4nm/dA7GGgWlAZkqm+/IuQpkIhvatTR8Z3PGX4anmDBNqZFIxWLtwryHnf5C0uWQf
tgvXLnDGnaXj+UMe16+ejBnNmNgcXPBYsuLHUUMzqfYOeyK3C7qa3law8dINPdWANl3+NkXtwY4q
FQy8YZsCW9HJvh1C7i+W5T7FnxJw6PNCbWS83gG4/LECCcQU2SB1sGOpb/eixIY4ruXnMRcQ9h2E
a+atNtb2AVjEB2grelX0cqEh4mteb1uKitiwRX2wL/d2GIQFwS8CTf39frHo1n8FRobjg5wA2Z4e
zbVZML3KMgSqrvC0xM3Ahwj3hS4k3jHBUyx9DCtImcqANM1yiceum7LYPkZe6dCrEjypN7XX5Fgm
tYRuNth3HgmKnCB5W5PsDHO/fsIFweWqahiLTik+P5RSHUAJ++KHHHkGi5f7ioJNU/7iwGD0duHL
0cjlf06u3K9olT32kpnus1LGdkDNwZUqV/u0qVqhDGbZhil5RlsVCG7FgUFjQfg7U65UeIL30y5m
r13AhaWORVFiwh+JUV1BMcm8/kTKbCcSSbiNRcBBx4pX8w+EjWsU5mH3a846O8GCE/Za1bhmFi1t
VrgJljytU6LtEMTuxnUiPlRv21FmV7tXsLrIL8NGZSIlGE46bFFNh52q4wofguokr+v9UL/Q+REZ
HvWDh3PCY7qnpvrspc6ezD3lK2Km291VwjGUc2jYs/cgLD2AgHttUEjJ9VHehFwNEu9KUssmo/Xe
I6/YPqaWx5KtwVZVsEVUP3YZD0zT3pg2jEtcHvAhmMR7t439cOeLe/pyY0kCUsMK33TZXY81EngH
LUtNeffjXqaJI2pYsnUjxDzyhGWBz4zHne9ldLYFXDGPmDU/RbPMKEqCApF7P4noCYIgSCp3pbSI
AVUIvPsx1mRiohNM49uFAHKoJ/C0/F3FT2Fjspx46ExIlullgUKmAUih+prekZT5Jj6CS7ZnYrW2
5YwrUqgnwgxNm0tOmqhSefRosNCK8uyUHEPOWPGYvCcJxRlHtA6MOz+b9F8UHUh99L0N1TmqHD09
emkkXD9bLLzIHTWSlDBB7jIbUz7GwvPi7PFCriSOBoeH8Xxhvw+SdOpYSSvHq3uzbUajXLxxE9U5
Iqv/3PDvhy2Ky8RMh+Pc43LB2liy5xP3ptU6syENIY8OQAnVTQbqSMCoNqa3V9zfJjhRoZ3oDVfX
3Gz6Sul11qhgRkdK+SbCZeIfm5kVeI4Fa3VVy39Da45Xmtof4gIu1h09ouMyjCWmRghA1Bx1WXmG
QC7/MJGnLxpqsoQY09CHTzHKOrIwlNhPAQesar9bIQoH5+1e5Z5Xq1xntZpfRmCc5hP+muLH3h8m
nj4QdBhFCxxYVxVF6rMkcw8/QWKQtO4EjpM/Yhh4zql8rrOuQuwR1tUDBidE5/fT3bmTm0IqeEQu
q5Gxjnt7AmzoaPwxaox0RhzJmCFlAlJXRfZZtGUVbnlF/Ub9ocfQToG/S+gSTnOZfGQ26YLTjDBc
SXtleSQP0hti0VNmogbRIsJNy+qoSBtdxiu4roHozOr2VjRkbDp6W+tH8rfXMBpk/b6+i0nV7qjB
hLKKucSafaA8aap4lj5sVqDIYnP4UQQIsfmkhvsPnJkeq6/A2qLdpHYRx301nZfc3LZIPWNtDc3m
9CP9Mosayj5VZeJuA2VBNsvwUsgPOyB7ftWJV8OAb+I4ZDyfhOci9nzDDgAo9SzXI9P5Ww8Gm539
Rb4l7G5hk8d8q6AzgKoOmVnTkEkodQIX8Qtu5FrTFz3D+nk6Q4W7TGix4rAgDdJqgsapzUXnYjji
2vcl8JRS0kI9ztiiG7Vv952uwVXk6y+zNF+EIaX2JsCGhUaQo32tUAaGTWqXlGdOef9Eq5g0qQZL
1Wdaq1GFiARBEdOeCXOZaAgpvGoLd5CI5xEyClhscK0htuiJdqKP2dEGgIXd4AAZF8CQtFH8pWQG
QVi+MV382l/9scu0keeDMCIxgEvu9WBPzWUAHeLvjkaaq/vtlF+hxJWRbgje7CmY68t2QiPGAfHu
z6FlqvcEXXYGdSMVQ3ZRNYtlK9pieanf4j5K9FWBTrJ6b7QoXpixn4xgX/X2KH/pUR9zrEjFZARi
KtPIWZ/bFHYCd4fdbTK+9Lv1e1JK4lPPqgzXj+57aKzVqXbPTH/fV3uvWVT71MNaRWtFtvjVxnBD
Am3YpNGN5dUhh/4y1dFtAoivCjvMqPwZvqjm7bnyKp5W95+PZ/1HTndSiijRfqG+GASL0CdZQrLq
ARHDDfaVn1qu7+Syc2yzgQ2pfFTt8zgbxEH8trClnw8uRHDp0a5aM27rBgb+mlo41w9NqHT/t0zF
8LKMqywEXeOGj/TTLHc6brMv1p1bugb+oA42btVPfmM5phu60cOUeKj467aTCt6yb1c/2cRuoy94
VCMit9vC+z+ey+P2HsUx9iCV02G5LN9CvgzpzYuIdzChY582NTI9dWfFNdZRxfZhUAVs62pjLgT/
urvf/esj2Cuvu5AaYMAW01W65OffjlCjyv7u1i9L0GqbpVInRi1mAOmP/IM2q4b8/GwseWaqeqqr
yiG+Lx3YWxZRoRBaL5nfKvnklI0fgBvV55zwmTgindlvpZPRiA3vkZjnZhYGftMwNFuJP2Nj4VP5
Rd91BxEkNac7ogzjV1s6fU/D/eKVgW4xbkoSRl5d49MGIyygb0CgXpM75YbPTe6ZojUEv9LhE+XH
lHcnYA3BV/RreteqRUG0eo/+6/4aW34y2AHWHZUN0OTZJjq1zRIQRa7p4zxWyuZ+h66sAJhAaDBV
Sy3d77VPhkRyPEywNsw68R02j8RNGfyL8FlJOnqcq3K1AvZVRuYdCO9sH/j5Gf2+Ik/PRsYfyv56
4DhHUVimQsKpOQog1HHXwIobQcUXViyR8cxtJCWepM9wZ0ABv9cH2G+XnswHp/rG91agh6wi8nDW
mAwAI3AV8529PWp4HyE3xsxrTz3M//Qr6g6yXrMAw6q69qLu1TTfq6zNZDZs65wuB8pTCLAhxwNF
Ik6miAaLZBnNHdsN+47/wWG8CKwhS97FEihEBYuy2Qas43OE+sfHgFy+CcRLH0r2kxZJ1Koc+YdD
5d9wKWom7n++tQ5UJJM5LqyglAIOhhlZObF/HxCLb3w8MoFkOOMIylAJv3LPA7eMdw5lAiMecmLJ
zUSowyLVv9ph+wtyEuMS/g46cJJ6h34zbax5RQMRY69/veGoB3OfrDYp4LEkqfgqzMfa3MqQIeSt
GmY7ryd7Y0UBQXG0LEMIvPj75AovZTTrm+zxQ6eIoA7bJ5Ok1MDlCveQtwyTvsVO22V1fHVi4fmJ
BRedglpkRfA2hUS6wlaQ7Bg4sIdaoqCtmPQ2iTCTDzGjOqoNxsBlqTJMIXjjP9qUrteUTrmhV5M6
2fqDocYzCWlH/ji9RafgngRdFhWLU19PFKFTE38wnhO35qEUOYZp9CMnRHKDuC9LUOCnWIh79M/8
76KIE6Vzkw2aSevi/lAWKROW9b+ma9iy34Ff0OLxxm1rYFEg3FtK0cAFiWSSeTU9laZ1e8vtOpoq
kHGg5TStU3fmvTMi5lMhpy4Yj1haHHddBPK4Tuh+O2RwjwyS8aANGxS0lFqsCnD+nPAToOMqk8T3
XzjUmG3zDXARWsC+IJJmSCjW8PBQKDyJUHJgCLyoEDkdc/cAB8siVOuYFqNR50dB7CCN3pqUo5iq
vdHy+gLuvfkEXVdhT3CuCgmgfRJ7k95OxX5Pn986FttTeQvA8KACDtTlKGc+yEzyPNfsxta+81Yu
/pCsgqUzT2I3XlDrpzJmxrW+S3Ru5A4UqTsFOnqT6AX9zPkLz3gMC4vSRuW+8xsBfJcS3vfhdq0V
P4fbYkDltWTu/SNKNAw8810pEaFf+pV4vWqtK8jqR/wzcjv0jaBrcjKE7rjgg+QcDjiUavTVylSg
29OaBgsHkWnLVf/RHlds32H0msQe6RrpN9ozcDSlc/10I+7/fHzeL2p5osZAKZjAcYWCg7AzZhhJ
UU3Czo0ctie4UXKybnymqAXlUXV/mD6XbWAa+jjJ0brh5hHIOPj6Bqjkgl/Nm8UnXW30J6D7iEPu
sqCGSt8xo8eh41Cd8A7QDJbCEwu4ChvgsPFKLeRpjrxwMMtI+XOQ/CXdP0Wn5RL9CFrFI+NgJK0T
/IVAKRvncl9k4q+PSIynEY0XyGxfoeS51vlV9YcIuYZwDhbsUyXeLXn5tzrYO2/bbrOhc/fEUwDj
fd5pyCGhkMhszXBK9WiL9UZOuhQGo4ouS6lcBRTbq8IthOlThYnD6m7ptW8j+PbMl3yNhKRZLKr1
A6K97BLQ91z4PayRx6DOC1hHpaIKKAWq3MdSfE4kM5oxVdpu3bhPRlyERtsVEkh334cL2b3+tem2
VYibA3+fLib9mChxKoJTic7LHkFNxYwSMGZH3dfIEbOFt8J0TsFum9r3QLiuNTSLg31uiI2oMArZ
aErdE9XV6f67BlvjjEAQOGrAIZ+g0CYvTW0Y9oiocHKO/nfyOKyjGvZJ5v+TZPgfzYh7T8B9v2Cr
xMYZNCiAxlAygPd7GtE39oLchfhIFz4VbGi6P2JRtDyWSE77GdIWA0oy5sLtjiPmk55Q7FAptKWX
XE7Xw0Uw4tFP9yEIqyNSwCJVhNbuxzwKMAR+t7g7Tll+v8KNRZseWJ7ydHGOxNbzlX6bBn7/tVZz
lOeelnOpHSLz5tyjQ60GBORg2iXzRX/JZ/iRA7YMWtW5KgSSmuuGKrZ+hCOtiIcrgjZBtoJ9NK7N
VabbQW1qZXL/aiD8IAC9pBpASkDtpxyr+FHUL/c5E2YnSMPGOQFHa61cfZXf3A/pKbf2tJlv2w7S
BHJA3x2E08RR5HRoQ2q1NHNL3iPoCEhsDak2L8Tvp7xRhw44VY5nVDBx3Re0ucLHdRnJJ9RpoU6i
ihB5AGOS20/+LpYCyX0JSJWyfGItks8GWecaJzCjbTLis3WkwPO8Yd8l25jBnN8CHVFCbfM7fIsW
izNambNJDTaV0EkMHD7FZHJYsrj4kbWx0MEMe5Of/mhtLg5JG2oioRT2CWTzcVJEL7Qb3J5wBL+F
Xt+UkrRnGTsvZJPjl+ffqylSqIL9MTm5lS1RNePNemyu0ZesCLpkXBn9n5PEkXUQgpB21QGrw2hE
0hHBTypwagecBCeOpodeUY8z80CubGci/aEqQIxG28gOoDAp01dBL1KWso7Ihc/uG17W8WP5/Ka2
UUI2+nDtjfTyZ4BWGtfjEo8XLCp507duErFWA9rrampC1W/SZz3VWw8FyVMxAfOIQRpG0HWMkL9B
SqBozlzyYkASup1kth/jtpE5JFje3Aob0XFJjXltoHlC6Ll1qMttxmPhH7cxP7hVYSW8+eZFitOr
+aer9ZdsqIrDMwK6t5FWhdcvinJ0+HfVtIJbZEx3QfGhj/R54OC7+n6K5Ev3SXjWWQu9r3b3YGOM
UzdLEyDef6ljzgkFPHxO9zed0YBW8jvs0qCvXSyuzaPlAVVf/b/ZbWjhdU6/ThhVcOL6tVP8/cQq
YwqPFKC+zlBRkZeBNUd8uF2wJoRJ9Fk4ve9O6BO7i4OcfVyfU5ojnKcMzUXl4OQ6xhvaiO2A+WWH
CnQkHnrG1sr4Kb2uVjD7UKOElNkTood3xb9ToEMEDBiLUikVNH1Z6EQHQbrSlfvSYgKvCadfpf2S
wP9K2IfNw6ihLDghkOnLmHrR/noXQNAdUkRnQV0q9rxOfaJ0eeiqJuyP0JrKc2ZguKGJQDclM9Rf
PJEtVcwhVLUtHPkumd9kqLRnVXDexoHCqdA45wrUiUJbg/YjErWuqxN0Xk91AkMm6D5kkqP6Khem
NjOfgCGwGlJ/JM9OM/W4tCTTpFImabUi6pwsULicC3ktZrk4VDpfBJaA88TarYuRROq5BuchxYaW
Qp/tdrTt+8SSA/FttWHtEQE/t+lwH/xChK92murQX1kW6xiIE5lX6z554blRUlnhOlqDGaPkURST
4VIHjhDNUeJ8/aH+EineceqQS6IYYpBE1uyJq5XU3VoAK+g2RJMRHohxJ7VP8HWdhGUumd+BjItX
y8XO2bjQfLxrFKXiekY4NFgYT7ArKlaI2SWz+TZeFNDawI7FZyHU6sYwBSXb8XOub3GkNuP8n8SC
PQAMp1SHcQQuLBBTQ1T49lzIdFtyfB9F7LUqFEAADW+3ID6evvdy5/ui2F8kikt3Hmlz4HP1Z8C5
NW2tzAjLwhaRCQnbJGD8JDGS4ypF47VHx1nhvnJeEqjFFPCM7uI+LU698Wdw/LzL+5rFptIt5E96
KVDXTefpbxyysyRdD/cv7XNcF0BpsE7Bl4yK+Q9x0qteNsWGG4AsgWw9FqACrEoXYX1/BIsw4TSh
flWS7/GsKLeJqRnlayBhaKRK4MAycSx9i1JZWQtBnKoKAJCjVJ01aWwCMTdjqLDqkRWBV26OT4l9
lq+iRX55vZi1J+Y7aU546Y60we3IJS5iK8GZkLoj+qtjb2qg2RmWSrMt2csSfL06SmmmMduCIBbb
lzZSKrxeiQT5wfqoksYUAuWnj93FuxQYUbjQ17iEUSKohD08e29pbrD6J990yzeHL5iSFO18D6mA
GN3nSu9xHOlizKVIn4PFm0KFp6jETMLYsTYUB9UXsBB2ZXmbwEPjZwh0qrYbsehkwQ+wD7E/OLwa
Of1NbMrPQbYBYdl+w7zW4VDNmg0vt8WI6ZTqhQYc/g1elY2++ZW7/3gaGr1ZPD8YPXG8XYC7dAvZ
TU8uCa61iZ27+9l5NKbJ/K2T1OmyLVMgTS9e5uP1b2eT+Pe5UjWj3ADSgFmaPwmMF/jsewMKtWE1
xxiYMXci5a/J8ctvkz7B6jiPmdOY8fs+zzGNSfxaDCqaLgWEuNjcfRutCRdlftUDs1Z8lk8bOSmO
yoJvEZoDOmI2pmfoLJiWDmNj5TwAYIVrE49pbY+DH8/16gL+EKAqSpJR+LQsukE7Qez4mcJujvUc
WMFF58HGCe3MiwhH+i0J51QUC4L/IVNot6WEnecr3uGp6pgKn+kpgTgXX70lHrx87AwGYrxpJUbI
fmHpfl9w7I6A3wFodjN/3zoGQnRKQOEln5dOPSU7gCxu7G+XrSS5VBQNoMn2ev9PgDn5FwUKn761
PR8CV5lzM4eH/rEbe/7UJKWo3VJ2soQju3TMptrMHHjA0TTdqppZVnAZLcGqRgkmpaU+AQKXC61C
i3ZD28d2g5D6E7DQ/Ze2yP5NWTKU9H8gPuDjbJgsWmgrLO09oL7G/DrnLpcH1b+OuuTkiJQi4jMK
OPlzR6+V4pTexKTbXDs/JJ5w9JqKj0NhEo+UDXwmVyEyLRYI42Cmi7/BKVfGaOe0E4xirfkubLWZ
Regy2a7sDjBMYNDhQ/nMZFbxuaAx5ro5DRG/iz+IYngQONnFGuE22RnI1pS6Y9v18v4y0SSu5O+W
aUNHKpQp2Qp8LbhFRFoy3dgMjrc3vomhdORqXU15+orcQS56qmw5gGyT+StqXS1/sQrS5iIwFrB2
FKvktOUOzItXr6K2YgJpJDF4Als7IE/5mKVLMIN2sxH55LfYXT4bVB+dwQcEMp4XP9663Opctu+i
67/FtCeoTrfbjCu7USocg10T0wT67kBCy6eFrkMczPKNop4nF6veyD7b/sMt1/Dq9UBwU6A/kcet
05LuU2ZRouLKYiCN1n0RqX0lphRiDM+AnombCpovTf15j2DMmhuwlpSyW15/exOlNC1FaqhM76qN
3Xg0dZOQH8QNhtHH7OHQpbP8RfDRNGID7h9M7X5YW2TiGnFtfD3ivBPqSUuqD8A+IJmwX0n5eKoD
ww6whV1JbgROBhrvzuBAWjYTilgPvrWhwsMEHq9r5fvqaAgqavHlYuO6YvT1nHv/6sYHfaX3kYqn
8cNkN7X8iZffnE20fmsxWYXzi+e4ELT5JC/rHH6+4oLVny3ONCBwYAm0NA5SEFcEFiPH16W3V57G
kjbTJF63Snsx4GKtNgzagGbaFkzyUBjc19t/QPG7kl+ZmJLvLRDL6PF9OukMyjc5VGyUaUdoQ8ya
OP472H/nO+GF3TRdt53fZeBy09rVcR/+2IgfzB8WzbPQRYT9flZsoR4Eicur86s91ATy4ntSjy1D
xINlnIq1IkNn5S6IEyrzR59EUA0n/MhM/c3z414IRxxhsJsSWZ5n+Q8kXrfUq7h4tGT2mKzReRQ2
Aw+WjjPww1AWpRRtIY9rpvxsWsopABH5ydHikIqSJ4vrTSDwXzCF4lv26FwukM9b+u+O3QENLkV+
XlsMf3BGE6NuVhOlk6hJF/JBBL02bHHJMNzi1ZQd3utxTizKewHS2W91Q+83J8F5o71/7jTmpr0k
h/cVv/Exoe5Kxt+/KkOe4T72Td0QzXHnYjwpb6G4USqM5ZCIs2muSjYQZNR4w1GpeMKnu2fp5835
0BJZjxBB70F4HICkkwP4v1F5BhJqgqH1ujRSIXW8hqCIEuEscMCEuCgchX9jouCQsJhRK0Jl3GNx
C5+iOW4kd5c5cGCg7Cgus/ZhGsG3Nye4FKkHxnoGjDXdc3wZrCvIN++EbVhYU1z4CO9l09vy4PIE
/4EFlVm2MjdUlZm0sV1PnLfDdrmQYpbpBvNF7tokWqVp3BjqX+Feg6GhEg8UYQxA3syJ/pN6V+FB
Tm5UweqpALO7RY+GFqsw3IE38uUJlvu/9qXEAuDpawHB2mZ5ySaNxi7mE8oajf8gdIyt6EsmCMQO
hyXRL1JGtPUKiL4lHAlHx3q4v82ZjHu2oBrvPRkmUxYZmBiW3Gr5dC57NjdjS+Gr6Xh4OdZH5bze
auR80UYR5m7Ez5E/gOFW+bWPq1xwHgpQ1dvZ3I0ne0tcWXvN+nkymwSplKfP9DdWlxRnJxmbRdsI
ayQf2B48AQXlf3qi8iGRf/55Eb8WVeiVbZUOHuAFGQBFvk+5QkPw6aeR6KbhRy/HXQpmhEFzhqZb
drjeSTSTIrQDDfopzCuHYGsZXfqspIHq+0kJO//fChT+7Ow5FE3qlBshZo8lwRjByX4PoodX3Wq2
A8k9Zs0RJdYvIplfEjzI78Fj6Gck2pknjpVyr/EHALKWQV5vpeJ7i8Q9hia4ror7PXF5TCngZnv8
XyybJiIPJntYUloTn7izqXrF34Mo1Lj+tH/hXA5hjQbWJc2YyleyJRmi6Y7j5cG+xMbN/cET6ZfP
NFvxcg8LOHNcUNBRl70mhiVXF04mOeM/8iFPfwOz9jgF9oPp0i/Vpkn0rxZdGZrM8vafKBY0oJvJ
aVW6XQgRHlltgI7gBjfuDZZpeQJ1848U5tzhDSJjLQRzyq9+Iy57Pjgsd8uSLpsIPv3XXIprNUX1
v4TfBLSu2x8J0MummXTx/IPR7QmXlb1HWsKrVdR4pkA+70klBn3LOEYouEQOkLO9Jsl5nd91F2f6
PO46Pi6oCAKMFe9EU/YsxDxfq+cHsHYTPlBM+1DQI0TWUPwFyEL0pXuYiYYydzxPy2HGU94JWePN
eyonWBaz/Xoi7zy9VK9ROdq6O1BplgD/mhz1iO+fcdAAGzn01e38BjjfBrCy2+oicadtZDRfFIC4
hho/qiu0CfzYXSAli6fMHiXiimV4jHHBsn0ccHQxS5q5vey1k7RvH5hZhsSgsHD6XfBCp0+ET5ns
SOSpZVPWWJmwB9lhuXQjklbZitS6lq61mDpupK/F8nhH9x4oncnGEib11hxIAwX8J2GUVk+zXMrS
9CgTvTibrodg4G31rAGeM6l9LUX8T29BiU3w4jwBjdxYhA3HJi51EIy3+5CZPsJAp/ZpUt4BZe0m
TAHZCLu5e2EPTq7AVqfng5SbKPa9biAlKgJNjLTtlg3nU3DIoDqJFakxQkXlV01n7/LQ6q2I0bvQ
53za4IF5F836bWbCTkbXbel2801y0uXWxWEv6wfweftoHhtN4xt9HApkHiHysrRc
`protect end_protected
