`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
A+UQmdgqnUGnZvePCu3e7W/GOD/tB173CoSBuCqm77AGlFJwUgwxjo3V8H2Un/Ly1uRI0XJ4Xif8
kn6XuM417A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LcD/V3YgF9zxqt7gN9YsVVfxHbSyx3nteYMZbIe+fFunCA3wg//cCLYoVclpwHDoYPiegwg4orEa
UclpAhEo1/uBFUukrvvN+fSkqD5vq1hPrHSuS1JZxVY/vSyixo8jZR0BFyQxSGtiX51b2PTZUPWH
1cCvJbg7rLmn46TzhWM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZjuyV72G4Q94JZ7xCuyUL4oBzU6oHuXhmatbMpzmnr9lDvZ9wn0nGSkg7ePzXFbcX+S2Kc46S96C
BMR5VB+4OJzW7Ms1U8J41rAqWXUCEyLlh4ZfK0i7UM0HMm1MoUEMkqH79bpqzBmWxO0wiNeGNyUh
8I7Mj1+OJBz7D/L2NoMnJGYkGI63f0t5Eqyp38qw4osaBs/5j3ryUsut/E2QB3lfgADEMMhUE1kj
ccz0V3YMjsuL+eGSiOS6pZvj60Xup+bVKQQC+gJSPGbKdtXDvmNAKS/t+/5dF0lrpQqfIzFulIC5
zKYnyCbWF76gMhncxxc75OWtnG2ISeQQAUUNGw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RDF0CxZoqLMbhcouSvutLMVlvoj9S85p/NTlio8SaCb6eg2dEY8gCirT1S7VPycCYS4b7pho22hU
Tb3U4v9aQYQTWMToAISqA9YejesKXGGeyntUCjuwv/weOmaBf7+NDTa9rRVnDFgb/bjTl6z8Y0q4
HSZjQuE3yXzQB1uDjaI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bitLnKRHSsenWN8pJX0zxngajTks62vUFKKyiIhvC3jqdQlhvx/WnSxkmRDOEO3lcNa+phrUig4h
4CC6o31Rc0JafOB0d6tWPn6CxwN4ej+e0ZiJ7OUcfTeVRZNpkEy8+RE2G2tnfncgAqVpMRF+dZdh
nN2Lqju9J5rDTsvipxWjgz1SOiGifpVq1r29zNmwLSrDA5fiAdYTTIgbvg5BnOnAZ6iRV4XlhCz+
mBuqtKYvxJmQ3MT8zVsVWESAsGeuDvkQEWWu5UJI+EibMCQ3V1i4Qv2fDNptsSLFucVmJ2TNxYRW
Mq8ztJVhicQGG7GNEPmz7PxCwkLSk2A+O8FbCw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 29312)
`protect data_block
AKTURxVcLNKTHL9NtGPgcANclX7BzFjXoP86cQWPi0/qLIZ1df6zEvE+bblDvyRp0tIewySl1DpM
Mc2qx9tNB4GcP/20aQGRWVfoq0r8YF91vQoFyiRrdrwHYkG60zq8ogPxQiQvC+5tCzr8lVmMmc21
x5RJ+x8MYVXfOc5bigc40aXTFsTQXsLBjuL8XSvAIw80xPwJh3OU7621zBkiN+4Uj78vKhYZITDJ
kZZoBTtTyKETavSWagJVQO+OCNtdUei13Ybnfo6AwGxitrw29+Z69PMfUmVlDJxx73XHKqcnAcb/
Z93bk9ARJydDB88E2Hod+VAFAwPzFamMcdIuwHvbK5aV40xRII8NstRAqnyeUF+pU9ST2NA45937
Pp4oLBXXxvyGlbXGGlO5PIFjRzOvonOw+l55NV1mNfRpdO+6Ep9REvSa/0juJ2/l0Q9ZvI0fJeZ9
52mqsRYP6JnGFxsJGAYAEmBLMN5f7y7gGC0bRIqM87YM+JCgPiwDq4azCcMcT5YbxlWKqa2605uJ
c4cCZ/AatJjgMpw9flDWFT6qaJruZdXb/AY3ptf9g69+fplABDui/vcIsVE0aMB8705z3f17puhg
fBbYpT4Gn+kPCK2ZdtP/Nv7cpIu2oR3cSsfWUoie6Qu4pJoqvMBdtIsBfoXbsJgl1gPqNQKi/vJ1
qLthGF1KTKg4ODfSPP0+9LBg18e/mQj2+S+aEBD+RyQfSMTJvEY4JUilShi6Lfz1TtBKr1DduAer
KwyOVCbQdVo+RGRhl6O3yQMYiGtGeGV5dNk/JT2UK0zw0xNP86cbXbEK4xJ3Tyl4ter34iBaOmSQ
Fqn0sKz3niukHv7Vb9l+EeZZ6csXVLTMoetlxl/AjsUXjbw1OvvE0t9vbqXHr77aVviuEWubbWsT
Ta2IFQEXEbX/WsA0prmODbmobLoDPiHM+0tCz3RONx9+YD8u0fuCgJvlsi9VoRE5RVzvB/dMxbh1
th013wt6/bDMuWn3ipRyVxzSMSJVUzdbmZd+Ezl9TvvgKnBEcE+6QO6YvP9lendR4xP4BALrXo/z
38k50Gzt/Vh3pawWZzAit5x1LGZl4KxVAfPzSYwNQHWDBhGZzT/SweQhc7MEFZRw3h+hmOYcOn6x
yTCxDnVoUgq1gAoN47Lpxq+moedy4t2Ws3igrRXxxhp7Xu+z2H8fCKdpJe2L0nGpeJJFcY07X90R
VCFMgMf3x5HV4J72iSc/0uMAin3kkrHIvt1ziyN/DnQjXFQXUBHe4g3JeQn62vGkxa9PfxnIoRD3
wSPTDGpJ6dik1dHK0VkL//LNYtZOpDFRhLX6n0mHw0z/5DhZ1pvboQN+wI2vWE7/yRCt6o82JuJo
UBqPbyPvIQ/NWOcXQnXRSvEP7oHxrc3R+yJroOQbBQBwM70ZkTx19Dt/OCLORGZh73dksQrMGDqA
rw37858K3u1ZaA1vbtVXT2eGKIt6GiSd1jAas9YLvLeoTkxQSoARarf1exyCymNHk/bKOc3Xy7wC
kLFZDL4P5nq6dHb2IWw+8o+fWGWPsY90MrNKVAPtuXYAK2p2JD2eEPausz588hvLZToAAjZ2ilbw
VB7IUVc7xI83NmapbY9YhumYj0XGKjfG/m7ZHIJC1N3fYJQImp7YvXgwEhCFlqnYpwgUIVya/VQ9
H2DJTii70Sbdzg2DKOW9lvheud6bxqHx+h9UdjdOEl7s/XNSvGK/eA/gElMJAJ82Ae/KsP+BrElm
26iQKxfQUcglYB+q0siK8NI0CbwgoPtO72gkP4cGKFuiS4ANONtVCFM4mQIxrj4HbpVp3ctsdMN9
KJyP4USJp0OMSCZb/C1bZAr1W3b4vqJGRrC9CSOSX14HZ8GALEysAc6mokAb17Nvjl7NjN4t3G/y
TLrqOTQoZDeOf3q/wXLceooyUgH4//L8uXu23qDlcDaweO+M7ltl3hyE63lvyTbGlJKRIlwqcpUX
i7KBJAloKhjyFcnvYmRarHd7uilmGeAmyPI2YRYUGY9UPq9OTys8XH2Vc1ZqjL1m7hnLPhf3wgg9
RemwiDKB7sYAv17BtgJTTT0Y/eKN6qL4vbPd86j2jAv3zls4Nbu3BXAnvI5MOmmLZ8M7ZaaemUnF
aBgs2czzM6+gj3+wIU/jXRj63RGFjMhjAFbx8mKoqOqW8JIpt5eTBcscg25e+B9fPfuj7SlFCTq4
CSCWGXE/Y17XP22cD18Bp6vlKVBLFADI8uv/mEs+rIkVv3FuXjkxNTpn8LAWyVO9rhH3AFpyvYBk
GzboK3MQIg/ZxLeOiwSb1QlmvhG/qbPc5SKvKuSRBFU6FZFezxXw7RuRY7Q7TkGGWOsdDA9pjXAV
lT932JSWRD/0iqxqjlmoQoJpiBuuQhCPFHu6vEoU4n15eFRp4wQMoTWh3QWJGaIFdQzG42j/qGz+
ZpEmrlSOPtszqqa6UfAj5jWEW7Kl1XNPDpHVI7/tqfPWqJb2fUds+nJsbHFZ/3WEs7M75NxZU2KW
at0oO8yv4Apk5+G2ta2LAV50FU1PrUooJP/uK1TKM5RHXwVsu4IDqmDU7UKWiQgDC1n7YQgM3qyU
7KuRymp2vSwgshDYsEtxbdEs2bTZuop7IC1tQILz/efZFRD8jpoZc/BT3rr97gPVuPLDt2Gi+pZk
dnV/MzY8dA6PI3ZleQqEnTSPjaG5OZR1MacL9ujZRBID4huwP1d1YSWGDucsP1f1B3O2U8YIhnOv
GP2q98RdF3e8x+HgUWht6WVBzIkichUpU3qojKxIUmkjlBW1mJoGenQqdPOLxW65ll0opdB8/jqp
Aa1DBGK6XHMo3LykLv8nJKjuym5510scn933PRfqLUS0bU1zSr3J96nMZ/N3k7vYzvBC/EXl1R9W
D3FeLRCfnk2vlgtGzIxSv/CvzXyM8zfZyhcXvrSQt5mQ1g8vteGQKJGN2XGUa9q1YVyIgiYwifGQ
GzM/El6v6errD6gEoSVVMiq9igW2hm+8NhjBNraM2fwG831g1ZVJCS+XoU2fVDqdSzRO0Md79JQd
yRh1xSjvIe/LLtWCvB5AXqArjWW1a7wc5Ndk05V7qj2xv6+PuTu13xFka6bNQtm5HRhR7sKJdoiR
0+FITReQDUeR8VdmJiGoXltEeJw3NpA4+F7zGMeagKYABiJEL/jQMb0p86JXPbZxGkQdVd5VWweO
/RWrWwi4D+XNzb470Of3Dl8/fjq0zTzCqeFw26wYFcGRU7OKdcL8ze6BD5ExMBvbYJ7v/q+0kGJv
3cg2FwCa/t3riVX0zrf041YDpyfaz+kGLiD6FlZ7wfnkkTE67t9MD02eQYD+wlCOlsmAcVEUTkhL
SGZxSYhUrjFd0I96nS3PVqcg2FhABGmznyb8dM1Fk8rD+wRCPw/oIXiY2ntkb//xq5Xev/z/cQUs
ydSfPsjHOc+95OFmgNdCHpkLCZxHhRiRAqqbocWc98VcMiPWh8Bbpsbhe5IaK3wXk2CZwyU4FQdU
v5tBP69GIIgLTWTiD6KvBtyGYDLVpgWqFJ5Ksx+EsOGVyeZ7FewLoI7RQU4nNS7YtZi3UV5+S31C
qRPXbS0fQoLfG+ltifJMZ74qvAIv9LgSitHZc5oFxEJMgKKEOBYnlDamkf+H+U0zQobO5dESugcg
dlc5x62G9EM1zQKtt7ZLEjqGOSY1UUZWzYboZ9Akv9hiwplfRzT/RhFfiQ2jKGMDNQ1iPONmilqP
dM2ED4X+J+zoU9KoNXElAV+8Da9vrketNZ/t7p3MHbJ0ZVPYe7EMxrqD4+39kKESBxW2mn/BMRaA
tn1eC9n6etTohV1iapDhHwmhjy7muod+R2uzEqhY/6Adb/w+EXYHV4fk3lyqD84+ya5JtJLBlv8h
ha4GhO8/JgQl3Omz1q4fI8EcpA0aq+hhoNMC+RJUODVj0ANZ9ZWWNlGTAuEIk6p4mrL77927xLXa
XT8YSxf8xrH00K6ivIiiGzu7r9bM7569zzH3AfE7ARy+QPaj/Wdevz00xj4G5o3P134kkuhMLCu1
Uh/Of60C24M5pVXFe/+othhURTF1RQvVRr4vON2PLGboGSa2tJrqAJwo5kmv8dpjs29Q5CXLeDlz
PQlYX+mZ+h4hCBdGmJTKKdMms5PepPOjOTkkKiQUto8QQhAazyPtWaTg0JD8dAOydzf07scrttzv
ipPfBkdUjzQ/k5+k5H+sUdo1r5GpHYM8tJIcXamFYMvT8W+yWAaClYSY5i6Wk/XhckaaYFoobcnC
QOprSeVZOgOKK3k9GczeFPS7hGKQUD/msBth+QAbvYYlaK3quyLC357eRTSWVPEyPRx8a0bBm0n8
t1XbuPjDl84OKh9EeayWZuxxOUoov7uhRMZJGfKt831cfdLc7HZ13s+5+/kIm0CWAp1bvr5dsihB
Khq5h+1qvVuX9k8C3WOnIgzD4A9k0tjS6xV+fGL+AwScgJRtW+eOH8b4JfiEU4jwd1bvYi7Q1Te+
kEmd7lG0uS/HMHxzBqhebUmJCe+bLe4o6e2H47nLbtoFX/hkOZkfNxqHnfv9RHs2kY1E5BMBNOSX
RWeecjtRQjQG/MIlMGWE/bBoZMx7TPofPPkzLWFzuyerN5QhgoWE3yfczXPqaZd1cgNMy9xR1pl7
3qE82NG00N9i4w7vcHY9+9aJXdCksg/i4NymEk4G41RWj4dvAnID2Al1xv4InvrjpuNBte+SYSzr
HasQS44xqjezutskGYy8Q1UuZW9UY2HW6dfNLZoj0fp7YLIiPPYPM05NKHELLwHVMBCaAm22upV+
9CsE276wrWBHniXXVFSQh40xnLDOh1VradS8p/T5IXFj93jM/ZqxMM1qpVGVfyhmiaJQ7WN3poBy
DYLNUHIrMMfqk14/tN1lvG/qyN6RnDUOlxRfcBdZwCHjNoxuLWNpm0f7yg3CB/Gy2UEK8kxC84Ep
6Kgt8rdgym6ODOfxQ065EwwbVfR0KR0SHcWoRcUkivmD4ozMURd+EmgXZ4Y2OgFj3zrCAVBn5UDT
g5iHh9DfuwxWtOH4Hi3ZFnzj8Wrv8zKv0bDLQlKmEOkecHaIH/TPlGJNiIMLMLKPufzRXRilcmCx
XGkldRs8xxamzCF2pDLwkyxmSDBvV23lzLjFMkF0c24JuDJXF+/Bputm3xWQt1lDDLAMot4yh9Bd
a81TQTCZf0wZykx94e1L1fuBGYb9nyJu1Ai2U2UdH0G9nU8uR0yZI27hDJ+t37JoFMEuudEYBo2B
7n0BVFlhWb0TwXDazYCtCkgjmEGw9xiIWiO/ZW0NscN6cdroYW64K9NlrOKx9dHcBbsmOOhYgG60
fOoRllxsvS2jB+KvQ2sT5snLSk3gMrcJkgR8L6Zhy3tCjs+2Y2ICPMu2gneOW3ZlulxBLQlV0DuF
/3jTE/X9oLs518cHC8R31aDwOy9Hhh3WCj4Ljd7LGb2HGD1JGejvduZUhT34m2Tqhjh40cxh3XA/
mgwhzujxUTpswNlsUnOmhXiU1eM5oplqXS51RCOqTo6tKRvOlpGUuRAMTn+m/cxuB8Y5lPS/dgdW
kjemtzLm3Fq3DesHRpiHGHsGQZokaXSZWQgDNr741kNAYcLTP82IbAsaBj00MtqIF8d+ZW/WW9FV
s1Y0Xa3YsiOl5iJZghx8Fwz8SIlep/0Fe2OeDxxohNl1CMq8XoUA/VWe0rR1iWBaPSoRQKuxExdC
RM8T5mx2V37rwMUbGyYJy2jVI+vzb+m6OJpe0BJEY2s+7w+p6DI3ScUA3b1SuCFlWM+Id+xfBED8
5x1bpw4855bdfaAZxUyqsY1m6TyodOhfL9L5qXtW+8xPQLOCfN/go3DZZ0cpADjfW81WCdx5km6/
XHX4UQtggYeclitgXpbMsHvtgK8aTvlT9gH+5OgTmVv7HdxDi6CNwHSd3V8T2tArLNRyfVHXl4h3
YI2p7N4m+FWn9FQIgDieXfQZ7Wi0elj1kXUNcogS2LURp2JFnKJb1wuFk6ds7AxopMVm5nzttARS
31aOtAYj8oJA10lUfgqBBEaZzDn4ya0rupT8ETXKwcIB31I2uGg50jwiiztc4rbqVm+2RwQ4Sea8
EuhjN4Yg7bHR5TaubFtIKi06r5cdxi9IjpMogZBIJX08byfDDSt6AURqM+d6ax7jqmD6ESJ93KAr
m12LyxFFGOIMWZXjFMZPN9AuFkFxhPtodhPJS70Z3owmrj7H2KNVNL/g5xDnsrMQDtnFNBLmuqXt
Xb+04n6FZXE1RDBdceZFlsXtHPPDn/oURgCnaudUcrzp4GPguF8Inyh3zuIloM+pKz9TnLcink1s
fxrxEkwGRMl1n+vSP0TTcVesRZBugwnYlYiFHfioknPUJ9JwcJ0ueevRkZTsTVt+WVgqVPqz/awq
4MKh/fkrmkJ9AUU1GVg0aCv8yGhq9zQuM/icifGdh/nP5J/RHRLwCNpeSexMasl/3j5RNf3hl+O/
WRufxcJyDBkjzHplXeussFegza23ABGhipyPQY13WLyWh5A7E9Carr+osEflLvGHSkOycE5VoJym
Z1FZoYZc0aB04hLQ3iNuuXEFBr1LYZ+XDEwZtz2874GaaNtkChhy03uxsv2qc7OC7iOEPb0kPmQf
SekH4dFJHXQsIjLtCImmZVsiKIeFA2t0sKQCy7/cSyKU2QufW/AaEJ3O3mccnt9oLFdbCRsW+QM/
/L7pq0cbrwCPdUp7Mr83Co/BdXRgfuVEOVXwKBBmMcrc1chW6BvOXN8cegQHdt2PWdVVBwVP4a3k
WwE5Xfi+asN56AbkznpF2rL6nPTxB4AVAmSx22b76BRvmurXnJHrvIAbO3OByA+df3Wzc9SPb5zu
qto6t20Dqek1FpHyDQub/ZC6gzMqn8XRKo4IQJcqUO9MxaFDpcyQkQOFUW/hL52bXDgzN15Wf9y8
pTYbNsWBvVjWDT9e9GYZaWQFPb/IChBC7veSJNgNMCUEA2iRcfkxtqXjGTq7IL4QuiAwRVq3EU3B
SJ6FafVwSQRd2IJROx+qlvE6z1IChZMbOP05H6LhnilZSlJCM6fBDrzjX4IRBj1UjursOr0zspBM
N16LhE+9WBK5qHNtZ29v10UvQuQVXXnF67ONukhiylWmndORwEYoZhESNI2+ZwLOItNpT0btyv3H
h0iJqTg/tgcJE/SIUaLcQ+xXQnUk5cjf939whUqysFA/rIG87jx/aoQH8fVxGpKT4IlGuxt1MQ9c
Q7a4cFFwdqH4XW50NEhF1aCcGMWBMOZmZnvefEHFxL8A/ysX5SOK3xyabM4pHQfwGPM7urDGruo7
EZXnedDIRtdp2amaC2pXSA8B+U5vAJ/uqAUu/lTNtw6W4wrX5vHfLS3fi//s2MqdtpzA39T3h3Wu
pURPFL/5ab6adW7JEvK89gMeNhZ15cqpkyXJ6fzbwzdFDX1rCiHC9eIyOOEoYPCeLnQr9ePstl4T
OKHtHoF8F7QuGuOqMPOny/98TtH4g2OAAAkg0wGQtOFylx2jWfMhzvn06ubMv+SNoO2L1RUpTbDx
zKTIetRlOAKUQQ2R+cnMggjozAR0to6CI521f/AM3zT4bcMIIpCXgrpSQzugsGvFb+8ks4Hsnbpg
tShx9jxnAzscWvklpAXJk86Xa2QfzmKdZiKK0sA+4HObLisqd+KIB/HfPeL15dSkL+NzB/5gTrsB
l0cBiIDZGww7H+nouYxOubGWVNWwxWw/N4155n1OA19tdxCsZCPHfqRtIPebMpxBwVEGC/2CrR8v
qzeGhfocR2IQGjdK6ySWblSgcGLYcQjlpcoZcxAcACY9TiDmWaW37I8OPnxVwY3PDgOxJPYSvyZ4
PZcPfnjYFStRUGyrJsdQxVbRVI+ApTU2H8A4+l/BYyfIsGvZBRH9UqhmDsYsBnh2wGi/DtDUmcdh
acV0yzw0eg5sS0CK0Ktt+pe9jRuZ+eD0vxlY9Q7YZ45tDUM6nUZMk4x8PnNnYLW3azgdwglIbldW
Fcrveu5WVwZYUJGYicBf8HV2RYrPHM2rUrvWrcvbQDdlrjRHD1I/0rvQfdO8xjwu2/2VdaiqC9gk
VYFg81ufkqzN9BsREtK0uOsRxd88Ia8rfJ4k2kSOeQQ13x4DJwJtOU7n0UpItYSdp3NbJiVBqFwu
sAYENteTbHBDlUik7HMBsCu4HwCEoQY3n645idmGwOIvD6TvgK5p9ZhtA8dWw0q1dKF6BFxyFYZX
xrAc5d98eOPy8dA/Xjv/hzAtWuSwalfjiKV/Bc5VaV6QHPZwswdwj6+LUxXY4dy9snBCngwXZGiY
IooabEjO8pZHCJvgdN4ioU/pldfpUF/tSZ9aVmRC4xmT6NBliZ46goxch2kd3OVw2nWidHQbN0ai
xuDJE4AnZBlETtujxzjBd+IbK806dfUrBVQSdOpQXtiqp2BEz3dQAwStanqYB2Cyqa598lgpojOT
zjx4kbKVSyymsHI+FsVlR7ssLcl8SNcwm9IagyNsQczeTFVCivnUqr9jcx003AiAX0XBp6nIqSFd
hPZ3AR1Bc2YQyQawL4IEfbwMpyI/FOe/n+Dz3bXmTB1ku7nwPQbn2KHcBfJOZBucjV8/jBlUYtcU
pOG72hjCF4JkFAAEm8I3YfsKqSd8CpwwgmXBoqUqdD8mTg8quegWnVBIcZuhpliyoHthxxHkRUPT
hAw5AJbmt8SncJUMQ1d13pM9CRDvRBAolZyNRK5adM4l2+Ia2JV/CJNGg1cQ/7pgE5oIDnNablwO
x/ZQSCzp/rRaijqV8svh2ttUYdPXeRAuQgOPgCXdUiAKsA3ZrPX0dh3ObPN1av9B86SP69UU1l6u
W8ftEcyXkOX7kn6AU9Ik7PcKI3gN0ayWdiI9BD8umJ4deGBQ9XWR373JpdbONMWahjDdpzAAp6SN
zp0GaltuZAhNCE8K0368MAhRZ3R5/6O9hmj4fKYj54mnge2Je/MS6Kvnm8l9JvZs+w5dtryBQ0E2
U2MsM/mI2zO8F6YK+kPh8h83rJJdShjGwypn9O3LOnFKlwwYpQCkavB5cVdpLinZGVG304unFaFK
iD4pMedStDScB/rMFNoW3XiFRdLWpkVWzPPkV7JFyT9JKMqzekDvC0VMPMpWEIfhBhBbbt0aZjjk
6LpozPsuIoCHQTj5kKAygjAuq7ZePITppVZlimaweXHeDjxiB33ugBYtJYw52Kk0JAtQE6krmHhZ
2p8KLPlZXXqZ3uwpR5hy3VnyezBg69yNOhz+UEfrmnRiwVAkcmn+jvi+AttUA+jYFZomlD+iupfp
85YzqUxH8+v0kRDQ3e1pgulfplWYSA8u/vJ7s1jRMQWt1FOHpHSIvrmVyjQnWLfYAnk1FUw6zfL7
NH3rIf+o+g7hOIQct6n9Xb/eDbmzeNQVDNBT85KFgXFL/fpF82ZReiaVzPWIvpLsOEEHOCZv9dK1
S1nFbabSGv3Rrf9+F2vPgy+F3NBNO9uWPKmSQIW4e1zPI5Hsgxvbvb0b/zAJ2Cx3Tn81I5wxUM7B
YfrCIbBXOqTJ4Pnh/5LmhydCmb0isIr7ZXaWw/ICoI1oO9chbrN39IYzjE/1vRUZ/bYXRNlL7Eh/
JsC3UQt62eUlqM1fhP5/WSSVN6UgDpjkH0hmvU2W/2X6PRuJAgBwGu1+lHLrMWAAbQQh8Wh8ypTF
c634BvkTGQ0W8HclEbAS5LDFWesSNl5/6QrcfXBP3Zji6te1V11UMGNGlzIy4L3AkaFU/FVx8xe+
lJIr42A9zPnHgoKI7wfeVl12dQ7Kt0t//wNhbnyenq2uTLTRReuuQw8QgmaUAmd3mGgTGFlRhMuk
LFzZTzlup1R/7ur7YXT1WnVkq6pw8MLlTMAmTsdL9urfjy9aZe4qITGaQ5yqM2Ri5F09yNimADXU
QRA+13PKkEKVZ39eZStlEcsZHa+0UiBtwzI6w+By+vOiv5VqpjN/wmdQtxGeinT/yjvInvJwr8Ou
7HrW1iKyHhTkLxaT/XggbxwXqKOHLXmWvCAnh64K7dt9x0QGPR2R8DMclzX4dnEmZZJMxgOog0rE
2WlEp/5+IIHcDwiAt8x/WeOUyWpicwSzieRAyBqVh0mztj0aMIxG6dGT3kmtynwC3q6wzGcYXTH7
YZEvOKB7X3FaJ316X3ng23Nv/fUsdRhnLriyUSSpewNWin7IpNopN9KUnf/49tgXVkh2/fz2gut5
6KesmVQggSNOexpjofTEcvF4bY+K8i6oXNo79OHsO5inAkhdg6S8TvnVYG21LBauFF+Ko5V7QWYu
n+lO7Lgba6LVrIjtf/0vxxLEXR0U6wmDtp5YR0eaY5nIz9B8HBiwWt2BdPQ7NMW/tVMpUDwRLk4q
R1JhveAgYqWvgeTKyjxKOVbsBdQMKgWpnd1ReL4EGqf3K4tar6hkyoIb/bNFkgvW7EDiE90TzrzB
g07X0qhfQkZPosHq5pAujeSUgju9WV0jEjC/hYahp8WbzteRl9g0RjuSkm6n/j13Xavrxin4R+R8
3GVumVKfWZ3Ppj4Ylaq+fUUr7DtUqs718Y8NID7uPT8RufVSMWiufVyJQQhsO7J+gsVD+hafSdzR
xhh8lRwUEPU5MM7TYOS6l2H0vddy2I5vQvGyJq1la2OuG6+xDq/wESjZCfJIaWFYRJ7yPyULb5FU
d4Fg9gaU2pK8slbI4FAkHnmDimCTKMWnWQSFKbscocsv0iwsa8aSIWUt2Xh1Qvt0yXQbPSPGj/Ol
ximyLA/GqMlNmn5oVS/GmFFxSMrGgXI2b5iU9eY6R5vg56EkNQ4X5a1KpRl7DRj6qfe7mP5K0Es4
tEsj+2n4K/I6OKQsZIV9llUwOwRdsG1w9zRodkXJLkcU+twVy+B7GZIN/VGYn5c/zaIStj2nQJrQ
OGCB2b9k8w8s8pAZJ35hzq3GnKLzD19s52ofW2cArCPfTjFPQStgx21iIhMZE50oRyqugUtzMPh/
dTLBi6f+U1olbZMVGbS8GRmqJqtwUtx9jP+td91uLxz3NoRz1lhbjegEU+Pf59t+NTILjOJlN3NH
6gwMj3UzmL+og2cWAFfqhalVG/Usi6gdqbkovOLl1xOJUT1RHYY75p22aNiXL0WEx2xhbgm5J+R9
5xht5VV0zgNA9MHJ0oXtLGL9o+UHXhz5b4LAqQnaa+5fahedFvUD5QZkNh8B1jnSzKbaxhuvKQI3
x33vpaBnIJDOivKwOycyeqntz0efAADVCxhW6NvPUDNAzomAhLMSwF4Cw8eX8BGKRYw1v+4U+VtD
5WY95eE8Qm9OrNVGohMdN4tcPeDFaR+EcYmRJ1djnoLX/sWf7PQO5LTXqANv4zaZ3GtkDHAtfSFr
Jlb2/SI/8dKoYpJYK+NivtK8MBF4yjt2SG6T++Sq7yXgS7934KsKmfK/bpYs2SR6pF0qJgURStk7
3R0KkcFD0fgzX5ywnXAUUMlHveyWf7AZsHePblXjE/kXYa0VepAkmcdK3pBgujz6mzCoDwU0hRUB
YIXCMN4Zdt6yCQ9CcRsvu9wpbRUhrMTaLtW2NleDc3P/cyA8ch5UHUYsW1z+9yhLPAGLPD8R+dEU
pNImucWfWnhy9ctJw4rJXJ71c4IwEyFcfskaAGHP93lW7Zlkw/MZZ5+kn8TW7EmqE6s49ysiQaH0
9XbZcYY1/HkfDAiF7Kzvvr4xmI8rMXceeFOjJO4E+6fXRYT4TYc8Hvszz+FUi1xzytJ0eE9e6UEK
Zl8dzm6cSyLC9g/LgUWzCw67K7EDDfZ1BCd+7xM4W5unlBVD+ZMWRpy4A1zlk7zLVQO01LwATj8Q
El/ZrYFBEWDrNjZ3Hqb3GD0mfxGwHnIL55gg+CaoqmHbnCuyCfB9DqUu7MlM96HZa+fK9ZhN5VCY
Ghb8dcC13MO5DH6NHo5lodh+4jmi4NUx0U4VvtqJfW7r2GMvpyzWo0YzpqDUTHYNvmG3p1OFmaIg
VswVNVica1tlB1if5B3XnlwRLTA+8p8/CGSo2K4e2iA940FdZMa7d7o6ISN+DW6Kk6reYTOjR0XX
0K1JoB/mMORMzfVisBFdNuF1m93zxYik4OF56DQIzczS15VZjYdgUaU59pE/E9B+XzcQTIy+jyX7
7Fw6Nze1iJM1i3/Ae5pdz6oDAU3kqEyLq1D6w4Nk1PaNdh1ZOOjHb/D4DE2UpQrTSeTbohWhXjze
iUEXnAqVT4MglSjtfqyqUE5LVo/XSPPJyZa4faK9d7MqQKIix+vIUGgz9OeRVCo+n3yA7IPwOOkD
up/p9do5TEaEMI9vT3+GlGLmHmWnjJRRnLQuQbO6//gywlFrCIKw8wabDISdyX65tI8LtbR1xvjY
yksikRveQZIWQVUhU8uMeXxQL9jUiYqHPNiPGSvJAPSs99S+hcMc5O8z5LBpvHi1ucynvr8Xhkku
PAiXEguQ56sejyPk5pCUlCq1YC3v+lEfTw7+WRM5DuGGpm0+EjmX/IggG/sCQT3c3V3Oxyll31bE
DQfeHjRsHcKgWL28X/VWo8lmkQVyDLALdsll0mx1ZF09cM9uze4+Af7NOZr1XcJ42avEKXpANwHQ
OAcZ0KltPcy6jMfQ94UXZi3XjrOf0ODUOo1E8DW1V/r/4QcyWY6jblv+X2i7kjkl1HCktwRxXdMe
Zp728Tj2DAK0Ehl0cAryq6wUr3a88xZXkIk5xw/On//ZLhsk63aPOUhvy4D+ZOufohtcrWTiYSzm
5qKLvij1GcxLSwF3u9YlOgt66NJ1+EIXlDwYu79tHhlOjJIXx1e5nr9xeYAerXM0o3yppJZsJSVc
VBJzDBJ3N/TOLB7RveNBw9OatjQ9a+McXfGzVjrVi2WSX3JAKSH2qsDAqchdolvXYWzwmvG1E7qY
kfcqydxYdZxVoaFRQQMaqH+CPxiLTor3Fz244qQUTzdS5izba3X6Ubz5aBb5CIJpcUMt0/35NfTK
Wk1aOHbw5fTGJhuHvELFsVC5JnEvnS910IRslIgqCEszoyIoHQTlGeSrrSWajT9ZH0NU/fO96whQ
sD3VdXBvb6uh0g2DBNWqbGiucFzrToi3l3/8o4JoGtf1d1XG5pkMTUzk/0IZ2uI6WQ8zCjgEoKsJ
EWsbz705TIHZdXQEKYEKPaJuGqY3M5eSAiHomxdXdUbP8M4XWZvdMDGuNsEmQCjAtZUFmxsQUc9R
GHAl6FL5sU8vIC8HXIWet24vh4nu1pNzopOGxijEimcfVnGrfbIXwgEWK99mNymvy3tCFofzESLP
THUSWWYHQeBafgXIlvIBJO7pZNpKKuMidwzRN+ZxljfkjoTwobkJ6X9H/wvaKU+qE3gXq7k3wqtb
ReY3UiWv//FDyNGn6PMu9Z1szSSw34Psf7DBZpHK6dhGrCT/VyRKojU3rkD6vavaYtUgok8WpoyB
mZMns3PEs0BQS0YKkgj+nCG6oh4h9pRZ/hEql9MOniu1UcxpyllfZv1K8qdsggnfS8APOVRwbOzo
xxUij/yWjpRzTPyqP732NX+TvM+8EQvCbQWwlzT9BAPE09R4s+JKHkP3OooGJl34FlENvQCJqqYo
jBsW5rmp9Wdzm3vaFYzAz8HThgjMOdIO43dfX1InrpFHDiOcntbowBdfe5PGUGzs34uE27h4pRsW
Krq5cwUVAHnR5oSGGlTagLVVofKg9dZLvwtpvKiXnhVQ20OaA8JOnhI7w7NDscuUNPX7ljx9CMxg
uMgtgMY2UO+Yk1UwkNwkgGZH3DfLhBx8pzWVYs04kjfxcVrCX5nlN5qm8kwpLRo5wx+eX7x88KIA
Xe7AUpcAYfZ0dmU0gJz7W0D19Gc6V+vgZoVxe89ZN/r/PAz5m272zOTc5tgNx07ILmDyMVuukTXN
L5/4OVXAEdOnf68x15RsMKHrfYYqKsLwke1DEx0f8kRJbB0QBcI5XPl2LLEjSzs9H1tDAcXG07Y+
RLAEz2rZs3LRBHEkLVVo5PQ4guxeG1P44e1KPtWJx7dYqwr4gVPfp0zpwSVJ3ptAfETON/7yVa0K
DEw/Ci793yzookTJ9lCfyAh/RlnfNhbFv06KXjYnJs+l0x2Bf1xYuT/4Qo3ZFLRhni86tx8W2v97
4bQaDHYvDLqQQx5yAZHLU/zs/7P1kmv8bPRH4saMm/gQXK6bmxxyZzgWLPBbepen8tTIpk2bsJcl
Sn5na4UzL3bJe3ykvdreEBJ+SbmcB0IIpc767Gb2PBFu4E8dP1l9HktpShkUPeZVQcZKpic82pfQ
Z2IApnFG5I9R4vK7nsfdq4TMWImRpGvzIa+92VtH50ACJNKpQRtFLwrdWcRutiqaR00CkGTCB4Vy
actPZqktiGEYxKDnkhb8rhCBcwHw48L8E80Jt9/V0sLPuM3pDk1WCQ2DtOigSMYa3rXu+mJf+tob
EvYlIQvSVeDDvEMjCZyy5s2q2F0vTBaSnL/WmBgxTNQpbbDVzqK0RqnXI735/RjsGFOQoWN63DRo
E/UzpCQoFk3A11GxK3K1NViQqe2Gqxcw+FezSEiXyXVj5DkYI3twBCJMlUuCCkonfi2fWdlrElKO
ioftTFqS4fCN5FbzJiH/DhP/SPFteQPMFvEk3NSbdyhJlFNncjDKCat1soxhqCAMpNJpIsf+o9RB
dPF/DGAEz2DB0t5X0nY8MHwyuNJkm/AG6cLwu6DYucdLJbCWf5wkBE1ArsWdgVeVj7cO8Yvw35rj
THEowdiMegXBxq/AIaEqpgsM4lTjMXWWKCCwzwwsw+SAILjlZMcIZpRkMaG+wvPOG3BYrBHUFU4l
y206rSpjH1o7vOknOLidhbhXSNMJingtH1VWm9MRdYZv59KSLJL69R6kVtUw7pZ9eJmeKFjfW1gf
3FusVXz2MHFVU4xLFVIdgwXXSPcHVu8zXocB9ueZve7e66ngFy2AarLt3rj/J6FQfNJEy+rpPe7R
bcybK+nDDg4/iBuV5uGOPuNYMnfd/2UWaYLRiHhH5gdRqbGKppsd4b+ZAdEo0zgc9a1a4xe3ypOO
1+EXWzx35PBjNK2xjN2qAuQqiDi1mCGK7f12ADT8JOHFVM2gB7Qi0jvqT2XB6T9qZScNxzwZDuff
lr0Qz6Q5+Xu9aKG6PgqP3HfUP2pRRkMywEThmiMOEc84T5UiWtBpYiblUaICeeldRvlO0b9ttc9e
Wcbv2xHBFIqaFmFDACfFGECjFXfsSF72gy/+MzF7oxrTBhxDjd3QphR5bvRg9814I+GabnJpo4HD
dceTYkpHnahPV9K6vhOteQroN8oixvKYSvh1eYXr/+1Auj8vcG0PXUDKItA3yRYlFFK98iJySaQn
Tck0T/q0iGRvSlEPJoi9LZJYMaIOh1uedjNek/VVOCHNcIEG+nH60XSYt286qOGj/U32vnDev6/F
CaBD+8Zqs7eW9qJdhbtmC6Jr3HRSGx/rdKEXUS/bfltOdpL9gcgbIF4nzP26+jtSEu/t/UJOga5A
qKn010VMeaUaeAdVzlpvtqfxhQft6f5Eb3Ai1Fz3k8ZcUw5/o8rIzkPOIreK8xlS7lBF/9uuY892
Ohn9FzdksTNk5csLKe41Q5ksAkBxFiSICYNCEvBBm6a37aBZ8xXcaFgRBmbVOonJ/gUx0lHSUe5N
D63EljgAukuGPBrbwVrdkGXSfvLwwKGvYxF1FOuHNmzXTXc1YcvYWsBzdryAJB15Mn0pR8f+48Bi
dTKDgEa6K6Kfov6ItjvpFH8gXmuygHBKFvvOscTTHxFU6OmF5fM+gaSLzbQ7VrQFXks9H5D6rRzM
vuMUIF75GunlZtJ7zFaJVePJNTByKRQ7le5tKZO/wLpi0bxbL3g6yftObpfts/I947w7CEFhUl7o
CK8M4n3MwXuu1mbvyDbSaJ5jfg1Ah3GeujRjaR/jBb7mdDuLDAUz2cxcmD4aXZuYl1Q4BwPn7t+B
6o1yxqbK2HYgdwIMQD8yag51eSvBS/ClZCqor0wkDrV+87Yedp4cUkCU/YSX08Sw5nAE5QJYWb5j
UlTJK7KVlyUKltV98VLaCkWB5RNZlimVP+Ghl4XJK5JHd2uPLUrBkBUN4PAW9cHrge6TqinfvY/K
ODrIkKcrYiOQT2oZxptsuFRsBLw3kmuvjDYLslR3VOJi3m+sgMFcSCWR+RWEgxNKGgCxf5RC5fPO
R7SjO+8jdxE/Jnpigzfb6vGJKxBvtSksHnD5URcUUI09k+BUGaXKfrfvoEyqQSjWLiYdULGJF55h
lYIXd+Hz2z3GCzHWg3j1W1btx3v2BjNFQ5e44ktzbKwYQjUJ6dpbJFXGxJMZPnP8UbYDBsZwHw/d
TiDAkuwdF/HzqBgHic2Ed+GVGyB5DK5qTc/e6fvGHValF3TLoAR40Gym/Akb8XCsUIpb/9OHWUSY
IEx07ldEbJfIfgLcgUSXUnTKFzCcrBnopC28kF9A5oNopwbCb3YmB8hOaztD8oPU5CYDdbgO8VZO
iA5Re0t2POF3wMPYqAPnSztEB1xMowhkHgRq8oVol31sJW8ztqF4ds0SYF93BiKGKopTTThmB/Hn
l4EXzJ9z9fki0FXSeMqE/C7z4qqMz2rlQX27xsoslxGpBQ4CAz2pPaUZ1HnVPNtjYWpJOMbXKD4O
CN2XNjagOJ58Q+YQAjELEtsL6aQoUHBM8WxDdn3uTObnR//27DMvA/LwGjXRSX5FQcXOBYf2BGU7
ukvaE+AJwEAuzWRRatRDcZc5rT2q+ekLDR0hhXz8AcwakJPw5hzJZMKqEF9K6oO1SIakLdJXt22o
6veLR+4YKHg6xuhgwN8uBaUnRt0b1fkF+6SIi7k1vQAMSzhdyudLFC2PUvDBSwWL+5aVj3piG5y8
jMGSfIVn390TwTdwz1ufBRMlxqPAHTJb2qImd66vmU7aOkqlBaKLt0HiCOMP0mQXmjaoDEBOXg75
u6WRmQiwwSN1FjwDug56elm/cXSLSm/2f/TakMdsMlJ2yV9FbrwzcyiG1O9v6tdAKBY7oWDkaktD
jbWOpd6453LMQjD19gL2OEUkIoDOUARi/RwbqW7L6cFHva13CZlpPSe983GjCbq9yZ5RofyFVQ/V
aKQ2SEtPnLH6ol8d75uEk9i2/B/9ifSwQ51yQXRtVVbr0LYpRr22BtK5HCmjhKwIUB+BoCK1V+sq
BPairMqYq/STSmkuhsTjL80zMT9P9yCkBFhi+1jq+FZKUQjXrXT4o42ixs0Vx2ofevBVN5p38U4c
xQ7sc2SIqq5xZI+YUNbuUp9z8qpc2cmbQoFUNEgjGarAeFBZm+Tj3bK8tY0x0oGFccCF3guJwhnH
LCGU+tSLFgDswah5NAYbMfhwyj29E6Adtsb6MtkL6n6VIHEiezuBZNFs2uUjW3bEUVfho5oMWK4I
oVTh1Wc3+ti+pBMg5p6xA1m/8cuJ2vUPu3a9rABghpJAdNTqEaAXgUAXTWlGaMwollXex5yWDR2W
j15zSrOBdJuhsklgzlKaHwC63Ke9T0Olcp/ivcMRf2N2tKjwTpejVfXiPKSAI8PE3lka2AJf9aqU
9u+G34stF6UfP16GYUgXFsacwz55rUCvQ9DAZC264jpi5B8TtJYPSrcGL0e7i7vt0irXkdIUlCF6
gVIGG9Gllx+BRZ9tB+HiSmE9CJYaonsSFCGaUdqDgW/api2juouv/KkFlDJRAwn8XujiAk23xPCP
cNQUqdn0q+P3oHtmng6w54AK8Tk0vbU4XbaPDNkPhHsXg6FYlKLqjPq8F5ENCHSeiXuwM92Y6u+J
FlXVAdkuqDFtuDTVLCiOknGOA3XQuOQs2fxCiHzmPYcgElBctkqamt4EWIVs2PrpX/XzEzk3K1Jm
blErR37HZZmtyKC1BYFDcn1vzY6B6WtcIhLTDUtym1etWr+TCrfvxgMq42h9zyEaSF5/v2QuSTVj
rzUbPb2/SJJlN2eOhSG4yW/aFpVxbPJyor+8QjZmMhcuGoKIZiI6NeisAkC7lz/uIVKvPLBB515Y
tyNpV/+IsVkRiU5lHC/oDf6qqKQtMnUD3HI9rKKsQ0HLqmCfrs77xQDpLMlzS7Li/Tunf2GM1yj8
jzMUzz6YIEErDuIzMWUvDXQ/kCsTZ8wz2C1lunkBhyH1OeFaCZ31GXoqziL1U70SukvdhUYVmjT+
JG+4i3VIJdqbqVr3cttxt8PmhvzDAJMlEZkPT37bbvVHzMypzbVyIwXcv18iSjNfYFed/rJmHAVO
fZJlqbQfc+4YcOQtXZqeIYJvNIPF+WK1ZPi9hAunBMgBui/q5SxdtA8/WRFGN2RIlRjh2LT9hxP5
8hpWPg7Sl365dDE07TFvwjkWMzMEdtX2QlReo3jE8Z4W8bPjpXSKY311l1KRJgiHuGmux5k4tyGM
trucf1R8JTm2arWfZ8bSYJyKC6Pjtsd0pSerXxxUwoMM/ljiBZx3IQmKtn6oA83bVtJI0mR9CqwT
Z2JVbrCZWxuPjIcSe1NypHhuIpJwccWAlVlpqMO9gk58fcUWW/rIUuF654KKtmWxklNTuqRUZ0wP
DPIc9WOmskvbmfb1d3TbqfBElc0UeysD1DlA0YWFZ0SYCPFt7CI+mVkKpklPB35G14e6W6xEOa9+
+PzSyIwvExVpKDa+1Gnf1LqtS3aeROc2EJNOpmFtTkrXdlzZqqkSlqOQWk4NaT/H0tuUPD1Q4V+C
8hKgqkHvDq/yudcXZXD8Gu3MQdRk8H51djNWIBthx4cpurC6x4h/0cKz2R3C8qzoOe2uTS3hKTdE
5HfJNCjyDGtTe+UH7ZLeMslkhYf/PQ1pyWYSzaZ2XzrEBegk9Jvo83c04864dZrwFIfSyULCv2a4
yPkYwh5JRYO4q6CwvbKhnqjyJCOh83A82CgDGtcqOZYRlBDfEpI3qiYgU6b7De+nuRNiQDNmmWRV
9FNA5O+dZhnuedVdP2C6izCYvmNGMcsHKePPr2bpWT4Jb663qSV2F+na/9gjAd9pfNxwzEW/XW5p
TzlTYDNO2Gsha+XenF/caB2E9us8GHbiXzURf8iG5E0qzkbHHtFQwZJhQiJhBm0MMjukKD9LbsKD
clNBPoVBoF0Gqsb983Tx4OsSmif8IZ/fAeM/fDjbqO5T4OQLrrsGevMqPZE0lJCFOjx+N/Pf9AqX
uR0tv/SZstualUGV80z60pk/UszwLU1ElY0GSoKK7NbTWdTghYtqbR+EtSe7sJhYSTbdzs2u8XqC
4+rUDHQf2MgzkF0SZRJnbDuVdGRow1lAP53nzGP3ahWTV/5VRUYWChXGrz3p7/tISvhmZrDwHF4r
3SEFBia2V19BA1rcK6LlaDR1FYxV9LaQZlNLqfAx+W0O3OKwPwdQj6I/PCpIGn8qXFX5wNinP/xZ
YWDhEzSgc2R9qSOfC3vOHVw30IJfLsX/JbEZWN7EPI2iRcgWx/6nhuGWolcRheWlp/RnV79Q8hWP
DmgQJaH6HvPLVEfMZZF+XFIAIAIO4geSl1DeIeeowK6dV2uUuPqAv55qDB9o860v8kmC+yUCYwPj
pa1HsGRBLtMor9CARmq9mhufhHEG9adbGITQxdK5kSiqQoRuflI5U7cJccC/Fw+n1tF3FqYP9c7M
Ej/rzWdTygc1nzRDD0lCaHWioTQXPzEFU8W11b/0SglCcavG/8SwfLnX3ik/tV2jUFyG0dg4Nd7M
w7PkMNErkiutn0LBujTadY9QI7YvvF8hSQLfpqz7D6LPyxHmJLmd7oA3fmkpIl5Fk1s8ZlKc+P+E
5wwgO2Ck4OwEgqvOOkzdSx7i5Vd8co1Nhggq53uFOoULehsTk2BJcvB8lvQBSQqet7VfkPkIcATt
WEx9XlFFQlTWu4lBJ2bJ4TZbwprTXh2Ge2TWsGjIk/eoUnIODdtTKhuiCfOZ1wpwzXGJE4XV2YNv
LyzZE+3eBi0O+Xrp1TZoIytgkE8PmvTqWyUOHkle6G9G0/RntWEYzz99ipmnD4p1sAZC9PPPw3tw
N6+HnClOBStBQMaptsbPpfCjBTgZP4VJePud/TKKnyyvrvOcj11jTv3ggkYseGaKMFYatIw3QMsn
vjsYj3LOZGVlzuC9dLx7YN+9EOIQn5DHDKbaUtlo/lak++5a6SAISQRrx5b1z/YnRVowl+AhtI6N
A0UP02/jr8lMXULLoYRTuTnbLqur4Icv9i3niQWaZhwzwDRqV+64TaR58soK9DrVs2C9MaB84qwr
fTOypdRpW09IfStOguWnLYOkMqS1MiPEQYLA4e+au/fuJtnraoZ0/traDVF8FttJ3+g8+WvUZctY
d0DjVoyRtDGKxzLsfsZA70tfvujqRCWSsC0r8pZWPtDdPKhSVypk3m7h5IdOqWopnwDIyYLHerj2
mEPQJ0SD5sqqZpO62GIkqCXd/KGSefenZJB4JYJiS2C0XrPrHCxkyPYQkD9KCXIgcupdCYtyR6U2
eW7Y3WWUlurUsMFyWvEJEgMni9n9dw092p9Cmba9uDioernRy02pgp2ZrKTqWnBIHsYOTKA4Y35d
f+/XbZco5rdZoJqEyNc5s877q4aPEAT9ZaKOlsruTDn0kPO4956btROMTKfCuKS4AiwqiOS18/DV
lkTPG+/wfEbzWPMVNkV5qHH4MoWFd3tdcL4YRJ7Ox2MNFNx47/eRK5aKm5pMNHAwVhO/O6rzjLeY
zU5xRYcqqAICu92tjuaLPs+RDMll7u0YJ7ZZqYzTfxm6/O89LBpXaN7cwGcEEJobD8qaAajiTwTb
TVPk4lr+lA7SWJfL6cG514B2Cjum5zVddynPsxBCgh0K8r48dH5rwtlqcw7cLC1cKqQhOH7OYehK
f2dQDIwYkuVG8FBTIOma6viRBRdF6Wp1S20HcLZIEv+csHWjWu/C1wl1YrejrtUBo55iI4x7T0HT
DysE8beFqbwE7rzvEWSd8QU7FuBXxhK6hWF63hdKasXHZs2eRlpYKfHDmE4jGin3xezB6AqYqYKK
jTGZz9dlFARAphoDT8wTnwuFLTWJ46JbuaP7dHAz6qgPyx6Z50gPhBqTOJ45eHqMEdC8FEYY20SN
9ErcuDh+zrbN1XcrAFzTWw289ZO+HHeVg3T4AZahDLdAt1q9Q6U7A9Hxnb4FcUY7Yd72hdro71oa
B0HfKNXm/9YwagwWNbU/A/QVCxh2AswUPVL8gSHpJLspfo1jNA2SVfArVRWqDIVtbA3AiCtdevB9
vviQcABg74yKBEglOHiLafWWHcgyE21Wwl2tW1GzXdYmFgOL7ngzbJ4niGFoBCEHWI9aRERqpnl0
IUI0UXWq4p9PJB6aZG8GeAD3dFcTy2eAOhsO+DN3h981RfWHdXn6/EDIicCHYsiDb8kP0WQXqfYo
fHRmSg1NOJeKG0pa/X7HQV515rfgmkOo9jpiqr61ZxWLcR4AY/D1g2xbII4zUQ42z+A4Ao81PbLB
B7ISF2ogT7mhZ0eZ7X1t3jkmWg0nnLbn1pp8GHT4ZH6A8LaMKuB3Zj0MmDWaQyRO/q6dJL7IiRRL
FIELZlJXTtncgMBnNu0wvS8qckAucDT8qdI9G2SH7dETxkZZiMYKsJjyH6Tt4kdvCvTdjg/WbZa6
pWfK4QjV3WapyuXxHMppfWceXzLAOnXGWvTppLMwULx3AyuXp1/vipURpyxeD2Emjvf5ibdNHeUw
2oArxpMzf3KD9faFCybK1RxB6IEOkW9dtFVt00M9jCmTp7/9n9+9c4UCx14jsd8sdLIF2KTA8vdx
PU18TWnM0ezxGGt1YqbXagmCleti4DOboNL9ezvvFnVwZaOSLBUP0fkbPAq20w2u8Z+trCypg+Ec
K/uBl4aj7MBlXXFvOqaCYX89tHAA2xu9dnCeS55aEWwm0oOVcAFg5oT/HrL53BlyuayDp8/uEjkG
ulu7N6grDCOd9uGWNCXlI12WVUKD7WEQNEJAeRpYkzNhG5S5Uylw6KAf9gaQVECvBuJoP+aabnC5
Kdeo1C4ItvjjlIUoa5KMbTDiqFKvXS/ByeRmlR3Lmlrw89bU9QayyKa3ekVifOIFnv5dWiNLFV96
qAzvrbteuVvgLXZSrW4mdrVVqrepuGSq9LMmwi4BaJJ+geVVvH/8rF9+Jm7GqoorFMUwfO3Kp87X
xaABSDCwT5YkMuL+1vor56SrhoUuwKxEmVTJ273B3l804XZEyUvlS9MCwq//IzBF6s2J0DODFbx7
egE2WTKwtWKZkhVU7Rq1eITmvwE6N3spU2A5MyxMaYpOYQ+4X+51RcQ5B8FgX6acLucY/wBBJa/r
Ip+0d8A63uT7mEmAbBmsNxzuTGW47dD6n/8iqIHlmT+qxz1mTlbnV9hW6OIYYL4jR8oLJjoNIs6E
O0Vcet/+q5hPp3q4z5xAqdABAlHcy7X2XwFaq3YxZektymZ3K2tB0UsM6Y+1gAKCc+Tn7aCVVM7t
8OWrfzEY9drS0rXO+JX7jecFYgboVM6p26zKuxaBFwhKlLuoz0N27cRq1AVLYjsbLMLoas5VjGGu
Kpm3eXO4EmZryMmCNWxPUn/udhjX1XVD2C3ck6JNO/u0OeqV9vdudtVOj+WoTxguxiTV0uvLWZcZ
1TJDAUonlqxg52ekuQnRdt0qtfsKNXAx+fl8qXkqlg1dYvvbG0S3WasE3Dxrmt4orJX1M7jn1VIL
vAXLuWAoyqV9BGVC5+E7PQ4fqnCTvErHkz3ltM8czaLjy7zilSjtAt7K2l8bxxZn0+wRV8XnNq57
Oq8wr21gxMnSUfXtPry+oZyGkA9qRrRJbX7Qjj1QGP/xfTzVMPMcpQJGFkE/0NwELogkdNSiTtlx
Pk2kV+FPnNOYZWaX4sxBwkjJJg18d0w7ynwNC4MwY2hy6P1paZUS/w3QI29mGmwx9r35evpw/Ak1
bibb0iXAejG68ZspuuPxS8BoaSIwYhBrZ7q1DgzE5APDeDCxjJ7ATlopterFMkxrOzwkz5TN2z9U
sd6fojWdw7WnpCPXHKy9znuhJZbYNTSf4mDJafoHLWX9oXASuwwgdGmW2pSlHksZ7hnromVHPjEq
R2xp6gBOsGbQBw6Zk0AnECOz+BlsNDhtKKBnpcY+/ScDHe1+4XpphWcPeRy0a7AtlHr/z4kygQrm
5xu5yNrtJSEvVMW31qZjrF4yTgznBu9/vXGpk4Po6Up/bjIFr3r5Ha/sc++3grbpeZ69Mz3Z60Dy
HmtFp0kRvQpW05Q1EscBAYgAeXutkkuipfUKACtsmVi4k/Jwqy89gGpbXYhp2/DFLvrHGKdLQxzZ
SUsJEAzITzR17t9/fCTMbNm5t1mIZv46Fg12RXcQx1esiC6IZR6e87czzWeZEJE5zWij06+u9JFH
FUkRihCSmfMiHOpScLufI18cgfbTH3Jk/z/BqbcWydnIea0T8scMJYIT9kyQxulpzXACgkEXHQ/e
0dQDxVMFCb3gwwLku1BI/e8ITiW3nzhU1GIgNV5/9mYryBWJZcUhEkpCWdywJhKLohnzfhEVlact
OisWMBWKyXvbBx5KdBMFb+jVPaDGUtMvMNjAltfouIq1YhGKS5PkE3vO3eKl2hP7fr8G2wHIL3vX
KMred3/u0yURfg8FH2p7W5nDxendHGecOANIUkOCegqcDkXGfRuApkKw6/zTtjzlglhA8Bi507Ci
7eYSIDtD42+wmu79WLWeygRYJnuDgMsV4PFjkepicypvhLdmpMbM68zXYvnSknayzSK5HcTG84ex
Bbp80QvJ6Lfk1bLM1kkKQrrJoR7buO/nYmuiYYlTI27hsDhCVTu++kh37ymmBHxJQ9pS5EnDHk4e
UMZF771M+IDx+BdvhqEShuqWssyXHGHmZsP2kK4E4FOdJH/yffy7Q7ZlFZnSVOEtbd/8SjOwVbT4
MdKKo2B/xmQrcH/nxzYfia2UXIdbwZBzyObUWH5vZWazJYWjZrqxlMHAkg5YU9QSYABogksZV+/P
H/fXx4jbqlWSx1D2dAzkRgiRh7xuNHuUcVcj1WULNZXo2z5aWQWmHRbeQ2Ppzcgvf6gZ/K/ZN8Rm
Ovn/qhsNw1Ludpq9bmIDrhPp1yDrNqrnmsWkb7WvUwvupTN57Lt/cIhgrHfP70PWoh6q7OXrICU6
C0Lbm3cnk4lxwncKJPE1QZDWg2p9vcqLu1m+pt7A5+0IGlUsN0OPI9Nt8TN0JlFFXS6RK4p+P+4r
JT5fENt3QsYrv+hN5QRqDtmxsuO0ytrx8vkKBsnGqc4mU4cdSw7yfHczSeqktREqHefg385XWKVJ
DSZvK5rtIT7Sp5UJtmM4H5LeOtiWuntMTfBv5PkaO/v/CaYKjhfGW2L0a0qOPOTgtmdFUFOvj+9l
13kg73VoQoqB87r7Pf/5r6lTvXuIWTNnkynnPPPoGBlww84xCXepcmvcfTfkwUpLKfnNbW73ndPc
KpbYfkFE1fTFVQo3heRTRNRj67XQtQ/IPhWF5riWEP0uOKegPfailFe0KaDlwCqevjT42kPwUKjK
d6AC9SQ5gAcW3Ugmr/jA0R0BvTd178UiNH8y6kJEsIPZQcU+lrGcMveeL3Jhx4Z7opa/pDEzt4qS
DjgEWrcxXs04FWjz7F+YT/uvaw4b9MRGwqgClazxx+5NpUqDnp9LJSP9TmwY01djgW2c4edyo3br
UoRrpsX8HFyLL+MKh66bcqvZ5VbWAYMgSKw5ZEao61mkjFsJaqGStM80WHHhquFPSpmrSNk0MrQy
wLhZElLCthkK0eyQaGUtiSl/IDXMDmGdLZAK92S7uHUdbgkjk8qiDL5HQa5sy+zcte/ZuRxBRvVs
QvesMOGwo7I5UaEEDKXPVwufqO/aZsH6yoWLQJrTMeSioc98ZnucUCnpLPrA09mGTvNUfkE2W4l0
c51kCDBwT/C2nRwvR/ob6vhv7f5j6mQUwJacodyIb17css4YM6DCvD8sMsXLBAgESu2cT2ayE+E2
YwcuzTSXM69nhIfdMGg6dzHUCJNLvRw2E08BqgFOdlZf8bNH+ZZB4xbnfChJHt2qZtVlVwP6ErwF
IJ4jXQhIfpSjaXOfb3e8ziYpEBEL7m50LbWMlyrFeAneN7iDl0+o/MYHC5FTCC4vv9ZnSyfP0xTK
mbhdWyjl2CM2ByujfjyL984HPCMUjOSonRk+M1t8jReVvfgJU+cNM2CzbOu/HhFhLE/ItBiplm8/
6QKJ3osTjBZLmyW8PI4OazdbiYMjVWyJN0Ydl36mOUZ8CIRpeqKebg/WSE8TQ5Wy6H4Ffym1Shc8
t/t3yBYZ6BRlK+tQTvwqUK7BrElM63o+Ag1L52j/WIh4gkJM7T5uTTYSy1j7v5g6z7Irx/xOWlMp
3EPK4LEUTkS4XnDJ2n8UpilRR2ZMjE4M5hmTg1VLeRG/XWIy4IoPGSj03QxV5txX95vrwZZIszpt
sASuECalBQO03K6oDoO35pdoVMNf2pTTZWmUmL0pgg28Xf251UFNh4gvvPT1M8PwvsaAZ97xL66F
6LZfM8Ww8l5udIdRCJMLPhXmakadoHWeLAyPyfF9npAR6ONg/Wjj985tUnr1xcKSy/W3duzK0nCb
Xq3rQPXIQ+dRQG/cIOaFMt2kIhvBX1algA9KqewlBLXF+f4L9ualQyLo2KgIGOXfWBYS+qmVtwFZ
2ZPNIZQCUr84wbjB7/2lwRS/xl6c66bxXYnhihOc1t2jSn48WQU3N7ux1Uda1O7s6UL8KKDJRNKG
9RyABQQaU6ENGR/4C4jEjPClOqgcoanB7gLGzYUMl19Nj/vghM/FHrVmbrGJ1DEXvf23eBjPT+/q
xi2NeSesEzwgEfluOE0PBM+2k0sCrlfPpnm/g37xS0s6a+k2uiLr17YjAPCcbXZwUqrMYFpnAP4H
IlX/prp/Ke8cSBHmL/uDkEZUSav7Tiq6oyGSpRTW19+QEJm+/QUziI7jrTbKth4WZVdlg9iaiA/b
febGRqoZYzW8LF4Ej0aqNtIvxF5zVtsvFiwtNB0DH95XP0ebjv3O6nytboBKqYncCA4vMXTUSf7V
dBLF7+nuw69fXfxKBy/g57dtE3dks3mtbc/2id6bZ73fLt4Mc5CvOhdtEavnfBXr6G6COVrVEEW9
r1s1a5NTnuM2irFJMo1OxHU+afjIPaFhgz4Rr2e5fXL0Z3nAEkK2YUCUmvxm5yTLlCYfLzrpIr27
qVImYfzdtjHbyh1k/qKXSYgyzIj74zHAwy244fbx7ytKeBOgjpRysiKv4UfpDz/ioUplEF/6ks4v
Tx6CZJERLWHo6q7XcN+F2yxTkB38oN12OBbu1gNSE6agtKNdbpFppOq52aVA3UDLT6Qpg/Gg6m3O
NG1Ey9D41k0JdmE5GjZHRwR9ndYWkfs6RRUtjSDIMklYSQa9V/b+NvmuoqhMnOB47WIFGvSOq5AX
lwrpKiCS9lD3DuDQhQD+9+kON9DMY4D3HrM0RH5HuiP6Kt4z/fG16+nkP9RIScEc4me881CR24f0
XCMVYnMoxQpJdq8905JBJX4XYXtbgDYke0Xm5GvBV6UUN3YgHXkAu80kaCjvJCV8NOTdOqt/qJmX
OvmD7PdbeOfT7DKcfvKI4kMgdHUNxMoTN5Lr6+0Uriy9m5nLzWAkxZiUVGC12maQ3dD5s8XCywoD
Hjg4ywDZ7Jz6X/g7bG7vNEP/tSMQc5/g43bbZZq8Th/qfbJuJBatwgpXVBJ3ywoQ5qu2xccfbmro
JtKe88+s4oR9+QoCkcP8oS7PNg+SGYqDyXRNHy/xXRprBjLxOm8uv16NWGMERHL61d3HsyvoDT2y
b9RdmIKj5pwQaEeBoxpf3d9gwDshKMwpvJtwBjrPFWdG3wESDD7QK/cY1+UQtZcn6RhCAP/dUaVZ
OYi/JyCSQIDb+KyDnV+VwkcRLKMb+EYkzcBhlzKeYRjmm/VSR1wG+wkxU150J4ebRtcjzMaolcp5
ygDYzuPrX0VbZMgbeHsgqIdDZdLX2vmqczwFZtc2bW2bqnuCIcEZtkIsph+EoDlzG6j79GcNnyIP
Cmp2u231vtAxW1EnEpN73pjQWhL2kI8yQox4/gTeGyMM90Ah21E3yixLc/rfjlD6/BSV+Ek2NePL
3SvvnSTixDOLj4EAW6wtsdpFQ+gYaIR8DwJLt3cMxZdnrnaQzmpTS0C0Q+cozdK5QT3vy+rvzxCP
Ig6sZihkJmtZoVUPmkAqBKyE0g6ERNVtiYclrqa/UtSqTBKcGOrjnro6tp73r3fmgbV447by4VAQ
Ba1xHQCr5d04pTX+t1ZJlphFyOfWb0c8GmaRA0LLvVzBQBQSXt29hdeP7ZXa+JHmNB2dobcygxSX
BSSxkdbo4yZ19ShRdCDQkUd1fudwGha0p8wc6op/rQUem2ZKz4iaW/1eIwwzTaDrQhIG9RzDdiiF
shM5MGTMck7d/stryKNROdlbHsDybPZn0nIMazhp9zLOVtfdKzZJV0V9+oUyrIJ7Gcu8035kmlBe
ntkoXwtp5dOslif66s4acK0UmsID8dKKKNOH04T+P4GCj0oZffPLWUTCEhzck9WYlD/P5JdzMoJC
qqOZ54RXMsN7JklrwxxDZJlFmjagevtTdfNKI/PWWmduChCkXvMuJxC82Pk3ugd2FmKd/jlEFVTf
aEzHKzJcAV9Y2HvZqe3gokOd7U5iuAn270/eMxV2hEsg3sjfKSp4/9y25Ejvib+uUqVtxsEJvtIh
NncWWWQYZYOoYPfxFNlQHv+jXcmfT25GK70TCYSYl7O16N5QGb4baEeT2UgZKGJo9Q2OUOvxciGX
5TyRqpRqvjFLxvemYmx04K7UDa9rArAeXTB3K40wayhSqD3iiJ9K7XnGUyIhL3qqCNNtSFrQFqEx
/19M4sXXP4wUJBZXNixeMXsrlXzS3KlFlwbX8kcsRry05NAltqqlTd2sfv7UGulk/662IX8iqBBc
j9TUQy2ccNF4v43GnicK2+9BgRDV+qmZ9rxGrcY58zBzP0z5TYc7EYWTbAnlMH10eYCAzM87srFB
w/uvnjFHaYI+cbVJXzAR8IeWvh5eH/JcROnaIIh1wTo123J0nL9tyHXjdKPiq0HIhWhhEQ3ddcgT
Il9c/PJtEWmyeuh7Yg5t+Qkw8VaLQGA+QnqP30/4wMrb6Qe/pXjKuZUZ0X16ltHi6uGTzhe0sdYi
PypjTLG6sHJ78w5UIk+os3Olf7y55Mig0dnlZDHx4fQNjJeWEO6w75Y1/FQ9a1DxpuyFMVU0L3HS
sa3SxFZRe46HyAhW9mYPQ7k7xPWrVflN3CRmzjTgU4vgL1RV7QF3fYlDWlpiqVGg8Zk/qiLxxrEL
fPY4WYw4ep7L+BU+D8rrHwAVR9qYkvFuVBkD7rSPT6Mp/zmvXbqNt9cnuUZs2FQK6opqg/W9kz5f
p4t8ko3PGnvvujT7B9P3Lw+o3MXSyLWVlUM/f2/gLbVx0S0aA7/eSUHNPFDgQoM5j7RahEFMPLBr
PCxlgTbVdBGM7ser3Ksye1WxZZp5JOT1jKDO/X+p2msVk3rfolATuTJY60Nfs4rWP9VdOba+ueBF
10ss9sIMd7ZQ7z8BCmba6rFVfj2teOoH7/6XGIaU5PkOO4ALBnN9awfSDlw1OxALUfvIB59Q9UiZ
+IdKVd/wr2Vfr1SXoX1hWePi7PMeNnUqFL3GXOeCCXoybZm37ZmUSvt2f7e5D8mjvD9alDTgm58G
ytPhnsm4TwL1vSjrWlfCU/IQea08kiHFwC05Jd2EOduO1D2nJcYfUi0a552NumSacENEpRc0Qk5i
r4PeM5mS+cW+3x8Cbv9LpUqNzasLCc1mUAK2LrbBgWOY6a/6rOdlASU+XQ0ni50zYrKVRms/VeWF
coXCX6/ALe00QEyQGIPCWdEmtbAQnQEM9EdCKb7da2IWT6kCZP+Dd8v1FxMThQxLbN0zhkPX4/4N
z5j/1+0D7a+F6mS1xQMWKDXwcFeMh4H+pG+zThrm8B76FAQ/15XJnEOk+QtwAFCQGgoQZV18eJEa
DNEmmTayBWLQXJ6stiOHYg3MyiuhsPQL/6DIsS6qVpHkv6aciCRAiwgyStoUeo9TxO90V6MTzp5Q
aEgRPEwup0CuW55nn5+1YCDdF0K0qW70yqQY3m0niNCYLof6fSkv3OcRuwTMxFUy89oTXe9a2lT5
JKVVr4ngd9h2f3fnp1DC/iyEeFfC0qPkEJxEsvagWwjwZnXOK7kskF/3WLfyMBTVwd75ioKM3YyT
AWdp1sK2ZvktpHwhHevXRdXzpEjIkLtEzHoVsQB3R0UNu+Gc+YVGCE7YK4yu8l7V0pgqQhyHyygU
Q3zse+zEWWUZL32tfp4WIhujxQkG60ZFZYpIGtrpdeG7YavBVJNh9SjfleDj9WLkcHkL7EelC7Kl
lfLaZrXxZbX2KNvpQ9XKqp6CneFS0rwWfW3HybblXCoNUnnK3Kpsht7lBVDT+WvpggiGsWv8aJR4
84tO7TDocQ7KCQoJ59fAh7a6v9G4iN0kM6jganBA7cKzz/GepZGGL2Y7lsLHaMtLsj4eWWt8GgLp
2Z3JNwNc3u+43kKaPmVGj7kk7AdGn8J+CTjtKfneo4bdOfxWoyCiDPXFdRNhGq2NiiPZY8indphj
V/eSXkPxlPTQ54jE4/EV19AyhcGfD5k4/N7OBT02+rWNv8wVLd/AAGavlqosuBdUWrwnCQ+b8Srw
CayV8umuaSQ2Wbis7Y1iv3fyab+Xh+XLLwQxcbRtZ58vcwwUNPZimbe7c5sR0NR9QA3TMOjJnLkl
8bJxEHUqgK7VlYMjUN3QO+jTDSzDSnsY08TzOxQCC/NEPb6DHFDQXc21pKtW00cS8sJmwNDW/QsC
VzkZrXqAedGZWa9imj+WTHb3uyaP4hp+d6mXI/5TSn1oN24F+iCvmV4dhxL4ynnSJDqzEPvTz+++
k2xqai1duR+zcWv21gBh2sXyluEI0eZlf7zwiaQXhAs5/6BIDkWgG6JNel/318mCsCGn71Hifwnz
MpPXL8i3CIIglAQlJ+42fdVJYOdc7unnZE9wA+8KwNbfk10DiNvNo5mEnQFLgpSZIyQ3gg7YzUaf
cLr4XGZTQHNVkm6QWcf5PKfD40ZJ1e7yGCE9iWde6vYE8agpcZ2Y+lcIinl3JCjwr+NngpVwH8ud
h0isc7AVVvHrL5+Rq0PogC6hh110est1UGE9Y+jQAes0eLv+G6obSGX5R1nU5bc0wt6xXbAhrkBS
TRRfkp4WuNRv2zgDvc7nLRmRkuonhDE/GVNNjKM1x2g98Nf1fbVxtJeQSg2WeE4lOi2OJw3Ktjmw
37RrHNJ+fLQ34w4RYcu3VHuvibhIoTvXBf+Iv62SDyFl3sEIB2i+D7Ab0eK5nGx/tB4hwLLm0Vf5
d0+IZ7GkxPZuciQWcetHTRA97hPpq3MzxNwUWNMwzZgBJSthvA8wCzbXhKo12QBcjH/28oD+8SlJ
mZriaTZoVdnbPhrqHKmJD1Rd5SJLKevHH2CbTZc7IR6a7mYfnXIZYYnyCdJ/HwKR9rsT2eBVKou0
W2WzXRFr99+GPXu4vwqWytcIIM5sAwDy5nbLk97unJ5PqzCtB1BuAwZVI7vJ+YwUEVUSJ0/AyPNp
nNsjJiwfknqqTYRypF7mkidVVwCY6A9rk7fLw0UXbFTV4JlNQ6Fd2GQJZS1F+4OW4rIyZYfzslOo
w+eG4lkJ2mDeowQO7QJ7biBaor+unZNu1sFeGlimcgczS5p/TXE2Jp/ZljP+5UvnILyf5eit7fOr
vVmn+0MSE7PoMc/OwEs37plecFUNV4GrYh2AdtDbdqNzRNhi2iqsnl39i8Vx8Oqh7X/y+/o4CBA+
DZyqjTDNKUZNzweaF8IxFMzPoZaryATvsY6M3+WSkgQtiulL3p5UHPw6ESzgqgzacBl8FnFhL8TT
7y7m9fZggIkSvo6DLtJKctqKDzrPbwpKeOR5MoIeqHgedIg7/cZkemQAp5irICta+7BpeoY5v0jS
+hG3sr/ZKEidusIdcj5t3LGLdLUPKSrzqNIVquB9a7QNwTj2UB/X/qfjYsogHs+vaxTa7Bw60AVc
w2gw34pMm5h46SUS0ttKu0BetHVlyP8m/L+N8WhfSM7IgANC3JH0xMJ4l6umMU1YFhOPR6Y3GqYu
j1DFnzzPVKCRoz8hYVlJZuFdKb/ujKO745YbU5pCfqTllvbUA4b1qEj5TWyvqzO8cBtmLQJergPR
uCXXUlqQRQ/KQwOtdjKf+CF/K//4SXXkvNGRUSWv/iCAyucXvSeBtWCoWID1lMp0aXtKaekMUfqW
bLatiMsemOcryUCsJvgkBTXhMsCFMOg+p8xH6qeIEtS0BDwmzNwdlTIYEIWy09hhlJlCESvhaJg2
I4OVgQSTzeCpAWgMpuvP3/iCuxVhGbYeTBs5LfBsgFWgH7uoGOgZcFAyiSNROaSijF0oVbn2Y/Jb
d70sKnY7KszDvC0LqujvAQ8bdabg654Nkteb32/sBwBeMnBbwBmKiwEGCP/Q7H3CcXMnrPSD3UOK
HLI2mIKA2F9lOTmJWqtSo9yalFuCCvyrzW2VdGAfeDXEzWJQAzVGDUDOx3Ueu2vDepTY2Zmzw9TG
20vrISXlO2VNdDKmMwVe7KL28Nw6+X1qo8n4sZNnWQNGIZUv3/06eW8MuTuUmVu3eRosSiPpyg+1
70kywSIgfr5mmBnBU0I0d/yWz9sycEEnAoqqmWVqRn6tLit0gfm3yQU7Lm5flk6hkhiSBl3qG3ea
mWjFImDAwxBxwCwxLCCCwmqzLK3hNW696IeIMU4EHyUZLxANXWExWZN/SOsmbQwJYin8dAKG6/bM
bnF39VADtCP0apG96gVO5mK6qjUqG3wzpkn+8RrJKr7rMLrsWjPKH2QuhCHGmFrnYk4CgHsFGJVU
ZGYO5aVVp2dTBoDFtnE1wTvgVajaJYIKAqYkOgWB4Kx/3z75gu7pGsLKAJ74WMfBzLjfQEpLd82+
9MsD57lEzxIMmKf7TVSuKjq+dMrSznqIMq9WtKo0UoW0T1Hd+wYIiGU+iyR5LZT+0KFL7xoSoetp
fgamzfHENyNSOh+xAyO4K4RV642cXOJmMYdSzmT3wNm1VICitoq2QnoYgEAII8AzJKox/BfAoN5d
pjSmeiB0701xvQIfbay0hoKefdinf64YeSCwf10T3oDQqMH4UxRnf3937Q0L+OUt/zZbX2hAkytT
4JI0Fz1VMbWmH1N8i01210LoE/m4XppDZl1bYBmzBrxqY3A8CNpZO6rGkOB4Ey2n2T41nRgBYkHM
jcYeGb2uXTgnbcB7gKaTeJJGs3lI93Sa5L7YMByv0gEq5y1QGTOQ97/mFsXmfT4dv5tfj+5dbnih
jJU8TLmMcMk/8rFy729NSoAHElmI20Q7kU2ZOHV2Y6M4aBDE5ko6uZMDV3tDw9P+3UvVB/3m6h8Y
Fl2pTmtaO0qKePOEDQt7wqfk2z42cmSqf98NstPJsQ68OnvylSA7qBNi901NPCuZB7O/k3Gg45S2
tZVqsv3kdpcZHh0T4cCaORGZoPIidvuGl3FEhJ2wGo0wcq/jslgQIhUTzqDhSKjWXNm+e1eudpa1
Sxc9twpUNzRt7c0PIdVYkCrTehuocDYIRKJu9eFVe/35lTp679voKxNNDPDe6ezp42/TKL/Cv2JS
+bTZvi2vTxQhl+dv0VJgW8w8Qs7Exq3njbqpSVP8TWdB/XL88OgloxuaCIPv/LeiN1ja1FtVHMXe
VvVN/HyLjKeULf0V2xqO2CLitUXcOq6HVJdandpI3706dWf4pn+6CUQoESYA2I3fOyk43n9tK75L
vAz7WvNbozyaYOkX+iWQmgVGHFQBdgRDyFvJyeBEsLinxdU5Q4GpEJ9PE2f3WjB2eN/MURmuLULp
CHpo6Fo9gJ4U9j5l7Zm6fXzwMxYOefcc5LEkj5K3AGS9d9as1UdH37sfGmOBJr+pyW+4XrmuZ6Ds
vBZZLg+wHXvaFOTRz2dTWrMJH7sSPB+tvDv8tn3WJhf4ez4j/SYI7ZuA6LBktGG6RiOdGcph/NGV
jMWBZkMiulW+6Via/N7xq6lCWFt7KYkIayljnKi7Jd5bU+5hqRLrHBoIvpPtRnftuam23kUBVpN2
11rCPSm7P/5B2pwC9V45wwWb1zKm7NWauNjnYmFuPNRvNW8ikAQoTDZNY8reKSIep0r3nmQhtxD1
gx8DfLyKswfRhEHXH0d40yr0+19C+Z6NlSCx7qDX4JBhqMwteni0ePxOmML9TgTsMMk/cQN9GE5b
MMV//m5SdrkkEgonmuwY9/69GtqOOiVAHu/3TiQQEPaMjNUAnsk5HJMp5C2SB9ZpHBuAWrYLzSOM
fKKHJB+m4rS/s5mnF+2HBOTzRG7NEzNX6sK4t7U9C8sLcjrISFH1CX7/9qYAl2DG5u/wNHLjIkj6
xZq/PHnuf5kEffQbC9nouIfT7I89TnvzSKVsS5PgjZyfeHgSxvn5KMjDDJf/G9Qpg6vJWi53nAlQ
oakW/Ts0rLNvUdARoYSeuNTAIUs4+lI2a2ASEleMtTATLyhnqC7WC6iLqFFq2zMAFT85D40vUD76
pFHhAph6adCsADlq8FqE5ZzUeBi1wMCwnUTtWaygmnMymMuAwwYFvb3Q7BpFN/XvL26dYZ7w4WkU
Qk08Uzvqq/SHQYhGakAkO0HEevl2ehFI0zLXgwI+UJtsyzLEYWx+NSRXfuBciv/T5/VSGET8CvLG
7anOzusVdZhs0GyUPEVLVXD++tt7yLiQofEyMXeyYrGnS0mDerVWxwgxFMKCjFC8ahY2kASl43Sm
KNInlOy1btSZmyrdXt6NNWrQVAVihon7mLUk9vyvNHFxf+3044bLeVZG8+1DMdAdUrD6l4CP5VYm
GAe2T9w3waFpuoiDELmPr/8/k8xcmkeAGsYriyRE9LfvQwWnc+o1R8FpWB8zRX/Ehb0HHkmDPI7Z
XHCaYZj9nqH/t6GJh1i/z3fgUCXASue0NTZQzq54115guHBEFkksMH1I0V8q3pUL4IRpc0kT2NqW
ieQXrO03PqqlAGUe5ee0Epd7t8TMisVyKqjccNLxWuxkMp4Pzu7SfF6g+2uMKMAQwJRZgSNd2Ebf
/MjE7ii+iUiDtUp8OxwDLyNfaWLfyzYhKt1W1NfsK+77USV+rRsm+OZFVtDxOrwPh2WDvfVJfxoU
UtN7RmBnz0uGcJb/vzoLAAE1U3egYsvuDcnsqJlqqfm970cvXkFNXo3eH7Eico8hdyjniQy2cgBc
WpyinZ0EMov7GXvH1PPjp85hATn9SNXz8sNsOrccdZ5iV9FgsQzQzEGUaxQ4tvNFZ53c3BvyTxB8
4qv1jMotomW7fG1ZoXaQUqeiOsbxCoPsPXw/AIOwCVZQcG2HHuVwKoEjt2pWh1kADO1GWHjYlCBl
9AZHNKo+ywMMy1bmBC3/mLX3vDdtxqqnVy0WmiTFUB/VLFjRrOzX0BDs1nx/BCsRU3zcjP3q4Znr
XfTNWDjlAI/twAbLNrvIwT6rg13J6eWstC2/6APWM8enZ49zXexdRikMJ5mcnwqvNMQuXzyj3Kyj
kMwktD0kF1etJmZrs/b0UbmtXHDylbf2Zfn/GHH5UPnGgcWs2ciLX/GNh9oRU7L4MR1BmVGt1QPb
Tn4cWVQjmetp2QABbI8U5onJt0sDe7J5HTY6BANuIdxvj+HSRjeRN2oDW7iOuUSE+UVzoaOVzaSR
t8Ee158znP0d+hD1myCikaopZ6wfUdtwYxRt0HY5aMpxJmlQbD890W4lFa6eQdqftfMrqN0FXIXb
oszoTKC+nVuDSXDSx8+V0m1wy4bdJZxmzR1UntI5CqnxA8JOIWf/dQdkYlSSQwwTXHh03/Fckm8v
OKSyo55S3keACRuroGvYCTh1ai71/afmRWZtSqoCn2UrA7I1hOuv70evDtXwvFUrubSJXjw0y6KJ
62x+HKhPqVNSjOHcobSlC9aVfS1IAtA+60eoVSv+9wMAZH2VYbHUjEtG2fjX0QDToSOQ62lalJiK
4lnYZiGHNbvsAjr0AIPHRiO9W6Uft0K5ytsMtRuGT9GKgrOvW3d1Qnrwpxy1sfV6hxlkrg+1YXSs
m862xb+cN9p/YEk5wFl3vYh2Hu5Rhe98jjI4Y8HMqCATGxmIatGL/eGeeN/CqKWAWxEbbhLZNDfg
xvxmdgT6pbiGjlFkhbg8J/RHACnj/a6SShaHLXaF1k8g/1Yi6CsOpJG8nikomRThHqC3TSYqgAop
3pDkDUm8jdDNcVVYcD30EBsSoOPCFJCmQD83tr5HQiN0PaEusduVS4ANp8Cr1r1GEzAxPTqlso+r
6QJaKCQOjY5+P1PxHAMy110uKCteopSxCF2pfbnwJ3MpYYzvi2nNSnPyDYAqgPiNVXSfgB7/LDai
czDWPBqy4kYrtG8RQ/OP/FeJ/Qb59kZ1naNhyGIijmhnw5D7s+dYJCGfQ0eGES/lHkd0YEIqWA3g
+NkyvuTzBDlSIgj6FXEfRc+OGdW7s8itoN4g2A7oNR68wz/Imhp2fIbgJpkMUgENirXmXizOACBy
BiqRgQLBbmCy96rgrQl+kr+qW50ezdl2ta2CTOJ8snMz+NvDNIjLtbF1EUBhNBkQq1Q6se1SQjDo
AbsvC7Bzke4cIOh3wf5074Pq2SGNk8mAUWNiQcWEygUXoJr83XXBa8IrLCh0iKdqZWDcjM/0EGfF
ChkYiK9JFZZeUhh7FkSmxK4BR9L/iBaozTN2bHJpdK+0RpHp+WAImwYqWYg7VV2vb65De/dds9BD
PoAT6tkwN/lk2D8cvLkCXL+eOYcQJoIjsBKzcbN2yr0p2irSuJke0LpFKa7rlSqLcDJHw4hDrRRE
QtB3bVQugbKnsZdaUkgSuGLwWaP10q+FsJ/F3WAA+rDLBRJ2stYwRNzwOHwGMpz+uHmrbn6mHPam
RsFa6AW6nuqBjizahWDoO49p65jvDQAHPeuB9WEazlM7nTTdKOanvtMPLsdq4IPiQB7OBF67s34U
dYOJkCbTtXE/+9OBzjNpfi52Zo7YNqwTHZ/HyJVW7k62MePGP6r+g4B01LGGSFhswqj0fwcKHgc+
QxyvVIXHin/H4hj8IimjdV1njNlsFhO7Xnvl8XVyBK6SloNyVWYa5IeQ6WSpHhiFGrkMgYbu8PZj
UfFdzhPmJDDLjkp87CaOf0nKPWBydmzaBVpn1ylpfaecyVPVDANfriL5OVnsImBjZ3GFeBAglU0Y
S51kDvsNtAno0Alb2UoaH2s2z7zIlld75/TxLhw/DMGWVc7Uar/7+SFRFCn4EngSgKuhwM6+ZjYi
OKgYIsybP+n69mzbWowLyWW9Bk/FYcsIyYNpuIzr5l+/Q5pvZ35PVWUuJXzSyYX2Fiwy/YF0aflJ
OHjz8OOk/kFifHzS6cjZuEaKaZhxdp1yd4GhQXuGvh7fUukVHbXnSq0DgkU/CQM80Gxos0bcSWew
dY2wtQvG2eA08Cm6k7Lla+TriHX2z3bAfZ1O/Asj233NOxoKvTQEGBoXVULDWYf5D45gn8PqEUN1
cPuF348BMS/RiuxCJsoO/AhQh53T6sm5EncvDS/YEKcl2CCndwegKG+fP2U1EaJy11nly6CV2x2r
Tx0RQ2hgOVOvTOnopeFeMLxNswvatKo2tEXOc9kEhwW2i9ZrUYb+Yn870aGEo1ph5xtpIR6w0TPl
FBVtO9tDw6jEZBAsoHUb2BhN3HqXvPWSUiLNrEwSUrZR/8HNypeaJeCmeiVYyA3CvC+fwMsClOHT
D/pegIiJFHmxwzXhOO1VQ8vsEAl7LHR504zCljZH2DO9SBrm2GX+g1Z5o4BZEAhqBD3+C7/om6L0
JfhC4QjSlkunR2MWvlLwuEcCRpvSKUSyEZ7KUWfFcf1y8ipAFh8fRQIfiQ78SG2AEIPzd3r4bIzS
dcC96DoYUdyL3FbZPF0BZuMJzAhTGKh54Bp5xV6bz9/SfjNchwHMTrdgrQRA6xTKWC2zwmmPkDRp
c/lEc4/PaUoeDw6SnOr4nGuUwm/nVv9HyYCyJHDpf9dBVtUTiycWDGIfKREETzcfxkVFeeWhE2gn
yPmZu4iQNkcHxci5Rqr/ib5j+lZMwdxtizMoeSjROvmd2J9PILf8QpiPqPReREiEQ5XTCIVB44uY
6Hau+Gt0Qb825lWQ3PG5PVdKymNzDYP+r9oXTNfv3uIPQ+1tOSVbkoFsviJwtebarRiVKUBPS4oW
ZNJHFAAs+64ILGiIVenyayunStimYLc5uawG8EYA/s0eLRhSJLBSAjoZXQuWCsWAYP4C4r5FggWN
ZV8Gn99bAsjfy40VTA4irgHr/tUB5hKJhsV7rsK2CasE3AuTW5lbj1zck7o5/0uIUrRVoJGTfFON
3nMHohqX/0NNt95zrGgDIVR1/g0CEPH2NDvavZ4jTrx7WV5PQGZ7TYPnFhTn5kvqs3BqIKHrs2YD
PRx4iEOux0wbnPqf+7bqAmpEJMkcaQZtYCYgaLjg1RCs2MCJRpGD41qerpl2vdgsnkm0Aa08fyZh
6Uv/6dPk7FCwBIiAAlqax06jxlOrRejis1nM6zfr65ozLYGcX+e0wto1Hai3RnL2opdRnDgLFlMp
6BrghBx8uHaRoQRmQFz/yCcNHAnjwO+lGUUHIXBXKBeLlqys6jisqokDOAKzb8N+AB4NIX8PmohL
zVgtQkkOfgC/55nTaX1oWgGYfXXS1WglcGXgRjrXb6KbxW72VsNbxxHnGEM0UwjMJ62hJMN0GOy2
sLTewGRy/dCOjXYxrsUOY0ELszY/gxPQePmDh6uBPyTATWNTooDCRh1Pac8dmClwqsHbWhEEgPYg
E04ijQNfCA7zHXV93ib76Rhv39O4w1v2/ze0zpls856rN7VsEewXtfFEr9X0V2R+GGEd3U0CYX9x
huHCNrBFXqjY+NSuzc45Hu+iWG6cxN1NbfmyrGTm+mXykYJ5Q8K3TpwR1GpZ+DsljT4cHH70/7RC
5UQ1AQk3/+kiuj8sjGgcRLaZ55bSFGB2oFRe/jSYer3t2VnipKTbTvgcwMtfQnDbCUVvDsKLS4UZ
1m2m/t1sx9QMTdmAQG21oxgADSwPo9rnZe4EIXNIwxII6Bc4wsqoMatY5iSvdWDX8H1IkJLiXXY2
nfZj6fhY9is6IOS17yPQeXW1xbYnFQy9LCIz67OFtT90ZJwIAfoUww7LOhmWKxuRXhN+bpnz9z+i
T9A82uxFwt8qoa7Uo/zFrpMktKxt19MU40MlcbNDh3rsKOQXEgCEdrxcgvkE80jbmWrA0m9bdC4r
FqH38BK9sbZqwXAKNwNdw/Od6DfzbTJwz9WJSkPqE2epb4RgXtAeyp7teRNU70lU2u/eUoIlF2Wp
KhX+1TCnJE5XBZIe/hjU3lJfnxvxyek06WZGQSYpxKI24KJvGgrU/CQSa1bqMGxv5JWZuhIfexpX
IJaxCzwzbES3AAXSXcDhvALjVFmpfSjiVWSrTdDdd/QLJ51fHbqENb1+GtgWEhTTlaeV+D/Hec/l
jDnaf2k5x8OvDd0LPf1s3BkwchGAGGAIiY9vzQ5kRWBN9yyQpAXDQuEXysSUS1/w0rFzYxpHzfi5
l4isErljSZKZkaxV0JLGDn8GGCLa0faI5M/Y87KDmcbpmd3XDwKlMy0Voh8DH+S9Zgp+wrarDIsP
i7rt5wI0dunQd+pBBXr0HU5Zqiznaw+KG6QO+lvas7SUSi76A1grDk4kbgabuVVv2QITpl2lBCg1
tG6XQl36FigPTGY4l3FikaCzelW9ZvB6t9GxXI9zk6siFVmDG5VEA9itOzRsjxiJK3ZFvajsYq7/
IXgzZFi/Dhpj56sHjGyYg16+MGuIAWEA54YSNCb2EvF305mH9KiLKBuQGSWvdV/FeP5LZl3Wf6JA
5szRbzfiUFWB1FmUXd7eVbafxzJMflntZH5riSaQadnnLcvHOSAc1V/JVSEn79neOS3fU2WMQdbn
ACpfA3gFt1a5m/knOYRcfttflsCpM8OR5AShznS7oeILYFaWbIW41FcCPgzZyHpAro1C2MuJwbhk
GjH5JFLRNa8CmHn8iv5kU4eCppgAj7jfe/nnYCp1m674vSTI7uuSm5rhKdKjKtjUxcrlmLzzzLg9
Dj2jzQNXZr9SElHbb5IICyzKs6seO4QD5D0P9eTMwKckKesh/4gYdT0s0PZGg5zgKmUAKHijrLXE
1f7jk7NICDbBSqnSiGc=
`protect end_protected
