`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GfDD68oytDsyjK9rJoAaNxe/H6p9+7lfJ2AkYo4c47rD+vP7w9Ettsm9s7B98wDsnyHRZ6+vhHKA
lNUHX9qKIw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hzJ4WCrRc8ohMB/GPkJq9t2Dc1PKouHzu1AfrIbb2XjAfoYKX/eaU1dH4jb8w/tkt3agRCukBrDQ
stv4GyZTM4/8X+obAnVLBDxlAB6DS7rd825mjfJTmmcANPqjJGv/ebUGd+YqcxYwhUF6fKcYaw+5
dGguJakCy+DWrYrQZRc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XBb/iY3aITy4MMgTd8RIgziBK+IiCaxdWeaiyZ/xIu2RXbLvdkAZm3M6/q/qU+DycRTT/x1r54sh
ybKTelHU/3HoT0oL2qpXoTkPxF/kLUw1BRR05V5rI4SAW6GRu9AuauwhIQYpDVsaSQe25Uon2BWD
I2nMCeLV+iurV8JVkHNKiCIGGv8+48nJoTmU5lkOZ34pA2HmoHS/hs0XRTOhjgt697urESDZoPc6
C3sMW9+A3+SlCjI4gox9wqUqv9AkX3m8oOGNEQpqM4Zez/z1Iy2X1DUlf0SlxZa2fP8qn1hJN/QY
2p7MXQv6XItMsiEt0qETAYXF6Eb+wdaLf0Liog==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hK7vhdcgENj5rjKLjfg9aXfkS49q3YirIharCVuLRJLw2tpWhJZ+39NU1bPOgtrpWbCwvAGBopKr
gV0ReFSx62w6BP3cFzQstdkOUkLWJl29iJtQg28016AkCU1sdXBNO5E0dPfXakjRQmGIUXzxE/Wg
O8rLbOA3/gGEukzAb8s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LmYu62TJuZFMbqefKd4M92eYdogAiJlu+88yB/xTs4rqvzNCmqEAbIiEXy98X4cdn/GRAfY4N9eo
a65aiAsfiwU5YEXvqPpqL/M7H+Q4LypM/+2Ky+JgcKIl3kG4pFRW+U4vvlvymA9pTCI9jJgHLMg9
PkktnEEvkOStY9W8Ybafayrie8UuGCnofxn5Ew1zPdtKfSp5wvafb+HX5IQNWAjn3RENAskBclYq
/TUUaeF9vS9wLjpxp8nHBATmDjzIAPWhtH3u3C5xxlAkDIVoxLTWsbAd0E9+tIAzeU08UJ4iS5pu
ZS13DhlejZ2wN+t102cpg6qo70h/HhIz4wIubQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5232)
`protect data_block
lnsCABYLB1q3geykGO7xS/Eh7TWxf78JSmoYCEegtt+WivhwVu48XwCGSprzctsMxxc85dvkQiZS
Yy3EDe/dJg2MITuVK3KhGMG0TZHKBdwtWZKZSaGB9BUF9Y6BOUI6hiwufGp/cb9ksc9opJE9JasP
lKMucNG8P6Xvu7vV3un8atCXJrRpACogVlU7IDYapPATAKfmViaNFo8+RCxx7QQ7qaUbKDzzC5bY
J/jxGT2G33+YskPJmSjOXL91flGMKFXBq6lf76b+inaMykfuqL+T4kR6FY41kJlG88ZMrpqGzdvW
4o/nDBZ39hcD76EEbPGW4iWtL3Majw08wL/gMl3HAmRXteeKSMyZmk1F05AwKRo74819/NKGGiNw
+UNhr0Ngg9iWgWk+mcnJVamm9FsIVAN2xVzJocdhKaEjYcFUGeVENQLHrv6D0v/E6dvlceqPTKH7
2WH0wdBuOsHRNrEgqmcUrfTQipAZ+Thi6bvfaPCUBHTq0R4LH/xWiBsbJS0AzZFSrSPnpcZZQgga
/jPO8vbD9K/ogpPcvvxC6FV7/ZaXwHP1UgNxZ1tDWK3BJ6CJo43uD9bDUytg6amxfAjLXuLf2y1i
UQpm1kFl9f4nbCnfpW3UbSe42J9DNMtm7keVAnKq74YOQE42geWDVTS9w2r02iFe8Ra0bkXWx4S6
lHSf2lNNmli1BvTEjZlaDGBk10i6KsOgA2Y6G7YT6J1B8BHSvjxJABFAUpFTE1gRlDGGHkkOW7v2
AcJrFrBEDan05mqv16KsHD3tqPLoicseDCQzaw30HUMEpdeS9RX+pVPCh/11C5XRqI1G70zS6EAj
Da2OW2qKBfeTH/wdUV28zWP/Ot/p9Wq7+V3StJeBRPFG2kmTTbzAMbKUh4QWQS31MCsqnM7en6pw
lGNz3pmRqt0KZwWeEh8Bzi4KF0/g3+TS+FROQ4xuVFLcvpZUqz6vnR71Lv852xwin4bYOawBL5my
gnmeYIJscT5ry13+Q61W35m5acHy37p+BHjaNyRGQFnKh9VpkaqJ0wQUEnkSzV746+0nLqhdiXGI
ZuuEourGebohxP+3ZwgzbBnXvJao7o7E5CMf5WV8q/1GZBBjNeSS1JfTaopb0C+TpsBvqLyunWhm
DFVQ3M/r+ir+RRhCYI3tPvubUechrtzCCKKT705P0z16O1UQTHjcImll+pAn53PiO2AR7o+pOYYa
bZOxhw6eQFEW2cJ8j2/W0ElYIeqI5LPM8pQbFreI7qVQDKtf+OI/gGHBlXlYs6SgNx1UEUQJ1nEd
5GP/3M3NRf7uBMDTr5CeJKuFtvUbE6LUovtc4vK+gvo4M0Kqk4Rinwk2g3cyDmqJ8VpC5Hh7DJhk
xWwu5He2xaVUYn1/IZ5VnIw1u9n0P9+g/Ui4UPprsxzaqjlao+4V+4LIEHrk6JdJ9juoQrdXz1AV
B9/DO4gvqNUWGInzqHBUrgoeCsNMxNB4OPKoqRm+4g9AiwWu5jzCUYCyVxCR05N8f9m+T13aq56L
AfaTwjvww/cMai/VnGOa0GucXb4R9HZ/YdUkMvWxnq+Avv8PdfrziJXEpNjtQwHyhZfqzD7rce/5
zjVHVLhpVSklUD1rPwBtMDRGIFC+skZMjIs4uBHGdseDSvuJiX2GckX9WKKwxs+7glCKIhV9TMzG
ir1V3ZXhwycVIJ+/iGS35COGTgfTnewPCOO/zHhePYz486y87+NozonnHaRATZHWk04nn4U5dYEH
FzXDp6AGcrgevhb4qRvKmurj9DWdZAqffdep325qtoqJrioKoC0WOZA8ThMKBCCVJVOVgBAeiTtV
hOxaOt9jPur//6nlBIyVxjCqcxbw3ErItte/crW2een3LZGpYq03KMOAmqDR52bkauBQolhCvO6L
DXQt9DZSBjWkR1unrwJvvBkZMsrk5A7gES/rx45PFfgMRs7PP1T8H9VVmATrQjD94WFuOewSDnzm
1BRGV8E69GlvXVuxlKd/XaeQWgVlqaSUwDf3Amc2xCefVyCkC7FgPlsP8WsW36PM+HYqTySKnT1W
QpbFkoXemyJzc8FNwn6knbI0KslG20p96lp7xbI2Pwgmbe3T3wMyfJ63i45seTH2kV2rwELqldsb
EBR8oHDOWRqnPpFUl2MR6od8xGdEPIxz/fzKkmXglOu7Nm/bX9t8fjszL+fQt7e6jP2KSlAesLOH
EDiMJsTDjHvaVT++u2JPAFu/xlwT7ZKa3c6cSHV0ZgQsnARX3D9TItLR5dvt9GfqDJ+mqcSqNZVN
Gs9uRUtGTHg3sR9DObD+hXCAaLzscjWYTWdJPODsTu7Y0KyFcuMDzkmHNMHniU3HbX5F3tL14cjf
KTWOtxtm5svt5dDLFTCOX8wuD7FfZCCL4Pd9tY+095NPau4e7xbb457m9NPtDOVL4RNxB1FTkQWi
Ihe98OezHhPre798JDjFYhptWVtMFlSs/fK2bsqafgmfQiNTCkYt/bnFfRXFH5oW3G8OVHVHk8ME
7NVFbb6ErSi1586sqj/r7eWQZEnWue2KdMpbA17IylkH7IWcrvRWkTWNsC5pcl9rk80SRJPlvFUT
cv4OgeihgfclH59K46x84DaAbooGFFHmbAj3pVnSLqkz+nSGz5YiorEFgYRalYw5ezK7aBK4OTt9
rdMetx7wkD29nIwjjUO9CkChDM5uVvFgD4ElEFz1p4X02gJmNMfiv5Wa2OzjICiNJxt8nzGEqZjE
XOZRZ9VwBjm6vXjyxhSH8qi+fKr4HrwV3G+G5gh/1DAJ+lUWIvAHoewNM7gJqI3Z8OgLbGAOqlEi
OnzcZnSIqzdRBMuFK6OmCmFVzF6eFTDp9RvAAUhr3MMxZc9MIlsa9iT/7kSgfmxCmL+zgKC7Gbp+
BeLCJP/E+dF2ocOluKYvCqj1NALSZI//SzBbXrXoM+oiYuY72O36mczBw/T6JuCp5+r5HWgJURio
Ein7gNGo6qnDji2OW4T4533ITkhsZZM9QaqkiRq7T4fcxsXgvQnuSWpd0EsK3uJw2XiRi3HaeZnk
rh87WQSI4RuMcu84RzCzi6lmLXJjqS+tnsIugVbxB5DoeFvwDCN2j3MdNXHffkX18yJad5sAo5GU
WYMpjFq8dxqaChFi5BQReqdfOKhCIO5HlNHlGdCM5fb1Rf48Tpxt3SSEuG+UA5mlRjJam6tHzqqC
UJWuT5dbTx/sPY+EqI4gFyuPrMR+CB8rhRlxMQT8Xo2Yn0iIzMe3bhDGbYBeATvOCdTcwSilrbs4
/wSkKqRr0TUpHLrNehcjRfFXsBaPcaOXWQCCjNAdbNAkN3Z6tbLgj32VZfqMLXSoyK9PCqP7SaxF
h8lNdFmIQxgarCUYjXNqzfANV0eqA6ZNhuhBkK14ceTWT3Sxo+2eoJ4v0XEFZ/mSP315EOsWXrj7
mqdmzcJ5yK5c2/e5hRXsk5WA/TqY75ymIFIYNyAO1HAALv+VgOOdXQdQnrPwb1KlxVN4idX5Hztj
qAX+SJgLqYxfNHn6V0r7etT41AFvJ22m5/bFmtxWrMBFo82ytuQtqYzLQVFcnJ0Zctm1afQFDxox
qVx5o193PQsB7bMg8MM24O5NFb5ICuNFGo9HF1TGCDtoKh0tqyk/X5BSyVRV9yNMAGCqrKXFtAet
5f4iBPeFOuOLNcE6z9WwjHtqz16AC0zmQCgVMYmtYue31eQamrzUANrpljEflyKPKOS4NgSW+00O
M15rlhVk8BIT6z1utsflK10Jz31F9+sXOAEu/o25EsntQjtXgdUWLiGhNswjJc25P4jXusFlFilF
rMDJTuA0PzdSLpJlgI9DyZuk83NsmpfHVgRBITPSRJQ7NOB7+xs62f4qHZNOpcmixu62D+YTAGrr
NHHKu0NMLrlRHBUrwwML+S9p3iU57P9FCV8AgrjEaAWCkTUsiyxZZAJ4TKXWqhkT5PVuKLx2rlaf
vCf4bj6jx76vIAjl1vysJ1d+/lVrHWoS9DcpIsV8xtyeNOFZ1+fqoY+VLCh0K8QQmfPw1gbJAk1/
LLzpnrAgkp2FM9qPybQSiCeSj7SoxegL0IQ63SR+2N8bZ0kLWkr/YIyXSXzCoF3cfLWX+yw05j1J
vn4ocw2hV8FiROYpxp+mc/gNNEUWiaxdgEYYbZ/bMttSQjYFqQ7C7UBQrJbjmZYDUAx3ZCRnuEAK
UiYR+2Do/IR1UIRgibPXEUVpzDLuWxPXhzMi7baythlWw13NvjivmRqVatFVHXIeKXp++h04ttnH
mwjdZ9RFdItov2NzpSz7ThyYZE6lqzsxJrdpY4WmIdoASsGUP0xYbXwky0lAOVGl94Iasuqgy/Yd
i5P6nchpkpTLGJsZexAyZl5OLma+3Q8yCfm3mLME/0KjjyNJaeCOoTVpMMIpcNNk8G2QUyvLLQvJ
NFVtj9BLWuq+Xhx7GQhRYdoe2OHdMIT+D5vRoGaa7iIKjsK9kK5s13G2k6ZCkbGGbt6fam/ZGgRq
E8LCV6hvfjdTlihY7PLzTBkPh1Jm9QwsjNX/LIibx8YdjmJjnqsu2Zob1yZakc+OziwvesuPuB0K
GpFm6MiqdiGbbCN5BOrxnOvp9j5k8QX7f8CXxBdCGmw2w6ywxmPOByuSKHU4ke9BTB5LKKkL0sms
/15DUW1u6YhXPkqE1QWJFIKsnN9NzcTLJ6ygH8wz3k8k94IQPfuttcZbbSBSCXU7z7peZv8LlKpy
l693mHLVmEsJKhom1VJ915an7PpYCjR1iVdtKWI7pi15vc8LrcatvzoX85oHlPlv/OxaV1MFxZz3
2TJ72PB3b1uHEb6a1JeibnhWAnKeQ1xn0gVaeby/WuQuPBQZZgqReV7T8NJiA1laTKQoJT/jc4fg
JkUuDsrSqZE0wgO61YRuTODpa+Y9ttJ+UtfQaRHw6fY+CGJbDQWNiO6J1l9f2Dj6PdeoKE2fnz1/
CO+ilBCCjBNpcBBJyTxK/Xn4xVO6ZaT53qao/WLu3Oe/+UnWmmcOU1oy5RMEkJibx3Ale2t/1qtf
5Oa0+DFF3VkIMlKsspDtD9OfP6FUvcT53lb0HRvDEQzT65icgpBOB2ef8NQZoS0s0eQLlsQsuv5o
c4dokRA1ENm5Wri/CBC5M9HHWfq9neNfwdW3TmjjbM1Hx0j7e7sQy7G3FVafLuzmf8reMxtPGhCi
C+j7hR1GdtJi2lMvB18KD8J3Q+0E4VzhX7RDNWs0scj2t2hQ2uL/L8xX4k0jBAnqO3i3Lh1dLXED
OUv9bEEUBZ0MjUEsHP3gSeHNydx1wUpqXmAxTUbopBAZz7ae/FqAEcEniqdQFRgx/kwlwijXqAEB
wAx3FvAKOdw3m3Yo20fU+fNFGFfJIY844JSuz0BOoroqa89dQXLzcvqkw9yO6vpJwr4axgo9Uax9
hH+1B18JrmX0HX96EFEmtYvP0fmsTdUYdBWR3EW5fLdpWLjbvrPZXRYRvbYu9oIZHO6IFvlh4TNz
YIWTacZqA2YYzOZ1pxH+YviFdCOAbwHgfwQpW/bY8ZPcOyldBsR7FitjAWtg1ZkGdFqczL9E2+ze
N269xzLCkp7uC/prnAVFE4NJa0/Fhh13Fw1by7FQ99WrvZZJEx3kzvac+sSOsfC5pEVDWjdcMf1H
H2QDF8sTBMIiX7wuO0er+ZJGBcYjqzk40iWRLmefr5HjwUO/4c+v59jwvdtBLn6Nqv/E6IxaKpz/
qtNyslCTReDMrk1NiupFv+iCd7qRKTEkMB/XDAxLRbGyRqXRJkF1i++5tscmU0IvPUi06G4aeXn7
mfxwzx5Z1Mpcmvp00gxGNfni68IpxqSJsVr1k3DA30kyTqhmKFaDidbsErSeJqPKp6pS7wPpGTVi
K4Nm+9m0/k6h8Rm+viX9Qrn/d9rj/kvQm4ILT7Zgy4sCnLKA3LfwPpp9Q/UGHKR8dPQgdH1DIK88
GzewH2196F6WF/SlD0Qb4E4XUY5aCcwhe6rtxTq7lyJtRsK9UV0i7lW+nweSFlkYrgwHy8Tppk/V
SFxF7Ny4HoO12PeHdtBSZKwKNEEDBEyiMMPctb5tI+mR0QI2MFkGcuWqzx7eHd4+J1lhDjYWGv1c
ImjFQlreHkrby+XTrwA1f0U/uPqvowfeyWOqp1r6Y+vuPvLezhgnbfNjk0GlKstQyT1ocrPKixCZ
ziNNTxKBaK1YTGmAXZFFPjegRfPnSR3OXHgT2ot+Ct7u1RRT1zOxlrRSZELUPlxHKy4zzFH6AHVn
xPgpKMXLkmf3S8PN2BCKldGqSqnTXxOmhFsvIpb6vQnvH07HFfLWhOaAy86JDtYODwROIDChz4EP
hdqHP4avNKFs57onvFy3ujKJ06u++5/+kNA87EKPfHeUiQDDY02ojTdesdZReZTEzBUYBhEAQHDn
qKjzIt3cDa/Q+FXFEp2u/QGksOXzkJ7H4ie0o/Tk5vAv8CdhIBk5EWFbaHQtkuhpL+z+v14Vzq4G
VnaiOYelXYSgnnXVDb5mGJINtVibpTqDIL7PaQrHd1sxHc2L6klMmqRUI0o1oZxfyALxatWZJD9y
5VTdWkVn7XvqMQQ6BGJVK2b7+h61KF6SmO5XpbDccmH/tHnITbtQxmXkOWi19cS1WkqIGSXW4s+1
EcJp9W0hdL9zCTjGOGYvPFMA4yFVS3Uu/9lxfvS2GexH7/B0OOOih05+k6ezTHj+cQdkfNJX8rHM
INLDqu6DiWUG6fc96wNzZGC4NcNGOCYXEVBWaKyAMwmJoxnJNrlOxyt+TFLea/RbmYKtmms+8QzF
cKyGZUSTtSgE5NNLL/gbAvp6FcWNpP4eo/sDN5XOz3OwPHX5RZObdSYZCpPP7v60DKGfaMX7MFOL
+5lXAKQRw/AChqHy/zBAcOfY1MuErl9eCJeOk0muS5Utc1Pcv7x/D/Lz+VUno6IfBRPVbisrqNOn
4gq6b30aJvMfsP//Zv0bNttlLlAzfi7izHHWsMKhuKx+OCboMpEM/H9ioup/
`protect end_protected
