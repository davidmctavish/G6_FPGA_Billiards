`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mqShA3L0xrr1CXM+0YZvvtaaRUJ1WqHYA1RkCJOxptKHHEZLZ2TgJlJnf3C7aYSPmzwHBPgrEZ4t
59sA5Y98ig==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsiAoOXS03LU5j+lvMIHiTAH/76YLmtmAHMzaEvrbpLRgWJdLPDvkZ2G4KrBYwycx6q0zyT9xham
NLNIS222OnRpye8y97Z4zPgF/k+fzoe9+Vs8CWpRHz8nk6+f6b0uArY2VEg5b7PPDlTlt6PsmkCi
T6ruBr09P7+uMq+TDm4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cdLiP/b6Cg3Rbajvmj8COjloYcjaYIzGNU4tOjn5Nj2i+hqW0uuYV/wb62Ban3cr1mK+DUGNcziO
81eRRbw0ZDX5lmoiIv25wRLqUlqPVQPhdS189inchZozOdz85xbDNO5FRT2jRyGIAgQI9vBlr6Iy
61XxNTzzT8zAGz7vaSrYNcmgmFfTuNhDKxvvi7Ayc6I1vRu7P4gbScFBa0WMMOrcLvYpnO/9nfiR
plrYmMPadMOYBckYY9NhM9TfVEfCFxm+qLVjb50vORqJwd6EIeub2L4WUJpFO4KRrkst0TJ5mqZL
Cpnlckg6l0srLlRyRThWFvuWbiMgAcHezzck6A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e9jlbS1OWz0ZIS4Verkx7Cp/oqMwNUuBPenxtOPRz7MMFBJZ7J0clStLHI1GtMjq25gVt6Y1lDPH
spzV//m1IH5JReHCGtvCxl9uUegxewzheDdOOL6yJEPGaCFIk9lHGqWBnF5uteUuswXTaUSnX9cD
1CtwOmmGvUOA7Dy5B1I=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YkT+wIHcljuI62r4ou0SHGK4tNN4pTAPncGz+/uG9RXJkJJkOwAy0QMgF998sE3bQskkqRitfALy
TGocAiE62Y/7v/NTKuWndGS8MGKgIi30t8b4B/pbdK0pyac2VMdGsZI40Jk5PPbMZMerhyLP8RnP
wNdCEZiEPw7IWzoYzJwMoE2oczEkviBY1Qx4AHm++6e/BXfpQdYo73RMqp9ybDmrX9k/xrDfe9hW
ydn8D+u1UetmVzbFjtSnGhOOyByAXmsM2T2WvDoiIodFPLVgpIVT3/MlHhFWWLxbJcdBitX7zcmm
jF/FfyufENdqG+S6cqog3/Ey8LLxEYRqY8vBvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15200)
`protect data_block
62u3Jmav3COHHV3CVY1SOc1Re3Gwsv2/fu4XrrTLj8zd/ah/f4mcbx510XsbXJYhhRgjkNw/450p
9LlBydJPdR0xf7A4wId1Pvq7cE9KWemSETo4nQGt+CJNHdwkUEiGBs2oIYKhAmdmlqvsQQGwRpq0
ZxCFuXIaZomK+hkm2xBKnB5LmwP8op7CTPvI4VKoE+7D+rWdRH6kiOQU32kHOUbDfoEQYeqloUQd
ztg+QGsLcEboMLd/wpzGX/Es4bqR7xEeqR8TT4SJhuay2ihF3WTOQDvpheK464yzWX3sX285m1R/
dkTG7buvDHyNvY+UAccg/aiI3QJFE8FrJWnb0QB0h3UE0+KHH/4iIB0colKbXuQvsFQCI1i6MQdd
Um0jdb0D+tnkxvX/Dz9MIwHBq64NlJwlB9odkZ/hNaE+8IHh9bfnEBkgyCeJSBP9H9v+l2iJlTvN
kzfhSPCYqq0vzUdP5ybZaXxOY7Z8iRaX+8Ybin73wvJmw/EQpWaq7mKH4F+Xkzy2m3nByYU7vLuz
kiB8uakZOw13/rfOfuYSdhkHSxdY5R+YOh/+v/UWHvLD+dj46c16WNEwm9HF9hevOivjprVUggNN
48RiS9cANNZud8C+vKl1wi0s/Am9bAe55IFEFP7eSv4FNrhghxxmttcfulkDJPJBF6igub/t3L2N
A3Fs4jS1l7AqS7zxOE3ISIwSv0uipCGlHXF8SMCrBhYCYyyuGEIoV5Oi0pVml12IZ12NnyI6366W
aOCBbY4YnUw21OKmQ64FKesO9sjqhxvOzGVoiz5eW5qfKn4Luktezfvu6VxaHSQrw+aKLhKcBrH4
Mxx6KIQ7Y1GVKLFVjNJuvmDia3dNo2Ma/filKAEYj3TqjS4ezy2tSB0zzOxHTH+oG2NJChTqZgRa
1BoPY5lWuRCx25xXEr4qw3MVBE0B9V3xx0bQySXkVNFE3UJlSwz2llUVPsqGjVDF0BWZoAZDy83x
ZlmXAz4F5YgKfJn9gxp66mWN+46nU9vzQ9UH61aPRkeD66Dojmu53DrYwtR/db7yaq0TaeVKrRwE
uYcc+zINQck8BfDCjc82pOfgQfe17wQ6zZDV7JW6FgfajqlKZyGM5/Vf+Iybi+gU+XmhI9pHYu+L
4tSsmslmB5S1O5vAW2Rdlgq9iieGm8eLXfh63m8rm0QIPNQIXquKAtaU1uJR9wd7I7grKmTRHiPt
avpROTFIT61uCYmMT/Xa/+XaGZJfaJ3Pkq2ocCGUbnAkEKpmrc/PytEMNVMW4Dbz3/etrHFnOwn7
kC2x4YswgIDR2dn8Hax5WkXMcGvp4o3+BQeLr9IA4/rpSg2UA1VlxAhnAMY0mB5DTCqE1wh0nLyf
zrmb3S4SKUvkp283B3eCyF5N5BRZT4NMLYGbMSW51GNpTVTGOia9rEsulYgFyG7BITz9qGm8UrzZ
iXKtcGqg1ccqfbEkQn2BpTV72Fu8xGp0VDtSMPT48fg8NPdOB/FUCZk+IXHLhdLrHaGoAqukmjj8
oZrO/8YixgYj6FlPGgoj9GOzuBzvyn/6ATSwyylUxyhEe6JlU21YQGocmJ8pd77ut6s63+7oh9bt
I2rVsH+8ZaUU+7VfY/AHE6f2AhHUoe6/w/sPpQn31hkeBsaXIKJkJ7O2NCUi3wYG6grAyWoCmTe3
+BuCq7XLUgt27jFWC+04aJhgYJb+8qJIXUPPWSOdYlk8qdhfRKmzV5xQULVm2yat+BTucViywTgp
Viv3012bJU3FKRupNrOLedVxYznpC/BSfrTDJBFzFASn+MmhF0De2lrsHa1lZPdv+65CuBjB8ZuD
DsiD4HkFNsWPVx7J+KKYN/eHJYMVAGv//5CFDxd6RtNzuhxI/WWu51WeknPZt7QFIlYXEPq1lSEp
ooxg5k85Hwe5hr0vhLQHY9B8sCuQSTgOlh9aLnc5yPAd0eDVGlPNbE4DLx1cZuRWA2zCNjq2oH/j
Hw7XUzVGRLzylUwVCQZJ6xqIVE1n6ltDReWwjhy4xq3IpamDzo2biEbS8rfAssRLxP3a6SA4tv4R
MBGIftVECrz5khPjYd8aESUAG4Q6c960UhyA4dSgEE64sl0sLD6nsOAUTZ9/17tMbt2N3NVnaf+I
tN79VVYy1VEhfVamaycvgedhrQGlvTLzdj/sZHBWPTmtf5JwRG9X/JPR0D/MnH9EhRsMyD/zzSvC
q88qlRL9zkjtR8L0XOO//9dXMObqIzMY5fFxmR5/+4FQJRedFx6hshQ8z340OX081zDBM8mf7A4O
CyUunzLVaaEuj6lHZk6SDCZneGnzyf9bRqFBO8ehxzJa7CnGVCd4USSIGvttdfFI+0m095EZK7QV
k01+Iqw90KiHnF10qy3yBEHNJm/+HloezH7pEskR5FHw3hQWy9ei+XzHG8mUAqqSHQJA5aZJ7CXG
UJj5EZGgOaftySoe4Y19Fv5gF/ZvQnmLMfSHVY/N46sRfQu2iKeXEwctC9wC8CUDxnf1ARUW7QJS
o8YEV+wvHfQG54BoVNrX+Y69/c65ga2ZCMxh7+o1bbq7f2oud4TUx0GKUPtNFT/tBeoSPt5oYWHC
HxDmKef4zx2jWkYeQDIx0gHnXbDUlaMPlvQunsr3C+S+NqkS1rdQU1dJZ53KoPZExEvEca21nBLP
K4uvZ97IMRQx+fkjApkh59njuFs6L5lYpaNEtRrvA5WkgKQX+ZBU8l11ceNS4JekISOjFRoHBAPx
Xe+aAcZAOFfmJIJgbrrfKxIlJTqLAzcizMhvrN9GkkA6Nm2ADB2jaN4vVbZn1ePWQ12PmaKcNf7c
rN8s6UPahPm/Mynl35rfBBhOA3a6z6P5ekXOiZ8YVtruVpz0LoCGN84M7v1aW9pMck1PnllMGe6j
T5vT19RcF2/B+tcp4i08idcAjCOcBGAgTc12enqoqGZuYBRE76BXQ3RhpuwVi8mVQSNxVnoCsO2R
MjiXxxngrBGZ2Esy+evsW7S1XIuTjZ79i9ayqXXKpMTEfRz8nIKi2c6SmAMh+RJkY1TIFWYF9D73
sz18WtfirbiG3i0XdsWdh2cyPmGNgcxL+Gox8kQrfmFwECtjgEiy5jh/4M49QFQb6ab5d9hS4J3S
bCo/mqkhptNIKImUU6tIkqfMOJYWvwAYE4Bb1wVzRChG/R0uOzPgTVSVDs4Co2joIar8CCyhFLVB
6XcgCYfpdNEMhPu5RRZRXy65x35lzwWZzzSmjQ753FFMROrm5Vs6aakop2pToTN3Gc91zyCtn6lM
XsWamhUzgQY8VJmOtbIgb6J6XBzyc9OT5h/8JMrC+LR+Y8VmZZEBIsQdlIbZ2P6Q+D+OHJmt7ftn
9QjFWYtWB9pT/n178GHY2b/NkD6YZg0HOwf5RzePvyTJ6nHpwumHukDYTqAXHFsyvLVrw/Wa9/QP
7FInl2xRMnASi3iC73nhLWwVWa6tWeLph4kSC3nkHR3WWSjcyKbZVjiIRnnWKrDJXcgQ1/Ok0Vpx
n46nT1drxzZTxQ1jH2ds3q2udZ3+w6TKFrGLrG326QPySuz3sJpPCbqWl7ohOkGP/5IXyCUHPZkl
56PmGTk40qfOQ+H4fLlqzNUVvcsilp88ZtdCjkM+vyxuoGfnraHd0iRqcjwSzBPRgT4ykLZS129s
SGHLln4ehyErRJEjl8543UUcmlLzpIiNQtiT/zfHTe/oaBWc7lZmJzQd3LyHV+ENDKGqqckMHVxZ
UhOrebLSCikvvWqLR45To2YrhlSYbgu0vsinb0mjN22BwrFBXyI88eh9/qsjKQTCt3pVzI6wcSJh
2R3NbaNJZuM8vkfuE6dhw7JWvrcIBF/VKLFtl4i7UkBzywB5qvFwxq13CkrKARh8zDYBn4KThujK
XHv74wPly/gLU2xFdsPx9KR3WoZldhNNEj+fstHSkcFlzkyof97abO+xxwLBTvftRliAHIlhErSA
dGJ8stlf8cBQW5d24X8DAn02uTHxltTvglzAzunwMhjK+Iw6EX1cx6hG+9Ws21Q38dEbtRMeiiUx
T7FFiFg9fAVnCGtOA1Swr1yXmuJEwTVIbAL8OSZk92QNRleB5vPis8usLwCEA/ceXnaZnsbE6qBj
mUSZg33dvFKh0Ux4IYlQbGkpLj1GxrU49vtMny57LVKgAxHjJZEhR9HQTR9ig9xmGRTU+aBIGhp5
rM+x3bEoeFwmELwYX9fCiDqS9uEyuNrfeep4m13DGl4XZUjvwiwV1Wkbl3mNv2YbuPC/jLvSAPbh
5DxpYPkh5eAJlI/WAZsvWNAFycF8m1tut08KjBbm84EgaCa1e5kYO0aT5CB3L1tiryUTL7cnavz8
5LHhIRhPVk2dQDNEkznbypKUESNkn9bGaUUNTRpMRCcGTdSI/nQ2X2O6cG+0s7mZTBK65FmeFHFG
52XS8gGTY9kEzxzR0SlFZVggUmHJC70oajCxwQFbbmpXVJjUnM9blTU7n26FnHu/aXUfpIxbNrLx
PdsUl0XE8GObPziPAhsSdsapgIweT33Qozx2xW0CnkJo5jcKzbHvQIccaueFOW/ZBoFF7uuOswMj
Iix7BOwntoB/Dh/CrqJZmrKJKd0oZ19l0FM5bPeB4eGDdbHyR76PL2NIuwE2+cWiHdOkYHmmncJq
INojKlUCU31G1siozszs8/uFFKL3P875JO/mlo1fBaLvC7C5CSW2owD9tCj0Eqk+KuOrgcHZQGG5
MWXLYD3oT2CvbJneoIeUuQbrFvA8WYBG7kPSQ1LjRLeLQ5gzMjyYf9aV95G565/tZz19YxVTkBfw
BpNoZ+ku0UqrPchiKrUoWRIhfnM4AvqVA4h4EIzyNfxBkEVG6PcFvWdW26EJ0P1QdmzAKsceVe8c
ytYptupHiFm8OdFVVFMQGBedqVQm12J9eQ8eauNBtkyKHTZES7ROh8+6ZLsErWYDa0/0/4AkN+GK
XLg+QJM1Im8v5Y5GrpmNM1wGTvQhBPJ0Lh4qwKlZF3z3x43UAZNeVFk80Ctbg1Z731aO6sKknNiL
R8aLi13ZIRnpkc/gQhOEkGPJNNqiNJLZBsxc+/E8W9irta28qVnuQxq7+MAAprfbk413ZD0x53Nq
690Yg3ePjCMoV5Aqp7JfXqXlANJnEacja59QD8Vext951s9ySWndySoVzfzlRE9P60scOpOxEKMl
8HKMVbgetd1/QHL8ofyEzn4XbQllGEWdqZdwDEzkEbNLWFNoTtX29xgJDXLZmoXjP8Auu2Kjm+Zk
Moum3aRgA+TzBPjrXMZhmgMhLaQgSqC6qOR0SW4eaFVSyFGogjkrORpVqLnAqB+PCOAApY+x2U+x
1j+LvvdaGLAKJCKacjUuz9n37IjjkEBpJOGqnrSgtD3YKSkMXw7e5pHDIh6gXlyG/hCYe+rqGjqm
z3O8vG4OqVYBLmr0s+0iomWyqJhS86QtD50ESLkG53D1k88COaxvmksRPLaJ/KMlYrpEVOCqUS1I
jgaybWSp/duNwZSQbjKUsRZ+CK3s2ZWkJNRZPG5RQlGOC+EUBZf/nb0dEiTRohlvAhvn6wKmJ4BT
lHR28QKnisHifpuTEQ/A8Xtz/VVuQdv+LzpJJBEWpTz9WluRauUl1QjU3H/dgDwMMZ+JPAlL62bP
8ytHOlWl6L2Ar4eq/b61hAT2COc2eWyVWK+9+Sb0vrh3EpNiPvEN2IUymu9svNWXVLd7QvZXN0ws
L5twHHeWU/o0v46dhNmG/aCHLwUPlO1Yo3m3VsqzXm7BIFndTGjU7IvNMDc0e/6pRr6CYsDUJc5m
zGnPiJ+scqHz1/8kpvk/Z065ZPEQ9jtbpm4+Ok+y5FkdgkzUqGv/XXatWKCDJ4efb/LuFwrwDFyI
sKprfLKE+8D/3d7MWecKwlCpgpt58u4eCOkMcKosQbQgihqIWDYS8R+k57gryd6UXBKBPWMqSMAB
X3BuJY3+nYPFDWgseho5MU6XOvnLRg24489ruiu6rMwP+Wa05zl86a69slkgJp+lGZJvQTfCME5B
BJZKFpYSv1zCgUgbEKpqeNvj/hXh9ygXmm37MdgFH0ES7/01e5D+J82YrGKnuWOZpuA6i7YcBlC6
Zhpmn1xPERWVf9NzUy93g5EGoVMm/wvYJEnQzH6m3XW87oh0fwtajl10vquMZELOBRUQulmAKfq0
jItg1L1WJgOLCHXtbAio92a3hdQfc77lsLQ7izwE0IdbAmCFqQxU09l/9+AV+fvhPk4saT3YejUQ
1n5CdRWvC6cFpl9sAJwWsHrK3t4rIv/LC9xOBDB36pe7PxDSKXvIRyLxwaqj3lJgTn6+dHg+WL+B
KiK+AbD4MVUCW7niYc2MeqlLOMwk0MxYui9xvvjWwVIcb5qfSZZxD1a5IxdrdT1La1ECt0gQVMm0
GTGhE1ZmyJEoacGC3VxZbcTWunIyPAhHAHyHiJo1OpDb8ThuCqWKZIXIeVz1zACfjyWhnUAygXK0
DQcoF5xdXBkQ7/czlHJSjXv1mdRWWf2rU+Y5S2SbauTtCo460YVA4qS5Ll4Vco0z2KksfJKKxZpe
KrpPENXWrPAJdm+/7GNgvKJp9FQ16LIfDbFIuKIw/5+Wl9UtZ5nGpsZHTm7M1uTdSw1gR0lJz5I+
bAOfvI+WyNP0oH0bql3tc8+Wk7EGmThcD7M9e1wZ9UKmL3dhl/4NWrlFEEb3H85op8IAqFDo0LCB
cWQPEqp8p/NGdoO+X83ZzXbf88JHec6rMcWsBi0G9fFNAyEgufs1HsqeiMOYUiXMS9WBrkhiBd7t
eml8dioyXm0wEVQ7juBHjrPT0fvbof89YiQX1GjKFXjcgSfWozqdcwfxv76Cx3776CDr/CUn400+
w1RAKqMdZ291hMVN1smo7iA8wOTsdxwFIR2AAiFGpVaVZ8LfSgd2HxmGrTgNN1NmfzFQ5KDgH7rd
ovqlyzNuwwOZfoZ7xPuADJNT4nTpYldx3sjLxMv3TV9F/x6z7P03YXWoGg4NGdpbeYKWI7qatnBw
vSDb002eTne4jNCvCcGwiUNyrCuX4sRbFOlJALdOhbuQNUhEBIRhQfucgCw0YfF+tItjpgt8d00f
LUuYrAOFN65Kccdaz0/nO0h31uQ5ErYwvCm+bseo6u/QyE89EhhYOnlJcfjs/UTaeB1dHsJTTa1n
3E9n16G2RsOCPf4i7+odL+JKKQ2DL+2QTfnfoVwDNiFn6lkvKAts3QUS3iJe5EFUM8y5f55k6uOP
yDS9t0QRUyYarEyS5KK1CUrVGqi60uE3UZxSzv7Le6JN0iO9XVw92ePU6PXZbMslDlvVZ55oKPXA
0gkDxh5Dlf0KdJW81MTd69+l3vUFwJ0XZOsbycdM/5cUf6buyc54hNSyQMu7iAXNLA8WT5SZIGvp
nwmIu/C8nTm4tdGNgCl5cABgJC7wWhngM+Wnfw5gvRUFxypETAy/MHntmLLb/AjvCIWihMoA1/5D
cYjlQBj7eBf/G3C8UCU3hpTdwwiTEzzq6mEVke7ed7bkKLzbQd3HqvWxRHEt1IGXGOxC7atqlwpO
T7dSw8tQZa2fYf6uNPugvJ4OTqjwBOwOhtxh3a3rn82WIsO8rrG5c3BUTRPZ2hZEVAkSt5XNg1JO
ufRPtEaIr8ugqPzBHx8/xJ2f/LDs/7wb4aLPcwnW4hlj8mcijrlAztf4SwY5dIL1wmj4B/KD3MLH
rRgpnAppFW6lAxpZpk0PhwPCfWovJ5NbfgsazJrLWYRf35XGmzjAW73Vdj0GUX088SvWRP+qvd65
V0wLEyZ7yRGutf0Q101MrrKuWncV79/HGLm67ySfNtAPbEY2eS9DWTQmhXPp47BMxEz5WAYhiB9/
B2LOUMaZ6gngsu3wQM/ro4Nlt8pQL4m+wFAWM7AhEsYMsJbvLt29nh7tDBSIKKyY9ItVuKS0rCGA
FmxAfLRxkAaBJOhiNW29UeIwD0ee+PKzp9pKy7209WQ+OA5Pfx9BYRbsrVIjGu6/way0x8IoGAIy
7WSOG4MvpvcGUiF1IkMy5hTULaZqrFq58e5+oYVrzHGbF6IRl+Q0CsoCY0sT3e0xO7I+eDvmy8Fq
c9Zf+d6A77drr0Zm32Xa9AC7DmHiXBMN+ztdxr7DSftNKBmcv6BXW7zzYJXfGA6BPOAe2VUef9B0
6VZc7zly9B9EtkyKw4T9yruTrc7Y0upHWPjxZOO8JUv5JWGDRDrRq5TzkBvTFicobb0aDdUUA5Y+
gOPT2AywdKYZKniwWic68rA0SNSAvTOZsIgCkGx3ZHeG6QZ/4ku1T8E9RngIXDCVFQT+mBCUPDFa
V0E4u9yrMWO37V6OdjuDfnnA+HtnylJ63nxbRydRLmoQqd2E0lMnZKTirJ9LFUYx3F2YtLL4+Kgl
2eV+NWWjBpdxOtfiW+z0yM0uNbbHD2OfLso9g1oBxnAIaj60BxLZyiMPvAQDF8FHypgx8hqTJ9rW
8tf9XtKdHRq9TFqLtudGiI6nsUUv9pmwNkUcoKFWag64BiliT3vMRYKVhQE9YbtMgg6gSRkQjY3o
/lMcA4vms3N85ZGyzUFMk5DFv4A2b6xLCOSqI9nVPdMcJQArSUV0UOUQGkejwA2sCWXXz7Iy1Vwd
7KM58Gb528tO7qpRZr4k//PCIXjDrry6lDJEavGb3vDYZ2PBIYCDhvwRJlRf7mDxA2MqwK20LDdq
mq/asJjB7wX62OxcFJtcC5YJGUJMUr4uHBwhqCrD3ZagrUyvyAgUKN+XaoeIuvMu4LTg7kM/9zxF
MGKazfboZrj2fVKt9jMQISDr3Th1iOGcQ1O4gwh3Rxb62RUVxGg1Vqlx1nPVpGEfsGcH8AZ7dCSY
6U5jmVpH948zlX/yiWa6oU/E3/CLassS8TBP2EgYTjsE1JYdPp4Grrf23hMLO/aRcHzJgC9qmeBa
9PsuUEkaD/L884tt3j9zbOQROBHCPequEVK4+icc2xo9Nqv9BVop5uWskydwM9CaoD9tcWHUc3VU
BHZkUm71VcmN94l4Vxcf5YKMdh6Pb9U5bDPTsd5d154f3Gj/iZDpRV9dA0mErpUsV/hq9xqb77Ts
63ksjtRqD5K2pB1VZDGjXo/xImM1jqYse0CUeV+IecSftBWRaJPPu1o3fwLsb7iHyZWklcjpi+zG
tiNUvpvQhLPIg4GomQZic8LCU9nY/HWs0qL5rZwite1GDHz5wlQSwXwmGIWeLWyeI8Ecpr0ZBkez
QvmYCC74MJVUJQg4T170cyFU//O/IuYSd0wHqJpYPpJGOnlcAe4U80ijK6AMTrQuEK4Qmw/alpl8
jur6sMEAkg7+g3MUP8T1M/5no45g4AqHFmmBKQNuNMxNgVgiv8I/yooZaIeAjGM2yyza+23P5juO
LIDE+9uDXV50X//L2bo0YsHyGfbNQqOXFlddu1jESzg8Aa39gxel70EtGBFyP+Xu3xTGWfHgI5c4
RazTViqm5C6y/ve0n1t+0jdPW3pFO7T0aJb26tUbHnhwAnYh0mCXFLdgktxe8jEoIPWoYUWgY5rQ
FNQdDnZtqpajRxCI6k1il90teF+314dM97m69caFgLgGcdso7AOSY6FfpPxDEUMu8pX46XS3Zg0/
cskKc6UxOj0hNhs5gDdovuxL3wLn/bHDXVEMSqyz4GUunZhcb9KPQUw6ROw1T9c/Bab48mpN9CoE
D1fubhyr/mg1jhjRF+Xkhn04Jibf+ul+sk0wMHNNTRxCz7x6eQ7iCdbngWiDkgpRjSVLLgoLf8u0
xU7rDRkLZik/nTey3dzSkfo4YUPaGDlv+2EYg18ZVF6bHnmxvf6qc+AXfLCq5PCjtJ5yZS9rZxjx
6WS6P8sgvp8cXrR28++go4omNUnSrtUNymShSTVGJfhgDJ+z857q8B47nD4VC9f7ACI5SzTw3qRW
NqUzJ10V2iEiJydi37PVFtvi4aBAV77p0EIrhCRxrSdBht5Wo5iYQ9hrMZ4EMKcL13PloYoKwK9W
0A2NKE0Fh6ZyYAltJC4AYu2UUerbVfWP5fv0u4c9EjuAcowgZikuJaNTTvzClTMhSmuEwI7nXd+M
W5y8Rh2483Kz7UMvcavVpPL07Aa8Fs/xpDuJJjAmpaQ9jpizTxSEGw3cD02b1l9t2KOhnTY9nccQ
vLKnD2yIhjMoikMzf+Uftddu9bMm5Uhf6byrswk33ignAlOIZe1+I/BslWE1eQhHI4eNRudODBC9
TkhRVpu3M35L+01ofdGtr53X4C6YJbbB3flfhMv1z/voghhcKclREXV6HCy+f7U1skoqN1OMkKpN
E/tGiDmUJL7iu/UostjWtSObVhxUPCL/jTwthURvRIDBP6Qr1nnt7lnBKqstf9OxCmwvCEZbBTqa
xmCzTFJXldnBRYmtKz0MP2/igEIN0ku9v6+3GEgPdt7lS03ZH+GAXQjgH8DRzW2Jx8UAdrVmf1QO
04aHnYYrzGWYJiaTBF5C3MW3hav3DbvHv5QB26U8mVGzyOj0LPuK/Plo2EINpJtYdnxs9hp6wZVZ
dDOWJkL0xA768dPgHlL6oS12lBvBuJK+9kRjm53k/w+LWnXesO1hdB1d6x+/WtxYTukh7ldiuPEj
n8vRVVDplMS6cGK55tOfu+64fPJDTRlGaruM0kCzX8XIKadsCp7y/6srj/T/YfKRvyUmcP/IAGn2
ZtLRBgEQIAfWnawCe1SLNL+iIZqkOctR+Ure+TYuum/tkgc2I6uYqUWVEHissiv/ASjMgWgB1a0W
XBuXwoXWU8TWOaGWrHgKk3JZMzznqKnLIyKEnplCuzf/8+/7RL6KhpQehY4quhtdq6biZNcTVH2e
nZNedENQ4EYWQCVcaVJhPjGVh5/E3zaT5bENjI94lAfU/JHfn9trbgWTzEx8s6KV+7S4oke3+5O3
/SvXOlqlqhi/pBFoG7AVlxsjUXQtNVCmO3+5pVh9C+0h4A8Kx0wYlCWAL7BrgQ63YZGeD3oHEFkb
jhEQDhcf/HDCZwGLIatBCihvaGqgdQYu++qAFyCjQaqaj+axpFWCxGX0MQq01A3F5X3NcVTyLrE+
CJx9J9ZBVPCGgDEfGSIgHL+rS34C4Knfgw/tBNOfkdf7Q30V5YgujI717eamCiPalP8fdEpgGCUw
aYxZPmBuxm1xURH7j2BY+yo+KGS/DsQYe9GCObwLZvksW5MVzmU9P7Tfgzu+YP/RXx0vtOmDtE9b
3wvy4OcRXLVWwBpejfiUhfT2c9u2zU2OadSe6IfhBn5h8QxZEikOVi/OkyE3zlwX5JuBO8f8njfT
aFp9oWLCrXtPxW9nDUMhdytR1jb/wNJiqYhJg1RGGoaEzLYjYRQr+ivECeV8Vvx8VtlQsE1/e0KM
SC4khtZApVW5Bwoi7aHx848CgxeV0eHU21OSUkXHBxDvChu1aYTgb577snc3jRb9hPMJy5Nqt94/
9UQCRVEUZl5u25GjvdbSu+dywy79Aq/IWhkM9mUlPzD/h1scTnEjo0qlvoesch/HM9KAXnL0MCEM
9Fra3V3XlVSIjuSES09/OOQU4n1kkyTIcF6w18rUjm0XDs0EsHd5k0RuNuw8E3XhIQ61iSG9QDFD
7JSNK7+sf8w+nSZ9G6u7g5y4oh9yIXutqnqpvxZKxV9uk6QI3QHDi0iFX9DzYLlDFUPmb56bGuVW
fUPdldZUyBuEEx527qdgEOYYOmY/L5Q01CUql/fN3eDZ4EjmsWOrNtIikThbq3hwfe76LD4xUaja
Q5Mm7pBQa29BYktY5u9RHo/Bzgh/xXlyI5fCJpOa9rXpT3Sq87qt0vBxlIrele3wh/lc2z+XySCr
HRCwuWx34b187wcraJXvcLlbpmJuwtw6kthJgOrXk/w2EzqTo2DajbtUha6mzME1yfCotoxxeb8X
b9E3goD4BczCm68khU32+QcAHyb9aF4lG/dNAlrSgB5jbVhJsWluNu7BP5B22855V+T0V0PIZ6hX
qz/eY3tA19rpgOJBlkfsUDTT+vE2t82MA60wR6os20E58T3dPjSuv+qRuynFhTXoCfe3m1i/AuVE
nfvQbPYZJh21mr9aMcay4ca9mKHn9vwA7nEl22L3EVN8qmwa/rg7sGPNiEF8KQ6xPEh/eav07q6G
AFXbSaQmYB8l7sbtTXqFkHn+pQc+o+4qcSmWIalHdmKynANK5zqMcX/q/txaPQSETUPrSZ4gCnOW
33lbPEffZUWR/l5v+MAyRby7/6ejTVJsA2/djEg+Xp61M/SkuwxDs0xEUqiBXB7GQgRhWj5t6Rk7
XJg0Ez5JCCvoa+FOFJPCWguin3bo8j6PdHKajms8+fmP5YvY6rE/s4bPth9+UxanJccm+Hg+5V5l
1eD+p/X5Os4HnOQ3E2HroJuXMwo5pD0rMc4d/Wf+3kmBLznTNlusGoqrx/DrjiIhZNMzotDs+ycB
8r6EnnAI9hA1LUeyZFUWqZ9pbipLiax76Sy6B1vMRER3BFmO8GWrzZ/Z59HmB2DAVUNn0BTuqIfb
JpJQrVnD+G+r5dMx9lp3XWTNku/so5e7LW0DkXGN7soIQ2DKwKoqk3YGAuGDIpHUYE69swcPU0h3
9ZqwxEzxb0DmAhxGe6T8HBMNtQhzSe3ltMZ+tjAQVRCQhEh7t0KPHo0saNrbzbmLHQIt/m9AYXuD
uBGK4qC7vybRT3iLeZ18CymzeQlgU+nJsiYFMZKdON1dOY96CEx9qqewpQHOHF+JH5gRd3xCAxn2
WMpyqWvsuCd6Df6IlC9zHYx92/9p7XOHmsJqxAhFOJD+KvT/RfcQ+6cG/BN204GQD7yz3qTSjXnh
7PtqCljFA1ZdR4R5qhfUjtQcXjbY63eQSpOkz3Yu/BrXMDSYoXpeWJjA0JrXKengh6TNg6MJMqUZ
vtWsZyRNb+IE3yszqarK1O0G7vVYZ/4eZcrbSmEFF177N37ZTBGaWF6C8XDCsIT55/8byxYV9hwi
1Z5RNWVj/NEWmcugm3xUrCsvFv36xf/2TwswcTs07qOax6RH+IHGKY/Huzz82p+FX6BPOnUi4L18
ebKAWtGtEkkL4YmllGFgYSot3MC4+lLai/z4pCOKE2FTkaw2/n3G3Z6F8Oumhar4NatyW93+a+8v
H6S40ShfExRuvSnFdYqVB3oSLHaz4z7O8HDLmIxvxURTIF7paQpBfmTnWgwLr+ju8XCMuaEdKiqX
zij9i/civ8GzcGSW+Y5Jbsy0BIaqt0OsYouFgdAvN/1Lwy1GnVf4m2wYxBnva7jZcXJI9bOdgODo
9LrRfJCsNBRDmH+kfUIl3j0ZxLJYNZnAFJL/RT8isCuFbgWZsNFSn9qW10CZqu4YmaoZLv3iPTpj
9IdYyqC9du7rMw+zSdMApB5Xl2FPRAFCRhfZCmpP7UaofDW/qR/By79ywSNT2VErTu2kM/XnzDX9
kBRtNxmUl9dvoRGZ1E8EC8Uvxi07Y71W4kShFVS1VRbKB8XXB1SpHo0hX8JtgUDXkEj/4nxujgqI
PC6vbnL6waI6KwWpj+UJcuA+F/icC1xTHaj5YfKu8vbZhDbMX4b42rIJ/tse2iO228kqApcl+b6i
f8nGL7F1PZfoBzEB/8OAkfeKr6qxHA1rSHNlcemFNsgJMFndI1/qngUvmKm2vvZ2FL+irWuc5+VD
crL+CyaXu+Ivpyy58wdaAraSW3lBytQ3yWMHGh1GUweFaps/V7JzLQyjTdCh7xixiNeUX/GzaFFM
RB2gKcY97kTCcCf+alW2qyBoDY+aXg5xE3ytNycS5hTjMJVSvx+oUgXY8qyrskfAtSKpvwDmI1AJ
UToMK2HCMZqe0+x2+AbxmBvLmaBL/K/C9+oIed+YdFTA6LrY+pKc1SddaTf3zYTFB6K7bvDcRU4B
G9pBcpmp+Kc4e6+Nv+GMrN0GFFyXxftV895uafbazhWTlmOv7jUOD4o+zn/wBHT6SaYbgoZmJPzs
hpKcSUItXR1RpFRsHWMqrP7IIonJACBBeZqHZ7tZfITJv1ueIoIqa1nvzj57CLmfTKAGA9Keb7uU
1gloHhroNoonAB/Sv1szSnQDb8ECx+unhIMc3O0D77liUcGX9xPp7vujPCbLa7rVt/fexB9CvS9I
2mlhJmxu6QtY/Dbm564+/IePNty2HW9pHzVu2apCNSvYCTlQLsb9Gvh2SrYJ4Kw4OZ0TNFmhpUpT
R82we/2x5GE8/2xS3oJfzcUCPwo+XfQ7UsXrm7AMuEzU+EW0dHOfpuY0TTV/pJKXO+8u7B0MkoJC
DmL2BBcaLKhCWxSd20x3i0WZsZanlZn75++aFXUCX1PubtwfNGoLPgfpcYwW4AeXZn0oSowXd5rZ
oTMS9XI5JA2T/9A+kv4kOoBtfBBLRJSTy6WSz/4gU7FlPuKbAlaxT1VbgKCuqck/KQEeJWtHDRY3
QSxQYnrlWn+H6wv0H1F/8L1uAPTOn8m+JSYH7CixpKDjYqdUFWQv7y5JE8owWpuGHu6qZnKgefWM
dqL3MRgNbZ8rapH2fAdQhOr5R0jAUCPGa/fw/PHl2vmf+iQf0ONg+2/enKGNrbeXGGiXrnl3M21/
xFrg6vl0y1Zs0fm0AjnXZ+vo6pWns9PMyoJ3qXWvTcar6mKf8RmcWfqHM923gCAqyb1mv89mb/l3
e93BqWYF7Bon2+aafoLJVYhOrKnGXnrCyfTWQOhelB2JJYYlxjpL0103ri/0NhLML0DuJmhXNpVQ
BDHajsc/NqUZ1fBIpDCqTyXg9Hi7u274w+qG002NmfSaE0unIGSZ/C7wuc3CBjso+g5rOjzbC1mz
Ed1IzxE1v8jwA102qoo0oSHhaQjNPQhuS4tjUATZptiUKRiWz0DYI2CyXHwr1700oDp0zWpB3Il9
h12h99b9BpQ5YfreI4HaNOwq/yIaymu4OC+DIGb75bqIvLWwWUWTXTSS4+sRX9zUGrLAFw8aAV2b
qTu7mgcN1Ceq3fCAoUouUY2EZsOfilVUoy8X42lq4Fr/M8gL5Q2rjkC69LhwrAyTm8jQDjLrSKcp
EdQ+H5VIFeco3SYrlv0U1MWYKMV0uG0uSKPNlspIjxxWYD8rskWuQxjdDC+rGTYHEw18Vzw+sled
MI7zMlrOT1iv4yUnZ5QmMA+KIXkJq1ECThbdJY6qMbXNqYNJHDE0cYHoDqVFI+ILf37P3cDTNM+Q
S08dl8YXbQ7Nc6bWEY9Fes/QDTnZ39CnYy5ILSJnVC0CHKnUfE/abAbCMeFeIGwikvOga5kOAHd4
SXTI8H1+Gt7iPHr+ggISXmf6EyVRynEE5ShUfZ5qv5K19xTylJmAzHJzS6u+gcgwnIX0v3CZaIUg
YRB/MnCrunQMeguoTk/rvRsugl27vJEnaG+CKrby1/U9jxzjc5Vm9i9h/P+A+A0wi2Qj78MfGEdI
/XPYAzUu3NcpOwsGxu5y/WiUi2nHhY0bNDF9gmxXnJxFwx6qommY7DShOR1Xckk4WHG6ATUjI2Je
5jDwQ2Gx5NZdJgZ9lQiEpXDt4cpUFhD0+/P3E08FBXP4k9EHzA1AN4HJAs323c+gRRBPdNwwft2A
aPbAyzRuO7cq6OeKMQstW16J1MzQKJUCh0UmBc4UcBOHZicJdaDcujQc01b3/w0V2/q2Z0Dqe08F
62mW/0BO6RMyXuJNIHkHHxS5GnlBpQegvBMihFzNFzze830YAM5x6XUI4pTC4vbpnVNAvDiS5gZd
IGRIM9Ebvt5nuyo2hx7YXH5Sow0LpT3az15KKgzozmAmpPm0F6m+1TmJ+pKRrVVBw8I1luKhF178
RfFYXUF2U1C7jSwzGxZXfFBHkqblFr08ezzkbQyVHjqJD1DF8nYTpR9pTnAeqkCStNrKAWrtPtfc
7G0/f4DnfBpY+vJ7fb8ELh9HNtA5nC+8F4bF1PBlF0Ezsa6aHWfy361CACgtPSzIZP6uMZ+JPw7j
eZ4j/LtImy5xl65TJSaCXJLnMPxDlyKgfqWnHdM8fhiIscLrwn7pUyhQwKoSeSbkUBAzwrUA3eri
peXWJn0isqmyYMHcXtFZ+LGOS/PNP0Vk/mWgLr6wec8RSAf5Js9J27PpIlQky0q7WeVTQRrmuZlH
rCV1bz/JcTqtSoEovZhlVIyizuyEEGBTSYde1fQX+WdAFM8YtNgCysSL9/z1tpzVUHoA57Ug9Inr
bAiWJ8kM9v8RO2KAAEWW1bQzQDlwBXvP1s4xYQGe6dVY/9MZV8tdKPKopeb0kXfTaJrNEK0/lEqL
qEMzDVEzAdVvK4gwCEHo2yfVPwa+JAsKRUtSeOYKmQ5mWO8IuDKWkMwyMAwKIFJHxex3tOLgDoo5
/2Ykj7tW3Y2RXvScAGieuQjqSUTGfSxh1UlUnWgmbHwwdYU+5m+JvmmG7PrniW+kpk7ePGzVf4B4
kgf6nYBtUWL6zc7rM25U/nKNjR8YgIClpC3jpCC85T38CXfceWjQhoGDGjjMl96o6he5vbop45ac
R7ciqXjaqaQRBV9QPG12OC5guUmTZwx+DUbJQ/e6HwYPmOx3Q6/cd59PtKyqLjmPNvnvLymfvY4l
f9Q+eFH5OMaZT1lMWoGx+yYWKmXMDEZiXDsfDZ0FDodzqaO9ajreeRYWCH+msqFF+L6wgaYwMI/C
bkt21OrQgoLo6DU+8xqOEHDORcZYn6H7RMLALxQP/abRF0UQgIpprbk43O1A8Jc2tBz3v/iChEkg
wxAdS1eIkb2LXg19et+Nf/ucUY07fDECpCVNZVT9vAHFFhISDFTOT4knLx1Kf83o3V+n8Ri0xfhf
spj+B3zz2D4ybq4kcZ/MV3TgiF+w/I70NxseLAWfmp3Vfmv1dPu3UTO58ksqlZteB2zJDTYQVd98
/7sU7ms83nHBJmvf2X7fty7f6rR9hU4kQIxJal2txd0hNXIu4SMUpd5XE9VwUkEe+KqPC3n+LJkf
PRJoOwyb9eenD/vMnEnTwQUrdeLCOQhq0mCF+uDgV3P0TpX/SIEv7cpqcicOTcO4Qm9RnT3gPzX3
K5xDweVge/uGnBiOoFtI7qtHiGiMBTK4ACv3jMqQE6C0jrvDKp2DNrJ0LXs8SRcak84lGnnSWiUH
/kteZq/dCYGmEuTikqJxhvmXQDg28S7rtxLoYbMY+h7wdMTOUhBb4NNNnB7pGJkF/qAO+2iV6crb
Zp05OMWouIqjw1WZpb/nkZkjJBVm5mXpXUKBinHN6pGPkSE9V0G1CbeI1zZ6g6S7izK8IUvCU0F7
iA9sa+gC2n+2tlIc4PMVH7n+Pyqfga+WfKNG0aPvuqOHeOpaq91m+EcsLtL2tN3u385U2LB1zBRo
J5Y94x0ZP9gczOZpB3JB6pJqn2Qk8XVuJLgbpR6MB1/qyjuH2L3Uo8hTOmCDHIOVzYKFTauqhD9j
eUHIYfu0rVtgQnHGouj6JPqvSU/oaQvEpiMSFokF8LjmQrEi5G1EpZAWidKT3deEvBeqX87zqAUM
12Tx0jd0ToLUGb93rV3m72nN+7bN6FOwCU8UN1ilKPz0pl2+m82IApHlwGO08UZ3DiHB0jG6y5WZ
TqIEwiMvSAouV99zu7uTFuIXxW3Kp7L96ehjt3pv2QJUwrdKhJJZdsMfvrP00iVrw7fgqNQW9hEc
nz2QNQayKpt51uh7X0XYN7SFeljUDXh9wOdypUuJkl0npsQNoljxuBeVXI136WRRfOBMjJLWA+1V
/HmXaV+t4tuVccx48aZZ73mHxE++C2J9AJpvDjK4FZhOhOzofIQpGEAnkkCjwlkfRMxlArR28CBL
xST4Y/d5w+FWpRuMpTHmyaPoREMNfAubJHmkNenOa9LVr4KLUndnfZ5qrKKe2uuaMzMoc2vjHrxM
BQmeR/iZAXQdGn3y3IuPXmdG5vlj5tsiHw41FU5iEgOyuxpnWLLtDjQF8B+AaGu69hc3Vka2PjjP
/kLVbFh0BxtFcs7buu/X51nBtRtOFr+Ld5V/trHP14aIjLkhjWNzZsYs7KGrkXWMJmYQc+1jbjkL
f2lzo6FBAd08K9QFRbYaE4S870SCXypjYuVSPOA/cG1jQ4fmjnLeh9JFImPTaBw0J3bmhFvlOXO/
IjcpPBy5Rg6IkYwWXbvRoJsTsxRlcURZq5zNRqS39M+CJmLvd9+EZ+Qlchq5LKQiMQqXOUk3dKQD
ylQpXoo4GCh5Kpc13okP6uwM1QWpx/wwkOfvOFOyvfYLtJ6agxklz8PTCAEo3psikSOKxzzJuJVE
PPCkLcZpXXX+OXUifPdYMJiJe4b0fxlkZSMAZh8na1tM7D0ORbMUtqctMKDgraZE8VVtCf9SHSGx
pgqcz5vAcPfEVOL6KEQ+nY3jMPMehmDqUjeQRYeaVKS5tkWv1hXJ17Ct5QdCdp0nsjD1WG8u3JaF
lkndsDDu9NqCcBkYVGZw86Gy8jifcIIOSKTOOskgd9+7tVfI+W6b0FTRxr5gRq/fxDOncRNKyAPz
Neo30KCC6aJ1rubYHR2AyyihPITH3dM90XLfX/MsBfjJeqprH0l7LHfUdT399fYFc+EnpkUjFtAl
Ve2Gr9zwNWQnL4raV/j2zaq6LYTFAfaqA4YGzD44ni0SSvJqdSsjrC+a46/8yKJ67stFNyfZkxVS
07jCdoj8+N7ZolKSyy5JY4Mq48R0jMFI6B1qRgCtOb4cimVILHhrp/umh9IUx7Q0TuvYEobDe4cK
73ROtdCPh50ZyY6pEQhGd0ZyUEH+cPn5Q+OfP9Xi9Sm3tRIMZtS6MVAfMZEOSCqcpnMP4j0S6uVD
J8LRKaupGnoY9tDzeZFX7CZ7t2hA69v7F5XAREfKC42S/YaGI3kcuRHOZEaRtM8TgQJ8UUUNTVf9
+oHRl41OigaI4ackC848IT6SwMKy0nTyvnwqKw5BqB2AwVP5TIhVWpwNMJVRJCYbZEZF60/N9hFW
JzEbj/GtKlCJyIFzT3v+KX5OxXYd0/XDa+53FleqYWrxtWTGaQRhMC1OUpMOzxPgMcpVSueKIImL
l98Io788w2uRqC2bFIETUSAM3CnvkkXY/Hfwb7hRHrJbrb85zGwujGrXsYfBMxQYwFwzj8vlrOlk
eud273fEfgBXWkqUalXvcHO3fzYdeWXdnPQxpsjSEF1ySR3SbGtX66lZhcJJSMW3DME55gNuh3uF
AZzyr3SQPs003B/5Q1AjJH+Armw9qC/j1Dgo/oBHj5q87fHluqBD95uJZl9u1Iy+DvqcGr5hWyP2
B0P7Md6fZFTPsSMJ9RCUYzJCwWSLv6Ingek6M+uFginHeyE0UMryLFinBE53TzlG2YB8WcwFnmoK
puLz08EqtSr4v9r6uiQR+AgatdV3C/L5OPD8ZeRAljZTIcUkbM7OAFllbVyUAU1a/rOUJrDMZE+X
56adRpjFJYKlNkHe74SqnO4cjbjjL6JUyY4DTuOvfNVhoYqMFNALL4axLysC437ZRzc77hGVdG/G
gG9DBXqqu19opDjjV096GYwIRDeV83F+TcyNjyYSMdYZ9Uwx6+U1rM46537joXgEyfZkjLNrcFof
HQXYKvea5W7s1mg6mId7SIBkCYvXSOgfqsDSnn3JZIQLlhEpFFjmWw8XQmuf/LxnAF3NQnKZDqqG
Q+x2RApJeEJPCdNhlm76gQINQSYRE8kVz1LMhrmBX2OHt0YcoG9ap2BrC5gfQWA7E4u3iW3vg/Qf
JCZuV3bECv1OxKA1tXJ6aEBuqyOEvjya9Kfezfi1fbqFlsgotl6dCbHmH/gAz/9YeQ6PYSZ+mUTj
22K60cKpLtPB3deLB7pcA63CrM40mVRqOwCV4CEu5ywfXn9wZB3mjXeQtubAcxPcGj7KzD91gk3z
cqJ7ijIMK/jg7jq7sVFy7pXZxAsPD88LX4UpPGK1haUIzq/AhHP/ngJISy/XekXjAJATtaqheuui
wpjOfbQxLsDS6dY7ED2YZCu+jQUwqItZ2DFUjmX7ofTwq8uapeIzQrQ75y4/Hy757WBBaAU3YZt5
GXwW6a+5UN3m5YIMxaMxW24t2f700JREBA001fvNnngkrElTwS30WM7NY+RGHP6CFURUm9RVNyHa
0VpR10ixApBFMB5aJGXR8hCkcJMmCj8tpkPZCkoBhGRKRNFjpDTdZ9WlQGHHLmwx9N8G/UozXN9L
0zRaF4O9Nk4LS2caLosywC5UfaFdpedcDNZRzNF2L9CfZEkxxDshJxCkPINjx8eD7caddG5BfKN1
p4WD2wFewp2CCAhCiab2D3mGXKZKd5QH0kCu6efHW59SpSNQY1yOZ7wp365nqEAw9K/AU3XVx35/
ix9QwOlOcQ08gGLZqk+DUmhqqb3a6bzk6IqxrT2QAY0Cw3ijhKI=
`protect end_protected
