`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPIim/zik83qF1bAgy6AN1G8KcbBgBForHAD6Q+9EDfPEHH6piR+6OWF0NU2yfFYzbcH3DA2skrx
vDJRZAj1Ig==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mTABHRrMPkm17gtYXKunPuFSfnng1BjQsQ0F3V11aM5fKjnYtLrdY4sS+tvU2FpTqZmP1Sa/Qiv9
3TMxHPo5BsNEav7oebaQoYKdYLXC7EdoJHMvv1obEmHUT5WtgO2a9Gt4HNpA6Et1ALUTU5uX231F
OuL4i9hXz04huZQGbAw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UB5iFriv5ddiFCKNaQdxkp8v9ixxJbRIOKYfF4H0oLazviBii8ZM9F9+sIvlflB9kFQHusHOvI+7
WQyaM/ua6Fbxe3fANfyIgRjSHwz6e8FK5Cxlb9TRSl5BQzj89NbXpbLop5FC5NkMOfPbsnsHxz8j
KOCe1cT6iCopOBp2fqgBbNx4HkGtFJMIK95Vcci5nys82V+Fwaqa+ahMa8U9ol4u77nwIjsUwhGs
ZVfgzJKp2Yc+1dCuHPUMJ+8f+L5Uh/hYAri7Iw4JyoIFZQV7V0I1XL8YIUPelZDqrgx3Y/gD635h
nsn8kLv7NUA0fF+AZcDsi7Eo7EsFSOB1CNmWKQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o02veAooeO9Ye9ltvalUYz4ljEBE2PlEJwaWMEgk7QbaUXh4VNkLRlVLc/5Jmm26c5DukaKPGsRb
UOd48KnfXlZyMyDI+FmaNAcDHsRNK0byS/ncmDRLdZY5bTVUgJ6prERuCSJxeW9eOPV0A+6JQ6A4
aCBY5V0+P7Re/G0UTF8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AC1vMV6byaT3/3Eo9C6NpeReUGL2DFlq+mO3Y+TMrEztydmLeH6v51+mHOER7Q09NDO+fxiiG57T
0pecla/PwpYXAXL272tashQQ/bH17t3IaOPNu6VvabwHBjdESRdtPlyE7mHAEVT6KK+t+/aQHy9u
aWdoB4pUCeCOGa7XWgITIgJuHiGRzFUaOzhRMenjcw39vjkRmaCt0BTsubNMOLX0CNBggoNes1te
/9I8D3aLp29Mr27AJfclsccMT3AGaNDYF/wD+ogr2GLcNANVSzn78PhWXcJ4vuZidM+efgQfk7r3
BfKjj/6KRLM1FI0piKx5Ivv8FrqXnKf/YU/rPA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22400)
`protect data_block
zQThjk7e7F+4fP0BoG5Wce87lE+i5EPaAgJogAfc3TV3/5mS0QsdYHk92HUpkWRz7Gu8ujMTvbKa
swzcyaw5UL0Nf2txJCxKvKmAGrmwqymZyZu6HQxZgSOvntAWNH8EpOs6VPQaS3k8yUd05cG2ZXgA
OCJfPb0EodSOCecKNgR8/bIWDHQt4fMWNi+JlZsA93M86Ta6ZA74W/PF++pF2KC4DyGzW4IZVH2w
5AueIgcUvEUPjb6XCEoVyjvNjTQGpo6NcY3gFNsCFizO0vH7SNhX87281qGmCBSSeIIo57DhsPP/
UxN00RTPST7I25DjKbQJy39Ue/DlDkvi31Mox4WgQg6cR290U0uIrZRbbL9Ooa3SJYFgqPuwz3qG
1p4EpwkAaoDjiOqaObZcrJhQEMEpIkTrKmmD3ROGzZWUaMNe2LgVtWel6vVZGVWcIhMjK7jU28+k
EBByjXlm9QxwwyIPIgOaqalGfvQdlG2ODsE37oE6tVIvNpPwil4KaawrwFBGOuf9hEDGUTPDr897
f14hcd6NFz/O/A7DvZiaad1jAxv3RuQB546ToSw/ovxAuVExI8XG/QoaIIg3BTBB3VoeqKSU2X5a
q1ikV5TRGw/Ufz7wc8TbfMNF3gZLHskvuo/KLLW9sREYJtICMNbm+GEYXWoSKWxst8B7LcIZ0kd7
Vmm1WOeeO8+hIGsFzLY/HSIVEM5ejGjrHVMrHnA2vHlR53qXcoy/unb4vu5Hkqj5meuUOr+W+wgz
QdTU9pG6PzKL+YRuV75PDhk4+iJ6dh08eiBVxRMO1gSu2fh5iTpzxNQnjbpg1tCSwxGohFqbnsth
DY35D1wgriafPCxaLA1Ai7KrZsnN5p4vKKjPfJaCt6UFXtnDurz/ddf+vuSsszDh/zNPAIej+Vgw
fi1r6LddU5LRTtF+8RG5FYZ5OgcqF4i/eiJOV5uSTVV0Z6XRTnLrHvAQjLjVhS/dSbhYf4UD7T75
7vnIUCCcRCNFkMMYNjAEA9D2pgPCR2iMKfEaK6cNOOX9XJeEpsWMrJudkqjKlSGvW6F2ihahqpaO
HzFri2IJnTLGw0Cv99sLxsF9QfP52xe9ktKfBafjcyZlt8WHCje2B5phA0VZbUCge3+3DURS8/N0
pX8LUFYcmDgsL3GRIw6Ys6UjAjfXI6PJqD00SkKu4oR1UAtYvTNyckFS7/6IOR5w2VBkiVdtVepa
rJefjB3HM6huv6S7V5lkdFi6s0K1hFfoOzNL2aqpAW2iDxkqUm8H04f3zI0ng8SxeDORevaJ1IaD
RJc3QIf5DYvLRSXvCSO/0yBLQLdbiSfCJBzHGAnW3Qlc0dnHl8hYIf5p8C17/LXyczWaKY8oZHWO
8yngefWUi5yT8nxt3Y19GHN4Ztj+/3KdzNHyS9gtGxB00Nc+Q190JdyLTf111VggKb5M/0jOk7I/
NpArV37Cdv2Jn+WHEkLrXUXApXHRb5h+pikecMm2K+yzHU4ItZ/x9/XlSno6j7qXcLk7KcrJfYYK
0JWBI6vW43d5+IkIAiQEJz3LVkVP/5Jjj5DWthSdc/3ghocioQqhcg+MSx57XRe3UO7MVnFM/+bR
Hx7BCpbZn4Riz4I6VfeEvFR3V5qywfj8m7YCe38J6qeBs2mdudkruxmNOhRbGqRNVpMR0rQLryIN
Xo2+F6g7Ka7O6DVbHce8dbR057vvmS7UU/p7O7VJAWxurTCn/izIpYuMxPKO17EeyGEMGs2uIyU4
I8c9dgRFif07PFKhXOUoO+yGJxHGKZ3NXmzuL3Kq25ynxZc4Gv8KQ+uVY8Y/JQ3iKNNDHB07afk+
G25BFNxR7cTn+TTNq2sgxBDRP850UHrb+DS5gACTiI9wXFelTBNSvUaBx81kCwNK37lETM3LKn/Z
wcq6gi15QYnJEqCywLn6TKhoL542dlb+mW0JxPFMPZrh2kQk0/uXgWjeDcPfEY6YcOam6qhJlGwQ
5l4Z2j/BVK159MYw9jcrFGrHvmRZZevermayBUBUrECasq2gb/3UaJVuwLgjoBKRy8bKXjq1fNlr
yfzLTDfL3tY1n1j/JngWQk8A/JDYS5n74HkKJof9kEBR2QlpE843w/nSs1Km+4lBgZ8P4Un9xNnW
MRnkVZVgjOUz/LK3SgnZRV98CfkFDRS4UClg49uEdUpf6dLiDfLlenglpYlNU/1+JlxWt8fJWepW
zQMv8USCYsgg4AItzJ+E7vE9bdjIgb5amdeoz1RBiR6JXgE/I7OpRk9X+aHQiHrLyBt1d8juHj+r
zFEkch2oPOXQHC68huCJy4y7gdl/TouWLEvv0AhiYkYdWnH/f1rAsMUrNOFPbK71OwKcq4zxyHOw
VuTVg+zbC9Uvw8Dh/aul3OO7TtJJVSIGOfTy4jD3a6qe4dNDebrNbBZ7JnnYarSer3OeKK8k9DzW
cHILV/hOKPxmej76br3ab5X3r5C+cmgV2aogaEkDTwdi+wokhDVFj5USns2XFZd7xs9bWXosgOGj
YspIecq4CDQwY5HSOl32SxC3fbExVLGAVC5H9psbaRMUe1WTusD2W6btKeO/o2LtaM4OGQLtT6Dk
C+pAlDof/mZ/Vfy3kCWDIyNtqbQ3QJ6pnhwZQLsqU8XmjfnDif3XuDifxq+H44PFatClKPCNkADa
IhuSvxBuLt2nC32Q2K9DgzANxQ3QhAIxp/Zw/RuZ/a1XRR46Wlk8AGeOlpDF/rtmG52ha++MDdOY
x1dXmL9xMpyGkpq+6sMY8jQpzIdp2jvOrz0ckqdgo458Qs3Dy8rviXUdwc3D2XdSdWnLVo47pjoA
ha5CWGSfLheM7Mq+NmxsLKryfFQWGAivuSKNGlc9XBN78VZPF/czcAOap+s12rD7yc2hO2eIwPys
LZ4S8jebx9uPhnVSQzHwTpqPmFdwelnikktBm2Cz34+IymAct3D2DxoO9TS4FeexZ+SK8HjpB0U5
ohuw0SUsht4hHDN6PlwZ0AhpZAil8LoOnRGvz5N1Hebf8cGsI0eu7CTU3fKZ7315nAq6SMOe88DD
Nats7JhED/tlWv9jVhecKhUxZqd+YkRMmcC5L5Bte9zLr5s1xcpHf9sMspoyjHa/Z0QUUAd0dQEK
CWXhZzHlsMo2GbGQa5+ANSk0SBMbdvKdJF/chqZ81MdcquLXJz2h6olaBcOgOIuyOywjo6YoihGP
UY7BTTxnvA3qxIC8GttBAt0r9ZGLUlGgxqMv1c7jkt2WuyLzg4mAaUncuKZLP6XYUKr5bdhmWVaN
rXy9JnxdF7DOn1aBfIYzFf6axJIzzQsZk7gZtWX1SdaqQ0mN6m1seAtlW/MqJyOojGphbbNcz0CD
hKdDrKNFoSg/BkvX/AM6mIe+qO6vwBJSDAmbdUEZkgESgtYG6RaQu751pAtkb4Hoqz4YfDVZ///b
lDp71IuLlWW6HldblwMkiBgjjUMoNav7vH2kn3+6ycRy5EgQ7+ceTeAYCzcfD2p/4ltvZR1vAxTa
bJL9ahFOpXExgID9fXeF61hu40VC/HMp8HJ+FvDBaKpktNlPNLT1ilhUE2b1X0d3CMiE/yf63BkW
x9/t4/zmGTx7jB5aJNfdT8/yeXLQJ6DltGhpWfGU37ZoLcmV15NSO4hgTLEGHzSyryotELxjx+/3
+cHsVgjnRGSbhXnJ+l2EgOoIuvcOXiRleMNu6h5Ytu3OKGPel2PgCtQmuG2Ed0uvls6M1/jHj4wn
b3rnRgKkKU0FZYYP6VAQGyCX6sH3At6y/CVRWqA7/dXtXt7RUoHl8LfZh/z58LUN3s/jHutetnCI
IC/8h2OOxqGRc99PZ4EAl6iQVjvsDUCv0E7amKq7wNAmiXKIu1p7aA36yjc8AEQcnajcv2kewD17
h4/YVKKtYcfruQgOGATpChkT/Si6kIZSM5pWgKAS9LBlWQH8W7Om6m5hI8lz4DdRB2UnmL26mY8R
bzyfqN8uUpIwkag9ZIwkQNpBGPu9hXR64Ck2qqWwVJl84vuWdLRoaZ8+QC6RXU77o0/5snCNg6xn
lQ2tlRao0j9/GlNLScBqc4WgHGo7J5QtydfNkdB1wsogpK1LpFlljpNtzhIKMSh36tzqUUB0t3Kx
St47pBkizGaFT6Va9djIIJKlVjWmvx8oEdSE7uvE6m2BjGyqPN3ZxmfGwVhgn1Dkw9HEewKExRyQ
ldVUXc7vdEMSY74RRETf/Dc4PN5Rb3AvYNVsfCV6IJAz9Mfc6Pq4+N3eICr75xIb8rcflR/f4PCP
PKQPfLDkWTWuPRqhBP7XjC6oEsXkvhnVx0zypcOlvnGJxo3vMDkY+MEkCHHFclXifEqq+MmiLKXC
m1scrd4ODZ4DKFP2rk1rDzm5qRjwEQEvYOp2GLZk/7h1/vx37ZVo6POeVQPNGOGRS4H4+rEfvdfk
GQjlN4LjU/KVoaVW4j62hyrHrnN5xTRSGAoD8SI+k1GLdQLrMUZWrdQFVbh5yv7fgXKGvdUYF0fK
MLZIqHFwP9Vi88yeouzQ/D+iRpOtGGux60PtuPpd3Bov90IEd73Vdj4YnP5AlqmjhuvSFux61ZPE
J53tEZ3PO+K0qFOIGzG0gJz9iZ68uqc3wuvYMd+xepWyvabZm83CBSD/0J4iXb+4h7jcNHT/5xJx
/ZfZF6u8XBZ34nois3xAmBfHvVW8Gjkj9GXMRWDheOprG1zVGCvlLvKZZE4e38aL4kwlxi9raHZt
HvH4akdt706+dIzTkgkVWq/2PH0xrb7f213khSJtkPDIXE7dGA9yGWx3lJ2rqs73MmTRelWYOEcN
dAapQUBetDL3u+hmOQNaT/oNOXqfJuHj5Vzrw9c/Pq6IwuIShBafcR7qBhoFfKFFZQcKXTDFU7eD
fklIikl05lO7kSCIjPstYDYjHtPzn++hR4bUyft+E/Z4xdwZNCoW7LrenEFry8OKHMPwgZEReCjc
C3VFxeS6h3TpbeL7XC4ElqE2YbKKqhTvxyTyEIJd6cZzdq4mlIYtNL7nMDY4KDtrpTCMlU6/lqQW
7uCAN8Wg0tg3+OkMIIB8kgmPlMV8ybwSdhjGYDV9Lo6TPRD7KK9vgyAgphAUy9JPD77hMbI/PGVP
H7NTTCJ2j2BUtQsJTvTeGVp+asRBaQeELtxKvwaflBkeNTAE/Nx+BY1BZFugcVszbsPL7RwPzMa/
nvuzdaYNnjAeNiZcSB9uxM6O/KxFWGbrTud5uJ5HQfIT2kEnc7glmgTqUDwFpAcIehaMa6iSTte+
EnmS4qIQzka0YN0x9YH2uJLWJSym30m2Z2wBv5jjuaItuPlS/o1KH0aBzEnVw1ByuukdjTwMWNPD
ZA2Cr9UJt9q88oT/j10o8A47o4azIJ4j+7IjTIBlaXK536lreJPu+AhpP1qvyvYnUy3LLCiECmBB
k+g4cT9X1/ImT9pnsQ8sJe3yEIu3OBMOD72p2QDWwa6eG540+IXVqtU7FOcSR6uzg6ZcOTTNz6OK
e1uqa0AGERqpiwwf79+ssHMe+wo9KYIFZ2cRfiI9ebjcMznWX9Xp9mN/k8kxzcxZDDNNNdJ5hk8w
ahpIHPuccyHhu3urtpHaRWeXCDhyziCuld8Gymc9rqSNLE9Mwil6Tsd9QH7XP5k/tNwgi+5GeFJG
g4zy0VzH3zdq7b1LT4rLeRFbeZgkX4rK99TZg3TG/c90L8B77rmpZuBuilUWf4Pp9VgHieGuzy/Z
UMteSadydj+e+BWmjJsYpEH5frYYtY75e2whxkU77mSlKhFBUQvVKVMRW//DKWKzP061xu5CJVlG
fnAcmmAlFno99FsO3VEgQndJTbQNF6QjJfJ+cMt2PybeXnCDnyhsxKPrbBa1ZwOqyhuotyJhazf0
cSEgo6cHPp/dwn57gnweNTiuarG0CxmKqUAbfTxjL/y/wNNqQHZKpeu9FzbG6Dg/JyWwEue/r2KA
XCIiqDXreS0efMQ1jazD97kc0YUdf9h1Rrp/fe+cG8lX05awD6kEkV3GSvsWfv/6ssb2ButLrk7w
fKzfOPprUTd1PM/MRPwovl/hFn9F3bDEmhNmsbFDkorEPCQJmsGEDhXUTPFD5CqxM+W/UzIeBPRU
L2d8zPhtXFir9aCQPwzL7EDJC4KUBh+tlMOzmmeH5cDz2/f2Trb8FAGEYZK2EkVVpz0heWO7iuQd
4RW57vi8tiveMRk4Wd1BgL/30RJwET71Z8i9J/2Y1oH/+bvBkwYjEOtijBvr8xriy5ReN1hDF90z
tSZgZK/M+UUb0Pgku9/YzUb/snktFmp9EH/X7Wle6E8oSe/mhgfEjJzJvmCuPVZhtk2YYI0Uqs/s
2/yaQt08WEKBCC07y3EsT3anJEPWzpD79y+TQZBwot4H2BXJ7Ziu1KSrh8fcAdtTUzijs5T05K3X
I5PdSfjOqu7eNJLFeTL7c3HTcQL1z0XU430yyXzc7I1kMaBPsK/0mTXsp3ffQSX9/2CEk4HHACa4
jpSKZI4kADjzHdCBSQomXrau/gLlHJ2khIWCWoHx+FSP2Y7HQGSbwqsT6X0lFpp7vNmY84gi0ait
DvK/Yey/z5ransX9/buwoO63GxLMUya1yvkP4kvct3cDduha0J5+DGuiFBmt3OeezBZ3SiKenhqC
OcCuz/qR7SvXcb9XJJZcf3mtd2OJfnbb14qrbxPZFqF33vbyr1pHLuNFISSQARJMJLc3bmMFNskt
EFL+VRFBL51vn77uKd1++7p9J8kGCmeuhEPdmAZlaIYtRT/Zq973LmJV26hF9TDGk2mngM5veHaQ
4C/b5pdt8hjzWRbaAnEz1Q3o9GDsG8nbVpAD6C0s5BMoPA7/M8SNaH+7mi/L0N0pRH8v/G+b+ssp
X1ATY/BVPv88DNDeo/moatpJ/+w6wA+93mPyKRwqaQJg1TvMkcy9I/ZEhKKLIJxs37VnhwtdhdYJ
q6+n8TfcmKbCk+o55W20DK3bG18kU1NrPEM2XpvjzRq5CG7Oxb0/hSROQO28nY/IvzTYH25EtEKD
TfxjiPaQfDS3Rp+6vljt9Ww64N2ZE9Txq+m8J3OWguHJ7r1040eSQKZpfelzWZLoKLFAqwfJcXRa
LraeZV/Xew0GYt47RYjro71q3yF3Gp0dgkIx5VVwqzmHboBZXO4KR/MdaoeEFhkgy8rNIjyercbc
yorvtZsqeVagBSaZIOwRSZ1BL3HdkJwzZwvGhc598V9F7ZJjGAEKVBJGA/OiscnZDBVIE373ocLG
p5xoWdfQ2dFO54QuY4z7J686XC12z7+Rc09xEKyqQKPDXkYz/RHFM73p972bJXBs1p4awuzVu1px
hdCR1q75ZK1ZXmIggsuxfLAuAFe0iN7XAAvbYG+Q6brJeqGAq5Ns7kl4ytPqJob/TZJu6IceCbLU
iYu02UOrNQeJTJHIMTDpDEzIDw/ggcb9mcVJ85nM32fCP2Z/orUEa3FV6BZJ0Hn5mv9KGMNRaGD7
UZ1JubeujhD5BeiE6ZVU5i99ymN4sOo4DdgvCUgvYh+X/MLZR3xjeP8DPG+QciHzl927IDT4syQm
KhMfU550l7SzGP68CZG/Tl1rcFLP27D+p8QQzd4iKj0e8xltYSMdnS9XEgxCVzPvpVcnfXWUoSLE
3WkqDcIQOc9wTHGZtmGRdwZKf0/LnNfHHPcKhOqGqWPi5dlcW43rzAn3Ar2Ho5W3QbAKZNaswhW7
qXUNApWMmorNmokWBcQ9UwDxvn+ne47i79yyD+V02TMrWO0xz7wMAimc8mX2SSO8b/8PmHJfamHV
iSSyHT2Fo6FlSPG0mMzOwmhc78dNTOlat0+1ewPpTbB71mNJB3bNkyNu/2NqJJMM3JNc/CRI4l+w
QU4TKtDZNSWqpf6yn/WPCrlOb/CVCiIsktRH3x5i0qs/MDD2+lv1CpxC7vJlBsKMnBh7tChEuuB7
n2ZwQ7nhvaklEq7Vb8YF82R8LxzNznhI9acECq0xERoZrICS4I3cJdUbAUZeP6oIOhBLVLcJg4Ew
mCd5V1nqFVnj/wsT8osra0RNGpMVBX6LpfFA1ynx/+73MpEVy9Zazd5VL7ob+z65ah1wurGvEL9Q
YCRIFmCt4m0D46NctVB5BmcdUNUv/daeiwPwipF1qI2Wc8HcUALcEtakNA3xZitOM1miAo2Qd5jV
W0A/IPzBgkECZhu5GIINsZ5R1tFc2nRkOZQxna/MvyB3ePXPqPSJKIALrqVMwRyJLPjjk1spH5lc
eEx2CxT11YOHlC2ktDTgvtrntkgNl7gFPv9Jo4YsHF4nTWaOLu1Uc+5iGRIOrWVFuqNjMOe3AJxL
bbuxTk/+riRWPhce2c01dsTXqggAMmZZ8B0xBhMH7IVh3HQ4ePC8K/VKmVEQyG/Rnnx3CfOeFSBl
9jeC08cKn2tzZFpWWHa/2nNEBFCh4HZtKBxHHYpWZ2aaY33Jna8ihRQJZc1f5mdT2bYDg88QsfEw
YDZjBbO5oEaKHBlooRDTd2yTqVLlD45b3OzaFdZ96psMmJLUTAzlXrYMcMbJ4drhjHcDLp/SV8Zv
pEGLjFUiHQWzl+sLlljj2MNHum5SQshDP/c2Ot1l5UdId4HjBGFYNCiCDh6bmLfGKswcErzrqQ5F
2BX3xRUv5c1N2s2+4wnt1UcSMDE+pzoLjuorB2RAnjUICcDygKBAittv8bY/TeuO/4028OfBgQMd
vXMStwEIx5nC2puBPqdXH8qjfB1Y28b6K8GxB9/1rBJ4Ih0FNWhfr3st/g63ec2bTArosLTxv/Uy
sDEApRTpGMlAZWbtuvHHVjINmhH3G0o250eHC5DH4QrTaSJyM/3BGnsUChpn8031O7UxMvgp/IQ7
tABTFkXwyTqJddQZYvTkCfoBJgEJtb6D85GHe2Gzo02/rqPPdkr6O0PliqyWNWguFqnNg4RPYbCS
ekMBF9AoI2htQndrObkLwKh2kHAyX/72ZX8OV5a+GCKdQJSag+GqlEiMXBklqYTyEKwInWmG4F8T
yPp5UNW5aaXwoaI4LKgjdZMKtcFIYnmPYk+HP2If/SFJ6Amqp6c0pbSA4NORJhB+cd05u+7/D+Aw
bKTnKqycSv4OXqLH5K7M7PXeZTzYKc6MHQv7fKWtyFP6akYbg7p2BNvgx6FRL333sxWqEkYW/OFN
804wQQuDDal1WMN5OYl+UCEmiRAK3KAqfWFFlkJG7hXJPTUkcDTjthf0vIuAzByli2w/0RhRi343
pPpVWAJsK3hnuKg99KuPBW53LBP4YDHYUoJlp9fBXJ4tvbS6TgU4tOGs2u2uCpFKa06R08XsC/gl
f5Ivad3BRYTuTOeI8/ZKQKj49/k9ggsuCv2UnRRgi+NavSSvodDKS+BGykdaYBFpUtDKdZYwb74b
D3Uze9MsYAs19ipjR70kohzLtzfnx3sdUL7LYIRHjGXYdJunDf6pEsP0Jrg7RlL/D7CDGRgYm1xf
YUC5b9a7bhEiytyzHBTaJ4zUc6uI3bfnG1bU2rpeZHO+bTyKWSRkPjp/IcT8alyrYo41PFAfZ1l4
5PpvjpUHl8XUCSdEdrSroojJ6q8l7M2n9YVvlbtB52088++W1tGQrb8toqS4TKT+rsp/MA/AM5Fp
PA252kFjpU+HOfUit3xtIT67+2Ec0UFpzj3gXmITXh0aqLUz/KsVkNVLTA93Wd4Z4JyYqcPpUAEA
Zx1e7Orp3wUzmaTXCXKC5D0Nx/fVP0quhXyO05r9AsfaPPWB7K8oVtUc2U916H/FSc3MIi7dvCrk
aIKAS6s4UOLTrsyp32AWGajxnJYyxcQikMZvaEr9y7rqpQIAoFyl8eXXBSCCI37Tob2jNaSC55sw
vjODwezwIxylDu8S/0Lojl22cD5TQFFnHWfFyBNhqc0q+sLx/d0IncIYW63D8AYWv+ETtepqDwHu
H+8M3KL8caxATHL7+w3EPldOMejKz8TlF2YDai7h6/k0s1QJZHDB/N988Bu3Ki4ZVD+GPqoZ6RP3
tyFWDFirQpx7IFXHwmNtbkIP7Cdyfi6qYmtbEakW3XJKi2Um6Oo2hhEe7jlSrzhOQLHhquZphFr7
/jC0Oln8swlgV9NjZaL+OrrHXXCtvScd/JiF5c/ErE08YryeCZzRsC58Q5O33Hg7dIsAjGBIgmPC
LRS9Es5GEpB7s2gb3vn2v/GmCffhUw8W2paTeEQtC7OowcVdJyFWoZREgu7zi6Rz9DbKfVny/Lfq
Nn+Q8PoZPoJ1evClUoRsgKRJIhLDvghZOZvIKh+GtrLYqQFTD3AtIg6hFkbiNIRu9quqhEMKt5jP
SfHSVSBwdRWQFTcWKOmVKFSGc2XTFbRxERPn3Ia/NVOy9jw85FKssf2JKDVyewoN9r4m4wcux/pG
Tc/JrFqofHAaeCKULOQm4mtwuZSLNqN4ckXxBY95+D9w9Ofb7023831kernX57IjHv9Ll25KIRy8
dBRapwPSOhR+rqn1evDCmjCZGqtlrH37Moc3B9+Cgi8iu2GOpskzGXYXqd2jq6njxyZGB9qxtrHi
+Ix+CLCP6JCTnyF5w/r4Kye0AlaOU+SMV2aH9uoIbBTdOUWmkqiu/fn++1uNnLr7euxs5SGAOGUg
KpDI3KSH5fRY+SDnUXWF46XUi1YF3R1/QVRY0vSTiTLxBsw7uVSp5IIPd44ZfnHVqGUKrLh5fGpM
J3u9h4TYMy4sNbCT1ShhxMi5Kc+wi7xLfBCBS49hVEEOxFM1kTE75AYAyO8ryhWzGaQH4iF1x4pD
06YsLpWQgsjcp8evC/9cC6St+h+lWvNJAcAeRejJ/uWiG+nFgmsBbDmz0MpS1lxQHsDbIOB1QF7+
IMEdBX6h03qU7cXlCqAVpwUKgRsMsv4fyqIk3vZ3yP+sor7gYIIE+O2Kg2cVbTKWmp4lMoHXPgBe
QKCSkqs8c8ImmE9NcGRl99jl2ZRtpjiyO/KFUFxyKcMMQPsoAPsdgLsOlFWDw2/xDwkmx0ZLq7M1
qML1zWvkS3bDR0RfWOCf2SN3BedoIulLvSiECoJyoayTrJyytcEWSeVUWJ1bySzV9+AeQlL9igam
+bxhMrF34kqdgfMjuAaGn3d2PLEUdSkwCRLS6C2NpUGoOAGFeWgfp8R7TNKXPllcaoTyTwibhEjZ
sgKY8R2L1RzfM2RG0Pv4eN4VyTpno8Nd9PXQeLjoO9Dpm5sPuFGctuag/VAZbK7otlhjlea2afZu
4grfWZxexKCdmIAc7hq3qTMakd0n2nx5ev6ylyjS+DZTAOsPiqdaIJHn65FOcFBhJJOtkhNbGcoU
j7d8UTwkPlzVzNdy2APczHWt+up3oTcJpsBuD64CYMf1KYXzEffsvgtzpo9rrqEJOSWza/WZYL00
GTCR01DAtepK8au7UHlRJE9HkrQcRFA9QL6qRCVfXYK1JVktJLErmb//OLeGpR7Oqe8Vp2ZvuTBX
LT/mGdlthq6GLe50ctPMAPWVUM9xiJZ69eAov2Hh7AhuXlXQWmo6ASpJ0OGMpYRwh5T+YPv71Pqy
+B1nCOSEPaPjAjQIoxj9BDzbkgg7q+C5Q0v46nN1q7P66Xt9M2MwWBKuQWJ5Oqv0b0FEMuu+Uxmo
M98cWCKFUnXQ9Sjm42njmryJompUCBnVWsPreCj8Ki517NdAT4fbdtSK6Nuj9DV1H/R/3qC9kj6P
bXwB/V1LUfKtzfZJkBBkIiu8xfDjYWX9eqWeem4zt4hD1ZCC8sSGfdUr7v8TL4tcnc+4e/5o7ZNT
WFAe2FqA6aB28nYK7shsS7KBSvnvYn7o+KxoZCH8ZjUEU0apUj1yZ6xHu3f7ER5TThzclFO1M62O
6RwTsVyAmHgU6iX0NaJZSJdDunxF1CTUNaeNmq2T361eKup91Gc3K9WrotkaFnqn8W0Ac42+fB6G
SMMLthyAP0xatckmdOWcGJbQCpSs87SEpMt740p8GB6tJyBCrNMHNmuDJrFSGJ09sHaOGc43Gmbf
iSmdy6ztxcOQ+oeGZebJ2GjkMPdRGWIXL9EQctgs15dnM+yIatHYJgAalCJSlEO1MLws2SsLinpZ
v8pJf6i7MXxxYwiD2ATeoc6Ms5bbYDWcWCOjOO+ZA6G7XUYrcLb+uQvqk00eIN08f3nTJOOXzdpV
d1SMTEcP5rqz5pRvSIeDUIV8FuVFOV7ufel1NAt2nTPXlBY74JR/xb4/gGuRaOTfpiu3YzwyCQuq
WGOTJP3WIwImao/q0zm+gaumsjnfZMH1E76hXf+AmHnGmwlDGTbwmwk6ecbTKYRE0Dco1LGoWaer
FRQg0RTjdBeo03L0W05xzUrddG0qtz3GOuwYnsDU8lX52L0mWI18EXRsZ5873xPpb7ctpLxEUpx0
ePvHOJQgxjr4tVt1ykLMt3z7kTqtUUgKU8OLlLFcu0IW2mghNQyBP72q6S1L23Wqvvh3pu98nylY
Maq5keZTXZn0SnEjNpSpJKss2YYP3BOaoD92blcYZJy8oANLoAv81Jym+ymoYAd0UwMLJdxAlRh8
66VDyvmCue0cj/iP45SIvSs4v0QMcQEEtWjgcJr/lnv0KefnY6G3F3vXpzOapOZ/gUpHhQKCX4TR
zsKTgbJLm3NzpSKjuRUFQN72EuGOGMX6a09TJ58KvSa3qLjArU0PviArzIPeb91/NC8l7k/+KSF4
LfRkEznHj8mbM/hjcuFvl88CZ8kAAGjNooZTcs/De9VKLyo79uk8sD6JuLzs9ijKqC5DQISt12jA
019Lrnol9vgXNvxfc1QOPVyzUISJ/ww/ZuTVu3Hqq4M6yzb0R/gT8lQSsTAxib3tj+l/hU57duZB
ubQjZvpCPEWpCBhdLk5kPo1s+iy36Nia6GHukqEZiJaMetdlvCm9mzxtuNoJ732PcUfVVX1l3uUp
EFq4tCDQKFx1Onse+0xkO6LjQT2idXW/HedUeEskgAeNF0Y61UCHFTcXlc1Wo75+Wkv9Dn8NJ/MV
OcDyr7KSEeWoQluBFn+VvhVNt7/XaM5XKYklneBD2KU061WyXJiHiKc4Xp9YrWKNEOT0FEU453h2
dh2KVNCLusqzXiv4u4sc7j1Fmyqj8iE4RsFriO8ZvMrV2Kqw7VQDuhxvqNySn3Y3GPnx0cbA5ZCs
9cGrONS/P/7+lJSzRPLFV9AYftBZW/0euY1ZzJYPyx5C1yFcIDqaao++U0nl4WEg3W2jHOqvB4W1
BbRbYxWwApY4dbPMxf7rbc/O0nhrDcWM+N9maP/l/jV7wgFAoiKTq7zJEJb5DoiHZ2v8uuPY75QB
BPX0PTJMbeDrBRrsdL3iQzs0q64VD6OrDPDYg4RxdX+FUc9VbVzMtcLQvXr7p0OfM4Gfj5tYwH3X
cPATBof7W51f5PGLC/YLt5vs0isaKrthI4MnWKv1bYVmM6lV7PBfLGBBJ7EN1eYtcM8aLUsFVewH
6koPElffnybQRQ7wEvJr+fH+2p5UUVMEUiZgqKnTPZPp+nBxtaT/dYpdySCL7RI+zmTbaQdOPNYk
8glfM+9YhbHklxJs2iPvoGk3a3EXxuJ3kaRApvJof4lXl/hEm656Md6zOkdnh9JRj1PtJhcLzDXR
xFOFgNshIiqKOTIOhyRKgsx5dMEwyvwHa0obuSIUZ9E86AXwLelWAN6lKrw9QME7O6iRQ8ycaTL5
QSlsFHMdSpds45AaNRkfQ9QVwTkVVDO6LO3+yTWBuAWtb8bvQYVjbHyZG0ik5w7sPFZeImI+Ggqz
VJ4i2ww8Wa1DdS/yHRj/j/7Z8uTRGVXkhRDLbjwCEjpBxVTaOr8pVuvfeJprJmgapdcn0PpJ8eA7
rgkSLXFka0MGveBoIi1iR604zJ5IIZYnMTcH1Ni/Ptg8/dxd2lLKHBWlC+rKCB4Vw54j0G+9mwqb
fcBhmPHuDvMDpCT/KCi0cD8NPTrMnxT2MLpyEptwuBCa3WZh96Ri8NPGM6UP57LZ9YmV6Hfuvvaa
M6i+JpA1ypdxqSObYcydCU6jmU18BOaQ54/rCI7nxZKPNkM7CpZAyrcGL7X1bo8mCzYngE3Lzzwt
Vzx6bWsf8RvOgdGmmE+clt5ASTRwOOZDPZ1EO1ofqyfKkNC17OJKc627Bcb4d1zxIAmionpX5Zkq
rDf+2Fk0AZEWqVedUmAzOSvN51DLZrFD6IhY3KMXgSROrO+slowF9UsyD8mO9qospdzvl9c47YHh
Qhtkl2NcXZE1MPcDoZm8FelGxvWNGMAOaVtOw55XhA/P7EbIrIzMOFzU+FgYFOf9qz6IGyLVWp2N
us5O4KYy+0bV33jZYv+yNa6vJN1HTkvhxeVjwJ3XVHq5iYcDkkLCAnTjqqlphiseYO7v5TqP83PS
PBBxbJ6/aklf7xXWV7nmltB+0c8QtRKev+xRRKj5bu9svgYi9l5NlVjzrlWurstFWKvbVMl+4pQO
/Fp3SGlNkW40XVwYjj4vO3uAF6F6yTHQOa79Rj85FDYdZS5B+ofsRcx3ayor9IAqD0HTQsVbCXtG
K/4mUIlznhXkr/9+3Fa6p1ggEN6lCcbzt+5vtOPx+tEZed4OyQp9+tWvRJLHzQ/TN7P2xfdrLfIs
rMzCzGerbHNhOwNsQfgyyWKx5ge8S7teZ8Mp7UniKSuUK8rZ6uUxfVwSK08cs1xTKUX8q0s+1hAi
rKuHU42tx71f7ZbSsNeLOJ8vil1cUC7JmRsvVqG9RlAImdYph/pqaXYE1oFqJaq7IGi1NjhTTSCF
kd8dgm26QxfVcGt3VdlEOTgipa3Q31KvGVVY7SYakAtgHijix8qjKsYjquk4q/B8Ox7qlywBuIVp
Jg5XEns8f8WdALMAkBX6mqZPlWHtdxcvkS5y7kBOfC+umlbihDtO47gluinYpQV+DNuBHL8RcgTU
bRMC+CWv9xaLitYNZhdpEm2ux2OtKzM0ag5jZGCzgPXuI9X6DahLDse9QzfieMsLsk/6yINZ5Jcy
xKzNTJ2rcsze2iAktGthO3cN60GmVL9FsIYL5RgjXfujJrd3htZg79bbhQLgitiPuKXjRl+uzXnb
beDrLizwFt40pbuwU/7UhR9t3u+Z174M/f3RWBaFSfknrze7k94igY3zgsD8fZlzwNmeMru522SM
/7mvkSg9+XAd4TfSqAfgZ2Cp1OR8uT+guPuSyp4pzMkG7P53ibHheeUI3jri23mJagQBB7VObuRS
18nahv3hN7mRirv8Yza8/5dakZ6DCFd7Da9ocBqjcXewCQVsJupp04Fxyotrg03z+yzL9FhDn621
770EN4X84KDBdRt6Fr8Z08x8MbVNU3+/fPUjVThSZ2Godc8+1fGC74pQEFo+qQfS+W62coZFnC74
nfkdXEYN4ubj/IjHkiNStzjz1pbeKA9oAbhQjGEc67RKGzn40qcqnanlSRowfSlQx//WVp0ck8e2
X4gye6XXQZW0rYbhQabZ8xt17IvjSrdgHy2vyoIkO/aOMhEhoSIEUUSGju6NyGupelNctW+2twUm
iMo0LjlGVhNMgyS8VukgFwsCrDH2wrpKkQaJWj9UbEGMxg8YQXSHyDB6CJ72bYUq7vNZnlkPqisE
E3iFeb9ay+dW9SHw1mWdED4/G+6XOLDCqnzZQGFeUKHk5tbf8hgvYPP2EdVsYrmOdNQIVriqKAjd
EkQQ5TwYmy5MMS3gWtwjLpl45me4opA5gLfu8xiUtph/WtRAFH/pvZAIKL5zH9urw9KlrgdJ9a51
WMmUly34fmB4dwN+478b4P6UGg+k5cemmgEKEKgCc8ASFUPg1FKN4rswicgmv7yt2naEVDedkbL8
YRBcR5rP9gFUbB82ukeb/q5Aq8YBqAqltGrRf2T6vnoicon2+dt9NUHE6iKl8UK6KB7GFp1vf3mo
9oi8AKKJvFPPbyGbpWR7sAAmdFDSpH9Iu5P6zpxLr+OkRnOWlmEkGrrdU8revAri28EN5B4qzuBm
5B7mnWVxANfieXmH1WB/MPbVK586m+XPnYBRKeKAR3lKMIoqwMNtELSlOwXXO6B+O72uq5G0VeEv
nK5c1/uXL0Z+ntMZmi/PHv5bp1kDLvXDXjhoAHPyMaiu5DrLGJAu2+Be9Wu40fRZfw52GdUcJzy5
W587Pti+9xgkEsRzked+JQEwVfjNZyH2u/qlmfL1rApwoxUgRgYLNtEFzEioFbOKffKpQqTPs3Yh
Mmec+6ToWY1adPeeSlNdfADfMqzdh0SDBLuKgrjXG2iFOUhQXPAIGVFI7h6zkmE5SzfCnA+gqyZG
b1PA7TWUltxe8bKJ8VdjJ1TrLXDI15cTyTL+Ad0vGsRU+zlOYFAXCBVrSrgCSmvkBO5O6hCOVPAm
2bg+f3AO2LcoV6ikndigxnFV3TRf/EhmKX6bmLclN6cT1P5DjGr/uggjdXsqinRSrkfuc8Y9Wh9z
kVQ0bE9BZhWnVfwmG1EGbaKJMgLWh1YmQlesamtmPh2Vj5UJPF17Ce0uPM4K94QP3J3nsYmEEd4E
sSAuR+8OY0zS+m7aYPJm29+g+pN5uYMRJx5f2+ln5ATNFbPtiUZCvovrdu0wQyUlPHYQ65GUdTgI
UVyU+KPwclwvmnwz5YYTg1fJtdMwp0H354lnaNdQBO0Qgo206mCGC52wSVSuVRSI839f4NURltJw
Gai91kDU/z3NuDC2kpeSyVV18ne/vGUZhYbiLG/39z95XPqxN6M1j3hZvTtsjXlFaG8S0JhTolJM
WaU16AEl7INtVZ36uWcAxOtKHbGP8DPWcWDkoDsVJfXEzlGNhhp+gXdCBZURy5OR188xEuAMg2zz
NDg6Ps41e4HnxItMPw8JBtjx2yLXS/XQzBmNyzXHy+XJVYjCkctyMvpiVUkIpyZxmvIWpfKM4JeI
ToTaHIgzrOJCmIhGhqA0AMM5+gggrPG4mlu9xRxzsqpHrI/PxWgrfg5Cl2fBZMsnJi10Q0YUvA18
m1VTWL0PAjCkJFYIHOj8+6aUDMDMvP5FmgnujDwXyz1K2b69BR0rVR/K6pn80N9au81JhzRK6CUN
ERsl7RPUTJom/JhhnAyH+IFbQFiNq0/DeMGI1n3CFs01QORJzPntthpr7+mRBKz0H3pVEOuzyxSn
qr6M07+fQ77dFVXdyTr9gsUkgS//4YTfgAjnKKy3DI7oxUhxNnyOsJXt2Deb/88APG2m/4vSfBAf
oPIS6pPrLbGmtQAkOCo+mj49F1uJ0c8d7PlFv1zJMnNHJqGq6t9Dgcf+ovjgUe02R6/M6CTfZDs/
7IaetAUyqceFBMFxiz3+CjiwYOIpVTnea4mkazeAuqqRi6VNKQJtaua1bAf1jWYu0+EnuCN9Duh4
8rKEcGfI/zY+ZWE3UKZJuW7+ynG6oIq5bmBeP/eL+DtEsFLGgbPBTP8bMFv/uj5G4bxEQSGljvmf
gWizhcgGrqgeGFFcXr4hCBLibxu1EFaMOt1UpedJN/sgPIFcy7Vd3aWgP+sVQ3rwbh6jkVG1G8yw
QzDCuX5zmoFb+QS1c+Pv7E2av37V3+kCOpjiOQ8Fp0q9o9VOFCXP9m3qhMl1NY+Apmf4uSXjLmSW
KB47lhpIpRNVbfg8x9k0oG4rcskDHhWXUtU5hhXVcVWNG9cY0FpjM6dqAlCp3Gdz6BpaE5DiXDxY
S3UalOhVG6KdU2dW6VVfsP93GPWioPv6ztk0QXK3w/MvlxMnnluiB+rl0pXwKniEozjqnJZb2Ifr
gxWCN1TFFWjEItF4qZQttWsSzfavjp6frsTEU99gOpHeaKBJlsVX2DYQFLbUkPDlror+fJr8pKm9
Aap7D5dcZN3SypjGKgDe5vst9ZdS8TF5hEhmqSt6UHEHWTAmgsW6mwvbRvgRSauyR3LwoJR7b/Oo
1sxAYiBjOt11gWY367aaGB794uP3a1Ng7sAiPgOjdZpPU6i+sw1dXzgEcUFLicTGxtv9Pqm8iKor
7fxQmEWqgBe3rcs//VMb7qtHrkKWwg6svF4FZ2MRykvwT+6DWYKQIFkVkf3cWyeuj3DkRc6WLcdm
WmHk3oJMm8sm9p9zCGk8gilG7SBA9r3g2GGZNqP04NcSZ63yRQymsmcC98uDMQQtpeOLHYzW/lcO
KxWXKjxCFPDmTrPvB9gcsZbhE6eWe+6EfqTmpptFNtecRwDwC2wI5Lb8f+L0h5mPxNedUWV5hR9g
S/5+6MawnPDEOns+m+1s+PRmNwz6NHC3qa95tV+Q5jujj56uWeEe9HtOmziaKSQXspRGaerahlVr
EB+9XrFVhSn3gynTeeEQZusVGkL+fgzE8nEfU79qXkxCFX0W1CYM+rxPepdN3R4fZ2luh0sJ4Qyy
fLOu+O+n2b7dL76W1zv6zX6CfxUrpyT5nBCWpEjZnPDnPHtO/Craxk829wv8X/S9QZYaG1P6Wj81
QDgwAb6NDC4NwBNJKFuexHFC4PvhYAsrIvduB7Y/muJbSnKW8V4W1abtCljMyJoa2FI6zIqbY7eS
DufuAO44OAvjMcXJ+T1L2TEb530IozahQRr7xRT5oi3X2CpZsQbTsk8f4a9uI5sipMZ/XbeWXhBL
Iqg/Kobs0PmxtXQdIpDPeWFBslAfN7gcYG1dJuN6Bgam/T8zsdI7rIAKO0FdIwNUV/1H7QXhXDUT
+xcxwc9kIYJDEDNnIy9yCBT/w9TiVvPFWsY2ZYLSWjH8deM36+FT5wyeoL8ZaFQPxauFLjgIbYkF
SasMtS1UyUWrPVT9fzlKXoWuguD0DBBrTXYIMh0Synl8vEgpjz9vfQi4tRZrnPjjNqkvgKkVMsmE
V950JWsph+F4lxsric7uAaS/cF1g4kJt5sVoUmy27cuU7vagNDRturOkiAzVL/NM0dLxKy1xUMrT
qLhp4MQ+Fw0wU2/Jq7o8kp7iFHYp+iB3iFNbAEclP1570yaD6ZfNNvrxEQKb2ZKWpCvYPsVHMVYm
n+I1z2r6xC/N34jiM2MayeLFh4r3iGRkTmh3fOUTgLlcbGQY5umtCpJtUywBsuBkryQQmlWduBCm
mh6wzUg+soS5gBqkcBRqrHKogeC9ovaAoCuGRQlnQpxBlxY4uFPL7nyYxh48WcDR8N9EDoyC5C1I
zZXYYJGoR/Z2VaMD0UaaRJ9M9xdLdsj/wBbbRiu2yLa8zLWMv3mujoMp0+pt9Mcso8H3Z7CEv3Hl
n2GFxYvfqhKyEbcnGp4j8UQC0pmruNk87Zh/LNKt6JP5qxdw57nvoNuKd354ReKpnH9Z6Z+j2gOI
m0ml7u9gVnCh82oBqTqh/8A6otHIA+n/51EIgKtjxObBN+PqIIocwmGUst+gfNSixQBsiwWu9IbA
4EFXTBxU/Fvh+9FbZE12uvPD1xHiig/R5ShXORdXoQc6clh1lbo7nY+1fkO2lt9vh9roc2EU2pNF
4p8STs38Kuu0VD5AGGiatxkQduGFXy7C/GL7ZXKw6qFtlycGp6h0tHPrvNFdaIe6kIs69nLitVyc
ahP+S+sSDkMWlE8TihqB7r0mIywcN6rDkOWIdvx5slKFOBnvoDklSF/8/sGJxT6DoT0g4r3djVhY
Uln4oV6wPnkKbzjSg0SciI31pM/gmXhTdv+F69yk44SyZ/uiprsQNCj/GKrtRuSPX0EFgkCV5ale
octOLzeFIDGBN5XD1rHg4To9v+4Pe8BtraA/x+VSn3NRQc7TyDiM3yUogoTWW/TGB3GeF7BIsdQq
a+C8Z1WjbhnEg76LW1rtG7AHc/K9cNEW4Zaxuhc9ketC7qTeAMtpBhLrkX4zUVEbo9RWykxl7zm/
ngTxUrl2aZojLrfkLqoUXRBfnj7zN5bmuDm/SzdewxnXmqmli1BtpXeFhTx/pZ/RhXy9apQQhBRu
pFOboS3FlGN54VEOMZ5YDpIe2AhVnuDia7SjWkXFWYnfl/S+xIxmi/r7JAk+O44lJ/bO3I0ZrEtO
ldYPPRqIjPSgb4gFHOXxCJ99pekpKfPtrjfAijef4rhxOiixvPUiNHHsjgY+WZRFBTNMxWKXixgM
lp5x4ccKdKZFS0+mqOBiq/ewn3h3QEg1AOL6lzZOXzMjauO3BzxCcYZoTY4EYPHPG4MstOqvjxgt
xTxv4uS7d3oPnbigUlxAQ2DimZKb4aWR1hy7wn9Oeme0SFfy6//lOg8V3gAp9Irp8MDROWlW1hal
HMZsMYvFW7q1ZrKgUhrj3MSrqzJPlf/EiTuHnE7IsNK8NgamVQwFGO5g1nyLcpqbnKBLBA6fYkQt
TOdGUDONRAHn1KHMjG5uEQox5mQ9XUQXynq64pwD06uCwud6koEIlLmL61vdG7dOQALDeB6Vz++J
ZDej5VhE1BFi2nSK75EiOjzm1s2KvAev2iCSzHYpgv7evOHzZSk4YOecq4YTMyucZvy3iJVHEbSV
vznNIgrpAWiever8Bqks74mkgR0E9Fm7/r3rzALDEXz2ELu5fe2857Z1qz8qyCHCyDV/jYl/yDSt
ka5MSjBah0yiNvTUva17rTg1cc1eSFHW215ouoGhCQkOBq1ZZrWd2gkY4POxFoeQAtFuYwdaqfTM
lZB2gpZHmrzJ7S2Cznz1rncSmJODESzZhu7SjlUhb2hsSRcRYWkuQ8/8Id9PH41GsW9Fl616MUHW
7XT3aYKw12FVgmPEGBjF8NWOI61qd2bAAhBu/UrAuojyrxZceG5N24REUKhv8637nNwiDqTuiEqL
1ZdTVMtFvFzIdYgto9QjzdXP4FnbphVGWNSq2lezOyiPAJvYTIPih2qW7Aesy3OEOkZ+9r9w5cTp
PQyNTQEX+7hrCUvcDdstte8RKuqTDZxwIngtrGRZOWy/lBZsL3Kqw5IcCJwQbA28pYsuD6XfRTDl
qDrGRN4IGAXk+NmrklaViCpU5cbKXHF65lFuV34WuwgKMsVaNzANQD82oRZ/cdd8KxnX3p6xO7yV
5zieh5QOca/1oVBCrsTijsxiMMjR9w79xvYO+27eTvoSmaSLrNczy0rMjtV67hynmtt59IZ9FPxK
eBl8Uu/L9Y30j8TiB+t3PgNA7hRzaThucr2GXeuU8ZB4UNkgdZsCmQV5oU8Xk1q3sBj82o4ygHUs
6HWbliHDWZLqYQLq/YBl4NwEV7x/5e80wmCMEsFFlg2REWiof+sPBd2sV2Xa1P10m7l52Q31Tv8n
A+tFqYnJ1DeGzyXJuVOtYjojEIPWfWOOVyqENGBRWdoZlib0nVQF5nUlRxmosOtgL06lpDx8ohv7
aW6jZCT4EZ6tcl+o7bBnfgRNctn+qXbYs00otiLbhB80esQrAebqrTwAeNB+YyuZ7WJDpfHEDDwo
XNFYUrw1imQdIOnsJgoDCQJamH1vRkdoBCPOkiTYJcKEozc+r2t46TaQzJXq7MH+cnjY7qP8ips4
QNeweg8iVpvtt9CUipYJXgPAS4VgarK4klrZCGkerpbdRIID4W8CGEeG4LgJNttfa2WZucJHjBqd
l4XuSf8IR6Of/qSYcpO5de8RjAkXYLyU5psx2ihYEzT1OMvhXzJ3L4XiZL9/4AzbUYP89mrug48I
86ZG+9EwcUZBVdtbPhe0UruaQ7qm3dnkQiK2/VsoMlvb+8svrHvtu1NlPhURF5afzMMWIPxrIgNg
N1yv+eHIXsUX3aft06xGeVTZfFBgSRnysr+9W0haur4AImudVGkjjQCnaoSTVFeBc+aOZccTCk0k
1s0Ox+l5koS99I2g3ihcq7QUAFvjn7D4k09j6bV2uaiX7bmBtCuRRmEvHyTP1xPxkqIjP71d7DCP
vlyqcge52bun5GD+Hi9vVDWckLzgLSItcUPnDTCLwV07O31cZZPOyBMgKXKE0jamSj1pl42gcLnj
qCUJKutHckMrny4k06znvxDB1qmmfjmpXeRtl9P1Xxcc8B27sNfZUsBG4iLRi0buc+2FRngvuHFv
5nBEyakbyeLxoyzoxcH5yQiaofWMuivS4hdPCjXUS2hUiEQILDgI+o/VS9SrPYYPJyoKaoWLjm8j
OtKQo0/RRN7z6/p7LwKfPe1gZJd2Mz1xCJGWoYBGHz7Bb33Of8lLml0CdiMU5NCwSbTjauxWcz4s
VBDaWrhksPq2ubPZMw1C5q2VpC22qGQNCIf+jYjsALfylm98xavTxd/Lj5zFAOYOyTa7snJo2M7/
yZMIJJWLvdStQl8DRSGtgOpjaN+TbNfowf2oSx7oWfYxlxG1u+nzTJbxQWAKFksJEXvHqmJ4aXGC
B92cDpV4UFBzcgWwxQsHzE224kCeWsKUhBXEAPEYJPYT7jMp2kMa1rjZ+JWAj66VVJn8q1eQbBvq
AA6I3aKsldYHQM5a1OW9EmAsjyfuVTj4ukzQYajnT5lhdQpsApA73oJ6v/B3EE+zQHTJL8wj8Fxb
DeYw0cJle4002Fmy2wkzu+iKeAv0KpsIkt7RodQr0WisWXohwjm1PUhLfkavbuymNSs0f9os+bb+
KfJm1CjrhJSpwxGxsuXsqZBhnRbSGbrgpzkeQ6dhsppVoRSFv1+mHgv3fzDKxBPzh8a1JJwapmBI
h3vLz3g4KUPfeMmp9Cvk6dHBtaqwFZqB7QUVkcA8Ql1Okv1eJdSTs9rt2jOM19tdKlP++UuBvq1m
MBvhJzQ0Ufb6nkXdaaqFVTm85Z8/fATLEORBscMh0751mrXB+Ade9Y4MCJF50DOFbX5yL3C5QlS9
Bape1dmcBCYvEetUgiT0rCF66mT8puxLDsZy4ZSSafxme6ccD53SpqZm676fNguyB1/MHoi24tFS
jm0q9wYgA3MOn22PnjZkdBj1UTqYQcOxNr4ZKRsTWrcPVISK2RvtD9dR9LiAgKeIuEHHasd27yVd
XFqjaqHp0kkfhnz98eaXjqWXN6RVI4jTgY+Y6llMjulD94pq58t4/zOhkxVlTFxwbeWmZjzVBv8v
gWui70ZQL2qGdUGp2cr6gN7Xz9M2NxyAxHiJPGOVSnWyRm495ipRx6Ci3O1wzEmF13sBxM9mjjsC
Eo4T88rgpc16TutyOCFDfLRIfroXQ+dcYSoek/qu/Xypa3UDEMHOtOa8P3Dd7snVFouXuB/7ZxwG
z8542/r83twqTcbDC6WL9UBFeIylUnMmiaW2ZyLHWz3u42bwLqqV5K6P0Lrz4EehaahVxrwSqksa
SmdI4fqhAOAKbtJd/Mmfs0XcPev/m0iC8NVsZVC+wEhv1XxqMxsxBwwiqpgDL3n5GBoK/duiCRfF
scMRcLo5kRl4TE6kPOOTarUeL1mRzaX55CVs6l1yB2MyAeEETTF7bqTYMjI61Gs7fRJXwSPJCNK+
PRvZDKaNkkDUgUdhap+QXjUmPKGR4joO+kGMqNH4ILE3RNnzp9YjyU8HWdSkKaYKWfLuPjaV+Wn3
R99Q/Y2thFuVvGN84S5DaMe3cW01f4EIf6VZvAC/F77Oe1WKMJu4JxBhz/DeN5X5kqU4z9h16+Dh
FtjneHiTkOCE39DsAITQZnd89ElpoGJYiN0Vwshd8UXZoFuS4rDOcJvER2Sx/SYQoevo12HGqWlD
n7EnCkADp4smB5qbJfznOVp4Li5oFvZCtMUJtM24s8yPv5Hz10s2+kV37WIdfjC+MhyfcsxAQKB5
dNE6lPhrmBuT4ZZA9ald/lK2Yc2Gs8Uzou7g17J1uuMhZOso80SIrDFThcKYHl2fQIYhvcKWE1eG
RNZ508m5cCRdVQ3PCG8ay2CXqm4Zmx4PqxG8thq+92sDbCW4lAcgJUmrehuu+9ia0+18KkjrsglI
PiEsy2v8FBqmIX5sTwvlb4xkAcvr4kSn/mT2Erag5BIsbGq4XQwBm5F7uIg7MHx4GZDEKmPFrRhQ
TaKYEucHM3N6NgwhH1pPtjGfhO+rV6ws43wvM96anTkHVH1Bb2juVrtEAvlWlIp4Dbw+sX2cIidN
yIPT9qWzvYjNaxm5nAfkx5xmd88DGbzU0PLJMw0yE+IWp6bOiGWjieAArPoaROvChgfb7Up4ULOZ
fAX2cMiMXybuBDOqMpH/mfBD1wAUyAlAzj5Y5fZXGs9+ukvYmVkpkSuK8itdP5d+yDORUc5Fz/Xv
tHMynx9brADXyIJtRdSGaeNl4rJlGHFQVojU2w/fg9MJ9I93Mtd/R8mya0FK5KWtoTIV27dNybX6
/+tXKWIZJsuykq97qyITw6oSxVTD9G3LiH5lUDMxavUXy9HZqsLXS0ract8yYW4jw24Q3vWl9xcz
3+Cc1zv2HWGQPYTQ5/bFsDDfLeBYL8tyRAMMNqg+XePAqiSKLVfXu6/ToNgLIYvZcZd09r2kLY5b
fvIniY78eN9CQpXG05wTsB7mgfU6BjVetVk4wCp5BGAM0yDIofNP7roz+1g3KrCN+Zo5qzN9ZVE1
ooeLKDIq8E6p9pexztFpy4hwIIdT2HPrj2zDcz00pwl+EZWFINqDW534+WIzTtOQytzrpZsplSGt
Jbs+MdFDPVvLOPgftzG3/WYbHcVCcREto1jpbuY5/mv8SZnzV5VYvikqqzWG9Xf+Os4hs91TWmmE
tbU59SkF12JX96hzfGgliq+itgfwE1e0VzHBeW7e4pzNP8psRWyzPPsK6JwgB+qEqqxbrYzafBI0
BfyIiSmFXsWtvK8VsVW9jtXThq+M6bt3QWG4rGV3d/Z9Qh3kQfavqiJzGAg7ycpR4nXagaiI/qqC
kDA+pJL1rczUgfGcz98Bch0Gp1or8XXh74yGE+3EuI9LCyBCJ6p4Jq9ZHQ9wIZtQFwwJPmOjaHzH
8fMApjq8YTm6paPfauGppk/6hNJ7D4INCV4zIxUbJ6lwELC1bxgjKMHEU3zstoRh9nftpCV9xWbo
QAUCWd0w8ADzGC4KZaPJLAQAsx4BnaWTJNxaKKm08doaT6PecBUWl1OsxhsKttdl3kO/TtcpahZX
rjADREaUFPasr5loyJ5fKiehtxmKBD+2e3g9/Wv26a0MHdF5HPwC13SazJcfwsmUM1b9p52538Vp
DD9EKjYOT3qelcc/5Rc2Ok/DV5xWQWd1UlWWFwx67SWcvB6jTz+hbyYuDyYusqQ4pTNhU3LEgkao
S6D/ygpgfoT+43IrD7TlCvYr7GqoEWZnAwM2ms/uKOqjHRn5l3C7WY4LJMlgkWPljZ7dVkuj4Elc
USQSigrGfFaLesLvJbvCKm7Nwa/1UIgNa53XCrud6mN+dXUoHXLdkIbnArbh0a6N4nni3fRnxftt
CvHsu/fsT9OJ7PK3hbh3AMioZPIl0E0PlY+Q71ng37LcV9HYdzsxxNM13THF2oqhzq22nIupdD0Z
JALe22HT0eUx7yXqDWo+3nhKBszro8h0QKvhY9oYyO23LWJVTKNmliDRhSOZ0CVEtgt5f8jeIqPG
2PZojMALJVOLh2hg2K+/N+1VI/IX8GYq+v/v+Uetj1+rkgDnNxUk9+i+hem32DhTEKsjd8yACI8f
v18il8FrEhExZebba7uC1ygGqE7J/7UjunlPssuDLvPWRRAyj9VrEMgl9jsZhTpEoL0HGyoH4UL8
RPqs8AcU3PcNI3b73hEHxKxZVxdB91++F1lPjJj8hA8am0iB6ASYAWz87QIvozakukqo1mSmGyy/
LMp1DHJFdkEsBqRiFEb+ANOR1fpKrbuBW6k7KMeJbc8WwoIGT60yyFkgZMj3GDDYNtoVSoBN9pIx
MgThtdUWZf8z1GjS3CMk/8kl0H4n+DkAnIQNoQsJvHnoBisUBMCLak1fEBlh1aUIlN07/2gWNZG3
eeIlKfB0GohYE/pk1YA4S4mZo/b59KmvpHMb7oyOajORlvjp13XbUQAE/eIBlQepitmZflVOT03I
zLFFYKq1XJl6uJvWTlsrP+RLH7Ko9BqTGW9vjVrh6tn+uJVrZLSemszwPI/tZ33em7mbFSvM5ZFH
E46HRsFgY+1bvDfp3qWMSUrSpb2ZFKjbyY53Hw4MfezdZpBHtrDZ6TTGGiiMKt4aLcvaqw/eC9Gu
t/4YDI1CSLwacJ9l+N2jxunjq8EMR5Y8bWiOrn3fiWUbY3UT/lNHOYyL0nMZc0rdmyecKHFa4b+Z
OsIXd2hrjPQQpjcH3zB4giUvAaS0xUSaGp/qsoeOucW86k9D6xGAjF64xtAfGiFcFHe3lbWO9Pt5
XesOb6Rb7Na5RhHd3SWxrr8bk6NZbdlkZvBng/rQzjYW33tN9Dj+Zy289d49xcDbc8inkkCcOQI2
i4B+CEfR/bPP59277t1d4y7T0yJHm3mnpriK6iwDBJ7t3NJipDgf3QM0xm5nXhSgzYHhB3KDSIYh
S788eeF5nL0gGW7UhI6OT66GsRszteoIDzlw3uV8TYz5AFhCAaQTw5/w03GconAh4V1ibCpNnvOP
oqgaVyCwccnX61tRnz95p6ei+VMFboQYNPGCn5Yive2rwk/wLPKhk8H0pQlIh9uvd89/ske1oD9p
vO+NO54UQSmfD9lnzPxh/OGX1Pss4eZ4hoyz3BGq8Kcs7aoFhbhtPUrof2/M+a9YWxr6vvtX8MZX
/lGYDenUhiAuGtxybOG0g7okQA6ZLFEpJSGH1yJ//L+8MBdkL2g0jdNXQXkLAI/bjHUkaHriB0ac
K5Ytja3eWHJG3qbOHqvBUzqA/YN4d9gDu+E5ZVvqTVgPZTd/8F+faXqF5v9ZwsINMmZMqQR6L8VZ
D2sOV5BMczjr1hM6cxu6XVikiK0lvrkmsl544iZUhi4eV0hiIMnQfT8dRF+WcvfbfBhLmSI1a2QP
thf6eg1WDrtRO2jZDj/fDO+AR5i660928+xwkDBJuQzPyvx0W5+3p67vHfsucLmHcxnGe6H35HUS
KtB5IWX7Ym+NDco/4mm/2VRUMjGXnXLNBNJVWiZMBZ3tuvHARM+z3AonaBYgqZqfH+Vb8kdScpA0
79dVuPLVIjLCGswPxbbnhVw2AX3cxKaq/EigUJW3ctzTZFIvfDSbhVIl2eH+r9QUVJr8j1uAT5Bz
zp3zp1CrBzmlbdWkJKnU2V9o6fB/riTkq4HVjTaZ7jM27sOCElgpRE2fItJ8OWTMj2WPFF6VeJsK
1PqQvLh/fPSwqt9CR6GiwlHkcSf145Ayvc/FRbwLcsMaaltrdQkA4eY6jA+SW7Apk+6gUIfWHXy9
ZJwBJkwZNC6qWUoy4a1OBgYjVKObl74EAo++JYwnrkn/MKvjFe6PQoQ2F7BjSa5eBl+zjNXWTAV6
eFJYC5QAu4EJCIYlCUfiF7dZjW4CrIm+boqPp1gwKePDjoNUxF8lecYzdnZZnuEPE4pCvqbq9mKM
AoPVJPegXR/wS0qm1TaP8Z9oqqdnbljWpsLR8mZaGwlLHj24S3N/NqvVF4W8JDwvpdd1GH7q47zQ
ezKx/qSGgLxIqKI69ijnORVNYMZDkc8XisopPXsSuW5VulwqHMhGeq9c0bjs7ItTTFMkz3yumaSS
FqBnaMt2UmiGSKgchgGm7rXBTYySW5mdvdf67QQ12qvkdYq1isICDfPC/4KwNFA8EMlumRCpXP3S
CaiT4+zliTm+m/Z+9LTih+95KgOZq0jrpWlVZrgCsF7Nmb4ghqQB45a1gFkk6fReMF2aImniV741
EOXywRbEIhVVdL6PdJNh6lHse7TXKbfiZl5vs0aBm9LPe2KrihfAHGAEr8rUNrwvdznuSxlQ7W15
3V3P6IiVOym4nJNJv2aTmpSX95WlXEGmdViOtZL/46niDY0bbBwyVJbcDLEOhhbS82iu5+qmaETk
tOCPejmvkC8XSk3/xKrcfGCjJ/gjxGVrEBD15z2Oi8l2MQg8OGyj+lmCvx+3T+BayeCcczAqI9vl
FKphsMOJUknmywt8NecplxZ0sy7XlxUCB0zK/DEqnbGdkyLb4t+bUAQDATLHk98bf17S2nW/AEwE
StZmnYnXhrmLkHS3+G4VBz9zbNXd4TuReZlujzCVo6itXT5tUQqrxLr/GwsG7PfCBS03je9p6gis
CcpUdZ9ZslfmaPiP2aoJY10QiPb2Xv0yonsmTvo/COjD9aU4+vw0rhDsSTDcHm5sspFROUD9Oqxd
IjlyiCMXToCjJ347C2VpVAo2btXK5akVoYIRepliSMdAcQD1+dmxTDVcEwrRrO0Hqxhae6pnkG9g
2AgfPZXQIPSzu88yJJw7mZNOXGgSqXnVsIY2Me7F5i40sz28fFknzv1igmY7/U50pF+lGWLVZahq
sMmRC31iwROFrO2XzSFEr7cnmas2m/dl6R2Lc2gMzBQEgfQiEmdAHBhL1SnlSndPGlr0U3LeYNGb
8/1trebEue/KUOLPTn0jEcSwK78c9usSY8d7FD2mzc1ZiqKG0Lrtea39Uv4Vtjt07tABSNGDM2Gj
bk69cA6JZJrmtWbiYsAYXMo7hbgDeFHBmBcpjreafcaSS5yqahgXLSPkM8LSdjpOnrZNycVEaXUh
g3WjObhfd1TEjFUInheQAmGru0GmJWuCM/5ehBYgbIOndSe18O5wGYqnjjbAVSJIP238jJ7g4bCc
DI/t2cK1+aXisQJ7PCvNoq3ep454t5aOcqAKaOqmkFCN8sF19+suXbkpfA2wA2+jMO984VOWV0K7
HaAqhku3AdV/4FbLjrqLkWCBmsK2k7uxB+dOT0ZPQW3jA47ndNVrBwpln3bgqGzAUIRhSZBulJcs
nw2JB93MiF52eD7OhCNZ/vexja2Ps2pf/yRN2kiGmQohzuWMBbPvkH40EUX4On3EvxYd4werzLQP
UHUxZkxVac1HqrId4dDLE4xDyWtEwpAbcUmSAt9SibCHKDftTLhaBw8tH3lpQfFrXThXBb2Bsemz
7hmDTK/t6aWUrSVK72PA0JZubqRzUhcuRfM2+P6Ymi5ChX5TSz5m+oRtJUTjBUyAOtiGtovgcNFe
4Dm0zm6ZDB2pEKEUtnpSaceMl73hn1IJd3tdH1fGi2uLJElwROsqIFDggX3vbcqkvFM4+j9kpnh1
Cs36oljYsMVOBtPrYWxvq0ShRmdQMgpETXB/vYawbnFv61qW8nIsTtw0FcB31QBSLnEJFk/DmRE4
pd3uooulCNlV269Bty/QQyonXUjOs+zlTua2CKlmQASr1RUife40wrZ7BwPLUCyK6EQN3kpsiEVF
qeydi/xVUhTEOLloxDTAw8NZYI4HAA3fFcX/QfgjjqLlhLzNdTGQf3YJgvcT+eMCUc9jqGw1YMsc
DzwA7fhycDfYlV2SkKNvu1x160GbBA2TxrBEibJ5591VHh429T5/yOSepj7ZIUeM5J735Gtgvc7u
KjYhOGvdGasA7mEZZQp+2cXtlOJc8EF5AJPiXn9a98tkdTU3xqmHAAGw8gWRYqrF4iJoLAdty8qL
dBziLLZfGL+d9PAs62/2PJlfUeFWAVgubnmJ20XF7006x97Brs25e7VuBWOGz0rhOZ9VnRJyaE7C
aF+S0wZ+JAInDtMwYfKoftsXtGSlG+HEvM/UKXdnCv1T6DnnY9U31vekyyFSNB7zBXPEpYRA+4Kf
5C0AuCyskkk4fRYh1aonrcbzAVr4OFnNGGbFm6HcQl3sbshCD6LWYSBHLGKBot+N9SCtnpv14BCE
vXNCdWVkOqX890ZfX+XWC58AEzDWYmDeURJUqlaMWPiSN6JkTmtPhirn531yBNO0d5eh8Sw5Ll1z
dFUGC5+TSb22j6GCGMD1bFuSjKxInj8gwMQbQtp2MQOEXzRPsiNmL5TwfejMR32fE/fKC1pdNRu7
qyyniD9muEiTj5thwO/wOWJBVg+s6DxH4JX2M9tawKncU/qHoB6sV1dRMZCPjnSXORj1fHhrFZ6f
uRGlLj6424C6EaMUOp2wnWjlNPoixVP2Crqy026EwL68Z2wrncUKjJCNeWhdbwhXfX3E2J2ntvr2
eB77Oie25Thjz8X9MO19sdJ3U0o5NUJV5ckjcLYRhnKJU2NdMC0ZAvDdHnCdJT+Dkq3+2ZJC0D9k
FB2rz3dI/y28zWYFc7ExaaeIvWLjxNzYbJHJ0y0h9ZQsdQ9xGiioyDw9T5pquOhzy23h9kXHT1o=
`protect end_protected
