`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KX3IK48HSUiQIxaP65FaQkvUKeHJSkOlKQWvWnmMjb4HRXbImMdI8j2J8lYcDFYNs4XloZPYhPjP
METnWd3Ajg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T+uhQxH37qnocrAAtX8NovMlyWO8oE7ivxMysBuXjeyLOEfQSQO739KM9gJ/VzHupmpS2hODT6id
bXdPcOhpCFx4Viu3ut7uuUHAsJjhngPMab6yXWIguF9eNBaR3X+ZUr2gPuHBTh/DpSnaM0AJs74M
z3lS1KB3le2pQnfU6r4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nal42/jMSZMZDSjlR0MRLrSSJscj1S0fXM7BYOpKQAb9rFfr3rwu9p+93wSd+Q4SQtZOD+oW2tFd
UK5xMnjnqkKNDm+3ZWV6+cR/5xVhm2duz7fRUq8cPcaAafkiuYMFQ8pN2m74Mxpo6qdRbIzIrj/S
xWttnxediPGmhsNFZ09nm3e4F2JFcZOfK+M5csOg4a/UKS3KflLNWtHzv9JUPU3dq4Ml3LkxQ92L
uyBA+4r+wZHn7h7ef0MzcZAYBKQK5xwYjvIxKzd+ckS2dinObDMecsFMFhNVQfwGWxN9WvoLs7Bu
L5qyRKvyuMI67CJTj2Di6aX3AuRxn7RIT+FrKA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n3PebuXzjUV2wLyXyMasMgoEM1euoL87B1q+eOR5v361Ufxy6eXXltkb1lGCtu7DdG5pGHzOtZlG
6FXx1swNQGZlb6gJXy1/WSsIUtn5wjtiYsUwLbfC4Z/r+5NHJEBSGzD4rioD4MesHKzBY0boXgLt
Y2GPksv769STEkdrt+s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IWEH64z45RV9mBVK5sqTzHWQQqYDK9RiVGfquW+h1rwrc15EbyLqVUZuGOVEHX3UkgMI1eEtnODO
DrD7oPyM55pkhzMkMAmjlAFPyPtrG7rqTesqiHIGLHhUax4Dv4clW5zeFufIS9xGilp0b5HrXBKc
47P8nzZCB3Lo4on9JLwFJR+1ufzAUNdROXYKu1F0r/GlsimRjQ+iwnCLycoVVFtTmZaDnAALVeqw
dRaloIG/DBJz8btLpbSS+dS+G65SunMUTrKDdDHkemK+bvPh12FN4phx6Pa6nWAZGt3q8CQ+IPH0
C3vickyhjN3H7WN6bA2nvWtItkAIfOpOX6xH5w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11712)
`protect data_block
jaCi5dUz45L0cVsfLklbIxeU7tBN4cjU8fy/cIPzPXAQHGEon/S3nb8tndg3PNxqzJnHTue30zmR
0taTi1GcKyh3attNVFRZa88Nm3ZZVct+boi+5xpVxZjHjA10qCuI9OWQupttIXzz2HTJGF93UirR
LjzvPKI6kIzBGbToj7HT6vl21MUHIqCeePrBgNZxjvWFaHNNG0RmwC/GWi6YvDBG6r5RZvRIKWC6
MzmwPjb/9coI5Qe7uMoy5EvUaItVSAyroxVllo6stOZYAXWDJWmaPC1k3UAXDtaUVu7JRxn64zal
3xpnF5t5X5mh/ByTiskjaJ6uqXFnp4a8qjPhH9pKi1Z4/uidaGDajk9buUdHzPttq0flFKPA3tfg
Bp50SPKjxY2sNw6JS+H5ljsCwIS7/Ga2kcJ7S537FZqqM2lj3OPxjnRKa4tZnuAqKoKNwlZjlGn3
/gT8KvsmwCDrspSAAP92OWqE3VLU6LPlxc3xPazLdCTytCQXQp4px/ZpgVBdOapPHwTFMNfs45Fc
92N7aN1IVE2lcFjWT+MX+0vrsWoDngPtb854bOTE/G0nBYT6flQj/9EFsaUWygrvRp51+KPo+yc3
O+Ox6s7vPVdSfeMoElXJovn9kdZEQGcXJf8OOD/zcZiEG0I+qn3VsEM5TdzZXM1yAie4EIh9uVuT
Js/js1WiE0n/H1e0oZewb3J2C2M4nU/lG8SjkwgyZgRSgEiH0kdWX0z8OuWBqGL3gUPApl6mpEN6
LjPHWueHH7uPVgkkF3Zj7ABryW2QsWXgyefMhusF3dbctekp9tPVF87bwIogtzUO3jglgYvPw4vn
BoLIgrp76IsGnDfB04N7YAxgqsWz5Sh/8a+k9+QWkHkfyzIf/qChca9Heop+6XUaF26c4yWhbf+P
6ywtoGiWaWXNeyxLBkFBCQUlzcND+uAXT03+wUnP6b5eCn7w/f/KziwAQ4ekX6Uemk3G6vxUh0wq
MjskOCIwpoQZNOMI2xX2wjUO7O94Bu7dSL5UMm8iJ6oMyQUWJ0uTZSJVWhXDYyOZPCEbm6etjJlh
toi6M6fl/BXbsulWpb1eW9oMEQM5TchQSZlNeeJ1n11l2Qv1JCJaO2SAei2hV0H3nNemarLnxxXH
21hNjzU5v1+9ODtdkN4cSA+elb7nkxAeYaoQMyp54WpUXt4HXdzDLm8d74cv3I7wl4ur2JOYXPo4
5F4HFd4SOmVbqnSzHMNhhsRhpC2AZyMu8r0jUC6EaiGRBcZ3zv/wBAZpvBMvI3fiVEsVDzNu7d+K
z53zBZmiIA5bz76YkFsu61RdvU6M0NpM6fRHBV2n3Mo84yqjxjPKR2AHyCubuTShNdDeY7PV0a3K
EI+jOEy+3xAyX+BwONZnTaDHIxIXgty33kC6u+GypQ2WS6GMxBr1lxZprtW6pa7oZgZWD0HRW8CW
kOjS5D43dVqN89aMXSGPywImvvISv4Pqwk0WaJPjUan2nvOj7UYRfgjCK4aVW49nyuD2OHMU0634
hbIFx3LUEqXfrF+JJE9qqSCrA5xZbvX8irmWKOJNbF2lrEXUSYtCKjhF60Li7zRlQn1sVeCot0xn
GIAdDwMroU0z4GQ3C21BsRFgG6TFaAR43K5oJR8lz9qjRgXuK7EBJvxuzxaWwCSJE3y/IWH3Bve3
vbvRpt7lt8hqIER99T+cGePqBZXtTXYlgBoH9QpSBs5mzAxBFd7FkhZ44zy2Kt/+9o8S/v27L6/l
bIgc8LeewStoO3aX3WsrZQSYctynsY/dukNLa7QmlVGAiresb8N5CisvnZt1SsvyfWC+gIv6SRic
RuizqtaFHID/NwWIlu+OASWwStafbBdIXhwIEvwqpdQX+8cvyQBLpAG1g4O4r1iTYsjq7lUpJIA1
BqRsnyV/WvAUD/LKoq3becm2IKtYtFU9NV6uTeFO8B4XSJC7/yt9YguVPs3OYHD7E7yKHnigpWuF
ZZjFoMpu5D+JNOAUVl9tg2L5JZVhwHEFgjfXw/iczQ4DECCJByWYUOJkB7SjbOgWkD9vxISFLW+v
aLqjFcgILavMYSmX+0GY2F/LT9Rlow3MZCinrR90u8vf7pR+bj7QVfctTg9oOF609GwvX3kO8ZcX
EOi2krg6SfKwVShm26Yz142MxqWfeGH3wsueAkra18Uldjt60vsHw5gAOJN2e53bdfPR6rrg44JJ
svealVequkhojuPsVJ2e0HI5OKSayBSoJLwR1JgnxiVJeePEA+ucdVa5IcpCztPVFqtmgjp+tNO3
8voZX/lQ7SE8XqHm41x0rvhxFDO+mCu2dEWHIo6wflXDirw40hiARz6oepKIwaR0jUMDcMQooxZU
FPsxzuMhFwkhpfe3n18QleFnPtnUu7z5UbgQpn8TZBZ+BEU25DZhTFzCmKe9CI/h0kJtXdUrtDx0
Ikc2mAoqrY0drB5YXcbQmN0VwF49rDjEh8vefRQzwQGA46LrbVCFcYVdrYv8SS8B+ERZyJhNTcJQ
FNSBCdSyUV9ADAOW1JJwDlLVwkSdY5dZBX2ZZoIZf+EV6yaaxzXNtNT/v+5z08oEpAIsI53ivJWC
3N6nx6m/XfgqEu7pmmGG4RsPJ6vcSsXkXh7ypLUytsYGz3YDWbnct7+SpxyavOuz4iVHox6AYLnM
koz34AadBaIqAjjkRALbuJSAwQnCUgcCTEXCUyDcVN3TPJmH3RfvN/jgI2yFriPXoxlUYpl+Ecvr
QStCucmpksu3XJBI9cSzE/9fZ5w4I6U9H04rWZw7eCpEzQIog8lB6SZALFjM4+89nbgoglOi3xkm
TJJXmRPH5O+PwTtOUGGU1t3Dna7ya4k6OylmA3zyOfJcvFNrYMRkhikWl4PRSRax8nqIUaGdXp2D
cByrM0iEgHld+JObvIRj+qTJBsFOy3cvBsPevOOEViQYXNzdxtDzbAdAjOr97dQ44eT0pGO9yggc
c5L0CVUpLPT6keNk630t1UjdXkHn0LayFgGYGfdVFWKg0E7Umn0MVqRM27cJrqlRg20PCSBZMilT
gbI2z5wGaiQRekDMz3o26kgFZ+T5W9FeUnoCFHVOiy00qImtPfFSLf1o7s7TibCtU9uw0mD9ydYP
eLb055w80B7wx/NOMgsqObbbYxLUY50IvCG319hjpi5kz8Kw53k0ga7P4YdOl54qyJrVZN/vpsph
6MzY7WJ/R0tgJlfBm66GJkB/8WoNKjAkA8QWG+8V4LRzcR/L+2Zv/CETEmNCRunJ76x45zc1FqZ6
q3JHYFOQgRlPom4JKyOlOhvFMQQ0AUBgfjJy4Njtob7eWyczWz/K0p67sAW2kLf2ww+as2YjaWJu
1B+mZZBh0gCs3Tn2GsOih4mU5BKGkqkJpR29rFHYo8SQm1j+3PD8xsXbioAx2lhOleY+Bq89PzR8
kx7EWto5aJi7gA9eWy1kwyoL6Dp7dBAwfbX8wjqGavEcoxvtyBwknrdQzeEehSNjPgMVbMY4E/sZ
NSETZ9pwSMhNAUP6mE6DGejFfFiGKosDmPt2tPlWz1Z2+GFzJ6gaPGVb77BvfVCjbZ95yRNSVd7J
vWNlEenWAP8W//jSSNr+9xCeszKY3i+wwKM5g4BCqJtZRjJhASP88NQrp/xAGuHZOYB2+t16ClEu
SZzjLVivsgIgKbghz3dy0L55+nwa+AxGBOGTmcP+xJHuJ9cPL84y39DVlJZMOo2XcN8zFJNa8E/G
bUG1wjI+aWPYitmy8rrhDmP34CkaYmWkjZq6/trqBPI6A0kWqyy01z65wMOSgbs1jCeE8zTpvywa
UeK4KCq/rhy8legf60CFpV77sndUi4jaWpPI7RbOq5jtoaRM5/2F11JwdQLdGWyeDuQDIemhlMtM
6bKExDGfI5LJYLdSKBTSjvONhFTpdHsvYnXhfs9965CYrdYAHYksWHh5JT3Isej4Ok8tKN3PpwNz
L87uJlK4VSqzu9IFLFS7F6GG2CNupgNRw+Ea5iVnTR4h8FmY6XqyO/ozBfLixx7EsS/rxgwwBnLx
oVotMixW7PQYnctKqV87Aq9DBRzjK/qK6mMeup37SvKfW38thZeOBzzO+fgSUFAel5EukhliUEYQ
AsPnEnHPiCdbSbI5qhGRBSN7Rd/Xzvv6ls+xGlOhzhVcj/6fKAheh9Ve6zzHj/7u6eFss803Fmei
u72KuTiOOlkifyPBDgx6c9qZ8LnF7P2EXgL1JkmTGesIg1B5DDZbMjTV+21GqskUN3uLJU7/exsF
oCWg6QsZTsjiDEihWJxkqTHmZU14DLsgIqzAOCJuP5j58YoFbXO7dRGnJWogHyeFZZAl6qK9y5Cu
4DrheEsUBlxg34/KSP5mG8i3INuDu8kxlnqJHs8JCd4LndorieGY+VcyqyYGsPShTzxnGYinWWJo
s3NRqEe3c7Wb7UdZy1prJw79xQHzrHbTvetfUL4SCQW2cXwryjERIIHI0vLsbzErBRb+3rouAftp
Njf28yoQn711n0ylokbArUjjJX1dAorXAfhegQw9eGyq2HSR5ZY4rjHjBfI3pBCVodfhE02SToBR
hElIMR4J1/FhzSDVs75FTL2Eh5kVwH2uc66pvAlPhDfolRCEP++gCgzkDAu/i63+Ykdo8jsl9gyx
QYrSpXMOIvHnruSLj2wydDZYa3AdRaFA7rkBTB3iGWEGdNHZUltUWyMCXaBHAvRrMlqKwes9gNtv
ppi3IVvKucRYjqankwqEH1KqR8lWaLIUlnqRrDpJ1zgsqZ0uy+cUwI2FQHHjGsXu3FJ+KNSLfywa
T5gMqGmemfAhcHuI9oPQe+CU5uzsOdRr9glTngI6QBsGB7kSCfSp1nVCPB17Sr/q1zM/cV0REvq7
bnUFQXAvOmfdLU282V6DU/o2/9bLKCsLqg6l1y7zyNuOc+6rOtv9IKVYimn1fGawFHYssRUC3qPP
RwWdGUUTmwnBRvWzVshrqvGpe1mU8I6vnYYqOVF7tf9y2p05jGolqmH1fq4efxV0hlaTbkQToGua
a36fe69X3KCKJxbGyRcgLe4TUr+if9oVzD5Ff8rY6vnIohyL02S2CZHs09YJHDxE14zEUfnVlrc2
rhVlSVEVYSWAqfgOFnVGHvXbr7F9PqqGsddFj200EDq1yDZxqOTAhCfpboY/TQKP1dLV8IbXtUGi
omXTNVz2/hEELX8nk8+qX9j3p8+90NkyV6uhiTiWuO9PSIFFSfhRrXzjwPc10I5BTbfeYl4Fek/H
3z/eBYWNLgGOERK/5zxU5xFKgm04rur7eKKWqzQ0GFtuRd4Urj4DAJUGWzbpe8inX+rGm5EMd0TH
fFMteaoengQlp2SSQdaqnR47yLJBai1A3xSgZ79GxR+ubjKBBKt9YhtahK8erJ4woTvj0JQp+3uy
HslA7BAOVbPVEsMv+/84hQ0gcWxSnWuFG800ho5jMkMnImsMgmvXxxLB9kM/y0EHOqjFsKYmNzQq
vxuU0V2kqQmQdAJaO0riENb63ITPYEIldLMb7dLoXOC4UwnIiDI61K03xeU3b67oR357In6JtOWT
spBg47NCUtlA0bI4KfLrjsJsgaAp7KMxJZCw6Nd+pSPjV7xdiMcWN2c5ZzjMfMj4XvaVWvS0OWA3
qSMZ/ASE16g6p1ZBrm6VeHe6RpXTCjgGG3nQgiCCmPqUg0kfWU++rB0f0GBycE7hT64K+V6JC3W3
N6DzRcwZPhRQ9KtoD7sXzk2s+9hqAVcs6efme6jJAUJM53eQoGFZZtWiA/1PZs1EGLowxP8O3WOA
+DwB1nEXUXtHGzfiSKYTK68SX3L5Np10h4fkpEEZZMO3P4o9gaZuHzIXydl3yKHCTgQNus6jZ1Cu
trODGrv1qLJLYemUW20gZN9g3LcPM2E/X7jTf4L0HWpmaN/KueOxkvgifETzvUJHUVstqmKeKHgw
ASAppIHZn2F7b1NujxX2wpsxvZ0YBad6yiJ8LEeLX4rD8Wxw59Uhi+ZdvUuY5N5P1AYazM35XBSS
7vSI3cqSPAxSrARZ4gG1mFz0hFSZVEjQNUMKLIq1+GPYMaHHar6NbU2kKhb1VndQfb14JaVNFn5L
Fpdgah+aNkS1TrdUenPo3g18LHuymxP/+4GYOqHu1IRgUmLzuBnnXSS/+u0TBnZhIlm86lh8MV0G
fdOs+dbvNqr4UU8SrkRZ/IWyljmcczBbrea3AQAdNeyPdHzRnik7bUQePhDA8lq5J5x/QBNMzZTK
8Mh0vAbDKWUyFauQysCses581xI+SbvlWy6+IMMpaK3c18S2fF5uNypoUk3BeEIG6qWjIFFvpDmP
TceSolgVhdz2wds9izYiUquEExDrJ768Jx06A3o9Vl7+lbV/YWHh45YQO0lqjczSeNfz3Knt4ZzK
7LmNuRgWS16UEoOomAa7nqYS9HhXltoGn5LRmcy7l5Y7DrhZSBrug8ulmbu2aVe7EuMYpQvVm3Uc
r4K3bEfBl1FYEFJY4nm0PtT1K70I01DWTu+rSB4GkzyBdgOh3hzDLNi8AK6dMVncPUMz/J61zbEW
82XFUSuqjC78CCmfjt3uPjjhUsQ0wmgEcHg5dczvXKSA1lXkJwbed1B18p/YMCyVxKkeDL3Zr2ct
UjNcozd5TFhX1/tIecJvKzIW4Gm77hertn6E2VVtS+MoNFbKzo9CK7+fMweDQsdaFjwE6zmKXTSY
x/aPaBhXLnVTKqJCLPikm5jrG/ownHoJ9uFARBE1tIkZdQKab4Mj8pvCp5mQKk0S0vB5pe3DcdyR
TFZImVVfZhaeo4QHl8sJiD6Y3k8abhqpH8giXssw9iaPbY+vK8pH/uKPyLRl6zld0z8vwSKBVmJ5
t0u5iVCasJHiFKNcoaCl2ivb/lgsqcN6eLJnVBwVir2YcXKs7qk4I/L5OOLYkLc1Lbyf+UDeq5dC
Mz1WPjwQgwEghuoGvIqY7jtEt7ijZIzjsGC9Uca1w96z6fKcOe/uQDMnbxW8b16zCG0xvEcQsji4
dgNuluH71lnQZQDT5ycTxwX41T3YsrOnBAWfbUIz41k2+QgBEPoRErPTIpjSKVs+BIOSvbFhaonL
L1jh1x3HETicS8rtXvWBzkq4NHOEUdKribF41oCfC+KGzGAPVSBunj51K5ePaT/WsBXrGOAwHAAn
9zCNnesug9CwZr56dMCDokF6crW2TdBUnofqtucCq+9mREA78SIv8g3+fGArO1LeMvDgTQgiCpYu
scFkAKviMApecDcF0t9FNWWaTjcp28JOUF8hJCGveXMkrCoOWOQIBnbs6jdpN7MgJbhGaa3KnPh2
YpmZdGG2m5P1sWKTuPsdr6DfB9P4q17eSlAVt3NHg+5E5zEqW/jtAncUjrLHef3Xwgztlx4/K76S
9yuW+3RKL4Sx9ljil3ebMTWOgzUtcWCcHy8fYq2VhE7bQqZVoaIlwJ0aY4tXDT7yvDS4bV23fW08
ln9FuXLzd6YSuUTq90WkhyzBrLPBW3THbK1Ljr+7FE/IloVx0WfpHPAfZjQR3KJqFPy/mny/UEXO
SRzE+gaqOQiP/Pd9toqKd76HFmW8SeI0GuyDNPQwacADa+dzoSvDwDVk7fPS6idiiGE2+ylPBv07
oQ01aFwB2U7/rSIB7WwV0fpa7O0nWfRt0W1nuWrX/MpHVq4X9Hihu7J9q+lOIv/Xlix1AUQn/g1a
TvT68W7uIABG/KpEVZUoopMyIAF2+YZ8c4W7fS1iUPo4KZVz4t4RaskXRaV0EBdgTeL0mZv6Ivob
74hjQAjASDgOZMFyOSpDnvqvn+GjVBb4zV+WofpqIKYi2+8qQMcMOAjLXksMXQ71CO/PADB1ByZr
n+Sff3vUxRBv7Z32gtjdRXFfmCfheyfaKkS17iz18ElqNw4u4Dm/VFLjDFEob/ZF1AJ4YHXtTAvS
cGT13PPNQLh+abYHH3IBcPf40fEFTQ0IwkmPdV5Evp88mRr7wYAPpE5fATnzh8SICcH6UTGzzF4n
m5MDTt7a3274xTifgzIkf1pr6rVeSws5BUbH8mZLktEK509fFJTbUvxDJLeLsfCuvsl+dper85Pt
jNuXevZpuMlt+LTnxlZtUIbLkG8q9jYuDQ5iLG3U2fcZwhKQnEdgPMlripLhwqDOMi74Jvh3WXfm
F6W/nwzUqVdyNz0ytQm0JLB8L2vgFgX5ESt9gUpUANHjBHQ/o49mUb7mnG511ncZIoUA1vDVamaP
2spAm9fS/q57mmfMfNSF+4J1xgbBaJvbejF6PY1RBAu1NIqeP4JHxWp8RFv5hHi4o8nM2T8Q4wcC
VS/HjtuZxl4lBsXM7p3X+YwSlE152ubcCddDnf62s2SsmTXnn8lQJR9hz9ODESVREQ6FI64N47xX
eJOrAS8wsY25rxa+TLNPyT8zx7gl3bbixjxk0XPEz0WKdg0aZMPiaXjaZyBUeEs874BF2T/NYWT3
/s2zVYLHCVwH7FmepgbA5E+LPUDJJRzwuhaYJ+UbNB0V2Lvb499v7bvUj00r6b2J9Z04KyCcYypf
NAgHoaHmpAovg18UBO6sw1hglu2ihpN8oTTxOBc9yC7EKC0yUT4kLjvd5yl7KXxQwfI+Mjc8Xjky
HTe8NUOwhZsNVl3MLuXbdOq7lC/xompx1/nSTdhU0iVCjwQNAzbIrjrmiOfyL3/mrtqbBsTZGeq6
x6UG0GAvVmpgL8bzxFt9lUFV4ZQk+suIe71pgAj2h30RHQdIhKiLYKx/iC8RwqdeNzaGXlfX05lG
WQ8VR+rqsggsoeTUfGxmeghSfGOLgCJ5dGe8CDHNGhB/84p3OHle3KzZr/g6vMkWoKxYX1g84U2R
FqasjIpLmvMTaxHmt8Ki1udjZoRBVGvP2Nv4oXuBe+5F/i8lxc6Dsi3wiUAU39byncH4rcFE8SVu
mkAGhgXC5k7hwaZ/ESd6F/V+3VMe9JovyRztERx58DY3XL4Pub9MUVaDeQ+jWHknJ7bUrIy1U9zo
GpAltQTdNKVc92QzodU6b/mwQjG6M2g3fQDxiSZTRFrmuU4zvZ8g1Dv3id9+nx8Jp3qUWvuNGs9X
y2lwSIM03UgdlDFXmi6tdBQiIMTJWdUFqSGzzDBZ3TEBd+YEAzCKmMJiNbg01CvD0xxOsAfihXO3
h1jInf/ZFCGBMbKMMq/HFN99OZE56S2B1LIy62qsk9Ty+IVmrdku7TVd3I6+OSdA6st3O0OIKSu5
r1PaNRER5erVt9ObVVAEYxqH5Ln04fa8wdqoBd022YFLczdL/jMly1TRTQuMhMSeaSs+Myg4p9Oe
T5glzaXpgl8KRJp99raTuhXTkKhsF0/UX4yqTSB4DnZks21O0GrKQiUPQzF8KpNW4ZDmUxFXCKF8
UA5eEVglF43LhI0QTUarMrZIMJdycieuNwwu7ZkgTmdFCi6E0farL3ssyV0i4deCkKINuUWvTESb
9+wTwtsHixeRik2FczzNiDH6t0P8SdvRr+QUEXYCgRnpfuAfbmLubJX2fPDSoOwBaFdoQ0X2yS/v
MwvUTWb1hNXiH5iFzYyK9dLz4kX6lpqycqwcvhqqmoXfjUelnAcmxD50fSNE6hriarKTds4GKMcL
pc2YlqTtaiKwRjXFZabBGw0XSuhzpOdJZSxXuvHN8vTt2VaKj6E0SfOFKDNA9pZKlTMQ9Y9kN5BW
7hwuMJCBllQcQLjQRHcr7DIKR7hySbtc94dpaURLITwi44hjI4HoHR/teCK2DVolB9Q0gpQmJ11A
Eav6Vlk15/wAEHZrkFdR05G4IX3hrnVUm8Jp+1srbYWmb/+k5jJcNPRK77Z0sWarBbRef2WXpFry
Li1QIlV6jAIqS/SqV3dyEhnuI8132Hdessa1YQk+UH9JSP97euFHmqSqdZz701KkkshJZ6acqvxR
Pwk023B5SoFdItY3ltWx5ouu6r70wNGxiE6AOOCZX5oUoklIeLIAKjcHl95c/XIkzBY2/zcyYB+X
W4V6Qxmg6fa4EwRGEQ2EA3XpAHFvGhJWQRsbo6eImgkklE2LA7caZJWXPIJhGVhcKevx90WGF9VQ
10iQ7rtt0e4BVIcntfnlkXZ1attdp09piD+t/znN1TmMFb5CQs8/FJcLKJb2iNBiPiF4ugCzM/E5
aZzHvhGQNkMOeptiyxj78TxxoakqUKO93NJWepPdgvIawvbqKDzCrOAyaEQlnMDO0drr9VBbOShq
w/joIrtvhsGwYcXiIGH/mvIKrbhd1Uj8VGw77sHnwYld9GZKmxWmyKVrnYFxUb/HneEhrMpRbu2x
Hv2wtD48l+a5DBkNL+nr9bqDhNE4B4gWaJFFIAzTe6fJsETo4jsD+JWn6KbAnUgiuz77Hm2DMcaq
mY8ayf28RqTN4R4bTri59yJwujhxDKBNJYr03JeInnwxFV1ftzsQXom1c8W5GBTf4UUeOu1VpOif
ozCO2mG7tySUf7EN87tEoQfC1VCCXCAsy1vLdP1JtahifJgidfNNefHWiL50VSKlYDZmXemKVfDG
iZf7v6ebmfFMNCm1E4LmY8yqD9QSppHRK7mP3xrDhtvzFAismM4AdHzA53eMDPG8kugnArhA5FEp
jTmiveeM3xt1fiRvPpJ4AUDRq+Fp+dMwwAHd2y9pf+m1ixF5JGk1RvDp3r+atkBeYROfVAXghREo
uDRnWQh3ZVsC8yvsv70FRm4Hx8ywJHCAe223kxInfuQFqm7DZBdmhM6Hp8CDOFuSGmLp4s24LTMT
Nb87cgKjltsGasjLsHBRKve4f0dZfWSARTZ8rHXbhsHIct+zkaQT2OPzJVjRjIV10EzwnYMs7kYj
H/59msiu3+GCYkHQEyIQgcrs62ExnDRP/ljlvpM96PhKahWbd7lOUoqwPun6tSqEaQKUfOu8utfu
ik07hYYG9bLzAhKMxDFNbVJ8WolxClbVvUeTyT8qZkd1vavIJWTSXYeYgXkSQTBY6AksnWteRB8+
oSggtC6X/gu/zYv0IE45O16rN53uWaOWaRTW45asns048upH3bF9VSnGsvsLAyMSwdF4mQgKcLDr
MMWyAoQzPp2QJQBtzc2H9E08OsFvFY00+6/ko9EHwQJN2tarX70aHWUJqwoogPmLCtjosgbgKKlN
XMOfSMDUxdQn3+5g/fMJavyPZoBoDF4H1vUhT6rYyNwyTx2gp2dlhkwXfOUQc/nNgd9Sdlg0QwX4
8O77AQ0H5Iody+X+3lUDEZstQ7iEVYYLhQg8AV+q1ffBofxDVODTWkq/Q03RM8K5zxLpO7+kyw5j
Azk9GIzANf81+/VqIHrDslTEfT46GoRL8cKB9FwIIfoiMoKOyjB2jZMe+DcSILTHsvUy0E+gr4np
7Onia3iiohNZD76BcU0FkvXBN5oWakoi3Uz1BDpXde62HnRGWjzkaR1FkxOUd+T1GZ+OHJIDlgqw
X+CEJcJlGiG6QCq4QLe2jIFsCHnS/0XDyLSE4UgOA+iboumz2Ejx6srM5WMyt8iC8sQK982D5Hke
REfgzCz0RY5UzoHWLc1rF9vaHDRMM9yG1etQeP8kkIjPzJvO/4VmsCqi5mps1TL1RQRPwGP0701U
bVtHZdldmVmfGRZr491GIVflzcjt0lyG4JzuOGV4Niof1lzVhc15M0gaDvAAcVkO7i83H/i6NtW3
ulLRjr6tK5iVeoJLxBCq5b5dN16oP9U0AtJ8t+eXQnHqCWJRxDrMcGsFyyRzGuivNlLvkw22xK37
uAeaJRgaqQhoElB/0jweafacASC4Yl2QjWFoE0qMOehN1WVWo6ZEVaKh5uvewmbzMo02ugVVHbzF
lq5xSIdRUswkpNpejKy2bz/VirN2WjRoQtSfMlPEmQk8MNKBVbKacwy+ZsakZFIzPD06Tyqj7AGj
UPatYTZDVI31DKttm3XLXK1hdlafiJ5C6MEm4XsTQq5XtWNqB1P2bUXPWZJH0elwIv5XdhuFFZ5w
QsiptY0jDCqxrN3f3DSIQsnDy8Hl7m5hXob0Wkq9MnyaXSlD7br4xTIp6D945/MJ8kZOcFGF7kGj
Y18ewyIMcMBmqTprS3pXetRagPX9PYwJuXOQQIqGBXVkZd2TSsxWfbx+ke1wxEOyR7xtJ+mj9olW
lp8ak8bY5JBwCRBRpO8irv+L9ZWHsBgE3hhnKoS62g2fVXjeEtZg9PgIcEoY8nYbHXbmTLfH9KP+
+cm5KKjeLjf7PiLmCygI2EDAMyZwXlcNfMQjosAWh+FMRXAMYIi833uQeNO+Y6C0wAdSaMe7QIeu
oHa1S6QMhLeBLL8OhuSdKBF8dxTa5WLfjW0lF8l3YZV5vkTX9uD2F9obyQWk1/MfmEIYuCcyLNTD
Up7Bsj+tDg9krc9TnqgrPXzpcUTkSUYNbup0MfBaBfNN1s1AMtm26GY9xKyxR/vd21oCpJTrL8Av
+lGBZud/HYPzsJ0vEz7sAY+fxNwUsYkr8keXMDU66XQHV1dupZOmLSzZCV33HTCoQvq19Ac7JGaZ
Kp3CYpqwvcAhbOKsvU/pFicmLDbG2D7f+lWOWzofcAda/bGo3QvTZ6R8JounoOXYawNrBRyjZGk/
/ecTIRPoqxom/n6g5sFti1Be30xJLpsaoMgvf62xsxhiHUGYnI2D8xl5FquQwVW7SjPsIa8e8hGV
HObqaStRKTpVhxDFnUGu1oDPnwhrocRFu1wy4/qjl3plX0x/RKZz7z/Ac9APiyCwSmjzSOYXtGXd
VtwtlDWzTajrSTqPUckjZOrwOEIedUao+7KeQdGSSMcSJI3Q0OcTNsNp5Wq+ql5QOES/KD/Dd2YU
/QFQbs/2C4xOVK8cDwpAS1FbgZF8qcfrLAfO6mptDQeJGAVWHEsnXskaiszvDKCWytg1jCb7JySt
qEH/gSP+FRtLF7ZdpgXlIIyJ7HNKLwegw21kRuB+Yr2YOTS/nSsuD7ZHM6lOiD/QmJTYXLz4oCy+
o8wkTpbndV5yoG0zGN2wWmzdJK97IkYSxD2Hgqfi1OiDnm3DsngMD8r+vPTps5kMZtVu6Y55+9tp
N7II3R0Z1aZxK1lhcJX2WoDnPI6Bo/3Wn82lmt73nouUue1XuR0SZTjV5gFd69eJ5fVqfDLE3giB
fIv49iG3+p/m1aG82H8U+On4on7cA2a7SiqNB6zeUZ+cmCqqPnjCFtmNpTiVLMrUYrfUQIms8QWW
uoij7jc6S39tOEcMzRRgTFyng1x2ulI5m5xn3shk0s4j1g/lncERHUfvCZeePo9/oDnjN2/v0235
xu6xNrXxNlA9V5JGlokEUWA+f1Q2krV/WtKLYehvLIDZEQx3GOdoBd/cYas6gVbL9TBR5eckXxHz
o5Kk6NKuCQ2w3m/GmXpwimeRjiJSZUn1GMwGIxe6QsQ9DE7lDESX02zTb3g+/ZoyZgdFZAf1Ypmx
/k+N+tI3yLql6yxyA35ALTX05HSAgEMyr+L07fJ4ahGz4L4bTBakebv44kuPPG5fe+l2eJI7culk
b0D32974QKOrPIdUXNHYki4v/MOemlY6Mux4rW1cfDQLgiHItvGfdQ3aObc+a6WlpbgiQlyM8VEP
EhT/JA9CZWoVKx/AD9An6//QTQQgcCkqDvaPxdNseDeVUoVywQ6Khh1v2W84BWDlEJibxB8G5uLM
AGe8c8Zpjo/d+jLkWIwr7rF2mNa4uCYTgFmYe9Jpa5M8gI2k5E4GpsdQsqd9L0WMx58Ccu26p5hY
uktZUMaPf3047Bv+jTf/jJVoL3LtlDZPO1KfWeSVGreV5C1aXPY6Y8v0qifP0OFCtu5lcrSiWnHY
cMWgFA8/tcoBsYsNQ85f80qTUxWnjLMW66qDc9aabi7J1nwyfSns+9SODTkYbkM0xDmUvQ/vqx7Y
aVpv3/TXTpxxe+DcCuX1fxHVttPNJ11iXGJYZmSChODO2f+sSZNw7OPbX6mm81NyYPpurCwhsVfr
Pn+DELnue/mt4FG4hMSYQILn7+skgS+d6PQ1B8s8wsKdxxx/5GYopYU4Fb2b/WD+WPZfDetvrt73
Rze3V0qZlixD2jXEmEfo+jTbXrU5bxnqMA/ZwrZ/dWVrXfr9VEihVp+6IBVB3hRu3vQKcehYM1Yn
+h4tUwOzrlm+M+QbzgMR4HEMg+iXeUuN5eZRHi/UMyOWu72ExOWkNMfckYS8v3jktzFLeW/dTEvw
55yjA5jMe60/bUIpDavTOiezBXBV3jiaPnoqVr/lSKHJf8RpVMUjQ8+P2foREE9bjwRe9xbLM8ps
aV9yxIEHA2ZlXK7gsVeupZzO7dchQapVCjPRHnZqhDuoxeIWpQXFcRY/9oTKqxINOxCQ34BW4sC9
a+kkmDOAs0sGqk5vlM+SPjdLSo7yic8+chLEjmc43j+5lwElUDhI6wX7YuVbFOFEEdHdJ6NKWJRg
Gk7YwaJoyd13i3RoM1POQoUWB+mj6rxn00oJEwj5HKk5nEfk6bJPI2kadmbfQVavfU13bzuszGjz
UF9V3TG8TB3i/Tpav8cnb+N/UYYjP7XFFMELQHZIB5kWVfj6JL8Oqzc9WNXfDOqfdr5/vtE6FjE1
uuU253O/PpdPv7TVEfeSdkFWvvdm63ihx51KXSbjG/9WZiAv2v2yRj13E4g4V+6wao64O97Ymx74
l2fbcB3QLoFEZRxWXAplP2pf9dPmM9drfPRovLkFw8Lokfht6ezedTwAJnR7+A9fzfp5LnCyrdsE
5sFeQk/FvkTI6m6MnAFF1KFDdWOJQUdpcPfs6EG8bzPobJDf4Uk52fo3fMDOq40wdtsP6uobAFyQ
BGxEZ2vYsr1dAm3J25Gh6gMJSUR4CebAiVImwc9vvfMWZ911r4d8HykJoOKgVy7RjAIqvxV1ySny
I1dv7Bhh3Td9Yu4wj6/p6jbJngoAJLovgzQnaBFt+WlcqwJOFOSoMHWKc9sLX95tQCcxfDMiBKOg
SKccJZRFrpsLju/yyAWVN0UB7HTuIsRFt0Yl6uaSSfkKrcblhqVHAd+lv/b+n31NyL0AyhmBL2c2
ptYmmM1GMQeCguFsHhwtZpbLIccyZLBjVuMhV7wITkvL3SE0jRLkDYrtamxl7X5vAz7ZQQLrjg3f
MHFhT2nJxrXoHMZgh3kFVBTGM5aQ+K1QV5VmvGwlxKsnqQLVBiojwkk3sYT2LZZ26EmKDM9BenRi
twrqoZ7SXrrmC05/JmwCfh6A67ylWRfpIqndD5iEnupPChZAr3t6jwDOZgftM/SEHn9ERxahA7wt
FP5VUrBGzO4toGXE2KrL8IGmT1VKmSKzx9PPqKlatPectagk2nlOgGiCeX2msAv4hH+lmI7xqtZN
avymIOmEh0IUV/kKwOW6aDfDQUL0MJf75LGw2oxm51TAkJg4F/VCurKQQwJFfFvTn9Si/we5ueLg
+YdT2/mlOojFLnGTszE4UWqZEeez1bnvhShJYicEydu1k29jWzRhWNdZnSVGM0t0UtSqrNpG16+v
XfkDEmTh3BlX5g/JeTHObu2m6XPbe2SdqLgTj11YvTgsvWMjxFoHGztS2nAC3dYTKhQCen7eM9SZ
WmQ9ms8nJ5jE6q0GHmipyfpbguDYpWdDVg82wU0IRGDxZuEJR7MKkX/2ATm0thLpi+y2PVPIrlwC
zbdjaYFY44szkD+JLxZoeszbi/ka5rXNs5Hg
`protect end_protected
