`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GVgRO7Dr/KsjnVa35ieIUqOl4nqUKmu8XsjgW4UckaPlmajxFL9W0N5oPN2UnA3cGV8L7ALNikVv
1kAPCg6Bvg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bkWq8f+reSrHy52xcAyiQE0oA2m9qup51X/HDFvssQqEzJrKhDENiv8uQSLbpPulVdR4ZmnTWeOs
v9PQfvYyDJxEX1pdb2tbbhp8NIfz7u/RByiC3xydeBPYUxtIWUZ6VrLYI6eYb7AFTUFRLXxKi+W7
MBjtq0jooJMKYMxl7JM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qxSPrd2yauidnrkqnXBq2SIFZuTeYt3LAMsh8r6iVDhFAL2qfddoX2Vq05FCdpzJ+SMOi+pD83+V
QjXo2qa+tlRjvW08+3DHtUfpiSuODST0ZMrvbSC6n69/T6AE285Ci/Gb+zeHtsgXQjctURZbqOi3
VIivc6V7135r6gfK+nJjwc0VQdmvkk7PV8FNU1lvgqM8hwofAj88v7DNMGHYw/aGeAMPGo+geiHi
4V31hVWpZAMEZZTc/IVAqhPIwqkRpu2OTe6n16i1V5xNvsdDhGcJ8b7wLBAqvMK6h7GrXKJ29gQ0
Kv9ldlCYdxvJDoLphfmorjKhXu5PnbLWtlyUeQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LtRBT5aRmHIdup+rQlBa3QhkBHtfBEOGSBQZQ7Bqj75D7A6uAv61byEeNKPc6Tay0oeO18s2zSJj
k9R/Ewl4KveqGLBBh5G/fatkgyS+hOfyBw9uY5MKsXu6IU4dKRPU536sbQ3kbGwV9WVZK6y9EEf2
cVYPT/DXNibgrYnm9y8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SkcYV9qXe13gJBvZWoWJgcZb0cO19U+qA+h6jHvcsXnyku1rL/E64GkomYdJtJ88v7BfAmT1Del5
+pdA91cCgMkIObztKiQHDDZGHZOVW1u65dpqje2LNOVc+gQZVnzcf/XKjl8tIUGQhYPlZzErMdCt
Q7F7rnsNtawtK9FRR/CF8w9ULwQ6nDTT7hgGyrHgUE9C4cgCNyuzdXdY8D1oxbn1Bpq9GP74ZCIY
4ivDWlnNOb8MMmNQKrHQnsxf2+RT+BgOdd7C0Vaj1u2aNzqpOl7iWm6Sh0ihvdePfXjjLbKVMeKr
b9SIP8OsFGOWkA0xNe8gZ9y14jW5yP6/BaIJGA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 448848)
`protect data_block
o3NtXHCO3r5Jzy/Z/xvOIfHtptNFHPkwFepo574zeFpSNaItLhfMKstxz2BRSwbUn2221X7kNWaP
TRM+El585lCF6TpazQGKiNl28PFHJiWjmgScFfEUDndfLgtudw940DnPLGVaIJolKWRua/SQ5uaI
W4mMZ0JtKdZNNkfV2rU3WtnC6kF/2KFU91eBxb5Upx9CY0hPUd/3s/AobH0hVAqRKOij2IIayeY2
cHNun14+T/QQSz4eADuzVwQ7ddH23NWUimmmaWkvuQSkiTE/nq55khr5xCrWgwNOoMuEXD2KvZNb
GKvvd7ithl+gHejd/ODqTgBi38yIs3yU9tO6WSQtBHF8LodPrSyQdK3sIxCOiJxJeMx7ypUHjqh1
bV+/YYnVoKtYzgl+d0Vjq3//npvETYyUBa3N+r+R5/EznMKg93jyNnu8j6w+6fPFvgZ+hIf0haC0
Rlpzk/TC8hIn+P6DaPbiFWtBmgmuLprmRwG7wtoGthBoBzeFfKnI96A573OEkvBS8SU9zGtJD70x
dunj/2kvmR0xumL+tDdsOIYxIhVrqTdcLlWf59O5WIBEUcgV/EpM6Dz/ffaJ0aSOCT1NvBrnLlZL
s74GKLXa+6jJ/3DL37iH+c1WjVfGRQg+NGa/HZwFPtKAo9xg6E7+2HLZCOf2Bl0ln5U0sb9KOFW7
/NHQBkz8hnUf49hMxksTbnWlfaXHmc0nv24RdaeoAkELl352EvI+X/xf/+CwzxHZNmfkbiwgINQa
PYtTRR5Yv1k6mJKO54KqSjGvB3vbf/1GX15GTn1Em0krjsKYSSi6ypkj6yk+VQKlBV7mjdc40S4p
bll1vzdXN3pC6tz0n0A/EPiX9ngA692NJdh9dBDUdxVxKB6Cy8kG2ZqgS5QcnL67VSLqYXODAx7n
qgrvcRlvaYkdFP3j78yqXX50dywV5OYCBgJaXlR3aSUzcihCkZ9QV0cxFnzZeD8JDBfLT/uSwtwx
7mf3fntDz52bJLs1HAWDc9OIBWvn7T03Du25FDTRBD+uLwi511gFLJT9YbIkL4xKI8sP/jEAj86k
7ioFtXCQMnpS/laoO0x02ptnHV7QYafL0V+psVAuFk5lzXiJfPoIMFy35AlvRnxoEkv+Vq2NlY3v
oRa22O9HkEaoezpFkm1N/T7iNBVT8Es1vGxsDnxKhGwJoJXIQBWIJgTx6r1vM3cL0VHs5moygbPr
q3t1ThuYAXk7RhS0BNpD7stKtYw+YlkqwHyTpWXqvP4hG2MwHJkFAChwlhFBBhV67gdEHpXTQSky
L/gvARaSN+xZlVcpcujqU67jEWpozfet7WMJ3x8U+mu+8Deu3AArIM9ZORVIfx70JURy38JbBpRz
V5YKA8HQswNzKyQlj1VMY2RDiBLIwOO9xZBHM8VL9Pdco6o1ylJ6BkhabGOCAz8owHoDAjZ5NjEu
GxUwZd1DmZjtqXholXb6XemARfOXXPF3rpZSe54PnN42jeuPqFxbAwYclMJQxvy7BOCcTdE/BJPp
fFocdbogPZwAcYQdo9WBdP5dRnyCFhOVH8PYcUOcPlvsrB9dc0d3X4zIy1L6XYWk3vRDdrpbcKV5
+k2nYhiq72Q4CFDp+bl3u/FHj06P4WWF1MAu6n2XzjAnziNp2nHnYlTRL69m2tzOSfxEzxZtgNSz
xgOpS9FIZzeQQMgUIU4XMuOaebmXIhAtDQXCokZdT65A4n7RuoIJG7ysf9FmFq3hi/Mt+6ej31+I
AO3rlR+XSpxwqZwh9tCnc4ALBojexDaZDADz0DOeohRLp1Ws9Ngo06oECbNEcPNCTyyiJWcvHcmZ
rYUJTom2fnikX/v32YXPw7PZdJb/lYNceV1tvYuKTQ8IeLodNM45X98uMn/njQFxURhjnZaqVoBD
QWOJzPiMIgHbAqwMnozA4J7TRusV8HRNueOt7+5L3M95JLRQfQPYAMt3tRRcrur03MUIasrgXf4I
2cX8Um5kMtepbE+Z0NM/t1lkGr7wbHEu+hGIA5QlNg0jLjwMWsrtuAtC1KOguQ/r4uBWbzXxgkx0
C3v8fkCVt7JQ4e5oJbfdeYQ4k4Cgfn0Fijv/TPTD0nCfB8vi0T3glvmMFjZZ8GHnwpfkRB0UNmwA
x00brk19z+VlpkSW61v5RyUErmlBGEp2gOJfe2IcDa4qM4oo2bhdVmflqF40OGi6IU7LaHy64b4m
RzooQd7O8KZ+wKlIEYSsfbzde8GhrdYk30QV3djZnshd3OaH9OBdgFieUr3pOYba/Ek2FfvLwmep
eaER4QiBpIPTaTNd3qgM0ByZztseERnN9tAy5ofxpjOVJtu8G3cIn4Gkkl4W6UictAWPLiLz2j/Q
vWZu29WQSRodNz69VcB0WUZqKuX/QgiIKpF0hOmmYZm8bI2AFXPVFiTYVpeWUTDWWYTZ33uB2P8w
8N5mIn2U+nPbMJ5W8yMC1gr15QJq0g4+X07FvhbsdbEGFYz7BtGZ5e4gRxgAcoRNxFGCs5yLBWle
TDn2IOmrOk+zFmdQ9NhHVTQu1niqeXAmJC8tLBFBUhRrhg8X6fIrZvXyzrqVTZT9K9i0QYBFZfYw
5bbPVrTvWFbvcYhkkIGEJNmeH/pFcX0UnrEhPd9VcxmN0JyJ7J3opNeD04GK8fDWF73MtZXJJf+z
cwPWSjAi0xopBHkmYU2GKPISyiQNuz9uzh7xXpuYRsG4QnHn5TCl04766tfRwn52vI6rzE4JBMau
WKJhYvUwMwkiQrhV9sgldn149wqFHG2boLcG+f1P+13nMA48GJWCIawQtFuAQou8rimmZwLJOrwv
6JOzSEZQbQf2vCAGuaG1Taoz/0d4omMsh1ZaJfyUTKySULuH9Wsz1fyd9fXMLJSbnAViv8ksRzQ6
HS8kze9R8vXj+Oi3f44oYy6kqrxQLWJ7WXSNYIFwWrPPLoVIfAi1bIb5VymbvjnFvwtzOkd0QUfx
03SShYLWGGw8Om+B1UaNVVJqsDuvqljdjqcDacZDveZwXgnIP4UrUsZr8pu1CERZUKLZA4WtH1dg
qDw1elrTC+AOUngNE5PjbjMG2oYBg2Hb3nE7n9xFTXKWbrdB1Rtu+RnRvwnFnsrcsQPPyrDeMrOW
o/SB6lYdSD0TqYEAxcnDgGLJ/NLcGG7Rm6wD+l8Rr5C82lNluyMMT20JmvChZmaDVzgw+9i4J0o0
h2IHOR27nlkjtWNML5NUyzaP2VqphvP3LWzjr7I75cRGKcCB0t4gCSulp3MX9h9eR3QTSFIFlUye
x73ylepumbxKwbuqmdOsXu5hsiM9HPL/pMUyTdfUlk2jxcdXmgCNUiFYPSsvoAyNQtFLT/FOQ4bE
sHWkyRT5q10mphZchge6sQW5xtzSKUdg8S0Om0cuLhq0iBNegvFszss5Wi6JblLyMN2BMFgBCuim
D1lTbvoLaQqgXHffc2wNvqBOqyntM/923LG/RWzpn1Z/qSCeC/UsQseCWrQtrZ7om67bFGl3mj/f
dAp0uMOXNfWAf3A2drOHQHtSe7TKNX1/5GZsl3nvFnZTkzfay8yw5p1SAqX4gGih4G8wa0bMlaz4
jvZFp9owjDCl5EsNPtgd/OK60PxpIKnNOLkVgdS32nM2OT6ovKYLy5+MAMYbsTbiJX1uGwddgBV+
u2GrIYO0Qefydc3KZhiYjFNO6S5owa8Ay0znhKFS3Yn8xR41WR0LnwHexccGkkilcDvZDLJZcgzR
RONgDuRldKRIkmjG+0dBLkXfWQdIupY+Pj2JCSdK+Beh/Hu51xrvKCHnr4LcPiWeSBRL9S9aK367
ayw6gytYG1IOc2xgd3N/PdhOW/YEeD2D3kS/norK9daTVRjOcznJXeEpeTKJCQBokC8Q8WK2fB7Y
1ph9NGw0ngvsUF3QFrKs1vk9uRY/KMN222eJ1H3i/WzP5hYMfk6NnJrlVOq2Cl1DwbgFXfVm2mnZ
0UDYiut1jMtAlXYGji6BkIOMUE75JQb4FVrVqVaG/iIcjbpUp8X16x9jQceKm53XhsJuXpNM+FaZ
VZprelQzr2sZbKe7w67PCsh/CrhFdexBS55iXUgpJHhRbq2ccf0GL803AU0sza/a29QktKMKWdUc
bkWAPJplX1vawh9JOm2lYb6SijF1pJW8F47mAg5tX8mfDGzL973rsXbIhEEcB5al7QKVSxGbTSfj
PHnD+VPz6iupUhfBaMCfUN9UsCzZjUpquJL2aEQJPmfAwBsPUNPivcu8aQJAEvIoqFBPcdxaqcbn
q0MvcRIwEnG1jSH0LoLj2TVusheuMr5PJMzt0oh8Nabspi70477mpTHxisWPAqC5k5MZCiI/tTH2
e6dIiiocYiUigm/G6CwQ2o0+Zju6NEOPCRCgGnqcdit5w97sdpbZ2nt8Bu18iYqItRRilWoMjEld
XY8hpiof+XCVW7ebPbaV6Sy/e+v1/PhLeSQ6BG+ENu6qboRdEEMINWc4ZxVppSRtARgajSZbgyS/
gJhaPMpfLyHjxMQiHkw3gcTCDUH1+XNyTIIGdd6CUNMUuxzyND1wMkV6aM3D6hwFeoUxny/9sZ+o
4bQUdIUot3CHEKrt9JrN6uZ9D7IPnzj/M9zSNwjuKweUw9kFyIXbEoFG8JIlGGdmxlimW6aa+Lrp
tKDbbTGzdThGl/kqSoKIO93SQwdJ7o9vwB/TB9eVITf9xGlKbrAJ8duPfADElw7ROdbK/Xk56gLV
rX5QtHhEG7fdqL/CXmybxcNHElEA2r1tl2Y8WZYACOGD0KBXpBhdAv7NHdEwsFLE/bHR7mxEmk0G
H9sM95VeZVOqgxLp4i9dj8Ytted/FCRT2Py9jxDqsUhSUToi7LAke8ptpOWW+y33+eqZd5z5Z8c4
5TofMUeDgwOl7p2Oc0SkJaR9lQ9UKikCHDqA50HEsVQmOG4wsBQFzzbEBtRnD/i6Jbn5mlkNT795
rUHclOaoR53WFonLYET94uPuid3jCmnKxJjdH/EghRReyNnOb+OfUpw7TQ2s0Y/vChHax7afJqpO
kabtbVyFKc6g7k3w5cYESK4VsbyP/cFYq86MSwEM50iab/jvP4fHl4TIP441Tlv3uoawuNlkGrZy
Ykn77F0H6s6JxmvmKWlvtN9Arj2tcGR/2O8qM8Gn6p/5dE6resx8I+qkVhOKngvEw5wUAnCTO3re
8JtI/7qsUig8AC8nfxDxGvH5VHGJvam1b8tFRO+yGSYnN0UKop+/B+SXdDFta35Vi9HKw5DSXxgQ
2VU+uU/Bv/f5Y6uu2aC9aJBXI7UQBsdJh4+1Tm093SNxAuyy/SzSZcG6ueHfnysA1a0NgKj7haWk
OCtFriZmGmqCHnMTbGkqg+4gnzaZDRTg/fmNR1PxTyk1D8H0wvDV+OMLF+CbvLxn6XBOfwMgHOU5
MT6hLJwWmAp0F38YW3MGNjt8VdgEBhishYgG8dHU+4hMIHW65BmLZKzBvmooDevu6kW9jvwelvdd
vi3mbfB3qMks/6QIDEH/efbDIw1q7Pl7pNoYAkRPkbJFXn0y6cTPa4YQCBGRlbNX/XPNi1hAznj7
1kTyYvzqdmiaQW58mYN1vo0yYQdwwLQpqA70XexAqHCbwns7CQRUZWhZnEd9DWIFI8D4B43oVdIQ
ujSgIKqeXT0EEvhmjOD8aft7+T7G+Z96SJZVHqw5DF0eA1PH0V9lXyYUW+mgroeaQWmSkxVxq0Go
5IVK6WQ17ss7Wt5JlEa/8l/w7Cai/D1YnsjSeMwqBHBG+p3Bgn/J+O/SHUeTiC/BARwjzhwGCP60
FsZhZayIBQv3sWo5YaVTyBJUCYCjN1AtrW6EFy0NkLLVqx/8mMTW0xv1mNf3lWv6fe7WTFlJpXIt
JLrw8yT9X+jXaksC7JEg+6yIjQr0ljJ2YO4lsgTjUfMqPYlC0OtyAbee7+eEeVlGH8OI84JEYcI+
8Y4sO33jfPPQAnfWk0uauMPcfTOmeF+JkSGm/GMUlANUBhVE79JPvVneRp8k8chYQyg984A/hR4p
EIcEdAV6ywJKormpMTB1WS2W7iPcUjD1fDxTYA5IB//OKhzSzoNI9KT8CUAz/Yekk2/LUKZ4cDLw
wuWRRa4AA1TTmZfe66xodjyXH7ayiXdfxTIDGwb6G/eX66a1Bnew+jtPSwv3ajezWumcax2q56Cb
vlDlQv7AXF7Kn3hxKteln0KvAZoXz7OWL5AdVyAFXUwCKqTWf48MbXy98LnuSSrS0q0LO8sbC3TZ
Z38kemjjW5+T+k8Hw2rffyh89mXSlWC8HM3WC2J3Yh6wgSS/EflbizmjhRyIdHZmuxv5O0jl3Sq/
6YA7q0cT8yL99o9gx6pBebLpVY/scA/F78YnE5STo8wg9cRJfoebotWCP9yJVzbC0V+pWt/hZXUU
vkjuFdrBJ4jbS7TYdmm6ybTvYbejNDLica+GDRZyF9CrCJV3rQ8rJX7EkDMiVrEGG1wmyUNE5XQM
bPWAGrqMKmucufqvpoiwmxLInUCBjasAG4VP95DkF/xCPL6j4lkSl+nx4uiH3SbMrdlOqJZ9bVeW
NpVYIN+K2xojUZbcUR+Ri/eyzcg4CVv7+BCzPAOv4ByLfz7hFPsVElk9KilYUyL+EaKM2kBFy2M1
T+FlFiGWV9LHv2sbqXY1f5BGydi4fLoWUXjiKc9XNMcAYnsTJRc8UUbA1nqBXifUkP5OBXgQHkCi
8eqc3O2MWBcY8x9VEQ2x3sfYT8q2K2kfygBrMYtJFOatNOGOP2TZnLpDFgnnNK7vJBC09+OZzA8S
BDlAP6xaf6ThlDN7rX3JS3ckUaI0mr6UcRUGADvzK6UYt+DjE1yfocS8GY6hQWU0pXRn2DD5voqS
licWJK5IN3ZY12FHUhhEILpQznrHdL91YUVU7hYwmssV9YKOq7QCKbroDQa0qqpjYhnkU7JYOEwL
K5HI46cgruEo3q+XyG0ugd0XxVugLbFpstsR1/1CRht5Nn1OAp7caCJhUrJHnAt70E0VXTZ34rMR
Xfg7V2HhwALfu9clUp2MazEvXf0oDPrBs7zswdgnkaoVO3OLYZ7Z2Xak5TfYwMrzewR9bvWXSBhv
lKCYFXvE0mSfsxbaxUmKzC/NFtfsjyYFKI5hBYb+1hLqM4fc0E3lDQFR6JK8Ps5RIadHRHYx7jek
qdbLBn/rl7wXNFPTzPuBvo78BaCchiyH5Z6+HYbL0lFxrRSqIxFOYy0AM6LNvdStFw06YZT+YmUq
evEoNB/Vbp1dTbxKoKo6IjlHzLa5X0Xf487f0a847i6tyatG1A8hI44AA9bE/5RWX79/ToETLDv+
4xAgSsOkzwN33qzhJ9yqDNBtbk9nP4xrqW5/A+nEB7nqu6ctoh8sO7VMsp0YXoOIrA6jk7NdrZpP
dZPK3TAr2LNiOT5yx0iwTrOiGZMS8J5Z+9Up8rKkYt1R5VwAAu23XQGON54LrjtTzv4wgnGn3b1Q
fxzQeumSDdR3bSybmEPzG59hw9ovC88o5JXL+7YOmhTYVsqnSFeGap9+t3zpTuqK2tzKo1j3Ju4S
595VKDnRvD0nGiuanCFoXEfK2aAWuO5zXwvjTGtQcQzSi+TDd3oYJh1QnIyA8h/ZTIFnYfKf8gZ8
iRuqu4bzcebC5fNrNlR+Y8yYXWa4K0RTFZ+s78G0ie7QsbOxEZI8rdkTdg52x60LkLxHG99oNcXt
IZL+Nh2lxhNdTkTrkOVntFXAz37Y9lbtpg0tpRW5tYeMBW0LMrzKx1hPm2ckzBdWMpdSD3l7Pezc
hDD0OT9SOJR6IoZLIga59NJQJlMl2h5SQ+x0JOCd04o0LGqNiU+qsEJVdPbRabzw7xxJa4InCft5
HvdZasP0XSlQkJC1uI+l0QJG7SKKD45GIR7aeATPrfAITSxC8qdzLQFATKHGiBPeNXp4rzwvttdU
apqnGqDk27BRVn6eJKk2OsfL2YqR6FWlj+vGjlY8KStG3WD6k464EyuQYx6MJpGqOtYKGqE2Rs1Y
OwVspa7WZxwXNlaczXA1tkIErt3nQJFg0pbP2s+lQ67s3k4RhaJPXGzbtG847jcMs3/mlQpajJog
Zi54HRD/5FDKptgoK4MTJni89FmU6VSyR88xvTwTM4AaDJPuH5Sv5SvbJZnBqGwBKGT0CJwmsIq4
lOBldt3ttDsmzDDpBSn+YVRD/J4X8RUGHksNH4RPXMU4lc8qo1DfAxTzZrZ0GLmZKnok0DetpkSU
YckEgxr0KAxMki1rKitmNNY6n04GjflglU6PydLtXDuslAfM8vuXZimNLnbC48J9rcDDRn6ulipU
gUWwCVSuYeWW81nJT4qTAeYpp3aKV+647bd6Pnw1z3y+1EXQ2s09P01aqCFRtdSsTvkpuEDoucWP
TIzmjIT3aGkRSGFQnkFDUNLab5UCLGn64y8YNc3g/cfF3W1syt+NBJtaRULDDIkDN8PN5MXSfhk7
XY/EpYeYxAej/L2YUtwvBQAYkI/qP6s7xa71U8PfNHjDCWC94k4ERtSccNkFyTLcXutKPmvBhahY
dQdQd64cD9sQqHPDgNtSeS8A125ThyfTrzDQalgbw0QzbsESJx5HF868ZSGioW8FXjvfeZJefQTl
D8hWRZEZI1EKYrIb3q7kJKNWcs5fOlBTXdY0lCpel74iYhCqr/k2oFm9EIRyl1hCa+O6hC6Y4HiM
2DjWWXdDrDz7yJ/EUUHvOehSY0yDp/XhpjSCdjREU0sj8/oB7R6oln7RiMip9KdVLbaE1tGAoxJE
rvoNCMEVswt75BUeL3z1tk+EIzVlBbBMyXuCnxrBM7aXmoXIA2Wf0DWoCA4P1dLbmEio/cARgX54
xZecAL7GSWIfPrspknuz04R2o1RUriWli0FLRv1f4JJtpKOfAEOHadgrpWZwYYc3xJXIbfyTX9G2
c3U/Ymg2bI+sf84iYoslnF+R9VVcMDL502cfhEReKXuc8pwNHYGEzJ3Y2ur20w5EDutlL40zUu0j
AoWC84VzxieEbE4hqjehLCNZ3LEzAmk/iLWExm7jET2hYHo49akWd+bwc10iCXIw6S4rA2rCoQTr
bTgtLOCt1iJi//+P+JpFWEFHTiY5JLaI5cLEYdHoPYIlnxsh3ylVDRvbkJm0WB/57bMIRStZHEzc
awbX9j4irEHTVxZdsqD2ot5Fs8cnYLNrmfgzpbHcd8OoHTtjsaokzVxqD+1IQuFL6e+BSJyZCa3g
1rnMHjeH0+1Pc1pvky2BLQbFNC+yShxzb/6CwXk6DxikedfNLFuZjydGMCxVHalc1rn/8Gwyfi0V
NdttS4jtCT5KOKGRzCVERogsFNFv0bJb/xCydkt4ccTo4CeQvDVi4nhQzvsb61JszxapWMDMY36+
MImVnnKUEjU9iC3Fsgzl9YutPnc/QJq5d2bCJXtYS8cXYDvv3ntPDl1fTmn77MQQJHkKs7zZMPTu
2np1+hbJxkzgz2AmAKfKPUq8k9Fp3fvoHrpinZ86nFmac8KUtYh8aK/1m3nFslFG3SJzlnwDdkzv
i4D/Z3Sgfz3SuuW4UrBfgJZ1yISV3PdA7Bsuu9Po4YrMjh2qnx5HfkP2e8tlCBNH+S18ME0EV8cD
WXWWa421D+rXqrEgH47ipo4X3uqJKOmTbX1E6XP5gOUuLhic18xoVB6fKG/OfjgFZDRQX37B+SZ7
w1xkLF6Xdv0wrTxnmHC4fVwAHjcB13uXRG/il/tzHIRrLR2NpzwTKwwwD25ihNUSjbVCG8guN9UU
+C7NAbGtBORETIE/fIVPNpaNvNJ5orpZDvc6fdg/gMMcfuf4crEj6IQIpuLoLiQbK2MU1tKVSpAX
jh/O9qSgb5xnPofrYF3z1V4IJ326fxYmvSCijPGwClMALGwaieUDTo5IAMyO7jW/Pni6KSfaGZjj
Aq6CwjXVx586uD6sSbYIZ39P6pVEMPw+anWqBOZy0Fpio5EcQ52cilyvj6iFqfE2Q49gn/CQnh6l
PTs8Y5sBnIw6e84QsJ5cveqlp4oK7C+N1YcpFlsYjc8T2KFwsa0MqVrxNKwTalV2sJVvgys95bqk
GsfP+JFb6BapkJrLA+h4WqDvMpItMg1IL2oGmyNjeTPDvTTfH3kQcVC/3Q2LIaJpFIFbjxii9F4V
M2+RRUMo8+nHExcV3k51O9omrU+8FeYeKDt3SQ9lORjCywkTueP6pTB0ykCML+Uj5VI1G17UDABv
EoI5LfdYOD/IiBNMFE6V58+yUH08K5DcMwu/W5GiiA7OeNKhHwVq/rvhs5+ae/FEGlGQY8Cg6LrE
w2GUATCnIwaVZJWj81/F1p/yDRmT41klaUuUu1EJ+BX9tsGxZiec0UzZLxjco0O1w/Tt+moThaib
ODXsuCDOAARL2e/MzrQgKjQwIW1BgNIR2I8cIr2n8uNGYuZgsOyFv99hjYlUoSXgJITofp40sOa5
1uE9YWPvFiLYhELfgZLAQNBY+5tFUpolNAqoVVLMbylNam5szzJxTk46jj6q0CbweOjDxEn7g30i
jIxUCIAP3OsMt92SfB34uKTKuR7/r7F8AVE/KsOGFv1ZuGgaXJgnhPrvf7FMqUXEbMXQWahLTodd
aAqk1TjFhD7wwbs5QKOf8fR66u+rcOSweH1cYeUHKnrpyaQQqAT6uR+Dn3JMkJ8TeUZS3K/EGswd
qH6gSrhvVz9SjyrRCDcFybCHEvgP0PjlaXpuhIJcS8uSgdeAHzTlIOjuqIioUfhvvYfw8T9QOTNR
NMdsDcLjgUZ+t8NwioZVz3KZ43KZcpL3+7dp0stuKJqoILUhdvxDwWjOeU1nFl4q0QEaWDZ6uYBW
dQwkp+TQqhHfFl+Ly7FDitZ9XXJM0F59HMRgxWt/0XBXW8MQ1KZOUfV1ygei3njkImf6cJ3h8iyY
O0RvBsRcR+Z8ZVYEVVCZT7s20qFB5NbjBameGn9t3kxwIRTOKivdpS6at7u21bLCUJpOODxWv8QD
l8S3XWThRy5RzVanQiKewHLD4vvxygIfIdpBQN9Z+x/WlgAqR7zlHn5C9d2opYT/2y+fWUv5uc9f
SADho4TpnoOuZOzxuJy4dL4tGoC0wLusuwQXDOpk9BbtVKVkLmamRTkEgykwyTF+wdumWaoc400+
pdh9cSTxPdoG6byEMasw/019aZbaR2gl3TIVD3d/UWxpH9GxlUxmSfogN0sWQKb1ju0Tnu4BlY1n
rnDIpuNneawK8NtEiroka83oodWd2xwlltqlK+9XjdxXWpkqo26VRtpu+6gj6y7av/5XLhSZdfBy
MD+V5MlN8lS2BVQ/KfOb+6RIW6AnM2macu8/TWq8o5B0rq98KZ1wCSekq2duJrYBk0K2IuS9kIXN
Nkgnt94OmChAZSujlygosP4cbYjUldVyakjgD5QrcjdSeT/8z8bFf1/in7SVvO8xJW/UHwWlCmbW
ubinHha1NG/tHt3ruZolj++/wJ3jjr/a1mtAlyNz4mesdhyP6t4hLC/iqsH+Mmzd9hZBoF4QIpqt
T7Oo+omMr6b7b3F00n/spvbVuYfnS5z/zPWNbVVgAWbRh5befMKktIgD4PYbjWFb5/8/Pppgi0KU
iofujX9ZTWipiAzHuGOjo0mCTY5iJ1gxESppAO3dt8zSUqcJmPy6dssCOffz5mbOMnID4gnUY6FI
M2aOMt1Tq1UAbmUHwfTnUBg+7K5Rn/GmH6LzNfh1duWIwioKb/FEeynetY2+lDfWbvdKKKJxdJZP
n7tgoPKjvG9HDkgWUAS5pCnvtif9CfbhB1QCCv0bnie4QQB1Xp7lAjGWnU4hM+pp1JxlqkPi8iIO
Ni8RPVhiP3NgSvrx09Z8WLGo9FgoeAEw/ev6s121FI+4CpHVKiY0upbOBP9vXdFNUjB1pNdCFqCJ
LsSt3+ME1F/0ni5z8K0XskZHmE5udruVARVPcmsRDRrXsyEmlhkWm8NloEAXmHXc7Hts2bVJ1EJz
KbENRkE9MgTJY5R0zYlt9p9cIX4e0+A79m2Q6XrRnFbbEAbM+vHaa2WQdpnWQB8pmQsNVt3cC+Yi
bjGjy8vM8JO1aHIPbHyRTrSehjXzEfzeDckTLSVNne1iEz84WVCLhWgTCpleZmE5Mw6WWL01xV93
iRxTjOFPC50g0hRNQOreh8TmYNcwmzsQB/h/evem9VyEsMIvoyfRs2/makDsXbkbo9/lnmVsxcpP
SrJnDByREngwd6lhBKyJvf3lp4wlniR3HmLLdIw+f2ZvPt709d5ElF/kjyZYDbnkAqnJy60ndevQ
wtr7tkpuxBzhz6Nr+hFYDhJntnlOftkIpE46nCsmSbngvT9FeGYvFgxOjjbkE54YvAH7RLwUFiDj
yHhnxzG8DFLTq0rMPDoMiIFxmb5NhArEOXkK04tz0GRssFeqhNhCXQdIHP6Y9TV3n5tBLvilY+su
oTFC1dpJ71HNp5H7enDPRKYL+NnPf/IuqWj72M/LyUBZrpndJQF1T5M3iIBa5N5s+I0DpBkQSX21
zwD4okt11OpFVrqXPDItmzvyxpYikH7RiMc8fDRuTj59CuZBJpkVmQ1N3/unNULjO+7C+PLQ+wvD
Q3xxvXon6VOB8TEwIbhsGVqkBke0md+JgMtB7sEG+RFb4mPz+ImyjZNFm3vSmSPrLNuDFeAkNAcS
VZzAp/sgIwZock7fFXuh/LWP1qkIL8qmzSbSy18GNH1fS7MG/F/zMbivzi112t0Luy87OjaVIWfV
J1JPeeROoq6JiLkITIm3JxjnNiFPrV4ZbFEleverQVafXqURuRYswqW87EDfp8ZkZet3UMTIw8aR
kKl5Era5Uqg5ygsRaHcrmoZQyZMrNqWnprR0gsuGesToNDgLXTtnOxZoCjy7guqyKmVTBmg7Btwz
eTM/9jOMGkND0y2S5jkvu4hcRYlTlqWqRysdYr2Gm4LeBbm4Fdg7yVUAjJ3nhSyWTyEaWtmwPsZe
r414QztobDLMeGbMy7dhmS615zwE0oc7xzlwQHQ7b9hSTxz+4CD2BZExATbdyNwde7g+CDMa1s3n
wnp9OOCAExQZz0bZtMNuQCVFDVIcRbMb3qXq6Cp//RT2jVDRZ1srGCplVmChTVDvWlvF/16DDh/f
9ZBEd+ObEvfWjiD2DB8akUxKCa8C6PnbWI6HJsBhW+jT+RnHn44321J5wdkKxQJzxZVcg7Bde3LR
9InUf56Uv26Avnm3R/oZD0lsiPLSgoImCSa4r1yNQ+RyIZ9eBAgfTZScWhmA2O9q4+FqDCiP/d7F
mPYO182Qdyu7mN+GXNPj+VUIP0SgCqZmoQh6MNrKizNdcYA0FzZN9GR0iV6OlKO1k0iaDNXn/ipc
vwdUIxBYSsojEiLBdg72Q2RypZmb9PHlnVFkbWVjDdkGmnRxbSOw7o/kx10Wv6Fny1ATNYxs9NMC
SBwjcPe9CPm4FrdJ9ce4WWeHAqddIrUtgHDZFtm8Si7+bkxnDC6W0S02vk2ovbQOe9Qn2j55sHwX
lNB1L88vE+zUzDSaT++W6CTNCSweX8ngQ4Up6iQMgJDbEFPfFCVnGl0W1R7eSvM5bfHBgxdDU0Cz
fepSW2YMnhbohghCi7xENyfjeYAaImFRk+af/GMDnmYWezc20q7jlPzME/eDkNSA0lyha3BKMIb8
np3rNXGvWRWpz47EaYJB5ZAksNiYUnTglcbeHOQGhlmNt/bJGYpGl1FQ8dKsryOFCHEma5PskFv6
2oed7iGZ8UFniD9oVsUTRrIo+fl/9v7gh8/SaMkhPn0WEVnYAjhy7JqYXuPIUgWMmDDDc+rQW1fR
amK0k1N1jU1zcHrdVrVKvPYdbesOkveOCtK2DOVit+hKFN+ntozjQIWcQsy8Q2eXUkN0t8ebcX56
i5+FztC8/5DizIBDbUnNCngjUrD502dj34/oDs84qERoBlKIDnwojnoI/ftJQCpNXvOZq0B2pa27
SRs8U4SLDJ1iN8qofHRgEw9tLRrSFsGxeE8nWOyMzzhOYGjTPDGlZbz02JWtJJzWi/m/2h+C7ioN
gwY0fWPYfN/8hxLgvq8YvfY6wpCKyGaYVnQx8AXAqe/E5256cTr4kvQrRp0fcbnCTMlmaphuQ5wG
qpeQRR02NErIjrXxZk8A6Q9HBZfAhC4yLqTKhhnPi3LaKmE7/zQb1yGl3O0ITVnir9puBYqyhWuY
Uvp6FcmAlgwKbDSxySfqsTm8EfPwT8Ai/0yaUeNDZuSVVOIVQm3R9OqX9WSxlGnx4TtwjaWCg3jD
ZepCUMHVYFqYOWbxn/P1towXP2H55wlASDEm2VK5bLiQZVHxILmdpXtKH+CJMwnYi9oXnWGUzLQa
yS6vtGnXQlWGzHqT0DKPFG2QkCa8o2NQbQktO0iB6yPnV1M8ToA6S97JP8N1ya0uq9dING6oALmY
NiWfiGtA8coQsk8gDNPOQoKyyPnsl5PSQdELlYUPuv5zGwoCL8QB5wwwQO7RzV2VJt0hN4L4Yjka
ngbkNeAwNpxIbDlLurgoh2PZeBunyAMqTrwdTnpyuwdiUSu0PBDR+6f/i3Z1f7/BYVNcobciHY10
+/oVDlImL0QjM0e9nLSVF1/LbibkQX2ufrynIPz2ZR0IZ5pQPkSpRbZGnlgLpKYMq0hOrl7Soe6H
KgIjm9rE9BR3Fi5YoUmZ8n8FS0g9tWBrvrC5q8cbU5Q/G/JwaC/SQkJ+eZosQ36DA9Vr1FN968pd
TJ3ouM3Kdk626BZUkEArCjOi7o30VBiF5TW1k/gWUw1SYWdc6Dxsd1tzdkEmIEy2dn0qc6QUDzhw
BKm4UtQvd6sm4fXuh79/yfxGfiYQHplqPsog0ZaoEGY2tkfdX5qldqJvakd63T3K7J5O9HsNU2g0
df9WbfDIjMXBUPk52qkGQBdD8jfbv/Y12bRiZPCUMwJ8BdDdioMyFM7DFx/vZdWtShCAhZFkoyiK
WeU3jwwHc20Ydreb3E1MkmzywSK3iXX6Zzvgmu1yiXpNB3sbuPj9KJ5eKCJGkEpH7gKRKZQ2FpvC
bYtQ1Wuk00IR1MfzDyYP0YhBfz4xTza3bImYvq/+pKoCWq8I40bpAziLZpcyWXnbOP2U0fQDtj4D
ttUaULpKOwopDhtc30ef0//wf5FBn9dI3NKkm5TqK3poq7f83MRcBgOe8Ryl8D/KN+ZzIMQEFsxY
yAIt0A2BiynX8BjFaqo49pFYStrRQkkWqxKm2sS2Gi5OtW7mrUc4RbnddjvCve8GUT/d8o2eKEIL
T1TgbwBxU9EbFoo6v4z1W0Gabb8PLuQVaO1KeDc379xHm8HWVndM59EoO+1S1JoxISnIAUTRPVkZ
up41dNaKHyF2CWaGBitey6q9SlFwkxoC86D4m3pDfbtRylqmJev7kF6v17ds7JIx49rg4TilRyY9
/k8bUluUTM+lRew/nk1edoCYyK9glxDxxbbJ5GewjdcYFoYwmoP2rmvViabJuUxepzz8vpXRf8CO
lMVMwi+ZkR3HT3/p8SS7MOxidqVkYoicUskA3ZqwfevZl1P9g7/GuHWBimXr7mOHRW8EfIpJoS4N
QSKlVajRRLZ7J1t9jLGjmATq5fgtsxsSmjZlbZutq3BOi1CFRS1/KbT2sjtdOFq11RW/zgIR5QXG
EwHaF04Emr+lYlwVe9zeUKOseU35bqQn1Ca3WmpvmtgH3xPCUlV4vaJ+nx+ZXA7TjbtiAfZBONv0
DZPC5w+K1SEwadQbLXrFpITw9axM3vZe7zuvtuRKk2iGYFTLR8rvXbQz25zaXsszwC6j7U0iqdUA
i0Y89bI92TuUuwsj6XYEDratRxRIc1fW+Ihfn4eAlKt0tNvxvLr/zFfkPnfxg758NijI/jJ1AFdp
5xeoPcZKqOspkoUFTGbRyzuMOC2Nl3mBA3590mUCwegNnQSAaZwW8AjHVyOI0ngjukyfHI5xHZei
stPh72dfk3TJTXPP3Qnr0jEgXJaNw5HNCo0ZXP/IjqDTz8yd9cdHOcU9WUBE19mkJFrY5qkkTnpO
nTipZKggfY7ivhqTEXLDBf+pGWrUbwOG5yJbgKB2BbbOJtvO6PFBf4MM3W31IoaGDBp5DDEyQyJ1
X/+wN/yIT2ggzpYhoJWTHiiYmMiUnbuFa/4VIVbyp8LXGrn7ddHuJ7m9/GT59ZYMRieCyzgRAHhs
y9sbvYWrZX9fSzq7xoWOx6MHpp1T+Or0oDd+ad3LEbZ7LiKNLbBt+nBY1FQ1jFge3rCKAkr/U0AH
bQRG46s7WhB3KnX3KZskoiZKCo1K9iF+kh3hmlyyuVdFmBsTR9DoJJD2kT+XLtu/2yc/OZkQJpJt
OOOEuvAh//lKEH/alngrham4RIXVx99j6NHNEs42vSPyVToXGeovTrjfEdK+aifyQW6CxI5rJUlH
g4HdB74EeMHTFEkM01GcLmdu4XN9M2MQ2K2iOd/KyQJdJhzKmu+vup9k6+YXbnfJpDR1PYZXCeBQ
qJDSWmntUdBpBDlMd4dTbdyHazLv4+SFERR3g6vVnw7ZcEz2zfrzgHCnZ9ZXri2gz3OvI6rUWafS
VW06S6w8qNPWRLH6ZQWXE6mskGCtHapA1FlF1bPiThJyKcewKE1ruBzkBZj6MRkH62BkKtiz0Xro
f+m62FVOZRmDKTB7Ky/eFoAej1/lLiiUgsQW2gJUZKvkasKnAIIxDgCiEVlWmj5qJhWRavxyRepn
c5S1ZPf1Kpfu69lQOEN7lnVrc9sVW/ivjpkodxXlmtCuao+cZJSusegDjIGS9tvOOkTGhYukuAwH
6pnbbnvMCAGh0SdAbAdtvx/V5UgqFnrEW5Tqq0494bSx6FLnLiB6TvdOTWEVv+EDDebS5y/E1tGs
qD6jhR22ygkwrXZAvTsCLkjEQXQf2vynjVb0LO4f+7pttfmLt4HBUUN8pv5JfARshaCZu6iKS+qV
UicGnLsWLDfCV/p7qA9eHQnYTTUrmkEfllRUsWlnDecrKDCEYrd7/5l7udhjvSdxUoBiAn41/s0i
Z+qpRwA3peduqgoPFg9DP9MHgdMkBXdcbmza0wIlTRsWbNPnPptW2o+vFXxATufJvEQC1SN1sguB
ROIZ0JgPNnUG3QwTlRo9/b4m1u/hERFwEQgLAooDA0sZ0MDDv/vhRfp0J2K2aFvGnDnnsZKVQh8y
AiMmTjcRSujZYIq08WDmHl0Id+gg0/H5cTB1ZagEH6UkG1ZJNekchriRcc6ycaUgUFX4nkL/qGQG
zE8Bg7J4kDPLRw1296RdaHNBq+wDr76OrTFh0c71jhEV0XbNTvbeWt+JE12fmZJtluMXnI+RSwyC
eK0Qfm1HsIXmN/RfDlfVq2lp3tbU54Prj2pnP6XqnjnbnbYghUpx8jS63uDaEcJ5soYy8UlY+knw
TnjuhFGUzdG54pBBGTNrzV6A4PRgpkCndJIc34fvgx6WbIwxpX7GWXzKolw9bRcdlLScjkB4GjAA
hzeQwddpsguNPjBUDc9VimI/4chSzNMp19+EdjVU8+Lvbb7PS8UiAbYbHP107n/pLlEm6buzaAww
UhMnm8u3fK9Z6opyeLa4lr6mnwPPrDPcgf8+vT2DL5Bcaxeptb4mGN6YZCj+U1ND1Cc11i0vOIVX
xgFwlGjTFHzbxxQ/cbB6CxNOWUCg2JspbjAH55P8tlGOvwwYKBcTwsswD40EEWR4xNf2ZKqxlpTC
EDy8S+6MMEPPAV7mrCbcfHYhNnq3iSL0tiB8SMFkkQX/Uxb29M4wVDG/ud89u77MYgSkKTLukIoi
k5w1LmnTzn+U2YCDCPAB+QNOWV3HD/5AhkQJwATuYMC8bOcXZsOFcBJD2O+LxN3xDCr/8969uszw
FyeHeabY+mngiDFHNfF0GKmWhnM2GEbyhP9xQ22iLgUN8/NCkYKZQeY3a48DYe+sXabXBMALPk7C
K6a3gjhTnQxG3E/5BUYI5i0lvdtfKdxCpXPCBqRkyHVV3riTu6zdwIu1NP3ICWtYDyWa5zH47kc1
rTHYGcsu4mrFRiJngZ0/oEJsN9L7FFDr45GOIFjMB7CChJG7oh83g6l9ILMiEJjg7hhl16DLzBDo
m5ZAGcl6//k8Gbbl9I6s6tg6CqE0uhmJhCkPxBxcGA5DvGT4w7ay51w/loYnwk1XfhxD9Z7zPg4+
Lw12e3BE+0Rl9isjsSMSB7pf4WZECwdecW2lz8h4cgSaMS4euZQ57hDq/r8b0lPwGrKahv4RIgyG
8/smCcUhRe4KvEIiMT/elH93b46iqINKrn7NJ9h0EwXul8c3sjrqJtu0zXbPtYYHP4RGY1YmhX5W
p1v1ZdJ9lnpfI3RqzLBCM9tT2AIhjKzd0ha2hm5uQyI23ngio95pe+0zozB9z0UDAZRH4xaFHmAs
HsbwicB6WcgX57AxfJgWNHkW1G941yKyxUvFwHiMj5QRCG0jPjl5ehXVFxBLz65b/OrhE/hbXChP
J0ZbWyqyl8PC3rbLC6vj9xXb+Pwsh4bsnLwzU8CYWGF3aw2p8woDniadhBv/TYQrF0/TxTlvB7J/
fZu9ALGhx1cNGbwhsv3dYoKkS83nWPilTH2MzY0/GWgBmcDPR0kwE34evN4GsSnurqRzFdjb0Oxk
ZCImOP6uCMTfWCPUc4Tvcdp+VWesxInsb1wK7JWzUvEWA5WrK7SYQnodQGyqywzsSgbtGMlLb3IQ
AA0deO8MUUGRHwy49C1rqTiKxPKjivTvgnqQZJlAusUQpEia7sQil1dyfPy781H1HaXMKQPEvx7x
ZN9FgQWg08T6xFFBiIjyJEJpBkaWZA0Q0uhSFjEDznA9PayV2u+RihHba1Z3NswCdFu8EW/0rdYi
5I9zLbM0outuACoEyDrl7f7GY4pWWp8L0VfHka2uT5PS1T5DPbNpCiQLKa+TUZ8mLMz0kOH59xik
Xm/ONkx/6KmCC6+otAeq9NSsadnoAHeewq1xwtAfFxQ5AXEhzSVeLY//VdTtuOm3rZ6IwyblQQL5
E9WOszI98KsubAUqVQ6lTocpdEuzk9HmlNigUJXQXspmHwSBsuHnLc9hj6Hk9aDn8KbxOpUtAAvn
6lZj3m5ol/oyXs7bJCikLNBgeKXM6OZIAmH4i7FTJ4tvNFwove2fCX5EVF4ZRuZEdxX3Mb/G/SgE
Njvcs1YEDox6zIve0mwxmsLff2ujrOvWzjw43Rnn0N1PZ4pNGLRfy1yb56hz5nI6q9ZuQR3O0n4o
s6ADNZPNWllYQm2jYLAD671XCVBMZ80ghNDhDomVDwFHUFvsAuXl63V4e9MZFOO+/gXYaxFAYiti
hN4GA58l5TPEEu5PrTyt0vOJ62QUknirlS/Lbd7rwDLwahQ8U2RidsbNIoP4Gh1exoz46KhRiBUg
Anbhjoo3FckQ8cX3St7WERWnqVO9VZHGSoC8isZxcJS7v7vlGJ7ouALfTnIuzfOm+AztfvNm0/DP
c3kgiirRDshNSnRhlx67qQYqwUv+5d5MNlsjb/8Yx6frlHf+AUswbsX8mohjaaHAFgyQ0vHIaArr
7yMRe5N1pbSbNmCWxQ1aInbq5VqHPxI7J9RAAdiXU5BivygWhVB9iTkssOooi45qfk9lZitQz3cd
ioBpKy/MhR330SpuqTnr+vmYI2AU3mSWNOPPL9FRieQFDw+UkpbqD9CpXGWcQ9seFzFMRoeHuvhZ
bEjqCPsUW61uqrxf9aQlD02USjSqFK1OWGFyJgdOpHgZVCD0Vw5EpwN0E3IYK54vuUJRdDti2kTU
biNiZtKv3xsDyhs938Fomt85b3pTrMMA0fvr7RPV1+1yGgbRYDioQaF00e1Qmrz/aJYPCvOLXYEw
iv9pm5OlZHLZsPUgbMua19T7W6B8vx7EThsUr+AFUCkZreT5i24pjphPgmfyCNXQmIhdFZ3DKG9w
5VtcXc3jlhiGVh1w4zomOflBA4RRmwkv0r1D0MW03wC7VdhW2GhRdpwTiv49Q+eYn9ZShrRg11pj
BShxe9EvSpp6SCqhBIQsVVftQk1C1EG1Au995Kgt1Zxv4S1hJ78fMpfN+BFinNL+0t/jlS3Tz5/b
pzc9AG90B90yQsqKPsXutJGzZ8Pc3gqXSAJP8AJEtVOqT4VOfXIsga0Qw0v04DR9DDvJXyuAd9Yx
ZMCvzht/CNiMoVoR6o4lffcWSdcc0EOg1Q4v9d6On83CXTpuazkbVyYvEi/Wg8287bYUDBb4Q/hF
x5LqO7iCSHuEIFjYZEdBvXajNKDnPygTdSuXYb8oKlO8hW6k5AFVbqWZpWwV7CAOLP1JTyitTbbb
3tDVCc4MhYKTotVf60tgq9eNCjD1AxwMb7Lke14nDNt3ONr50Oa+OKPzHCTS2/hYzSuQXxay6sOP
vn4eyPiiit8ezAODaVPXsNH8jxoajvbuqXTunicrkanx6PY/rvdT7eyCEXolsbusppMgEMKSYQq5
3gkPRBy5aqNgdfX0Cg7iXJuNB9/FBQg9XJkL8yrnd/V0jJsfSaoJlInVyMo9y1s7V0psfAzp7uwQ
H9vMM6qKkkVPOBbeYapSsMRz6ECnne3xqT5I3/Z4pcNAsXOZ8o0b+HH9JrxxfqQAqv7v1oFuJmLf
6jFSSpD0BeR9pgwAqSSZCcLk/9TXcC9b4EqKftMYjtyF7bqR3rVxrP2ep9j96tyvLHaZPWRcyP7F
SCEPn1OiLcaike9Y/J/ojfT9Y0pkLJW18ghgwXG1hPMD+sA4pKMe/V1SmYTlLuDLaLmWN5GheE4j
wzCBAyAnfHD0hTbwMoYip2luPKp0M4NMswQ4KgXE7zg80WM/hVBmk3qDcVp1f8CKGywqKlAyTFsq
l4ltUKjnpSs2/51nGyk4EPnz4luZKwGLa65AHa8K8W0j+b6zuyxRYkmyxuc1rQBpUqzTxLSUTynV
GG8slcrafGa6PBQBCDrxc1BAsSjrLtZyOGPSKQDzt6WUsTBYSxemLNvp4fOgf0I9QpogzJsJApax
vmKQEUQMIkpSonCSdZczIFkIRPslg8rRO19PHfEf4ULvrxne9WMiADDUBjluO+KM0ozYUNRZGS8x
iEUiWIJuZ3fB5rItTlqtmLFS2gfnztG6CkbeLoPP3iMtLL5u2xGv3MK6RNxQVtL0b7zosVNBy1U/
NJFp1WivVi+OkfNR5R1hKp7fcF27fWm60JM3kjHk7LClTzongQT+PEoEuUANt19X18Qotxak5cHF
0iGx9hMbjfAi+W0RS/w6VtDjLlN1rrjtSjrqQ8KIiBTwmAwyD7L7alXo3yw07U7p3nEqO+bTDJ06
DI1/C4lsyk3W8RlT+vygDOvFamznyMqoR1DE+K0inacx/4G3VFLSQ6cHF8bL15K0+dVTHUCozTru
70WOh4R1TsZWs9kQQzU3GWAArfA32I88fxtVWDcsr0RqAA05u+Ig2VWPU6M1XBS7kL9pfkeGdWJX
6tJplD1dQ/rfiy/yPh5RdLDb8R7e8K3temcuUVWiQNwxqFscZBYM/WZB93L+NcxPoUehXTc1otwh
dVux925wgUBBTeYUPxeIeanATCnN5N9bUau/rFpO7SA/Kq74gWfhddm7XSfdulP0GmBxqmUDOH0D
agl/ws3Gib6BTheSn0vT5j7x886pEenxwaWTSL84E04ioXpDHTXsn55uoNnQCVQprhFKkm+BotN6
3BTHazhJ4txPOdjk4vqNzUyaojHN8MpQ73ig75hXVmBSyq8IfFjyUpk1G2gTaP4Sa0BKcQkH5Mvv
1M3CKWyWv4F0lx2+dOXdO5myYkX1Q84FRAjV/oFItKcDLvzKDhBXlWBModGr5KlpFxYbQvWMErpl
111hOCR3TUPxYFvTGdOXAfDtToCR+pCl7j61SQegx3v8g91sI+GcQE67LF8ySJVlyuEKuph7vD+w
UyC+wMv+g7O6a9OFFkcylGY0Io4HcsX/TQM6AT4yA3Qgki5Lme5cgER3zKDgYuJbS8YaNYtFEAOD
r5vxA0AmyzwEWM7PoMwMESQ1mJxHRnpElHk4+SOQ/3bgDcajMppaZe44a3yuQQ4LFbJTTOSgBNkK
Zy65tn0hRb3PQ6H4oBGLfui42XwLijcTsm+c3LjRyoVZsAAEaiBqw3zo7WccX0IPDOFrrBmcIDRQ
O0Ir/QSmj27BJPOix5xkGbRQ5Q94pso1e+lR/eoMRe/mvMghPVoz0ZWdHbzFKLnumMbOrBGzwWhO
ApvY80GX0v9TJuOp8cnHZRef45Wslhfu0DJ3ywelqcqt0TtcXYdQdB44St76EsVr4H9ZTBX/GnPj
KxACFX2xUQ/MWIUZ6X4X1I+VbX5+4BJYJgSKygOWQCHkmr5iAU9z4oWe9vWF5WJWkfysSrr98Zxu
ICz0Y9g7dh7m8SL5KBJ7Wt/MOmP+mDSN5uDErm+t3ekpGyFudFWfGpTzELgb63H5zCFeWEOZSNoC
JN4AWfqn1fmpfdEgHmLN5IVC75Z8JPHCED0+0gmLz9eZlwEF6d6V2DdWOdI7ZXDfyCW+6nGPWDjC
JDRfX/XShrFprFdUVs5C4u3CQmrpl+TLj12QRvG3vrD6+ZmoOpQPYGUQQQbAvBClmQv0EdEVQCtB
pxafc/RpRijqcDctFjcDGWCk+C8fjXS9eGvOurLrHRj38b1mD8Ec4eAr5qH16jMPMIEne+wBnAbc
TtfwsPcC4EmpiUIq5R+jbtL+ut0TS/dU7IypJxOVPxDIGZvm2PPvkMnPzrESQoSr9CYOlFS4rfQT
APmLYhm6WCjH0ChU32fN/AlE+jtNDTsMdqiByN3d7bf8q96t8HBBmkGhRHAPFjtae5KVENlD8h9N
bDGwrbHVW1xVtZPhMlWVWbQMKeqWqDRmY6r3qD5fDVQAye3yobbasof1l0QAbW0idXJ+XtCuSven
ukst8ycO83TGZXnRs9MMxupVu4mtelW06E/TyTQe6aWoT9yEDj3XMMwwAwbzOK+8wnJmKQl3to7h
tsBKwEk0XDYiNafaaJsq6+OoACKhdLhgskXf8wCYS+Cgge/snRHbpE/cRsrMQxy+VctCYsAtdHXl
+V18P9qT97VLOhAVzLhfiLjULrIp+LSQjAPig4PYRPX3T6HH0RD7yPF1UQJNzaiekupt6Z3y0CXt
eywxEQZdy+1qJRzblONzylfY/F1Hyi/qh2VqOygjfRTMUj1XU78VbWjdBQPV+DWII127dWmlpZqU
YzIuKSjmMWJmiHetkzSx8/NoyfqFakU8NDr0XbYaJNQWr46qZU1e6ve16whXCmv/cDLVjQSTu4YY
Lz9ecWCzY/vdsQ8GE6/faCk2Pb+Zucle8dOsrIUpFX4TVygbG44hzN2NCsbvcWiKehF34p2ftl2z
W4fq5/5y5zXFYzuTtdHIq5dJl18agR9WHel7uIJHAm/8lOjO9D6sx8RE3AajdZsBw991e3SIXRz1
dj6CSq0gxXydb+5WFi1tUHjHp5Cr8wlLAUb3J/k8MdMMj+sYbu4rZgysLdlu6kNvzOLGmNz2Cq9A
sCOg/C0FCWbIkmBOEymLWsCysqO9EXr+eRWE0C1EWgrd6E/5fphUYUPSZPEolYzcMuvOXS+adME2
9bglInd4qO+ce1H3Rypl5uOFvjwcS7rwZUCeU+XGN4C3xzhluwh0wl3ASyuNt037y8cLiDJWcrCJ
Llk7MVXSiapVloY9DRTzF7/2qI2XrAfzDnKjQwFMFkzhw3npQEkETTv/EPboUZpY1rLWkq3LVoz6
l3f/RFqY5FvXDx1qKVomEdw6o9gVRP716/dufD+Vk/xXJFN5Fw1PQk32ilp0c0wxR6OsoGXoE/E/
ExdoXBGeScAKJl2N8wv3f6SlQ/nvb0sb6rMcLseHtMNVHRurdo/DoYPSSRxT6tF/9AQd11ZIEr3z
tN88FFtZd8qRi+TyHiReoytAUmQH9Q2VKlPtCjAyR2OoU50yPXvxXBA41vSseByc9nisRNCd0o8O
Uy6YowT+yDoWeCehh5pBrYms4IIcNAZXqpGeKbu+TqEYV0dyJq0qD7cC6z+4SqifI71FaHNTeliC
Cp4wu2HLxdi6hiH+5YPOQFBH5TQKsfo5woQqQ7e6NlR9Z9JkLWtlLjE4qT9R6boXx72zDLAEMdbX
b06yyAgb2vaC6Cep6eyf6xQ7R99DK2cm7dpuOQRxCxuLnHC3LI7uNj3fosZXnUk+5d/AnJMt2VtB
9gNbkitATZCUg+H2tG0DBTcJLCdOHkzsvk9LqosSt4b8MdI5qftSNsMw1ZOu/uvbZxV3UKpFxbp3
EqpVMSgP7B1mgaDQUySHTc4ZWsyXUgOwCUd9r39KKEuXOba4WLFeRcsHPUhJq7InPcumxOlAhwV5
SNC92EpT/OjEHr/Vs2lERKL63zZlYoYcs0uU6STa4IU3Ac97k5ch2rCxeQ8kzpn3wJdd+kTZfkvB
b8K0p8dbghtgoay0Yq3jR43b1ottCUrBI9D2gTFrZb4YV+n16sL4XF6E/+DkqyEKxMaLjR30Qjrs
mxg2VAAbQp3L5X314IjGQ4+eZ+PYX0FKbtErvWpQNy7zTF7+Vh2QqfRX97exCnTPMIK/+5WgXi95
k7FtRWUzHfa2I2YWvvPkMFXSDV9murFgTfL4UTzHhFmIwNBjRlj43aEwsOK2jxDeTNMjPUhr6pMk
N9qdj+0GcYQj7o8RduSh+eDa1WKBVW4YVTlHkevkl19W872n832ZqZNPLGAneYSVvx4zXhqS+pVI
Xum8Y3orzBOjH/SWs4u7r4LyDfDV725ZjDlIGLVP6Ikdl2gS2XnUENEizwvYO7eJCFpCK38USKxk
FxvuWVlMYnXJf9TBFNa5Ysz+mUcGPmhhbEG6MIdECOkDl/j3c9M9PNG83IxmPn7kK0n1SnE3Xtan
qidJU5ME5EQHt2i4t2LllUYl48QW8cOiug78qByOrOlwlE1TRQ/kFd2w+RG2+R5JojezazogCwi4
JGc73iGoN7SVWLUh8XWTPJfp207SSiPq0TZAHvy9DMzjqqLcMtTpuhyQUoGhodppqD7h50URyZho
9fHJ0CgfQNCMPLY+OiAM3/Ym6QYFYowB0vVhgx9XG3erKjGmFL7sp0FRa+a2K0wnC1xgf+Y1X9jv
DMxJXdMpqoUsXQ6Gz43OpwC8Ug2aoLeqpwT9EIh4loRhMkoAXqGmvArsMmjNzWHP0e649DXTnhWG
IG/cpWIoeYHtUECCKuFkV6VrcZ/trFTfelni/yQt0cGTdHt+BbEOZdBcXlmPKIts/eGUAc7vKVS8
DbKhd7mAbW4ydiHu45ZE+XiNrtkUoFihjxV5pU5lt+lIPLnHQWZthIvilJ7//mWkoHtkSCs1H88d
f6VVeY13cJlYHLgYmPTQgLkk5JeXzpHF2VdfQse0yREpIobIpzWf21X/SufLihjznKDDT78USM3v
TXDu8tb6qAOE+uhOE6TT1rLiNHNd379EvPt3QB+euxNlriqDenwP6srVeeluz3ulQjz4svMfCsSK
xgaRK8Ti7hLEz6tbjLPOjoy9/+qbD+hf6xkMnklBJL5RmkKcAobx7JXY0Oy/10Zv6iDWd6cMvI5N
vEv8EKVO1O5etg7QX8p43vVIUrqgCelsrYkfQtDMyKQC8VNRgykMERPLdNsI8T9JvKYGYftGNpSa
cdLtRsjX1hB9t6WFHeRHyahJ401cQDy8npioe/kDVfH1j3unnpAFiwqN5556LE22KQGDMmrmyLYb
KYX/P2bveWEELTHgHPluTJHSONXMnwQuKY3oHuY7aAZEIPhhZSCyDbNwrHyjhtWkyiWWqwGG7O2v
G8LNFvaSOqqK8Vqn1F+ws9N7Uous7L4V13i7OzHInaRfa6sceRaJ2BWOL+70LssWYRv5lXZnTtz4
Kqrdc5mRChQpf1Y9gSpOUjKqhRJPRRCDEopXInQlpYGnS+2L+DCKyWLdKJnLLPWykedmCHPIwLfL
vDtRrxhVLQWXdPSMAIqY1rv4JQ/yMu3xc5ALDa2Gtl+U4wMrgy6Eug8UkWgzUJ9vBliL641PdFzS
+yvjkeG6lLlnOQAgSLP8thXBryy7CPNJqwjBcGXoDiUSuh6rI7VwO8bOda7KzftTJ26oVy9IBdvL
RRLoePqE7/Ad0cUKljthy6yTbdh7RmZ7W4jgxxuJCD8MCPoIcLkZUew9HtxwpXfUwNVEFIhWHRrx
nZ3OrZ2mzzVcko1UniW6fDt8LJjo4Z2jZ/ZgVrwmARuW0NG/xYouY0jCA7NXbMP/9cqNJbCrUQXx
jVW2lOyIhK8WDhKbZch5c1gDc6XiejjmQ1skyHBU0/n9ngn1PrhwD8MpFUPCn4jihGy934wIfmXK
2rFviDMWg9Shaj126F81hoe9xUwfyemYrnm9VakBG9gz4o4XUCpRlFH5UYQnaVrqnT7hh/NsIjH7
HBWjWIrBNpbWhu2vi2StotJ9P/KdSGj3msb9hvpW7h1QMHPKmFI6TCOivfS9+zUCQqlmr6cUi9yz
3cotGBBcKD3CEKd/Fl5ymiLlaByw55ocwR8PBsYNEH8/YYULYSOTKsPmGP/3bYFz6OAEK9AY+RXM
6BMRWQcdNUreuWVUnpbX8KgMIfDTnwgXb1W+qc6x/biJ2iRUfPZN4IvAbAVwUF99dlCjRvQYc1Ib
J4xp40Hx4vSIZ1gk0r/EHVb6FP3D41np6LyMEvkpMVdJNONXfNzFIijzn7rU+iMAUP8N+v70r7o9
lUGINp5rhw5scEjLBlyk6/j99ZxI3/DPjdZ8Dt5DTZFcYmzozvfPDIzkNAG4eTeEbIm/OyW37Sym
xSUbgRSEySjtwYJjF1LN4fq2yHppNEnd+bIOONfPHqUea1J7haw3bg32ASvZSw5caDiSaQzOiW/r
y18pKM5i/RtBs+Q/awm+nirnfeDWuO+8TQJVLDO/QOAczuBWXjVmDxwi2XuXjiXQfx9hbPbn/+oM
JekQu6CB5VCMm7kn0dBKz6bTX4gkmOx5tC9I9baKF6JexdqCJzjLPKQXgJa/HP1onnGL6t3E4t5w
estnRjkA5hiH9Q5OpdqGHPd1qDXwbuZXvZ37SMDyGABZScVhWADVVUSRKMNQQ8yIkv/xLYCT7PHv
Ba3TQnj5S08hIqDQ6yBoOlPztHFew5dM9QPEyeJZcHgbI5My42mPDYYEg4RBCN/QWOmKyoNrA/uX
JviMoFxzuF7WCizXEcFONkosR45YpeAE8GVm2EIMsYDVU4/sX1/8y99aaN73xeCrRKNLmmWSbENT
wV1EFgK0OdsfGrtPCPiMQe7CuuCfwi4ItTHOQgrCxlOPENW4sxPjYFfrazqvU/AcjVQ4l8kE4Hl9
W2TQEtXjss4ezCZgU59hVBce2YR7lB1sPLqrjog4L3y4L9LePbwWzcvpY8e8Z7jtNJZv+l22kZRc
wVy3Id5r0fyA85fuz5QgCKOZI9TwEM1yJu+KLcGsai51oGZQQpFQY9Jswf6ZL6UfW31XGqk3eqr0
zmdr9pVH7JiYwYzdjMCfXqJCYX5xST4N6OizPx9vOeg79e4h5wIO6E1TevxUkxT1v/SSFSVERwaS
f5TNBNBwgaypXLcbXfpBqdGQQFyPYBU05D4KB3k7EHnYJ/5XyTvkuKFsb2HRXvg/VImC6pb5I9ZD
uJ3HRXGnF6kwvYcWuLwOyGpWwfzphm9T6oUzy2jwEWPu8+ieRyAJl6TGd5Q/ULCnYwE/D3lyhrbu
v2ECImkF+5h3W7TAa563kniffRvqQ6+t43FLsbfdtqjDzuNd7J16fqnpqFKwREBjaCjceaz/vef7
fZ00DAafguKERZGJX1jz7fz1tzfIKmg3PVG0v47Nc3U6BJaxzadaUGEEsDFohwAm2h09+zgn8VZP
gTCYNwZuBfQtxeyaXzGVKryBvhECeW0SVQatOTDArnWXlbk27bc6iQ5sKAZyS1yRA+duaw6Nry+z
H8QXEuyYsXAgSSFt7rRJMqAcSLnKVgDJI8jX0LNk73BnJ+SY6Yl2z0V26hwvCRkeSyLGgafV14z2
hRmVLVkqIztpsSZsEzkzUSsH5nIndNePABFRcNBJg25SVNCI6sRGW7v3mvKIp0S4COtdoxNFAcY9
OVRuIbFrfxTle827eHeEmY6x0DvUpcPHt46h9utU8e1q6eSDUySCwNl88Yu16vvYKdRzCtYkith9
24mJmn3g4L+zqhZtniZrc0Ka2UuZu7G+GTevKvAJrFCiGQ6Y6HZZVb8TdX83NhX5GSOoX7MHVk/V
gO8bBKDM2kRfBNknArJxPxbRZM9xSqYGcP51SPIs+dMfkmG4I+Ra3/auR505tvs/5qNTxAdV0xGi
7O4sc7OYFL5MugGGfW4cjkSjz4J5N4RYV0bhbfXG/sPYwH0OFKMtUQ6buYVVKDs2zEBsvpXXj+dF
XNg3TVnEEVqK+Yd8jJeg7lT3lIWv0b5hzEBDDWgHp2nEKKTDW/egxfq2qBiCXaz/ouHGnBQcaMYB
Oj2gsEdvUx5fxs5BH0TyJkyo31pbLmsqbuNif3e92JlsGuN0BHwXAMeU5wK5LI/g7mHAmc/a+l/M
kwGLAmX8d4H/m/kMXr+QAz+4xiI++rx6UN4rt2IpQPNKeFfnY+0x8yIo21+vzwfm5qNRyKBD8fWz
XKd/w4uE/4IMACo1CIFbBDfDx9Xb3jq7jmjQjK76r9uJ2R7jPqza/3AOO3XVIseffyZf7pN1th4r
RMkTQzkxl9qWKNUs/uHdFykjdaaaDHjWxOXhM/PRs+28LXf58/GSpBr80tNPTC6Rf67yNDg7I8oH
/rtCfiVUwleusNSOb5hT7HG4Ill0cJsNKoDTPuDNpdyFX1CAHkbVghCapElLONCMdEU5N5BKTaCs
VIZx20ILyfi2a3LdO2YIJoIXI0JAyxjHP8lWiZr9roQCB6FVUD+WfSAfj7DHEU55xMAsfAXMhNx2
SoFGzDjwDUc2PTZQT6+GLxg5UybhVb3M6Co9qfCj4wEwWk3GbhmW3CQnB1wkY1tlKX7UyDXzvyhn
bluLObc6ZgiD53TVwa6wfaPQkoALW1Fl3DB++vIMDH5GDFK6/xMVWLBpS8mwFAIAK71wgfl3n1RY
bamnz1gFvHO7RxyLpP+6NhwDjeuWc0rgX1S1+jcrqBTBxUmsyawHWnC2wCWbiVnA0/EUU0FpuFpJ
VE53xzn+9gT9ADBz7Kt0J03VUBO/MnwC1e1WkkwISAmQjMLx/eOT6ZrzyJl2B1wDBQfI9Yrwn8cF
RoTONGVmVwNpzOfKwE919KO3+TcNsxtXwvV7wfsKth+SZ3qbJ8H9kLxOVQpFFCi0s144z9QD4bUZ
7y36SFR2CqEeOMqCgHwZHxkTmNUcM0kfEU/t29k25XO6EPRsOKsNGuyyXgsG+ICmGHi8qFboeiLs
YCcOac7MsKiKCexIuXaVMWlm311zp44i5cBRfYV2MuAcwAunZzVoomKgSFb5CDh1qH1Ev0mzidRr
0V+rTKt0xcvfzBE8MSQzIqkBaCt0AiXf/OutNd3j2jP4VGnJ2rgp7DWkk7sETUPUQLZARUn2MxxO
mc/08QuGrfs2L0hfkSkt04QO/Y/8uRlsWyYQOiLK5DBSR7psO3YEphGloXW/uMQm15jMLw+6pg3E
BlzHA10pOvW38ztQ2ILhIxw1jXdStd3otzU1IvInEf393kbWrAiI58ZXOg21MgUrNuLBt/96A6gj
hC0PHQDEsGrW1ctxyQrQR5xVXdiXUWvyuwnIoIzVC50n31pvE7p/bILh8P1DPfpszQTzHhPwqf5x
9cN0GcyihUAFRaVtoiRZFldEYLrWPQJwSQRbNu/I/VpQkBAb1HcHIk8qCIW6V3m6KQPL7fFePZXv
X6oIv6Nf72wOF/dITh/oHki899j5EhpVNM+6gryeJ6yOy2yH0/YFuwu2T09QTL+rnJjvSAEbc24q
SmNW45JdKtxXA0uS7wsr1nyQ/Kb+KeTCSYFOtK54iiRTko+QV52MjZKX0GT1t6OtVQRo2hCWe0Ch
rIQFQFLgzxyQSTkGgTHfX2l+Bb0tJuonWMfh05gtJaI+fKDaepJc1LtBZIhG3T3mAXnxQdxDsmUM
MC4NnpqZrg6MxZ49Mykio5LYykJgtqcSXmxssmUs89PfJJTRm6uRcO71S2aAHP1WQUKvEO84lHvC
1Oc/SsKVxVh+a45shUS44VH7stkOE/ANyd7oM4b1Um5NmeVlGE/8Pbv4g48YdOWQSNufCgplURpj
lMd6NFgiA0Y1SjB89nyAIFTBZ154roBgeDI2Me42VPiwuzG8OFPtU4MHGElwozeXF6eJtCIZxIgP
of55U/768+792Hzl6idMhOTnAdbVencxYV3M8WPKGbmryvIwNeGCxnOVu9HW6L+b4Ttxh2c/YTXv
fi/4MmpT0Z7bSW/P9AdnpL0yK2scBmL/5bTX8jMP7fh5yDnzdXXjOIqFQ33qCsvdYWYWaCIsxFNe
1R20/e8AZderKDmZ6PCCKEmpdZJJbg5WCkXA662XQwp+3jj2EwyOw8qVJumwYQEGoBArp3pUV4RY
AgiwojB8p3ezSqcjUdwAvKkyGJpTnn2Xajud+jsohzKY0M5iJxXWYyYIkzAjHO5DQhuroT63/bWm
sIZf92eLt+Qsklm0wScv9FdsXZG9qEaUVeXq1grAGFje1uX472QG3kCVs/XURKqTzpP/L5UoeHhN
t5u8LJ3BGzxqdLc1vZ8iW0deQ0iyXil8n0/NdhXPWFw2XPi+I9APsleSc0OuYqKf8TxiN9DeLKbT
NHktsYAwnjnIA4y47Lwrz5RqyxOITtf9t7ASKN6u4Ct12S1FUhebRDCsuypt6AC3pHuMpGy953lk
QDE/OnZV3brrYL/5t4LyySvUZ/IW8OqglexrVX+JQ4lOgz01DxZZJ7y0leAlRRM8S5qzsglH0aXu
99KgzTUJzb+ZAsXfRncs4iCW/UeGMvM8BlYnMhtYivbz/rMgN9BDgKxZTkO58vH0Xq4aHdGgfC5L
J2DrP7sW/GePMVH6UmVNnLGXu+PIrjGiy5tfsUSWSWy8KBg7C0LHeSD7qZX19JTb9N1qEnTazhRf
Mr/ZNFeY5cwlEC3xKNPA+jk3h9w69vzmwEg+RtJMANBFdD0aqEuLEVFnsKrJYV9sR5OoMvGDNWYw
uMICSDJ1wu5eIu/zTeCz1sSBfNINOP341ji6TGnWWUODOrcgNtayWytFPsrSHxY/ApEUc4Rax9Wy
WuJBvcqx4HM0GNj1BW+spKYbp/Rep9QOrbJymV2fwnD1jeX+gHQqK+HwC9LVqQ2w+gbjSj4ETOYd
G0I49+98l0S9NZ2C3UexQaHBKARnkhpdfrOxSWs6D7vyicT+VlAnQkHc9qgdE72KKQUrvHJB9Wor
hTSJe2cbte/GTz3ZtrsvrsBYkB8MIlER8Y6t3T/yp7jcghuGrytjqxKfotjORaP8k6XiBuTMqpQo
0NwAFwsYgLhMBJRzZeCySIgfo0FK4PMTII6zz1/quv5t39NyNjzjDRnhCe3un/vW8CDBklG8zitv
fVDRg/RUuwvPkXRF7/gKb214HPj3688c7MOiP1n4vp2xnZRNt8BnxrYAuySV/270+sixzy51sPHm
N+KfQ3INtSyB3qGN+zn41YoZwbq3GzdamRz32AzeDkE242OMopGLQxXdF59Bq/C3Z9OTYlePByms
rKEjNu0KQnMtvEkUirdEw1NxaHk1z+SAINgVNatyXoyIMu+aKMT3ZvyeLwTNbRryDXioReMN8ubZ
+ErCSSSyN1HX1yh3XJ1pvNkiOmCJ769rvQgMqLtGCqhXrTitidRgFJjondNa5QUm+7VCYgmIjLH0
loATY/KbfdMpWOIf9tjkTGAjcXxhUYNMd+3IW0HrWpKdK6kA/QD2Liq7gpsjdRtU2PnZE/JR4Qt9
/na/qjnQXVf1lEXNW23+bamjuXwRDmmozIANXMiUeVfIN5phfmJAwZ5N6FrpYjYQ3d2oqjMJVVWG
Wp/RvFCc1zl8S1uWjBzJb7ADik7omYPlHHV3cVbPcRW+yVtSkbLQU7InSKynxv+XMSCoYnKhWDmb
rgrVHWMxLqXuGMVsXp4F7+W+R6M5tvGZCCITugxZzRY9IQcei9oI93EsjsAzF1R8gTnQarDG8G6J
143yUA5ry8Smtwt/WIqRDTw5TTh0eWYEoy1HHt36c50xiXBLvsfbXhV/9/TNqoTC3WTNG7SFIafN
RlaPgwUW0Td0ARHE0Zirysz5wbjND/C1rqhklhY5gdEqoNanHIKqMZ0KtDtx/T99xJgp8FaNccfM
iydjaPEtA1M1NyySS7JGU2gAiil6bbcxYcrIFcSnoc2Bq2Mg5YnLA8LpzoSBkqQgv03PYIbmW4Fd
Jd+3kTku9f5PEg1ydQhzQ2n5mvqIM1001I/9o5qPVGPhze2XG+eBELvB46FfSCD78uXOkqcW6jEP
Ez1PdRTXo3bsd8a1sLLyQGaInVAAb26Hujj3EDJqtbvLeDG85d91Bp9432MvbWzsMTzyXI12wN/N
RdoBmPvfnMlmB+fKcrF7HkDc+xM7i14uzTFsEccTcoYzh/gncwIBoDiKEX3JXn5TYXVdQEGItwAU
sOQ0OCODOKbSeLl6+ViAWUSXRvS/+GZwQ/sUnMIFuvCGj0sD8ePtuQ1qyj8T4N3xH++X6FIjPQty
kZWrHnpjdfDhPwHxfg3nZjYQaGI2859P8DtpHbpn6sMhyT5oj+XKrEFmS7u3cud1GGc8ae+GRgjN
1k2aqHMr9D8VxwnsO1F2WKgiT+crt9N1UMB7riffzk6tVOmSqqjen0Q9aizrL61Xj4MqzTUypCD9
gWtLPXjRASrOVansfHZduYuKz/D84gqsiQdTy6DckjC/EsXRyg8uZFTxEX28OnYu51W4nhpdGZ01
Ll1AysXgYoxeCnkCI74GQLY38UMuYsenD4rrojTB3oBe3e1wzfqUM0NemMvXYGFf1cbuuK6mufzL
rf+PXS1sY4LNhij/sfgfhiwD8pz2CGqxN/G5r16ZxLLVl4YMLVoTZ6ZH1nsE0l6PrpjbGZ3Tu05M
saLG3likwgbbKwubTN4pR58vbODiYWuSd36SlYWdTBhhCtcmQZTQbAY7SARr/QoXH+C3QAxEHeBQ
n/huzcdgN/msNaQ+Y5yhMlfqxDC0d0FRQjzGPCknrzxX3xoPKNoEexfVJGgpTvyWbjiS/JpqbDLG
oDSRaOEt44jZ5P4mMyJlCMTKEhFCSNWJWNrpNeuUI4JmkqLB15Fq5GUPAN9wAyvUXc4Oemoxxaf2
EcIyDce9lbYAvP0Yws8ja/hLhYR3AQrikwheynw2v3W/fKmk5afuZnQ2brcG72rMM2jYxK3k2Icr
QxO9AnNloVO/MtCWbtA2PQf+Vse+NZZSpW763WGqEKAzdctNk93E7mp2MWFdWRdWImCmtKzHOm+c
kHCZ9N0sl+BilSszh1sz7gcDmCSN/BGpWxVROK/rPPsIufXd41m7M+IQp37qZYh5Mnm7rJh5dG5L
9jdz/iIATCoqvpCDQqYprNDPFpRaI3wcYePXaPQGDBhVmoKeF+zvZMx4JU2iT5cSFiXDW5Z3JH+c
m4sSJ/QHh4IyU6HWH1aPmonITj3i2yT4qdHKA8wWNsTKnIJ5iElr9tHTFEzW931steRZ8sj1mmNl
qD+nLaDTxVkemu8Uoo2AL5lUu4AuCC3PiGEd3NrluowlClghmnsLgfw8N7ShAF2nj34kqwuwWTKY
B/glDwCWmz/rKTOYZrWnnRpMXtB7CXKCLn4QBa6RSY5/Sm/UAxBsHB4bd1jY+Eje79GOAvJGXQ/P
efLs+MQjAqrQerqh85rBrZGcVlxfkuB22Uw5rSZ+koPVX21wYeFOFvYbdV9ioT+HNEN0c1kbiCAc
3h8rnOSGOdtVGr7k9kpcMBF3FF0XImFVT4j4LtX1IBmv0qQbLfagDG7S2ywwpkKL8cCRiFliJ4/I
Gst8cB0CyfY/tesR903PgkrzzYpiadc3IdnqgQNHYMzQh5dn5JqgPn+RFz2Sg4TNpyet2yORZLXz
x/2P7saCF4kT5rgUXYOKI1/YbM7mI6nHSouxExACswDHoi51WUtBVix8ukNTnKVZQOBiHa/kY+27
9Orfzq/JpsZ7CxTPOP2Jwbagz4pMjDaCjoYGZy8V1JJuQEYfxVbA4mi0vDCPwdbT05h0/RXPRs9L
qDKIYoSbPwEw20B8jOD2dfmbkXqK+kYk5nTVmw9r/nBeljTLEIL0x/FTkv27sIdoQB/mEsp/Na6o
rJ6op47GMPumE4AsQR4g6qnn55Svq2o8MF9jx0WcGjFc7oEjzaArcdjXkmyz3lIj1BSSivxn22z1
yv/DQ8dP95pfMh+9KFVyV/oJ9ifXX9bX0mA1S1tYr09kxaWCtk6833ydfbAjAeeZnUvz1ClE5SAF
Z3oPK98VBa9y3TNTDhuZ4/EDTY0HgAMbKftr2DoKvN+4FrED4p191xqoTp/mAyqm39pXTAhtOfyx
9hbgZcX1ne48h6LPJ8WcfEvx1lpfpVSVN9v3+ZD/txCFRLhtBEUkpEtUYzTESSvIEqsA6PP3DRv3
lXJQN2VJlZ6PcsrYtmBlKWLKbZ+48ZYKteJ56BZ33ctEZOzeHI9HbzG+0swt4lHOaBDcEqjLUnBz
HaG14L1kBqJNJlNStHKmBNa3RtXuJnhZ7zVWF477L4wwivx2kdmb1J1iXUYlomKLcvjuTCudTOro
GolBdlxkdyCBCC6CzvwhPP7wQcO6HOXDqknqsMW5JvWrgbTkryajwDr2ucpde4vwa/KsDN3X5tmB
CslU17+j9AI7tTtIWj4EwcEHcCBlX9W1+NxWu9y0KAQ+ap6xOsDKV0mxjrf+PeHVb2qnb3QqLutP
9dcveipggYqaNN2ajLzE3XzrAGQTZu/JfTu6Xx9piCEjM+vM3wJMbxXASXS9bBFY+syRFF8ViiJN
hgipICljbMcWWlDgKEQT+dD1Wmdiwk2YsSAiPsO54VoVNNjplfmrrdZz7tehMahtoKqaBj4xBFo0
8Ku31IZr4dArnibhQhkN/v4mYydarKnOXmxKqVUhXV72pfQzW+G5vDMcJxF4mgW6ob7gXIXtKH4m
dUJI5bETuG8Uq2SejdoJT8tZJsCspgi+mqL9JFzcS2KF5xGdGIsyRfMin42Cs+pduy1BOvy8ah0E
pVLgtHz2jFM45qlBYkLZ2jug7Tmo6nxnhsxbwX8/qC3KM/2WFIlmhggJ5jspOiolLFvjpU3VlztN
X899mV3U0pKHMT6QIzHrlYB1G5RMf39eibNyN4+3wqyFsfG8n6efCVlIBpGC7rQzGDV4IGGNMC1s
jD4CsbFFQzLaWY4re96QZeOpbBuz9sq3eVXQzcXpIOq3h5bf2Cdd4khYMvqp8SnOE+2iILjx2Dby
K+6rZtmojGDpr9Zo+zORvO3BKkvURqe/gDPAy+eHSin+CrUmRTGm5eA+yAUxXmcYLviODB5a6g6l
i/3crdq3DnG+ScX+LnMVVKEEIR6U6gPMVWIrabuZ8mKOFF5e1WKFBezQYQDMkZZPLyLFDcaBnd0C
/crY/BpHr8Q3bCb6wBzVUVbOs08CaYJp8QThtlfdM4t+cpWIHwFQM7+dl+Q9ikowrYxBuNE+UJ+V
oK1MKxIIVTHxAOQLx/37E3Ye1i0+Zk+z0i//FrqzcXjgkVGYL5WNz6vXhCgKNrgRFpTKaA3HGWAi
BTzWLkz+kk3e2pVhKKlLfHF2WnXmeuHr6Qgo1x3EiNtENrFaYZA8Kark328csAsB2FwJ97AWusds
3CI2B48SbH1/ALC3fDpijVXHXE6zVYkNz6QFFmpEqSLvIidbIAySRBUhY4DvlXV4Py9ybhGUFfM8
wcgCdCgNfrJMUlYHoG/MApaEIy+s6yFvNnnJiWsU9jxBbO+eqkC3mC5EVqednvH+YCYiNw4hJi2x
5HongKnXaT49j3SkVU3Iv9zoh1UU4GYXzqu9sYZlLUb8BG7C/nYcDzCk4RYu4Hkz3HULielz4b12
85zVK4ZDnrwKlkBQNh7ctGw2NR7pSm3D1NN4RLszKPTw22m7t06yIDTZhpuGNh9zFymYGDacaHXj
G8Fw2tmsggjlLPCgQ6zrB+liq7darNk8U4Rdb9vew2tjy2NM93/8hCamJBm9OUmkTPrFuxbpeHj8
VtB8ToM90re6xmil5Rn8Yqp4DAlcQjH6iDS6XmVSFkSy9iGC9EEkmtxBsHrA0sMuG/p4INj2MXY1
uoOvwj9QnJI60v9y18xaPKv0BaEatzoJ+y3AvH8/bC1Q+WLEp9Gd6QW35AyJezL54FfolCGaiihw
9RMcwwtXcV+q0q3G5ZLI87DMmCMl6cJvDUXxQmo2UH6ov+bTjtgva4F9tOM7snYlFQd8QIRio9UX
jIpQSu+yp5JhMxeIAhiZ3GJslVKeEHHYi9mTn39zAyhaRezSjm7/jBTYsmHmdeTXfyGm0Ga1JNM9
tFTeBZIEp0osFmDudBkUUD1zpv+Hr6R36s7i4f0Igw8U/5QLNs4gz3lOKc/J3o4xG+C3q0EUme+f
LbTRP73WNjBklu7dW25n14J2jXVyjOyiYgL25P1gruBKNw76+9O+xej+aZhtHyaeVhaHk6AQN8Ib
oPvfnUukmQ+/Tf8itNyAStL+s2w5Nbi4oLlD+TfLh7KgCju3wss6TSXXZbBLCSTve6r1Et+o6Kk3
mpRqMB010rNuMiZNS3sKBY5H5EDUluGEuHjAitCfXpxv82z7AK4qAF0rbIpJwMLJpvs/cT3J+GQa
zLIASX6dt0BkU7WYx7TdGinsfP9BwHVy3SDxiUswSi76JCXRCr+2TiZd+51kdgls6ahRToKfwNJ+
FxssZvIMvRrDUlEX6xQ+wEC/tXDzd3wKdvqfFxE3yrzVfyrW2VD1dMm0NK+8BTXqwRmBFD3hL/rO
SiCXL1Ayt8Or1EOKMWC6iz9rr7s+WOcx4j3zK5YFP5bkQMbavoh6LsKlTyedZNiepWDf5KSdJF4E
RePAjQObsk98Fh7UOUYVV0HJdcgxHem1GGxqF2PdT0jYjqpHJQYbzj/untpQgDLsOUl9qRnVQrZ8
IQBk0RA6yOVDKp9k2aYORbcCVtEO1SkWhoM09GeeWkRKyfUjeRrtIdBMVrvexyyXNIo/3tlG8g4y
Sc9sokiIaIFhkZPoUBaTMdoHls578WcNwofdgdg/O4mS+xh+wubxRdEndGx6G7dwcenEAFZ74u+k
tv7KfDC4apPfuN43U3+g9eUOmxl5+T/Zny2VvZ3pYCiijTVC5wjPqrNEzKNSSITK3eDoaWu7I/l5
w4fbVrDbpdCoCtv0DxZvp2S49WMTnni9QhlA55QVx5g9smpbAkJN6JGARv6j/xxPPnvjs4/NHrRc
APdcQ21V1gXxVoYoQPiNEV+bnAFPYlKyFLmGn7d6I1jnjkeKk+zWsZLei1r6AXFBqTPWEOKhtIUg
rGhCJjObZFvUhp1kVOTFX96DVHAeoS6jXD/VuTCGtEKtnWpHEpzqbsBRx8FFxVU25wUzjwBhSTXo
Pym5NB+gvOxH4mbu15NAcDT53vGK1KN4h77b4orsVg1/Ozv+bGv7gyg+C/l557OODYl4Wopjrr4f
PI6++3xmBgzkM5MtQJmtI4CoPXSUh2cnarha4S2wx/+yKwpdbqzHf2Gq4tt3jsVB2mgfVQmVznHh
aJnPnKj2wZjFhPiuUCQ4+TDm1EQ+isbx52cNbLhI/iCvuEpeFDh3FxueNoOf6ZRW/79p4PH2irot
IwbD0LxO6GbGVsFDafn1XASDDpTZIjDRf4XpDABijj9G99tpSndV6zhT9cs5CdvGOcaGxyu8ZQGp
rtcAdb7mk5+BTCGnfu0xUHx16rzoJXw64lMHg8U5K4d85S9SLgQEbtFciaJgWjx15pjxMb6V6D5u
TECj1UAklF1XKg4Y13IXp7PiWw56Lm1CY21KAPpPt4WvH39TAKnxH6K3LNbv6khbk/DnZQGpwc+u
+Gk8k4L5Af75nPOp5Im9DAgBQsWLsPEG7I8L34UuU0f/BxZSAfnQZCkWMCLJkBtfkrfYKlOW9OW3
Jtw4YRm5xaSqn2rClrhiQ69tjJc4w793+l2UzIxc4IjrP9WYaBdVIuxxxafjlPuqHjam1Zh85PGx
Bd6nUpoLKRa4RyB0BiuoqpLBCGgB3422AAogtUcIHJ+k/lhh9rGOQxFkGI4hPez60yUB53LGBP4P
hl5FYaS3L2m8qs+glHcb1DfMjK01/O7z+PWRvqcEgZwXsm3VG7nfuZXaIU7UzWteR10Sa7o1pd7e
CVYpmsW+VzDPujOlb8BBroqDlEK8CWVCmDDSahUFdSL3ETQjP7zQkwEZEqYphiu+42qjLgrO6AQE
rzHe/qacyEYCgf0g5ynpJ18Q/al40GTSPt4WjAks1Po4JjZoyavBY2bcQGVphgPWPDm+DsUGhZsr
QDJzc5iIVVqHVc6cLy8zm9Z/wfPlkDpYy9df7topjSGO+k3U85YLT/UojC37lS1v67ZrWKpHSShF
ck7kBpa2/rdO655R/Znrb8zGG9ykhHK8mak+uopXK8XROb15se7PmscE/Sxs0vbvhswNhK1fE+Gp
rDSXmo4Dvy/aj5nGXL4HzFNYdKdqzkRwLZEK4Bx7XfSl2PtIB6T5T9AD2Bi++ou4Z+uc0owvmNlq
H2KHnQYFDZvvxj/rQ3Awn1JXfMon1P7HjiWPvb8Ra2hlTPaWOVO6Tz3lHZFyGM6AGokl4Ct//LaN
sl38frQaJ7vX0opyNMZMhykjnm1QlAr9dZv1oHPSxpHwMKVc/mMys11QPy1g4SkBLYgJoHOFZbyf
L8soQONNksNgQYNlYbdPv6l8bsOoBUMQ2dbZi6BPSOtI5w+RpYVsAq4vEYzVvnDzti1ZjqcQB0hA
EiL5yQyfaMQ46mrfBVTUr+IQ4TJnhe7GuyfzYMQHvJ0kAnBnnYMzyHDG8kxWxPrfu8p9a3eBBcAQ
sqpS2i7VAU1d5QmL0/aQw74RQeVsecLZ77DKg4LE0GnePia4FFdSuS+dXkzvImZGboGZXuYAR7rp
5pUniBTxMPiWrnQ4V4lOjZ3RLJTMRpPbdryLIn35QTxDzpkK9HfKjT3+WbBBVNCaKjxKozeFlAQE
+Kf7mSnALGExhG09rQzhKkFF/c34N/daimp1W7QN3ADU/NkWfLDBwzdU5jKc+xrNH68UnUqL5Cwe
mMIGOc89aBA7YP822ikFX/fAOnVdAmjlfiVDSUGiX+qgI7tm6GQqoM7MraOYfVLvcjtlRAAfr3LO
yiPuB0KYa+wZ8dOB4KW7SOiPhjrXo1n7ZgK3N9aCCp8AmDQ0NWbI8dy9FYsupInJG/308rcgUB7e
QrUL0BQrwQlwfpSujwfnnvOQjK7MnKlXkSwvmmXlIyZWmOadTz9z5ecd9TIX9nFUu4DYnze81CFz
JxEa7YI33mI4OtHrN1DMNsMfNG3Yh2YXHuJIcqM8r3Lzw5rHYpb7t/8gDjnyCDzDqWqv0hjfzTCn
TRzRE+R/i8UBFA2cigk1s0iO/PlTES+soFC6uX3yL91aLyw7RWUDtRxQzWUdbQ6A6fgmUKwpzwfy
lKdpKgLqeAMBTDobCBhSx8/7qOBuxGZyTdyBfcrlhsomzKID5x16L9TVoqFIQGqq+5kSwS1m0fCD
v7iDb2uZVqegxofQI+LxT5UHSFbHlUiegh7dI/IvOOGtHdTv43vjMm8pmxgFBQM1ozOPxR8tdACU
CZF3v6TOl6kXW0+vZ17Hd6IxjzEUKuE7hjDh1XYoNf6j1rsHX2bwkXKsMToI0W1gVAlw1zABxmUX
40Aj5aAtYe9HoDLI01sKAPiY/1i9egV2OTWA8G5ovZxC6mEx+CP7mUPqBGAVNU3epgmZZrhnAwJn
JWstYC5z/sQ1VuwGsjmyoVU48BxxEHzgFpfuZkOZPegeBaF8ZjI0J5C2aFoRI//nTm75RHc2lH52
ML0X7zFkRa2GFdcBBrcf5UCp6VYqs+lE92xunccuFFaeU8fMh52f9B8wc0c0p4uhSeoVJZRHoUH8
eXWrsgc0yA0z98wYF9z6iONNuYtKZER+TFSvmWysMZ0SneauzdKJCQgriejfTfaoqyPIDCHL00Gr
vCPf/QL6iVxFRl3BR3t7npopvVyTHoTT6kd2EE7OmZZjU2dgPZ9DaPphpNRYnD+iW0poqfFfXrtK
xx7uPotj/0WBdNzgVBbu4BCHoetSbFTjUnuJKm4nPxhzDD4MDUS4GSMrA0cD/AH15Q8JSudISERy
ftCKuW1/LgIE81yUBffkBC6CU26BxgPey0D2ADmlS3EKwIhy3+0Gyu02pj7MaZGeV9Nv+opiZhL1
2D+O2eMUHpzs1Cy6APHCvLJiz4wVQ9n1Vyt9O+9e42HHvN+XeWXr+o67yvxHRYoUldcl7wD8kV+P
NqNBHSHIfaJdY3FTD8+VXsu0N/zNsZ3gJP4FLij4cC8uildMIV5K7R/tCzQOSluubW45y7lHfgiL
t5+cz2OeekGgevqay+orxwPv5466THDdWztpKX1/MPIyStFR4W5Rz9AVGxXiXXmQEIDUwsdafkI2
BV3BK+8bhm1XodIAPds8V33SwtfTSsp1NjFvdEttLDo7gIrqgWJD1VhETIQNC5CsNpySSuHWbxCC
PQo79VwbX4N5f3ls+qQRuRBst81iSpuYZiHpIiaiQHyMdN+8P/Js9ZklPMih4DtxaeKLy3b7Dbpq
WJmAhT6NYcvpcno9qY3MJjHQgSWUbJIqWQAeKa5zNn61KX1YLv3XhejVI6GyYgyvCoStcCpDuaZ9
vTqLIagp4fc815UgM6ZbYJ6v6j+fviq+9IkeH93pntKdbcjpRo/HrDsXOKq6PDdHyqALDQ0ZzCai
o110+3BiliiX11qG33Lv5fzI74QxMvdkmZ1rG7Tvnvdgchtc/zhGT+bnk2iNLPa7Yj/3WMLHCJGm
xUJmr6sLeUOzOX++UsEQcDD/kJE8womD5oy9doWCAGINisej84cA1EnCVWGWzryAKINZim/87r27
EozAy49XXmLBnztdUOyniyISbk/k1+KOA9wTRljSpG0W2yvetnA1GJbLjGUKZxCkHYBiDURNGbvn
6kBV3if/oh9Pccj0xUw+eTWi4NB+87++NOErMq37DPJXAEGHGqvYKU2sqO2gOlT6QPKZuaafX+6C
rJbuinKyX9DpFu/H+wyj9Q+7oIQAmgnLcigKgkR2J+VxUx0iUpohEheYscH6qOaDrx5wqcPzvj6W
FULyUI1AwxHf2ALtfaKkHsXVw5Gfn372hiOdkzOoRgHDRxY/pOcyQYuNUHM4E1/zH2HpRrbRwzBx
6P0GKW8ldWj5bFhW772pqXL4QAopcW6XscD+ho/+kfSinLeCDhgc+5Zdkenf06c5iA/dbGnZiirx
D5Dr7gLZSRMxet2+QqQ1hvYkf1x6VzHXOziRi+FSjDVqYZr8Nf1zfe85HVqQJTd8r6WjXB0gOIrW
9nYYzke5qzMuS04Mg4FMOWKJqvDTCALrl3GxJ+/EoVuUK1r+77ECkz01isPc432GiXS7BxNss2Xp
YbGOeRnVVimyp6MiFEL8VFxln2Bmeoh6bx1lb9wzweBFT7tRXm+az/Qu4oudGH8Z7vC7pZ3kGHil
cteTns5MW6324TXl5TDaFlsB+JCFJu/JGAN/tpspEAL1sqfWuVC3IsjPGDUzxqNzQcmrKw6XGEEm
DOWZbXswRSCn5OOtswjMX/ltC4giIfYRVnkov70ETYDJG0XKJ/Ou922dAQUwEg2XrWROS4DOPxGT
TiVkD/GFMarE4/4GMm02g/GYYWvA0Z2+m5DEQ6b/MNW3WP5VeSkOrM7sde5egl87LkE7YDelqh6W
YLHc+QbtoNuJ8ClwVGdffNO5mR+2ioAoo3QTcH4eQhKyZe5LAnEPu1MXKD7fR0ZmuadirTgyaDrU
UG056h0thXGD2X269EFJZR5z8B9qx5f1vuD4s96ptqVD79v0+QsUkUHC3eKd4+fe83jEgUfs/PCK
MRm3IaBEKW5kYVs3MyUZwFPnuW9AeQ/ZpDsyLvVaYUqsK4DeVUPi/r5s9nIzenUUaHduH9kNq6QC
Xb4JxwfTmCXqnKKHdNI7h0C7qrm8cmk7Wu9nQYoZ0TsEPvVTj3SQlHXTKfCKk7B+K0kN6u0BTAmh
blOaxZdNVCVz1Yb3gypbhD2ShCto7H7WKRJ3cE4dXanTFuSmpWyv1YLFYpUodkBTKR77veznsN2F
+5ijA7y6otsH609Zhd6xt7oot+a6qLVxvFiwXDb2z1oY+ywQIFmVWSCk+rILoBrXed0qD4CpCyFi
QTDkeDQ69CSOg4S4Rehs5Et94ewDhkd/tSr2Ad39tzq4Qh0OtJ/odKBlUquZrypejot5wXjq5yJk
k/HBOshl3vi7DiQeXkbwMSpfOq/pAK4sdXnEL9jm4HIqu59Flx9bPWSX2BNNFJTldWlwBsv+UNAj
1uVFmYxrRFCn96Lzr3E0dtpX2navzoFW49XhS9rRonDN88DnXT+YJf2evU5HtQBq/k0Hrrk+fQhV
yxpxIJQ24aO+dblOF60dDbJLznEEHSwaRuRicRrV1k9BDTQhKxHndmZWodE3SBQHzBY8QEm5XZn6
DsF7qtu2pdtI4f3jh1bT5ol1SlrHjeAUY5URf+G1AVTz0HzGfxR4r+TaU5F9FXlJlfeiFvqmiGLb
JsxTOV9KwuuyQHemn2qsqwVfXNGhJ5D+Aro7PRwfsTY5OqVfBmVAu3igQWqzV6nn/Yh5SExOI00r
NJaqkqQSQk6/EyoaVLCdnwmi1BnfFzAfVrHcVg47wurZ8cbEbZwRnV/QUFRdmsxkDeMGlhTu1Yjo
r5r8VguV1BezlNOdfBQJxOcpWhgZZxt6Vlc51B4GokjlLaSWxG1DTjY6TsvAZtawAKP2v5p14Reb
XugxNuC/RlEzcf6kBQIlCIIeNpCPsS7Sdn78fw1ozRqKOwPo9FXfPKZY7zQuBcS1AHmbjfevJoWX
9EEFt1MVJV/rqPCax4/Wnhm2K3SZj8i875llWQeci71Y1Q7ugMKgm8YT5c6vVb0Aj2lWO7p366H7
KD07xGz0Zu6H2Kw11U1AyCIXoYuPORIEZD+IHzvxtfQqKdg17GmdkE10o9sHIzonMG2o8PYx5DYW
zGUbx7a8NOMUlkXtHAqu7l3TUjBNQObT9DZ3jMoVyIrfpRE+U4UHSYUMTC53BCmz/nBHzcdoDN2v
YqlQR4nZcULF4L6cFcLGuAW/AD6pfNFgPmFmVJsMlo2RX9cioM1cPfWMweeWuKa5XrnVUbqyV2Me
XdNFdLYiInkWAZiVG6NQNAlcLCClj+G7c7ktkqN7+IQrYJzjovo5Tou3u0WtLUfxUrjrTM9YbABy
Sq53QFHPF+X3w3O1oY82xEeTAghhYndJ6Gin/xD5pYc5GFW8x4KrmO85tXmL6L2YsrtRUTWMbLJg
tSgRCETlTtEOHW+lVWGOXVZ/cKCYuC9Mf5AfKcbqvhbIcmwhqP7Rrl8VsG7V9YC+graKnmEeIsm5
rdPGnaD4Gt6OhcEZohi5ubQCYcKfZNaH2CSrhVzpIZpRUoxU6Ygy5HDgxCQxpsp0jeZn0qmWMX2K
QH20fEqrcgRQBqAB5Q0A6VERbBX0UtMxnUtiZzrsi7OiCT7sUeikpvwpBzmvpFT4HKxhh727h8GW
foxhzMYk0hipFbRQI82DNBRB0P8Mlh9HC8zFqH7unHfUu06LtCGbWWUMlPrYOeV4djCssA+14BHG
G9fcInW3FidQChoAMZxafomvVb3bCK6GNaEOrVHQaodFT9Ys6l6dppOi6a7O6AiZd0DCaIsRPW8V
AVurJJoarWu+iqnexxsGwPAaCWkEApVnzEkfVscOTdmzTfCGBJViLqC2iww7UOuB+qrkuAN4lsq4
N4qUqfPJseP6gb2QEig5ehzCLR2VcIBL0opbz23YABXMQmOdTMkwhBAUnD+7+P++j9BDJx8og9r0
Zud43uCEcvhcC63nphwUoiboqp1DYtGqG6z7oXjFUu2AeJuPt3Vk74OIalnENaHx9udP9lYOxP5D
fc+Aexe05YBBDSkXYQ+tAJRlco1ObCV64Q9JJ2DEk4em3+6ejqUGnhpio28A/z85oAEuKRf3eKOr
2df+y0zBoZAstRcUs5laWdepLaJV/J186+NIiRsGt5OYbRo9uqe1Dk7DxL9RyRhUKjt0rgWpr+Ls
9dLUzdjcVfCpcK4eu0lVwPq2QAlM1BBai4XSLHnYjtPZx/ZN56PKKbDnviZ9qv0QYAjobtxZC1il
QaetgaSkVK3Qt7fTrtKFvkeUgpmtmiQdjUuSrpwHh8p1oJLuyWVWlkwNX/mbPjUbjHDu8M6134fc
QLJZ8hUiUTJhzTZMSyyv+q4Li2bZVx9+dNxzHiDMyLm/DhEoFuvZP3xC/IPzmKnGdGhR9j7oCbAb
Iygo2V+lOh+Gw8DaxzRUXsIEiT2fewfhLwLPQF9JhF50uDwc2yIzJWOOP5jvQjhjP8ZoeulLAN9d
RbJ6x6eq48Yj31K6BfbXzD2wUO9z/l8hyIQ0wq7rSgfgPuZZuxFv27ChkVACn2MeJPw349lYASGk
FZ2gzPrvYKBN12YsCP9xSqdMMC9Dq7Mqc3Z5H00jHfvFl5ChTyyMPZAQRyOFaL25RgVjag1h2n6/
NTqqq/bdKbODWcAERkDu4XDZncD9b9irShbrr+kLKlrDVffP+yP3yMoUDQSjYsRWb/xTjvfMqYnf
wDIF2tVQuuFO/kGlsmA3gKlZvOsx8nmruZoxlmfv3IV3yn//egxnNzwHChyARmfgcv3rRPLdemfi
QiyQbBMMSZQsxT5vW0U4eY3dWZPt3rBk2TEHnYEUYBoq4GEFVMUgszAICY0BIbFHBwBkpTG1nGvD
pEFNXObkEbvvu2wilA2pvX4NPiEwENZ+dZAd6q/7d1XWroaS7KaQW6/uxfywXbOZhHAZr5gGy8XU
SkhCx7mTPskoDEqvoVi44PhagM1ktk1R1exMxh6366ITEXDsygpMR83qy+QK2igxX8j9hjIgLxK9
gU4+uBzuRH/dRZpSjA5hokXubNFx6q+P2evJ8uTpnB8Wd5XF9PyAY7L3pazS7cFxgyZ2dG/Eses9
m5OzaNe3KQ1TdCnSNKCuwiQxjxgnfw2iz47Pz7oqtwsGeADERg3MwPfFqu/2vy3qGh/G40S1xMyd
DpBMziY4FEMvCgmk8hQswNLUF+CdwLLuCdDF8vWs32oBTamVvST/XY0tOp+gpCd2OxUz+W8TKZrT
tkVVBe3XmomkFneQSp7o5YTt6urndBTkynPRsB4vw7axkq+6MwFd6AAuvSFa57/dH/yJWp2Xu1Uw
vHE8NhdXw4lQg1gcmwt5UeMw6SooHtIROWVpDTc8sm+MbXw3vvL0HcauwMKtamSEWJXAOGH7UN3G
Dfpq2Wuel90vMpPgn1rNhdxJ1gVdGa02auxiEEvcRWx1hTK8KVxJAGrYbPN+FMHIl71QGeAMSEJp
PhTTtMQzZIKZLQcQbpxaUogVKZD6uXaG3qaT/SneNw82pDYMQmQ4wIaC5TYxCPZgvF8S9dPj0igj
y+IOqePxouApOsxgbiRh5FwaRT3LbVuF8FxgdZIhsz4csHY7YfL88lc3wyFrw5L/y1+SmRxa/+ES
c7QzhnglCxcXH67cAgwx9i1sDmSnZLtlDPvHlMWxIibAgxJnx8C7/ZBClPR1JPLS80QfCMDJLoY3
y3uUlh2HmDqDOB4B1z1CyTkEMNfKjvA+ERwPp/VuSz2FK8c0iCbSo7TSaaGR4WMDt7DNuCB7/SeF
WctXwGG+U4Q03Pe+74s3tJJqckSSGtwNumcTHQidl50ae49VzD8G31Ff+4AJBA9dbGEELTihMdi8
oq/SwHI25ycGe5+/05BtU9484yzUpfd0tfaBQuNZX2E9mO2nwhorpa8FcHC5N30IDu0Ow3dvx16n
7cAPZkzkJDQQs4W26Z1GkiK78acDpIN1YHNorFBJJi1dtypjMRgVCxiNtFq1H1b8eMcAdIJrSMfN
2Lt57EGoBEJEcDsgefJgGz/u6uNjzQ4u60u0cVHgJQOYims24A0P6CQJywBdH/6OP6Pto6vS0wWK
uCfW95DFnsCiokkPCtOdPDjKFMqTbPUtdYQ8Ewmey66P8YlMpD0oQqW/+AcyM3Tp94Q/rRtH6baZ
vcDAq8WfIHEpkcPpPwBCaJb4KIXOZys20vR1ZTDKCXyOQqCnCcPVVvk4elzvdetaXXiMkO+I6POX
jBInAoTNy2Q6uYDe0KCctOV9d0ukbTRV4WTZQLwcVdazuTbtHjeAcSr/SE628qka26N+XudkZX/p
S4sQJucarD+xywgoUMhKsXi8xWhr4aDxu84Ex0kQVKSspaOvUdXNzRyh5f/3KTZBtSzXyUUYmaNJ
0TIn7IHQji0q55SsPe6VYjTlhCSvt7hoU3w16k4//QMwDaS/l1ruFCjeM5rt4VPSGxiySt3YjFjE
cVPHJPbQXAxBfgkCBaP5eROmSvrwJNDNwrD+zttsQ8E8g9BFXptIHQOiEhH77UkmCn+nHJsSPMJQ
ztL+5PWP1epiwRcS0xRv8GmlgxjZSwnVbx7PLO9nn3VNiwHhssICKu4tbSBDn1/dAihJPRaEsdj8
2z1BRgDbr4vDxGc3SjVBABkGt4EVv9Uayd+ENecQLhGg6UTxRKLOk6YRqTZJFPXuntwYfs3lZSV2
m0yirueVbqvgOfzvpyMRL/cQPYyrwFuc/enAo7qss+HBpDk7nv1thzJ+7u1PXbHR/kcnRHDNBGfz
hFLpOeDGeGsiaj1lIGa8ltuBTC2qjPT+aP/VXOW/oZgw5LX0fyqu4Wk1n1cEv4oZ2fzj9CUDlnYZ
e/jIF8ICnyoSIBhJM2h2E3pyk2PCxvuPxMLqS/XfJMmY4mVfX8RMxQvWxn31UUKepNuPTF4LE5EA
aLloTtpGLxbSfXx8xquttXsT/ZH3r4oh0arta6+cOYRGoI0m0/smwcDM6jEQyFtu3oyjcpD3/b/g
Ae7ys/XXXhjSz2/nour/E5zipwLXpAZkaqPJFFo2oLuvIw3o9BkSafnRfrL8z/aDtgrySm+0N7Fu
0eaFgfnDkD4abZf9wRhDls6haFXvLRSsGyTHKx7VgBf0VT56I4JqRcA76k+7Ukzeie+WmeZLKGl4
zlxlAR+TtD7EpshmYjtwSWSmj03vjAq3sHdX2RKfUqLaEpSMhN8HtziI3Hk+YdH4VeT068Wl8a6+
XWGiSc/NfB8dLeEbIZw6q9sdtAOfnCts5AnwoIHNyTfmmsfQoxUOijcSR0tKm17Cq3m3pg842/2W
I1mtUf7ysj71JOyWJPTxQqVgMiIkX60b+GngbiathkjgAZyzycmtgospRGBEaILTYio74/xe5SUB
oIo6162SyqPXG/CsCML6eNVEPSI7s8is64cGsKGvyCWv3kmWdF2dUqLzdQ1gvOzy1nkD1DajRus1
btMrPysPIopv6FgKfsEp/IsVwyfsJp+YUqmsyWSE/MOkPjoiMidT8nRN1BVop78wLUuJWZIETtUu
xDOjczLwaW/bnpLpS7zEjvJq1hdloE9i9Io4gJBvm96NqamJkzVVs7u8mYdcFyhoPjgThgWUmKpY
cmZ5klErb1IWnqNw/jNVPM2TtbkPCPc6BtPOcbsSzHII5EpjpJFq0yx7dUcjE7hm0eu4epsUgEHn
m3BaIJON126tUUfpcAPdkIWxbG//7XkYl/uBSzwO8tDxtuhqqm9tDrMmA47jF9CAaTulT0ntRvWV
aimN4scN9r5OSnjHFeJ2z9pnUkYoj5bfrE1/XI61yj4ODVTBEBZS+UKouOu2+UitJfakKrwP0JOi
6FZLoyd7+BVPnM9W4sHSgM7k947bAiowQTCF9vcbSMF7yZRcCq+EUujV32K4ss4gSrvk8W3A8S/l
po6XOyGVutkmSoOdIwferM/ooui0hogm2Twa3s8qL4CsXgG6f/QMJsaUFLzeUVDoXvjrIYvZ9DZK
q6lKtqCXRpWGrvTZJbKiZG/IbZOATe2D/kdAD8ot+oSSN4Tgl9Bezmve4IpNJgH8MNw5N+XrZWc4
L3dP2kxeTwFa2ljHLAPAdvkvWrlPRDl6OWuFyGxqioQR76/Ix3RluEsqqfTPUX744lCcj0wG/KOQ
+q/DR6GFUiNcxEyue9xvmLQrhC+2y3IiEQmehqMSVz23zNm13wMvOAav9inCixAhrmiLaEV/khG/
BuDneWoy5gi5JwGU7q1e9vA4BBkDrYQ0bfNoxomuNXyO4C9NLM130mhgOOCEDSuMa7bTUpzlihbg
NhAuigV4mGJeoSRaleBnowPsDCExbWBPabbf3K/7Zddcc2un8NIo8OirT6FZF9XmwD/c8eX4Exin
YpHB7Dxrj/LNqr4k7C0dGtbmb3CycNluQakmA0LtUcSA5R0QKNMSfb/SuRnSDvICzekU6kZWZTfj
mWO0T6DlJs185L9ovKTN6/HSTATRlnGVIYEPY8BG3BarpwwR+k95e+IXG75UlWfmsEzNwX8jFApJ
ZAl1rWiyAq78EhDsqPi6/9QoD6MpCEJvQ11WKe6/BBc0oGSrp/SI6v1fuou2nli/WsGT6J9oAcG5
P5xPl1BlfNqOWbO/uYEvXDmajNEEcCwP8lUWB+k1xfTHRypm1icqp2LiZb3yznUsIEvfADVYq/mW
KaUXpUcbAYohs+fRJzhhwRTL9RaGIxX1K9MDkokSeERrkK4UNXvMzvUZC5liMOeVGbaTt8o3pTAR
4/5+sKPEltWJn7FyFb5gzkOETVM/oVWWDg4iigIKRGfKnMH/ognbHYoPtN4BC9EOmnKhfXgPu+GB
XhCEL3OU9ecDRYG2/bXl/mlF/N3JBF3SV/Z9YtUjiv7190mEmIaX3Q1grJYrPOOmq9OXxQCC31Z2
gTbI3yxFSqNL8m4+9SFC7ZLZP+ZnwTAyg2jV4v+PSpNyMxv3mEx9m0+mxxvwQiGRWYXaiYXT14gT
EVTNLtRVfx3+sDaMpww6veo8jK6yMtO0ir0nKi7D9fhybazmGM4q3KE/TI9QX7aWURxy5cAAV5dS
UirgLB6WFq/8pDhBXuInasrqZLQTfnZEMvacQj349ie6DuwqMENf0PT0Q9W/W/CSXe97dWufcKyn
laoM+MP6ezFamJX8A5evSkoEOUST4zal/O0wFmvpQ3XIhSBkgda5ZnLnvVLszFNIWzIgFkjPPpkU
tz5tMGHS9ILQenaHTqH/ScIpdhC0h/R6iAK3d0ugzAKda38P7x3nRXV7HCCZYGWje+jgxxqtmot4
mTb5JNpI3+ZZY9Bym+3RN1TLk6RIj22MFTZKaNB2+31LmOa5DpnTRSzlNpTtBI/KzsIQ1HXYzw3v
zAQT7TFsOw/beAMB5RgRqYHp9SC5xkUQYgR6YSa5QtUqgz5AUTbnOwveIVeZyNbc4AavopdfXvIo
d5uUsOR4Q7qMoV5d/71kptHn3fl+K+I3j8poE9tUJNv7+pL9tSC0yQV8VKUO1FbdmIQ97lSQCwrA
x+2u2bhcuMXkjc1dzy7kEvkDGGHgPa32VLDF3u4aervzUQfKJ7fN0a29OFMnYkkF6lri93s3Eemj
5b4ME7nhOf+x1IHqXcmUM/XVQsKZ3Ldegtrkum8+GgsrPXyCmiVVnvIje6BjnF1fRJ/XUPxdIVFl
NW2DiBGHde6uUs9UYm61ZQzrH+y3KsiPzvxlwN/xDb2XuTT3xS4B7asU6t0u/ZaesjkQI4pgFrfD
jBSeuxXjxUXX+mfR0RYM0LBrmelKazIj9wY6B6rpSpEX5Sw/V+y++bqJ0P3rTVGmujX76Ec5JeH7
kMnF54Q110pXqB18XAgLVQpNHsDltGsBBSsGasMoOwoXPUU0f9TdrgKMnlPEkD+QgZrujfkqADVw
UosbLxZz5hyjI8oDgZEh0TIVP2sSvJpbpK3cpip/fZAyZmbDzMUAtEY3B1yx1g1UB+yWtXqR7Y7U
bxht268+pZ1HSrKorkIXqbGO/eZHTIvqAKxkrE1X2yhPznj52sjaeBbT5VwiR/ejGGi/XJra5kh+
YVZ9dHFa7RRn66uXqgQuBy6Rt0IN88QyJDPDLeUzEuiXoT6rP2QgtY4lMwlBGo0O/aZ72dLJTdhm
XFTzIH6anmZ0ToGgq667pzEXw2HLyQjEdPZ8mHNPK2d8zozb45OUqdkDWO627jTDBB+FQcxDz7xX
eQh5tsYJxtsodNYTKquwrlUHntGXSlouiSvXZb0aKOLpu/NmQWgF+Cu2Df08rCqa23+IDX4xsz3h
77ceUnvX/HaIX3edRrRNBUuDsjq6EdnMhYdpCsyEY0wFPEok3I5rQ8zNwEEkjqWYerp38UzSLQeM
KyK2aDLNgvEMdfrZHsGq+IOJHTi06Asei82/aSZ4NtcJYNsEaa6TnjWCwyJybLEYPznvRUUv/PiY
JVcTQ7rsmixTdyOjkRgkruprc2fW/SbYK6TKAsakFzkPuR05cO256tTdLFNJWt4HG794H9qbU6lO
caymqDKPF3+vE3xzZa051r45q6KvS4rwehdW9ev1fNTT4ji3MKT4B20rvC0zTI4bCo+tHLvXoAe0
jcTBvvjvg/bZZ6O9EMXuuJhRBB+gOW6EPeciQEiZ/kV31rN55Bq2FylzCzBqtg2+7dD3Vp0iAgBk
bcrSM22usG/wDoFXMR1yME1oxxqFRRPlTXr9IxwkRfxf0PWYOBZxV6HQmdXy5X7fmR56D+gZ2jNq
FXAi7emaLxfe6phi6uef1ghDCQz6a26cIL3OroahPE1twEa7zyotwoo+SGIvK7o5kxx2S/a1oqln
tJhakAAqsJVFZFbUPhPfCUA1H/I5NAc/EROZxycOe15svbRPrWq4PjnlU5oKd2FNfJBM8ahd2X3y
AXUWrknGwkxUuvWdFasW9mAGm3A3Ws/N5l358qXfNy/42jqdHY+SfzdDGfnwrkN4xb2WajK03t3X
Fe57TADH/QPS/0/Et1nB6mAFT5qwEFjT9NTaZmnZYhP7Gz8KtFpqkn67tOW9w9PevwlqMh0ZOmG2
HUSG3Ag9QMrDJYwmok/Qja8rMa/2l1SFTzJugieS1ynp+NIYOoHo+9VRyGMq0ImziJF/G6xb3J95
4DusXFa4Qmh05JgPUUxetGgmSz5Q0j/dM844qoQsOdsRk0+XxcNk3bvKy38CbpMktwD2+66reLvF
q0IRLYzfatvCqMF7wMxys6BzHvk079lbgE3DUYsdFAqVyANSaBfHADLi/Abo+WRH6/6JyWHAvlvi
kBxRHUJYUy/i14xbWJTbkzUOKYBXNRqT31yz8M7LBiXTWgZhz8A4lF35mE7T9y6hYWDZ6xDJs8A7
DgEpmJFUs2nWpAI2qEjXZvoMzVw2ZEV+LA1AwQqIUoCDlMSxzRxBT2iRiRbAr145AA12B5ltnxns
nWph5B4KUL+qRB22urfRuazRsw2tL3pSlJLJjt6lUfSVK75uDLRtbv6FO90f/HaQPvx03chFiYTm
aNEoxAujJm4e2SJ94A465qpC0wlsL8e/XzQv6HA8XgpH0qjWSlZ2mdgJCbo/gfzb6mcGu10atJ0p
1QkZcxDr3n9BYIliPqVlC3aqZLdfHmQXQDMd/VH/9zizI/AFnNgZeh8tv6GMXoRgy7XTgqVqT1g6
9HTgWTpW6wypCBgtTVp5HxU53C6ifmhilW55KEIL3JB2b8FB4ENomJOJD/um6NYJxK89ier1Jx0+
jMUoyugeiIbgbD5FuobK8Xr03WWYQWJaZGPKaYqnYL1hLk0Hfbn9Vabz1oBZZiZzV5SNxfAAWuOk
rz69p9nu+1gu4sYDaa5y8iGjp/LLO7UZyhwAhGLVfvqj2FCnCx2KM+YjrVTwfVBfV6kHjfE7qIL0
Yqp8TlNnAH9VIuLAy9pGTba62H87N/6ExRFM8b5+NsHhu79Dh0HPXiEGuXDuVU9/Ps5FY28qLNPG
ZOoBldQDGChO0aBUjG6qS3/QVnqwo4r+2tRLilrzgleV9H/5CbML9vbG+x0m0XbtEJeO5Shc1kVU
7OuGIJ+Npvt440S5OA4d8TJBuOtSv2lQ68eduU5dOuNQuS/TRm7R1w3cpOpFlh7FgmG9WUiu248O
lijy654hNJIytYwov6cGvtUNU+rboDR941cXtf1rS0xlBHCK39WDfzp96Ph9ERd78LEXJBDMSvhm
ydk4u15eTVHH+zKSGsHmSDCkmcwyrNVmag40ob0Z0jWlx2bZrB+FHo2fcYUPMTlj9cLG1qJEsVtf
7u21PKS8T8MGpxqZnPwDY50nASV3uHxXlFsZNcMXa47TR0AP/4DoYkb4tE/Nb+CJA4G92wdME7y1
abcam9AmxyoviRri4F8PNv7mA6GwxfExyv/qw3cVhfZPbV/5Gjiy6WcYlN3tXPm9io+MRK9+f0aq
01wYFY2P3GGltUbr7HYMojlX8DD6/N86z9GHM4+HWj5He6PzCCZX8ASanUVr2wF1nWlLcNynQ94C
0nh4r7sCqiabLR5ATG+yF1MhPztS3pQyK1eeuJkJ350VwzFNPln205YZY5kEwa5D25EjipoOsNv3
aA71f5autMfAz35nMQ4p/d2zZfYMS187ZxqIRBkDUKRcovdDUjnmt1Hia48xM1NDr6u2c2pi2qoa
F/q3euTlPVk0JO69tkizo8NQQZcCqVor9TtrpgM6kNG1NZEW5j2RvKd5GFdo6UD3+gSLg4xsugSM
unvZxaSAYe3bvFg3at+4caZaOffUX2UEPpfzw6kSZAXKpYJSEqt40RJ+AzODnAVvOqMEc09134sX
1yWpqOOb6mgMyJpoTxgre1FgsJSYtFDcFjcfLLx5IpDx31CV6Xl7viNJOSDbTUinFK1XrwXRPPr3
ph4H4FItUitpaR3CfI5MhLkX63LG8PjMv3518/D0Bo2m1Ok+N4O+Anp/Ox2qCOnzK7H/bc6QX9XD
nQD0P1tKppFliT+1w5sqBMhSb7CCFLcSlmn/WeKFxF/N+kQElKm/hi/TO6zoSiVkUv402EwXNPJT
3QgIPBED1v9Fi39SNQbCbLPlptMhplx1ArIKOuOpwCM/cLVchq42O5HJixV3RX87om4mh2c9iwHS
tq+atMEiPaHgU/+Y/uA56vQL6kFU68EVdqTfVGDFOQlLBOi49HDsVegOKYaxAqTCmE7qvvTeqBsL
t0zpdo9iOYZYqiwzA4AaQkfGT3Scyzu5MqsdLPQw12YJsB/tABWGkbWe+r39gDTWZaA8UPyWp9td
Wz1jtJVH+O6jo6nCv6AGIoTrlZfgtlTgs78VG25fOcrY6NlSCtQAU52bBWpovfj1sELivbBYvBEE
A9y51OVu4KqjgZP4V6LMKUij/QrT0GXjMVoB4V56K2jy3lcnnvuPKW7KYeBxwjw92xKRloDR2FxV
rOlZCcIo7MLuPCbDg65NFm6CO2iPYRs2dttfQsB7wbgl+PybVA/9MkD6gaA8Q44PevgaG5xUyNTp
33BSeWgVJXFFVm+vKiY28x1BWCM6C8XeMVBF7susAHu6nIKtQBgmrSdxV7W1gwHHn0tmO9lkY8Dk
B10m81APqFke9yACuF2RIcYNv86VAvzYWQ/ECRzjvmwCnNKoDihwGYQyYFGi+HLJG6vQvFNedwBL
RutduYgdm4ahShsVkIo7BmQBTwulZyM89XPDjsWojnIZvse6kJp/hcw+pTWAGX8Ioic+8zpEur/A
+pJLnNQMWTDk1Cvuy7cmyYiQ6MzkUSkrnaZEIP0bX11E+VcTIBR2ZOu5J40ZATn02X6zWnVmkRDs
U0mVm6o9GqtEHFuEVmDmNLcBX2G711Cf/ZoZh/sQPpjrVBbQ+Ii6PcsEch0sJvlb0C3YxpPBZCaV
RUhUlXDdOHznC6BBugWUXhhYBZGXsSgC8u6Caj4nD1lYeqceORiFLdrZdheqf36E/P/ZftQcvMnN
sJMs3HTtgEmqSM5YVcjAEToqt4Vu74Wbo21J/TPHZZLqdNgoYntbBHH4jpbI1jhjwjQ8GhXjTuZd
N6e44Q1Su8WfhrMEscT7KW0/ni5E1pfmdBsEdWF5DcTx9CWocH7MFdSD4xvAxZwYtsDrVoNkoT8P
+6rpsScpHBRXo+6McRbLktyHpG/cJr0vGLRviHhR2u2n0XyxdY/XVdQgx/52e7fiOhz41KivhfPK
j2rjBOoMIxrhuxF2itqzun9CK7hVU8CanS7h/KhJ//t6z9tZVtvRepBzCUwGP0Ox6FhX8IR+yg2Z
8jcGt+fm9zoZ5T5+OIKp9zinmPlj18ol7ZdNFJidxXN30MtFapd/VoEeJu1tjBXhkghlvwtFf95v
EZoNKJZ8RSqsQlo3mfMD19/fmq/6xlZth85ufKBhNscFTrl+yJGYDk0WRublLP2OthcG9l9PGrCd
uJto6ehwkqp5PAXUMWFZEnd35ygPQ/86AOqttUX4ZVV6jRvuZgP1E93DoVQptW+Y5d1lm0Uv3Nn9
E6F9UYpb3i3m3kn4PHW91svDGgqzbXyj96RLdFif8smD6BMStttWT7jlF+AUkoYYGijJSCDFnWGT
hcBuXVyXgukJt4+HAQ1DL70kxuShykSNeUmuRH3qgpviyrbLcppwTF3D0zl6fltD8c8+ASE4JP8F
9nfkUsb3/ZPnEL/9M8dPBWmEAl3gRR1rQ/fqSlD9PWqJxcZtkbtRLwBxkzYm1ot9G5TGzZ7NZzXN
hvauUrtJDrtbVPLX3xgJe7GWWdYkNfLn8FEdJCoyJQ89bDbkt4VmQyX1eTpvdOR5AZkCBoQe/mRD
HoW+yLN9AT/P08beEgG/DKHWC+eKEYm1lkG5hJ+ZiWwXwK2e7Hoc+ppWv7isaqI5+Uc8tdDz5w6p
0Wp2UpzaFS0Ui6f51EtN4Q+B4x0TqwGoKJMPdbRUJF1mhiLf9SzgAOKYjmqaO+bj45JFYwN1/TFD
rK7EGZl0nhDzFvoBwDMvCx8E6qCCKpf9Hi3Xq7TWhObEdIxaMB4Ks5Xj7iOF2scNkMbxmH4zm4vO
dG/zf1ocgEAK3Lpz3h4SeR6SXU4UCinlgHgBW7yqFSqNSGkzZvasZXiS3XLzbKWmQsbLgepQGf25
MMpVmSPbhSvD/fuL95sHPwfByh8l+BzWS9R43Bot/L2gqIfzGr1bURClSF+4bA/MIM4y/uKm4Pt4
YsYVWllUj5JiK4duZAnlEP/Vo//lK3y7qGaVFWtwYd4P4ccJTVY7qnBYqswQfm9dGpOUU+dJeIHz
fSWbqsWr6OZ9EysKB8pBcDTFiOF/HTf9TB/XByHKJNBzxHoW/2EV4kYVmJ9THEIUPLpiZo6RKaQT
dx6kkbor3B77jwIquKTfzGK80TAwSsXa0xaerod1sbdPrGrMbc2kI03UACwp766NgnJLAPeHdtw7
w5P2bcwNqQrePwuXvYjwa/tKCWkVJ4lksdDGJUGPx/KsbB5T/b5xAy2bniVY6IaY8ir9G3PEc5zR
kuEk/3u4WZHaBeByorEssPtbbP+ekB2jHBVIG3jwugeDYQ2uLI4bXnjgFF8UMtLGJyx9HgQt2dGA
9/TL/FDsZfONPORkRi6tzbt7PhNN+Iptt/UmuPsT2oE3zlhDDGGe4pZWP0/bnZ9Ji011qZQu33O0
6Xi0/CUqhkl7ErcR69jdVzv/GIcxQ7vt1Yy+FYX5ksgyUoprMYFcLTSfc75iqHinUTVlj40h9qTD
B1sZgXRS4k1PoFaPFjrNrneuFh9CPuBoEvDHygYfa4zANFvVF6KZCjxozR92pL+RVlBxUkBIY6fO
SegjHGalbmDmH5Yo5UQEeSKdUFDUANytzMTUBprd5OjyY8c4a4LPYDZpLIGYnaB0lQaymorNB5q5
mnsTM9d9gdpTnyQGeEqPCqmrrgbBVc0kdAPDpRoato7oQtU7/g2HZv6pGdCdEid9hie+w8zRRegj
fd4/3kPqIqW9pKCAwtzKL24GRAFgREw3oqi0sCxBA7VyjqIaiIJNzol1yPLwKmQRqGabFiFTQ7r0
aoeC5t8mejTdW3DeHd3K+b1VB2xIRlaLddDdjtDhLZddTaTzSR4ts/XryPpsYCGsdcdKj10xs4EO
GC5h03oHUsmkCnCjsgqgsqsfOKJiochhw82F8SKMSgJCPpTsoCxFiCcFZUE57iKFgwpuEWYVj3c6
4GPHnbUjFDQYfFzG80gL0GjXsZJ1UNo7G9SzweICFpZ32wQZuCPtLiGNZbqc0ZEPywsQ+1+v7M22
3tYcURH2RA8yp0H0LvZoyqJ9+HfNgbXsylN9uskHLtUziwEK/QhPvXzXA5AcGjgCWc2GzStxLAhC
0z2LNr7RU3gheYnuXDr4BODxjGMhQ98sduewlm307K/lWaFX+86/Yh6iWrUU+dKX4WFEIWBdbhuC
tjiZtuzOuT7n82ERY+7Xe400dsSVHDaMG7pFYuhS773UlI9ccKGID5rbrIVqDCSCbviJvVyYe01z
wCKq0q4SaR4EE2LgAinFA0Y6TL4qOWQOsLHG81RSrCCPlfY3/U2LQHXHWWFvxMQZyXlZSSi35VTz
BVhA8gtAROv6Q8+V4Rq+4HmQY0cfCH3bsd0rgQ2jh4dqDPtLv21oGHc513FzpLjMVArLGSvoQWng
qqEZOXWsXumV+2ACN8u0kl19L7j6dbB1aF2pNw1e5ABx4OkLLgNnJdcrgiCHRea8Jfr2eB+Q0JvA
yDjeds/aWTfc42zINwPvievq/NdO6YVUFQFtGu7RuOH/ifxGQ7bG234RHD9/PSd5txfENGY2B1oO
Far5LKhsxefxuyt3YDUii2Ub+M0tswwVrvGMwdGcNLV2z9dAhUYTd3IDPk7R5QvGM1b/jc37X+Lv
+2+cegnwibHnSMC0Tuves9cVrbL4BlEZeqgU+CYWOdqZJE98PdnN85XMRkY6xY0rBXV9KBTHQQks
GNxXyTxmBUvZQ+o2nvj8FPJe/HzSEt5IzKr0+IbShZNOL/1mQZQGj9sNLP+T0hUSc1NP+xknk0b/
PzIuP8Csa9ONtxXvzP4E08OSY+l8v2ZTJcQk+mlFXeXi72XZcwjXQwNsmrNjfnLiXhPntyo2li/1
jY4dTPbLTV/R1RXvllF2LfT3Jzl5NZKmdmoQOVOAcFhdF86ZhjERB3+4YuPCkUYYNUiHBmKiaE1O
c9VODx1lS0ufkfnoqWKNzg3oW+VxqYU3G3YCHlEROUtBwui3+0ZXZRWJdYyv4w3NSCXIQstTFcTK
eIx4pUH7vETYOsLA2gdsg0OulmNl+s988OQmiKJ5QGkRnOKt5LlTaAeS9YCEFBempPJcDRplflfQ
lIT1qmvHDVcoITDqJexYfPjkV8QbQGXEH3Ek75qhyXa6VtnkIKrT1ZE0ho+xzH6SKzR8ihifjq6j
0SZhsb4RzHyds92AaZI+4qbRONIV8mkYNwCCPX7VBs6LuFst2IVWgcAOgC6jbOx0yaSjk2VkgG0E
GBbva15pY7HhX9cEMgsFEuNXG5CD2SzmXjetBD5DrxYcVx4XDcnb4pbI6fW+J7gtVIbLIhIKsfyZ
MC1VyZ1CfJS2QvGbQGWoo311RNMI2ngqmpyav+8QSln80sjwV3Qki7ChO23erW0wbVGWFX+HweQ8
D+uN3iAFB4ujz0pXM4IXV+xKvk6dnkWIqpS5ekEAL9Sgf8ENcXUj67m4IFFUWCArjfH2Qp0eRvYl
ZBQ7ZyzwmKcO5uPkoE0SlC0p2csq1zZMtgKbVzbxeLYm0/+FDHE4HOcFfS9Nrq9WrowQ4+JRIFUD
snQUQkVGbkZ/D6ddhz5KyeSCFXggUScp5jHWKs87g90NuCYZE1SY0ge6Ifw4uiHtlbxre+4WoA8d
/Qw/tOFDsel3zFHhBAhxut3YVwVHtdi4gU9vjpDOFiHH55HsYlEB39k8u8/8MO7GRlXbTmO2ZJNu
eVeIMAaep1QDaDRTZpROhQDc6XLfgwrbLtvrnT0F+VTaZ3119P1npfte93vIyOCS7D/T/1+aEnon
Mf/joXdpoBMHYf0AVe0Z1kyOObibw0qUX9pMSnL2X+6VhWFeDdBn9tY1zfZla8u1IQ438vcCcGDa
5DAnNL+dRTmkqFOwJK8uMm3/EXV7cNGguZuwIx4hSw2IGGimug59OFOsrfEwsmZbE43Q/LigQGXL
95bWlLi00ICV5nGGsJ4kAZYrcnF42jWL0XXJVqPnKEDzODkcfv7Y3XszJkZXGr2M+P3LHDs3GIqI
Q4UvN1A3EmsmMr70Ij8S3mFnJ8tIOHOai24xAGrJT0bb/zzEB55PfqLJjqjIKqA4kcr7tnRnGkG7
4AKjRI9S8D/nmSHPYOTZyvaqbjNYWL/xLKZWstTGATRaYVTrBTPSVMcAp2HvTAOryksd+94C+mIk
94boziOVkvW43s5dcdkloX8KSzIrCkijJKrrZFFnl7jDe/4LOcZDXFsGz7W+2IUMNDk8pS7tleJ3
mwJUs3fqt622J/n0/rcYIHhhinKPrHoRFvSFdGNAzNhdhZcf/1K55PL6AfcBGeL/LyB9vO11ZC2U
+1vnV10LrfRn8xIrkBLU0gFQL8Ia9nNuO54tFMY3hIvqMsERTgtoqLRUGyd+XYYAtCpwAs6RjB3j
m2/mw55vvU2CUMidPMLpaCpeyBbnTe8Y4i4e/nrC+FoAYjjbzZTrdB5A4RDdGuvPVJ+LdwM94UWn
nV456k3+muDMxMnuSdqaENUqxiE6OsFy0pFz3hKSL5LbYs1MJ79+aN7IzsaMM+0S9UjctUKmXrxH
PxA79RdfMKCp3V0tgi9KdduMz09C2N5+vnJ/1BpSOviyYmn6ows0LigbpFnfv+4nZ1c/fNn2wsRF
7GJtxu0mZghss3lkoDv2p5Vi89+HaOCf6cv72wrGz0YMKtXfmEtPluPFkxEAll+b/RdTTXrzvD+R
jYONbF8bpmQLk/hT9h1Ct7YM6hsk+bvIkedRq8zQ2FjmKgTRjlba2c5S9VXIX0ewmfYvelgSAsG8
Yz7FKY08a7TcHNtZzyQzc1hzRXAJaZ/9VGQ2KJVtPV/Q8ZFst/do1eQ5freR8X3bYOj9mCupaob7
TGAk14rjR5LfMECwE6iAfnGGggdKv3CgALudmIH/gxfx5dQxrVFVW9CISsPEB8c3Np6Qf3NuzVD/
nEWDi1bT+/e+Kq9XTc2E8ttKkkLc4L6turOu6h31C1uRAwncPmt00dAZznte14/AXJpJSCS1ttB+
Cuo6Ty3tMwZOBVhBGliWkFQbwYkGmeMivJFVflRaWmkjEzT7Cj3JNLlYbONjHtoAAEL82tNpn57z
Z/39SKSYgTxiw+6DzXYiFOgZ4BXqFQfNq2lgtVIXQ1uW2BFZFWceY09bh044vQHdAQvPdw2zkB2g
dbz7dMDO5SPtd5YU4ZLIS3c03ePSzC45hvgM8o1URjQvD0tVK6LaOElAEiaiKPoNncu4F/CRLGZb
Ed+a9OzStHJT4lme0Jb70DcHED8GPCjy0IQh8fa1QVlhDh5bgG/WGJvNDLuUcHgTztedJP03y91M
ElkxT0EJdfE9NG2a/ekYqJTemDY+qBLGT+HkPNkLqB+eCqmAjTzDkdRFUpK9M6VIwxVqnpSTmgRn
EftcOgqvlzzVg45gB6EeROPGht/kZsnzryx1um28aBT7LywubGI6VjfVwrIr/R+xDdACcIyS4o2F
K0rL/d7BKseIKKfjRnxiiY6jzdJiz6LzFB8/dqKIfNyK22CO8DQIkFo6/E4uKubhFo4DMmBn5tNl
Mn9+9sjFI1MtRNOBoJXFZdi7jNOjKuKvgYIf8xl1T7uzQw/1JExuE+0G6CGdhktxbxhxdRIfWtjI
2zzLvviIBVNrudbLe8p/uc+2a8U8sb03dOlSKizUtuPPit+LiDRjZTRGw0tkxTsP6j+6JCMFkbKM
wzkoCBwQsNsjItPrIWBTL/ZFASPJOze/oRt2oSx54tzom/ouGE5zosSzNr4OO2U6hOVwhx41zkUo
zgNcBf7RvOnBI3HBUHLrvl/P2aq9mvqPaBJqDQjNw3/xJLVuKSTSPqufsb4qqK2SuS3JElIL0/SO
GMSoTAleUUbrY42F2U45NjoLfAaxBbHgO13dykEosxA/XCq6E0MQevsf47a04WNciz6M9a3SRYZ0
6koprPPxSerQxT7BmDNLuVWgqqw0g1KTqrfnVztPIm1eqlGS5M0uEigRk5MvJjBDceeDcVZG5goi
hQMeTIjNDKg3WuF/1txuIng9/GvK8tvnVUX8JxaYO7Y9eb2JiZaP25XZIf5GUkdK7OJCguUjWk3E
7iSgA51QrPW9Vdrs5cx9AOm9eCID+IloT0NDhvP6p2LKYIVj6TsuknP6yOyWkGodkTjMpnyqDnHQ
j3aziMHjwjxNVaygikd0SbWveK1fezvEu6QleqheOTgjo2P/EKBjYYIHoCthc2/scG+sb0hsdz2B
oL76aBVpWts6lte2GuXm8WHy0se84kPgmZNrW6ujxz2HmpVwQdkiwrpvzkP+GaAz+xDVzLCrEKt4
8wBL6mDj10nus7xdyJpB3+kcoFaqXnSgWIRL9YbSb14kiYwLhAX0v8KaYEwQG8G3qaoxbNGi0q8V
hZkoAfryIw6o/nB3mTo7Gg3NDJPJgrj+0KlAXYl1jFc3wZ1lmGEvipJm5krkvv3uWpmfMjAbmSQl
2fN2Po99BhwVKPCCOamYFAJE34g4TCtO5JULqapQJU4dHs0/GrP2bGnr9ZNNn/XzMcvvbhTlIis2
CJmrIoynno0AYh+FiLK4MpUhPFUeIQY5CCgQAdWy7h105Wl3WmFzuPwl4/R3RmLMykdED0dQWUpj
DzcL+3WI+17J32iEPZrVeY3Ptq+1wnluAUyC2lzHKELLfVwkkCPplmkyqrNwvPRuXexzdKf1ZSA0
UAbypwOeL9xhQ3a+FDiG9dpSTAbMizor/dY2bYexMjobdAAE+x+sRPyyHKUIWNDaI4GAN/1j/0Pe
BmR6Puir3lPSKq9MmQthNpQCdsVmYYLcu7XRRXIoPBtAgx72mC4lW1R0FBvXEOT8fabTMX2m2hyI
pheWNKmcNGEvAnrVxQ8PJoCfdaAiUj4AVKMP+7W6vrE2sObfhIgfW8g+7/fBBlhCaoq1QyteOwOq
+5PKrvnma8EygCAcrp6fN+1VLVSae6yc28HHB5aqO/kjbZz66Dwd1QFuw94riH/jZZfNNErIf9bs
SIX5xM2TKtFlzDpnLsmY4lQO8ZF3EWRf8q+m70EM6xphqaL0aR/gpY+Jl6G7yBkwv2iqiy4U96mT
PW7b3WpTlNMs/XeNVq+ivHGufH2vGud7NBqceif7mRRKi6KiNTRP15C81UeQtV4uOssy1LxLfXkR
R7VX55jvx7qugWQ3+Vbq9mwuI4oO65uZ3YcpklqftUlijjOIRwF7OO+FIOylVXv6PMh7LdjuW6gv
3gKKKrH2CG8ffHZJuxGeUnFQhu4vC9YCU9Mng2DZU5BM8G5ACQW12hz9t57NhOFDveL3e2TlA/iq
WdgfAW9DZs/dS5Jo/9m6Q2ii1NQlcNniQ1usKIWmsPKEanrFuIovngJSituqlOMQLBxG1/JFpPFA
2FDMHd+Ha+IYZE1Ka6wVgJD+NYfgRNwcl0RlzOV3eb1RtJx9ODwyog0bjgS1v6eohZqFsbCgPmWo
xPI+9sAeU7iCExQA0Kxe2uUOdwpdbQkTecepBk/5Ml5O0ESs1NQ5dnc/z2a+7IGJb1FGW0OMdiza
Bk40J5hDiZW6YNZujtNePHRtWxHVr8H8C2YErzlavtE2OaJ0DgOApWvtc40uUsTkn4Acp/lE5gno
cPOGVx48yYCXZNbg0eAImJae5hFkemHG92NAatQZhnAWrJoKHzfniz+Y8jf0jdgg5POp7JbrDotD
wycOEUIaRbnYjxQtTH2QX4QcRV/wkTe6mTC+Gf7QUFtu9guCfC8SKGGnOOhUVfaaXGB/8gZ+QrG2
Lsoe1p6asvtWbyXKCBEd9fmX2vOVuzYiRkUZKRED6we38mkAk3oqt1symrvtZb6gx7Ll29R+Hwm1
fPTUmbB0D+3cSsrldriQ2L1wL3nsvQ3xsDynmycRCWWNDLq0oBObLSAi2hukU+wkk/0yQ5cyKGou
bVi3wLtSJ04zxqhsPLecyluFvWoZwHdxHrhqsntligKqpkhhKt0Bm8jeo7F2O3MkHOxxarE2/k3R
4BYvYtJMlYGvwhA/3Jz9A28HXYaNTm6fAvgxLqAM48mpK8SQfwch/X97ZraCG44OmdemY7t0K8Yh
wXLHQp3Y0KGnPCvj7j/XtYBdWgU0WAaRbZ/n/hxh6YYBiUSTXNfgCtogSR8ajFfFghY8vnWEROKT
NdrsbQ9yfCbmt1M4Phh+JOQluUxzyQhfi1bXUZi95lQ+hBR4ziiRvlWxJx0o/f7gTYpf7VeN2y5t
ykKhx0z5pP/1SzZFt6mnBmUjkE8wEktT8EVvCCmfSKuV9cLluxOM6BIvULnf7nODtOfLjplneUmp
Mz4ihz0b8zPtryOKix3536VkPPpEu8ThO/PPAuts7CU9QGjKJ6Woo+suxr88J7ksw6TXlujioqXG
BFJ7hMSDXG8fVC0l+aPTmJXiQQ+5fmiGpppP4CjIn0C2wJUTAcKodNRbdkwQbL+l4sP50Xrm6oHm
nyWFzHgF0u6fqh4N0beS67qCpQNEeBE86uV87Jsm7MKngxjVIg8aw22EVvSdY71z1GnfCk2kzBym
r9Zqr3/mY0SPItr5QMfSHwAQeO5T7rPn7RZsQIaj1gQn2q/6W4sdA6hbR02j0k30q5+lrkNaf5Zf
h7aHabgTMX0PwBTluvFVnJKYCBwFfGOdK1S1ln51LMd/b31ZaXBkOGjS0QWVMjoKm/96m8NQmUPs
62iKzhb6D5VAUgxnh562gZGIXZCtFnIt7aJytCcBTJQst7VAgfIgB/FeQluotle49hqQiADXXr2l
etfnPRHzJ4Y1YWsVoXWSPCaSVusW4GIFudahpshNiwAhki17R6MpaAxLjXtgJNS3+IQTNb8TxfJf
s8IxNrGKsCaN5lX1IiL6/RgTXuesFGabMq693tGn+LmznnS9KttS5h2vU4eo8E7n4E07Xwj91aRU
5ZAMCoB6TEy56xk1GNvHDZqmlMi32U6hHWVGwv8NhkCFTIbfHiaGK8XQtnx5TjvHGRgqnHyfFa5C
gx5SGcDqLWGQXchhd+xZjXEvg7oWJMA9U+RfAn6+PNccjM8LnBDp1BgK9SSrD0Lgsoc+g7WrWBvu
D4vENGYMWwCwAa8vYKB1XdGabsdWYpBjbDXl/m0gGs63cX3yKVmDHMowCccIO1IxOZOOYb7n7Ggi
dM3HzMLG8npgglvwvTtZ8kLxaCJdJQZ+hMRJWbTZIbAlWeFUg6NfmO7Kf+JU+i8Naf/3oLyD077m
ddz3GijMGOdTzitV2jwqsXsDQP/hC0iFL23d3W+mxR1Pbb8poOVREzqlOK+fNg8/XBPXKtALF4AV
TnFAWr3e+5M0ZiEmLARawXxl/cYPVO6Lj03YXpZre314Wa5U5UYYeH8hruoel5nVoPD+XkBgMGAB
8Ko21crMSOGXTMOaLEQhsHbKBjtj4qMVANt9eYf6OM+dT33VglHOTrFC3WeWgcw6yFKXbvLmgMhW
pgUA8gdE0zpjGWLDBPXlJa5rqgmA77IoABX06eCQI9NL6/DcqsrPYVp47Uo/bZfWOMoiQLVrD7i/
sja1w6lQVgsnr7Smmgq9mibwmld9x1ziYeKrRxncaqDz/yCekNh9WXMnC1aTXjiV2iFBdYV+3tcm
vk1UBeXb4Hkpc1UcHEJBbqMbztf/2OEBWxbcatOGy93lFbPFSUtmUY8DMtjGpjSoBRanmHdWbjoa
AHgJ96Nl5ZuzaEWWqb92jJZR5mMB1pI+SqxAUtzYU20JurGSvUXDSnKc6btJNROP9dxSEo2EO/+0
inGq3sm8Dnx787UCplI15BquKcaK5VHv+P73oSacQiGsKHWAkmf2wBnf/ee9pyrGwk3z1zW5qZQ7
v81Xm8ZW7oCdDUfbuNELerNwOMOFXm2+noR4IZpYAq4ElyW7suFiwPJDtzIvhinjjKD/2KkK+51b
vJw1Qjxes8POzM4uAX1r+8Qmyn9yWPqe8aZc1O9A4CfBCEs0OybOV4t4rR9r4tZ3w76wO+WMot21
JhTSO1JfY0GmD+qdALEKoO9Bm8DSLiTnwWdnTT/mG62kxDPE2FR0vrTsMSaj9YJSTwLTnjvb2TPw
gDjp1vvwL/8pPg9zt8qSj6rlTYIK2KpWrAk9BEjzFgPxEqZdzsKWXsHhjS+sXS3suYAvNYl3c16K
oR98VEX1BHrLVsluD5w3Ww78skKfBDibQa+f/98JQRVE32aAowtYKU5hBa8Zs8tShta++8tnYBYr
zgaeZfGBKXzipGafxjThNEc5NQ3dcyHQKDG8M4xZQW0FZ4qN7yH3atN8NMYAiDRWH4L/2GCcVGnB
zVr+2VL5xxxRM472wPFTBmGDe3fMZqB72jHmZvmY3IWQ2Ko6Nn3PUtl5LQzVJnQXnE1P1CefDO9f
uQKXCmX7TS8mnj+bsEds7Rg+e6PiGBsFBVrv/CcmdyIBdZFpzx4BxKIJw1gnEJVOwnMNHC0iBCDw
3ImJ06McjzFi6AhEjhU/XZVVmi5FaRrcQi3+HqLtiKDIcFLNd9+gAIrvpfEfjt/v3tceC7WmUJPw
jNcG84Gl/QC81JBZ5A25wAmUr3s5VwIyFUabCW11DHeW+Pg82dND7b7pCX5IygQsEF6ZrF5xus66
xMvIPKsf8zrq9jjBOGzqueCMfCmCulaXTG9SB6NeNbuxZrxZuBZlq3WEiDy1VkhXfymlVbb+iFzF
j1EYxlvzua9fh4xxDrGLTM9oLBx3ZsDJRKK5MpqnBpfZh//cmrvKt6k0Uz98f9Gc3kVX/+op1J+h
aB1olrMMFQNSxbNjAJqeochU6pi0n+2PI4qRK9MEALpnZNRzQQmIRI67inmx7ak6IuynovYq+H3x
9od5/w85/183EdNaJPhebLIStQk87Y8jj6Vqd9lEruiXu5TLwHmDFMBhZMO7Yxf+WxRwJe/KCWZ2
ZsHV7u/gAvDdvMe41whVPHmEshM6hBTa/rKh8B6Ov6mNy5S2l6AZ1u5Kb2kN7Xm02GPXrjIh+BQy
17Zw4wPonukxspHumyf8I9wLmWltH5rVhlx3NY8zgqdCJGPE5yucFvpgBBggoOlNX2jqt5WQTJY9
R0Fp/zr0gTYPcdK7+h90TI47QR7dMHDOzrOyTHV75pqmDjrykF6NTLK/M3rZt6JvtOubSDu34PXA
DhNuGHBsbfQ3IRdyRqfe3c4BIsMxbfNMwZb6cZEqXgimlOJ9YF5IGj80HzGjh4REFHEz2viAIoVi
DLWtmAKtbGZbdYw2zZp+5S/nZ+RV4DoRcnIrLdYSlD9SxZUsWaklykbdtfu4auFc221LAaj92Ovh
tAADq9vVk/dZRN+GNHA2xEkkojGt3EuwSeIDVMxUIqKPMJ6bVzm7TicBwSbrmegO6rHx+E8sZYAm
Usv4cKCVbV3+xGWaObr8uF5P3f/PHcdWThEF3ywZ/YJU4qVdK95K5Asx7IWHN4a1WdCdkEJP7byL
SBlZsBLUZBw+o+OTFDeCyBPOd3pmokotXZJwcH1fR4QuPeOxiZgHJoRHxFA3IfvVCMPGzkcL28Bh
Rsy8eYIBrGjy9V4TPDHq9X95zOLgjbT/Yoqq72aIcbzZViy/m5L5z1Mw4SmBdrYLCq00zsILAd3M
gHfvTaOiiDhmQlHCt9jt6XXTQAfSJ1kRH6h/emZR/uMskVDXm7ri2mZqoYbGyyNaJM8RStIudSJ/
HvAjsx7km4SZnqM/k+0QiW6bxdzFarHDLhquQgHf9rn4fyula7LG7Ln+V7d2Q6P7SDtZJzDgGiMc
/duNju8Q4T+pLj0gx/kje3VbTiRlAdsQwDm8/rvKw4+6b62dNw/81KQs4C55NrdRSHL0FLptSVvG
vvWrbdY8IIhJ22lgIt1sx2HEWYqg5bhodPoW8Q/2A0gNCBQ5I5u55+p7M0kHE3DrZ32UX0FRjcEA
JAbaoa+31Gut3G/Y1q5EHkg7HVDGGcWYJ2vCbtPdAGYWPKP51mCAtxSyW1/4swhvhtavuq3xyZUz
RSkAJ62D0sDJYZoz12tJElrBJu/iXSlq6Uv/TnEInZ063FgOuDr2nn5umTk5pypviPrxzFC4wl5D
2zt0Ddx/BMYCDAhZa0FhtGFd9Q6VfEP7Y2FZIwym2R6BWIbuI72rqDY9Wf/LDxgS19PyQcomQJtU
azpfCDNUuISDVy7bfN7Lr4wkCHgnjNItF/P8l789hyWWQdCYYsI93vQ9fqf1AfRGHx5Bzf0X1PEt
wxKzp4AfoB3DI3meCnnnZ2sp9VP8TeiwpoZpzSxSi8bqYF6W8ERiuwg81T7ugAdvHcOg110YrNTn
k9d32dtIlaQimeRsMoovM1Kx8mlYDc/PP7wXMRG/ORFX1t/iu5+JZ1YulMRCIe6raAdFMuegAtD5
6rK8q3kVsfIHp6iFMYVES5LpAmNYucF1Ub+0058I5EzUmhTC3QN8vPA54CL6E6LrymjitLuMu8FS
Aq5gdlNM7QroZQLkjV3QmnokS8xI6qALqv7LIaidXE5fvkZNnYacJRZFjeBus+z8zLczq+AI7kEU
/cazpv+Dnckabv9k+J6R0pmaw7mpOFdDTl1wd8AVqMZJBGaNv81QTGZWaXQ3jxloJAe6XdlFwLgz
YR6hX3uDy499beNNMHfnhjnsIP7J5BhbmYoFjtzFMjAExzoMVWwbxyk3hdUGr10GGE1Cb6tkHNOq
PPG2yHc7k1bzoIEcE5MkJ+240asDX8JggOocQ2JEQ7OIr7n+Yg93gBLSLYib/A7cQ4uFihKjL3oX
93KBHwwavB4Z9Me+xHaHPQxPIp7R9pM7foyRFywVkNmRbZG7i0J/yRJJJ2Ciekw+f99xw4Kv0LiK
A1k73ZurLtQfOROnwN6HapsAY3fufv/lbVGTWwHnfbHsVUtD47/y+AvO+J1lZt0wRZo8o4Oufv48
LpOQejGg5+wVyyvJyxsQJ1z9A6kwWIwcBEyJki37o7FppJeTpHx1p1bdQllX4bkejc0fTj/HyuZz
TGPxhyH7ikg57VFFv3L/ys7VL2qEt33sPnajqMQrgqNx1XWXtkMr0MFmLcnN5LHCzi0v3kcl/lwf
LJ52weFFT827Jpdm0cYjV3KkcQCz5pVo6gQHW+2AHkFPzpWhbIYKSOb339oneI2Lhop0duACx59x
+SGVMUIxaHNUqnMI6brbHW33ZZRfV7DT5slU4vi15JDe9J02uSSOrktz0Dc3E1jXvcdC+pxjk7l+
U2nSuUlG5DO2mNnO/+5tO1H1il9fmOl8fA4pFYTOAJmMZv6l4qsHFcVHThqViPYxs0vRWHYrj2l8
X7fByAmQ3IvUxiDQPQAgrcGJbLWFdVK9Z5kjPGvqW3VnDZuTbG3FSfmMekcM7JUGUBH+fsfvLKUw
505X+BRmZX3+1+w4AEzZyCIA3OHNH/70N/tok+3v9fwetQHqUWsLKF4jQjFzZblGQoeBD0Zdhcs+
V33c+f2Gl+ES8Y11fvxuW7mvX2x9XmxUGAj+wq+0NwhJrUJiNBurNv7g1ur7VVArMTwBPSpzdHu/
CcO79hvxEOtWK6BY6Pns1pbObaUfAWkMUh1f1srjClt+OimQONj61dKuIWYSeOzarDXya+WepfX0
3dH3aQYgquWbj6Pwtj3wIE9sdjPniU1G8Dvi8h+h12c/Cqit/Oue4xa0ldbIskwmYbBaIVL2A8QG
EOKJS3X/3dxm3h1bw2scxgWoOj8MRlwCtT6filZ5WNnfcHRkmKjaM/warqFmUe7SMnXHR+8rSJyk
IalcWO6SpHZzwlND0tj4IY0btVy/qwcFRMkiHOcu/31oMA+xAwaYuAggh9cV/MnFZGGLcP0uDkbJ
scHvKA43N9GLElk6Oj0Gfhsehwkbx3RXX4wnODOxMEvikQEgegtQRCEBsz6TmYDal6j+PE0eyXXT
VfTJBdjtw9YcT3m5SGjhzqTpxc4Yh87bTenPRyjyzmHsbv914WTPgCRF/ga0SwRrxfyqn04VWC+e
1BDAO4w84Gr6DsVvZmfs1u4Wm4C/9to6BoE+vostcWI7pNfhmTlzs0o+LSwbYOoWxIuZbhD+uORo
GMrv0UJd1QPF84gyvXvLIrstEYi8Zpkm4xdyyJwA7mD+MxxBVMievgHNyMlERwRK0K4TFtNFWFo2
XQe4ehqz2yKQDtWNGFFYynTXvVHirMiyaUyLSXk7qBU1pKMbsjMWE/OI+DDqohor3GYg9RfmLBtL
krj6sNCE072QIxSKFJcH6+PWbw+RT0/jICWrG6zyk2d72XpMEoG6rIgso6XI9NG6nxXDqvaIVtn5
j7UhVctu7pmIiS0ddAnHUyFjexwFpQoiOUSzC8M7LhGqARRUhN9A9pGe0XX56Iu2cMQ/ZvmaNhd9
AAjfWRZYkfiOMTKcq5A64QQieHFS8mkoSyFXWPbp0nQ340uuxXBaldnGnBOpWmCWeBfisuidmd1/
D4xMp1tcz2AyTOG+yNjjC30syKV7lR/pD8bAIv3IHPYvYcMHVpFE3bxv/NPMktKEQUbE3KqXblaW
Ub8h+yF5Y7W5U7TtSdgfdQfXeuBJet/bX2NCsQJs00/r0eRmSoa/LgzETEQiijEyHTHEzoa3jSqx
mkDb58eeborI6Ja59arzG9ZsSdlyNBN6XOwNVDbqIs39Vd7mKSV8ktDgDV+JPZhCAjTKF0poJJ+G
7oAZZ2VtF/MArV2H5jsgylxx6/Hsy+6Arofyx+v2/wJmwVRP4Qly0LuQJcbBDCDjLcC5zQ27/lZ9
WR3nH5+Tf5FIMZ7IgnyBiQMnhn3hUzF8tSd0sfmD2bKNmEv3xHg5XjZN1NHNItb2TVV/Ew8ZFY2N
LfH7CJsp5wbi0+o+1ofpQk8gBVVEtMURIxKyxNmV77rDTYmRv8mU6MPMQaTViEWo3jKXbhCtxzx1
U/wK0C21+J1iD9gFbvXqgKcscHkaL+9ECK6YmUHa6ZDnJHMYu7c4kpgA35TgNaoAHfPlz1w1wy0h
rYAa2CxH2qJMh8rZP1nhQMO/ZCP0F4tljQsZ2QK59NgsRG6BzR7QBrBJ9um8d9NkCiDqekTffi67
70t7CcGNIFh4A0Ys1RnP2bwPuH27ysKQz3GlUf1rljg/vzCplabYVs4cN+W8r69oQVuUxScsTuxj
pwOahLgi7mMEYFzTeXcYSmBQDrdI5RoyXlbCqk6AqF4lehY+OBp88xR+zOxUlSPZb/+B27G2swsd
pjgPkTN0BCQfjzxP6iHqCNzPYIrpuDyPJ4UBMFXXVbpV6HNqAZPA76ti3uNvdsgsGlq+YJQzqt+O
SdKK8IuBq8nbsiuJxrh7xk38toW2LMX5rn/odcnBcDp7v2K8jkxjI/t1hhZ9zAd85efs/Zw8Z13k
15af7Q4w/Bo5TmKnEqYZWRXFjySCALPwhHx5MxrVCjXQkZnCfVrO7yfsnPWZzNKPqiqu71CjzO24
YBJsxApcB6cQ2Vu1bRipikZUdLeZJq1khcM0PYfqaVTSUi4QdMSfHEnz2oLVS9cQVJVOB1hpEiKS
teNsUDYZQGEEHCZS6JPJ4pLYjUBK4WYY3K9zbZM5PQurG/RrsiiWif/ADmmVVJEhpavzN0XC9iYA
/qLhrJiVYchYO//m1SaEqmt3A4gGvqtgebKAbuE1y8Y/sbl0KcOGKMpfHxsTfgScw53RTbRs9mqY
072nL1K305qShcPpGDR9m5ua9vq4QcYE2dxGmHlr7ilTxiv35xMY/ZbPM2N7JQyRO14iRkQOXkF9
Xt88ffuW1EJjtqnAWkbaH9zFIk9uvW6JU+iK/zJzeWsBpuLY/RRSuKlv53ZQWvE2EixjcyWgIovl
US8kg90BD3Z7m6cjz18rH7pBvSy5MRMDBjOrZJ1MQCerG5eFBo5wfwL0AE2x22oQAwMOQocH11ao
IEvgvziI70A5ZRYXCfXo8Uv5LqcjJTM4NH07XyrcLEkz/RAI+EeDMTmXrfkhsW2XFc1YYWYy/2e3
hqestcJQp1NHc+IF0U1jlmy07ap59DgrBpv0uQMTV/hDetfu5kGWalbUjLlD9/aJo4E3zIOselo1
9adToMTtiKiTBD9Rh6mRur7i7pFL/7ltKNJCkB7m/MQBzvfH9I1yVU78kEfrTjqOv4DT0K3IhT9x
TGnFwkpq9YGa4/VFqrFaMP8UeR2bN94yLiqY0j9MlxMy1NZBWkPDFjMdGxkghZ4LgdqCtPhD2Fqp
WK3O3yRW9dMdBWOqmf+AqdvUaZbKhAzwdo5VoEKmoLZ7Wp6j+CHGAIO/5lViM+wcgNjA8Bik7Yr4
CkDjRPbuVlQDECx9E2KnpCHwHIZ2UUQpqt06hXPQeA26E1cquOn8zP5vYKgIijRyW3Fu5itBkoJY
5JZObzmojnvkC1q7jYzokrFUUYVJEalFMrd+FcWxIIUOOHzdqZMU2kAITrJ9ildbYaMR5UYXCU+I
wnDuL64UMBHQqsDDuP88OgkASyaP8/H/X/gMfVXdBzZZU1OEw6cXkxQibXz10acNavUhQxuiCUSU
5RbHdhaqqBt+XeFSubeTCzMdQW55X0UyyN5yotdcSho+rzqUWrX9O92a8TRuSsUOYHkOceyEpoMw
jCt2FYVft+cCLRGWg3CIPizTQbB+5IYwKeFJ+Y1tAHiBjpB/L5U8Wkdbjq9gIooC5NysbYA6OsTJ
gIRWMDiTOlYhU1kj6QtQhQb31tMYToz+KTHmRxy+5EU2BKXcjhglNA0H5v3vVvm0GDpeCqu4ElO+
Xejx10DQFnIdV9W4TrvgNaYcnDxiXbf2H3OQh0bZ7gcLmbrBhZ/NJx/yc7C4EieDr1w6ybxikRRX
J4B/wMB8G3N1KzkA/k6CiO04cfPR9XKSuL67oMeb4gkER/qkb/ME7V2mm0U+q6W+UIXg1GlHOEKs
1X/kuT9DP+zcCsyDPpw/QHnieO0vJzblO/WFSYmf77ezp5pAZAavKPLiHmtfJl1FPH9c8zZOMay7
1hy98JFm6nh0u+CA91MPyISAMJFRY0IWTAMf0W0BM9iDiyx/FJd0IULMLc+nZJkESi649zVvkirM
F17Ny/hQ4TiOfxFiFaTAQIbyIglQ3WSNfoPw6KITKgrSbrtjuH9o4vxbIRK5zHBeMFe/zS5mfVol
M51rNqgmEKrR17U6bIAu6bQmfZQ/gHYmfuClG4buchsWCDKf7GrirDmd9gg/JdaZtHJBbP5CV3zs
STu8sv5r44hL6FA1qF9HQ8QRqBU2SADbK7lLzuEB2NsR3vfoUOSnF9W7OIE8uvj8qzbcd3Pw3WA/
INQY4NOj+d4RMBvcC5w+WiJdxx3eqKHma6yw1gS47PCXPYR6do4wP4fJSLXUq9fB8euFUljtBtxT
DbHAx/72f+mje9cFTEVb3IfzOAiAvJUhgHxSyhFQ8aKyPt/RMHCt4k1luBF8Jsiy2x97yCbc9S9G
ERDi2289oxJysV2nFFn+aTuZwFjCkZjX8+X1spsHxa3NyYBcn2kE1uwM3eXtn6BQSSlrkx8sp+fO
bgI2PsgWtuiI963mXPoTvyhRdR2OjZxaNRO0gLzqwr6YsdAIH92NMtv+5VTZv1K/9P3xFVFMWHNa
9/F84Kx39N2MjXisYNwp1odTcMo5FUu2CammErjzxqgwOW+MoU97j/y4Byw1fEjBv8yU2Se/G1Ue
AVrHIyXPA9qaVGypwvNbwRz2TBR+J32QOQPtHZ9QGlvrm5jSfDfInmk0khYhu06aedpJfHTFb9dX
nUcfDCNQLP6c2+Dg3aFR0nP9Q7/kPvCEchbb7KhCCEcfochSCkkMRZaHUBxYBFo4o1RiCpuP/bBv
4g805J3zDUEmt9cRzVYGNwCGMyTrqwGLraOkSU3ObjiPpzKoj6ima2U78Dgv7KC3FFE6dVvnYS4Y
WQBoPr4BoJqwp21JVx2dMbXoYeipe3FkfR/j49pWYs+0m2T9xfiUj+a707tpfDI9R45Fc3/bT030
s96/PqbdEtin6GA/DV15KFCw9jRjq3DS0cEvZqm1V1Q6RlpHdKubTU0SelecTU2WA1/MgBmp5bvw
Yq4UPjVd1L6TjYnndCFF5Wrg4qXa2Usy80xNuoCsHUluG/Zqd+oHeHXlJcE8JPHrTq4l8Dta/PwR
kBs4g6DFizMzjXpB06T61kwFamCV4nv1joW7QTpkH9w1Szd34m00lEi8mY48r/2wNGZ5VLPNHPyR
2KvBJpGeS3hvMz0EUnsKchHKO25f2SOh4z6RoMj3QEST8fheSf1ZhISj76hazZ7OHSAJh5UjGOy+
itgFLwM41mEXYSGaiGcnxNHqV/kO3R9L3Rv7eMqYvdgvhacQteMNN/qErcW1HP6X7IFEigg4WCum
bbhw8DYU4eTLkkkTBi/GxDZcrIvGmeL3T/CA2pxN24dX4T5g7n9wRiPsDW7ycyMm/HHpNUDvTGaO
t1H0HnxPg89Fc8PVjPrNqKvKj/8jpGD4MILEY8+NPr31QexmsXLHvQN5v/UzkilS+nZ4t5VDL2ju
cndP69dWHst4MAy+PzvzKP+gwG/vy4sV6UxZaHPuqWN72Sza44u/f/mL4+YMPPS9P6tgYP8C9Or0
Ma3cN9A9psPB5azbLv0xWFJnBc5Xcw865+cwUGDU1vspAYPg/wyqXlSr/dBD3fT3jsnJYOsgJCMa
iNBuReNJaAN7sSI7JWsIRTXONTqbxKrykiBCP82OTclZfoOVkT3yEmfOAlgpsFXVX1KpLG5C9nke
8EnTLbxIftl+Om035k2ssHwtD2YDIQXFls+GDNqTbQUtmH6x54UIwGURE/wTaqVEMKMG9UGNcvxo
jVKVru2gAp8coVWpkkMFPZ8LsZhl7DX4oA2XxBSsN1T8edCihS+rjCjIQFnHG8RR0qq1JT28/PEK
M38HW5a1P6WXxpYkpL5NnY10+NUWk/wF+JEmRoWHcbqcx1l6f8TnOwXQ6TwhLQQW46LEObnztwTb
LZSwIOdNeELvw4AbvsGV5olq9Oj/igOtqYv2KDtSILe8b21sG6U+LIC1qSG1VtQjagAb/+WTAk61
hzBVuNuZuisoGXK38gb5IXdkTzdh514W3GZVcS1e90lu6MpyVQg5c3g0xWmXMSolBdV4IUCDIJdy
jBLHXVD3ydstDaLERTI+8UbwSs64gMGmA9mEp8VzuWs4a7oY8cCHLOi48DfxckFQHgAdzz9VhNlK
c+9cjZC7bq+mPSS4keFUiz/mjAbwTXAs9zbmqrgskX/QXtQbun68jYVbFPBE8OTiqVfrjzkSHP0i
1DVxGlWNHkFr67ZYCmsnLadRNWUwBrdvu52J35rndDZTC8eo1bz3Lj6SMGmLwoFdsZuME4JcGjdZ
Ujryr5IcAF9/6bOAM6Y3QXggPS4oN8nBziN+KslAE+S+dJrin5nVpHJr368qQaFWpz60qnuZeG39
A4dFO270nrNVMbdotSb7zY1UcyFIv6qzEGygBDEmiwc/btAAjMuxCbzyD2vK5X07tSlNX1aO3d5+
dPB8ALOyPvIVm9rOd+R4W7pF0lKQypUYqMXGb+GWsc0Tssyzec8HoB4ySJpB3EPjoS2KlNgdfxoV
jKv3OW19hG8nlliLxcVCcxc/a0NN3+K/56Q2LN3zZcv+7bxNNKv68XnzwCEel3guNS4SWN69Tujj
mcCAM4maBvUiHFUHThQZwD5/Dn+CFTNp5++AF43jxP3332Pv1Ep3rQLvnZsE8c97Bv5EorYDTyPA
Bb6tUPa1urTasBMa6nYFARRw5NenrNhZYxngmyjTMM9NL9BpHAIULpmdwUuLiGMVQq4enprddKdV
O3NDzylXISTx9al9Ke+X9Uysj3nJZhap4/gx/KoJ7+JL9X6DHbzjRE6Hhr+HuDskRWBl3oeCCxaT
1TKJ4WL9vkmVgVlHNY4hgk2YdVep+FDHhCOdNzhcZ188A9rfNcvfPuDtp84jAKVGsXGbL8GpY4Yg
qUVfhdkoVrBEEvMBIBZpONnv9vb2Yoxt0Zmh+aUN4+TO7LuRJf1jWvPrnxLaw1ciB8fHt5ZVbywv
8ihGn8L+P6+qb2DHeFjsJQnOklDMCxDbLJN5PSN8LdICHYbmTYuXQe0phIkx5f3gZIr+SJCp+vxE
DE36DcTSz58KgSnGnT8k5Ikgr5CpGPoU0Ar5SEwhHUguYJ7OW4jdM55y7ya1pHBOi+FeSGiH/Aji
aUpgtBg4Ug97wSrdCJVOWD9eROQUX46jtf/Khz3XdZM1T0xD0hbiIRXNERZHWqnDaoerWQT/HdKj
lNu18Jr6Gmh2Att3WY8EsGGyUQkKpigFtOpmh0IFkBriN/wWA2Jw0s88THOkrCcCWBvBub3n9TAk
F0p/IebbkSXSm7C7bScctJVo3HAqpBSp7wAGOU4pv+hxudHlaXr0Wb9UAYJo7+LrYcx1OOw6z250
RQbFTKhD7FYj+9GvCxHZ0VsxXnSI7DlaLyP4SDBZxfzLfcScctp18W6p7pwdbqEJWNvR8gceFioe
e93MHYI6A+5SF5wlEWegwvVJMqVtKfVfsz3cdDYUxlIvQkKbPyd7P2TfpdGemnSIm1IA/7zplxQF
7uySQeyAZyDZsTqBckg7embPqF6y7zxhEEc0CBshUa3k3prcTnBppzUg8p4EfggPla+087DdEy0z
RJBjOaxUeUm0ulbR1YPDhoYwybpAjNvkYk8L19uL0iQfW0SEIeORFDpnOfhc60R8YKxJ05tfwH7W
G3M45ixIK0WXHM7llsj4zQ4yeo08/i346so2UazhWu3XvLI3/4R3hN/Sw/fnUsMfUlu1UAihiu7c
pnTPeHVRHnX09vWtdgT9l3DXfYM+At0K7g0vl+le5NS24wv2C94CPBxm5z8CiySoqPH9RfdV7YcR
R2Ns7wGH3MHK+xpOiCN5CU2w71Hm9CKqL96CaQx/M4sBuZrSoIQy5WXS/4b/3i2hTvJHqiOtQpXn
tRZbKCIGpOI3Dlp6ALTOHTBly2kzWtTqcL0eFLpcX0vElOcjfSVNaWFiaZvjNutvQHTLmi4c3fLb
BuLsTsrsrQus3jK8MGJvv721fnthXaUi+SKNZlQMQv7QCkl5kdRHh8X+MHksF5ch2s5F2mJUvnVr
/lPykWg6CDQjy//v+UCqC64XqG2bwGcg8P390JlxszqLRM9jyiQPMdnjqcg4afDfWImPh+wlVYLU
CFuxv4uezvb1zZdRkrb0CuPdssN43uwkkAeV3axX7C8xDPX+4zd5nOlx94noMGu065oO3gqNO6Gq
dbo46YCna70QRMMIVmiBGAu9xlc3WWK7Zx5abA7B5AitHrfaFM5aIsKjB7xAN/E9U4tyF4Slq2o9
A6X55oJ4S2tEBm2TCtnwb47OWtGra+KFuATaFKQRsyAVJZEuQ99JSbxZGico2AeogCk1azAc+1r/
ZJL6K3n4O2uZ3Zck+V6zYiZPR2n5sZtBHsYn0bLJQNCvNq0PqXqVNlIamqG4tlyPVPJWX+S554SK
8taJpYemVB/wigq/WHogeh5yKPa/soYpy/p4LEb+3xad3svP6KN/vbR4qbkZAflmZ3W2ohyD45jc
tZqbab8WkD5tVkgDVhXk8jRpnlS9icXp0ehuALYtyiuY6Iodq0sw0mRmuKoK25EvTyLri+PVhA8Q
myl97vDB8z+PECkQ6wgOiZsDrhG5upVZNMmFQaRFDQ5LIydLAo4/OalUOjlKnRAC7BLyiv+Wn8pq
NNl2VVUCBXqxfTfqyMEKyBRWL5E1GoveknHs1lJzEHBk1B03QAaWsk8H3SPVok7L8+vEQLwgffcQ
lDemDCUE5Ui3yYZYcjEBJUi+6arjvLeUsVWtEjBMahv+dV1eRMglRRz8ZNY7CCLBn8w91FB0ns9v
cub5c7DAzjmgrACx2DsCszBiH/1FXh13qZLPWjhPdYDEhKXVJLqcD4nFIPiz5staz3BsorhH05WJ
l7u3yIJITXma9RV8b8GwchLSxT/XNwnTm+pz5l0tapikgOWS9HIGtiu3WZAMum3pDDigVMLRc3ki
W1o/8NdTNheCNT2+RlcVkuOPO7oTdw8i9xFQtGmtPqJbtCHEzqSrlyXLGfBIOGt0x54lV5YySjvD
SG95U1dfb8XhCvsU+H1j1v0v9waZyyQmn28MajEx4YwfqBX8NEW4PNZhQMmu+59rKWzOcI94r6RF
ZRCBY5Lj6yWaXBW67uA8gfZBf+dx5oOhIFJQKFF6vo7JaQliVhWLOw4p8O6qcASBgcnlnBS8dM3z
Rgf6pD1GMWdpIjJgwWX42qxDQonG5zd4n11JgZkF896NoSIJIdGptAmjuDt+8DUfQoH0+hkMBxGl
MuphVDAjuGt0hktdH1sVzhnHLG8ZkQNjs7OHOXZltf1YEaLutwsLCcofLZfzTtedKTd0usauBzx+
t9g+RUmarq+6nViyvVJVH1AVDF/CwSncqm9eKfCOvC8zYl8ZoQncRuYhkyIgHL4oQxo5L0xiCZzy
duCrgyQaErE0lUjTp2YJNYd3gDKLBDIhbxJso8avf+D+ObhX3K0DLY1lDoWUIE5vNicgdYvXHcIZ
/oOiQN8SasLpe8RUvU4xOjXG3zbXNGxeAu1K1/66EtxU+iq4ZnQx+xQh5ueGQaM7I+b6hHijgGkc
8nXPtkpKzkOh0KAVhws/6b0CF0C2bulCrkV5yYp4zpfW358F62tL/MYKqjcAQu+PAqWVPucO2isa
jEOvoI55gCMvq5FUjw8eY9pshzoMQDGe3soEVKdfcqHs4mo992Gqjlh3qF6GD95Lr5faG3fVBgx5
tfC21D9fJsdVUou9jqvB9SuvUfNiHUVHb+n8h7L4VNJWtBFx1FHdBUUR4eF2r9Lt/ArgIO9v1HYS
/+fWZD0ZB5dGredpcUUD1SLS5IFwYDTOCioIAFQ2SiZgA8v7yT3wFL6pEx7OXF7Nnh/3n0cdaM/6
j0plRCmEyMefIEkowkLro9tzl2+6EWkvl23K7HETAebxukXQalw1alCVxsNRShYsQw5+6ZfYNtP+
3d+2OEpCfuk+pVQ7VfBDHVfX6Wok6CN574U6dIhl6BQgveTbL9hUYP6K9TvAcxAJW/jrYqOByI/C
Agaa7fGnlYXYx9NpSSB07xEa0ohgINTdHoa3Pn77AwBYLjx3XrrvNZJR3tRj1CGsoSGHSgTsqn1y
Ogf7Luyb4rCprpYt0EpTGK738O41yw/jJzRWTW3mWvcX6PWsqYgFIZl1EmS/9sWy+bByOyIBomDk
BiGq1fmy7rGjsFhMllMKUM+xTNuh6RgbqxfzVeEuVr6Ay5KK/9ijvcy+6M+MvkxRKHFMmQEbsZJq
CXw4DUxm73K+vChm/a1BQxW5TmFSSRC4DHJWLXCA7NNhLrI1bbemXeoR36QCsyeSJj57SA6Pk2s8
VPYe5KRbWKPT0dHMdPoxbHzYWYbNqebF2s+6c8RH6wnwXMElJa/FuJH9AVdmDZeGlTTTjD56DyhR
wWQ76jfCr+cfnfOsp4t01QVJcKIXdafIDUxLU05Lo02M++x/48HehdKFh2pi1TBJHHL3KDk6dz/t
nbT/NfLDf2SknAdeo2JsOlPRL5zOiMy4wEU9nVX1tBgzO8sYKcsT48qwt1BzL+OJALlX4l2gLceD
OBusbq92c0f6dEWHdt5WpXR/f7RE2YGeoXYE8oh6I5IkdaH9J8e5GE7M4CzD52wS2RocptrrBKdU
kNlqLLxhu2uj8Z0aKGHOAbhHx9l3nRNSTo/uO8ao4n3MV9nEraCA/gSgMHTApeTFCnVpmkjpjPsN
+rnWl7q/NVHWA4StE+UsGi6bFfX7W5WHDoghl+E+hsgq/sw6cr02vW4Yy2FV3tUEPQ9KCG+CPUZt
D2zrKBQ1fw9DnelpQ8OFSNGryBYarDtfRUX0pFpRga1/lo4LctzTj+oWAKGei+BcqTvpt3iULrOd
vIsNYzsAVFTmVKGOtsZ+5c/ZfdZeXjilC+QXGpsc9ORDwrIZdlI204esHjioCcpYJMZYp5QyAOCN
zXoGoejQDS0WloTl3KkgR6+uBOy7UJTukBt3RANq/HIOzJlZ2q99qj4Hy8sYMy1jzMlttXQtrUR/
pPkLLSRqt4lDcR0U4pi2kD9mF1lX5Tz6cY0vpRtoUp//Jk9v7xtCw4Sk9b7mALhzMDbEOQ2C0uOF
/P5Hnr10e4IzIIXnNoyRMvSB5VWVM7zoAWhAs8SCfvJkJ8n4cW0F8+CDj6T+e8YDOUuVShOl67r4
Wgcoq4USS6zmTngepkPYRroEZ6fiuK6mALnys3vvp/z72oYKdZcfp1IPipIWbM8ZkPGEURlS7v57
DtB5fYvdYXjqoQ7MLxylEfRqqZjz1YnMzxTHrwfdZX4KpEqikkVHwQYilMHTyuANZOg/LXBUwh+H
4I1k2IEuAhBrN9uQv5cWUk/YdyKTanjJFF6MRNzB5JlzdFbrH6y8bUfhC3xMoLnl7pDI37aBZMHy
TiiulO83h+Mzevi66S2QlIPOiB+7GeywahY2s8iGAFAb0MqjYZ+BtPTXyZTpycXaWmf/1cOxPCqO
q2XIdcpONJTq1KnpTTpWQsxCtNMFFt0ZZyaLx0RuA8bMLN6AwM1b7f8zcnTJF0tKkhx69qsVToOS
Z6ovDUJrhRE2D5w4Z5OGiRNdfHHg2ZMrYJPXUG4cugDdCIA+CQpS/nTh/5TEpZ64vin5uWXqPBqA
1WUeewCf1sB8F8R1oHQjbMHK2QGirnWb+aZhau7ZtIIU5zO+8u+qYgasXG/D44zwR26kueLo2Q27
J3I2kendwhGXrZzYiJb95cLdc/xI4KGTcWCcbXD35xl5tKZN6nk+yNX4hejMVQA2f902S5hy6Fg/
662wFnEj2KDnGfuPpgbuSwpNs3QFM3rHOZ7a5c3G/Va1m9liOYul1Y4dny29RBeMPsNII1ITKj9N
XZOu6hQmgJGrLqYmZo0W2HRMVW5YdQH0VXGCx6laDDn7KExqQkOMpoYNO9JjZcLOyGIuuW92v31R
87T5Wumw/XQoJLtnbXifwF9vkvfy78p34u8i2X8WY0UVsTgsCtQCnaQqfMY9SzFX/cJaR35suF74
EhhpDIKmDJCcGNssgV5SFrBMnzVKsgwtyKg2Xk4oUFvEmzkxeylwL8w76RR7D33eSakOatg9LnLq
/52JOIEn29OJgO64CtuZfmtnMKuZeDiz4h9+uveRP+x23t2CHRsdAQ2XWz1dS3BNuwl9rYCJiD7S
M7d7pkBMeJ/cxJlSMGF/n7lcP7AI7Bwzwxcnwn/WHqOWzxKpuBhlVn/H7mfh4TY1caQ9cKNmaDjX
3SHRCCbqVRjNEZ0yw914gbAJsOUX7ZJ79aAKlQ9b90AfTvpTrUQ4cbf0P0lO02dckSbdGUisHw6q
p93ljTFs6+kz/rxUt7x4Q4NBUHV23o4lzSZIJElfgwdTQyQwgwyU10vBeh2tZGdENRjuzBb867jy
bby5xyIAxgroPz24QwmDFMPEj9RvuCItc8+8uX+OHXB4aiLvaCRVWRJk89USyZ4KBU8vCw/FcKQG
UKKanMIvezWyoqWa1HLmSNNIuqj03WqICI1GsBRu3oJlsLosO3rq7FgKRzuLUHbegggtLL8Nzy5a
/vkkeu9dZcf/bun6bHOmdCLyk0ebs7hhtFQNcYNLz8ZcqHi7b6kMHV7DJmiicez6YPqQ7lRUD87Q
Eh5Ub5U1G15/YBptgLgYt9UnvWZeq9sAuJMU6nZ/g458F7kGTD15VELbLQ+N4VTpzL0d6/E01Hyw
MPHMHLfHKBKEY/irD59koPlKQOL3r30XLz2+KcLSlZhkpSVJNUGVsl8peDnkxiv8wtmuaPR6FXzZ
8LnAyB0drlA6QI4jJ4f3fPZTPRskDu6TEGXApIU/zVF8lkmhJHbgujiFXwtmrEvyLER5hCIeTsG5
8ullcSKP7MP4Ipdos8+BfPkNdw3aeGjFhX5AL49+hCbiR//vVFD1Yxg36GfKYPSaqaj1pjvAneD7
lVwdMb7DdpaVsCU8tvrzYTZvpmhOoCvB9KZyf2uzF6cs/7/PVxZcR/55eSZfH2PVxEynVeM/TZW0
kAT4CWyKyqnCqN7+cTdksf/rVaNcYLlrMI6Tp/cS1d54r2lKxNCP8ylPRrTslQBQnx3PtYKSPjWN
iHPQqHXlqiId3hX+OgyV7o/JexC+13ztgC61WQafr2E32PGpVin4S8P6yZeID5fSxWmWaQ38mvNe
Qf3eVlTzDZaGSrp5+yrr1BPtjJGl7E6yej4c2y8uW20GqOmcOFAJdmRrK0mjVjdddb88PnrKLgFy
kYHf1uDHXs40evtxtPM9+5Kvm74fKAI24kuLfF6bS4T2/VNoL1Tubl65VNjSEiMrLFhf4olmgGHS
LxZE1IoIo2WqOL8ABju5K5xKqOvHn14gc0OsWUTplZ9soIu5brA7D/82Jr8+z/y66y78EN12mJKQ
yGdsnBMMXQdgZ9iyRdyYi0ZRgv5fQQTcK4doBAN8yEkaOBjNuKiVraKDElEgMO8KQoGpYH58kRgH
wepyVbP38v3vVzgRy6YWTlqtG36cMMd/BW2EfJS7/BZLTltWe9zToOj1Hci8ABIPX+PBMXzAdGkp
pWgf0Opu1H2ls3Ig0JCPnhcCbfLfGG0T9d165g5tIEKAWfo2Qo6DE8Uh9un5QJNsoaEujm0z9zPQ
N9ypQswBNtIHpLoW+vIN5cxQNT4VqmdP9XEAuBhPhsKQc7nUg7rncVb/9c2FfwTt4JZxlrkVgpVI
B+wd9jLl9ctha7bBmHD9R3BGV+MWJGnGisUXkslRCXZKMyII8hXbKM56tMEgrSGp/JlJgyt7OtYX
SZj7qWa8RvSPm5nf9IEZzfwhtJq92Ms59fPMtxrPUKVqkUJDHUU93eD3FS5FpYIDOFRBaD9IpXoF
lmQqsij67P5DFPDxhK5bEU6c6uvb1L6r616tTlsYi6E4spZLmi37MDERdDFT4GEPoNFkXZXHArgq
K/xmBWUTXR7UxdzPRGZ/iXFCS04F34crQQ2uxtqr8NuXc6vdRiXaYezNAXBbKPWQ+EFTAoymlbaL
sw+RghaX+aJMH3ashFpa4rEsrKxKaOJd6sXKg20vFoyHYYiCvNdiGAIXi6JrCaWj88dsSfzR++b8
jJxKHZWadMTkjsHFRGwFAtf43nU4y3MqRDZn05jEKnJ5XIA4+mO4vunVX70APqICSGXcnYH2096T
BN9+CCieDYJT2nfrY+RYh+xpPCkAX1opunqioSUfyKfj961pLYMBKyLEVPGRR/nL0TfS4P1zwK5W
kS80hnzhGxMGi2UGMZZ1t0gE0N4LbANfUD7XNnDtZN1+emtKmFrd89AF48xSsFbMkpvhIYkVaDc/
WejJOH5564JYsueAOQfAAwNxpnjzLVbMnpit25bmHwyuYBNE5Uj3x5NX5+RcakeoojMq4oxsVriJ
FJAC8pn5wwRQkPgbNJ1D6QYoKYMGrH9lG+vX5qdY6sttrNf+sKX62cUC17PMC9QBgmg/VTRtjhG4
mzJjkFnV0ZTLJhzEO/ZXWB9Z560NQhE1tLsSOmGBAc8dqhXrb6s3jM6hxoGEJlrLvoXy4Zge2x3o
FsKVbDzX5Tn2vsg5bsr5IRGtv6LbV3fSWAoWAo+OYzFK9zqYxpaw3HoD9yjtXzmWK8vC4+mLmtFM
qUbCRIs+aZUjMAXP+lm+jhrWds7jM5F+djc1DIKrrTpnveh2X4fcvZQHhRRyohiuVa2FB+5Jo/ik
OLIB8hCsVFEfHy0ZHf/SyGqTdT0ZrcS4hLrwZ0iWCQJ6uRG5qAAqxF0lZ2z1JFDrZnWoOFULax2I
SN1zBVCUKmgyRPzxeokevE+EnH1mDO4CcJaguicaOJH2IE8kPhfeuma/7eZ2t+GAA7aHC5ZwVI1+
c+JpDVZA/thB3Z4Cb85waQITkfayF1SPYURtr7ZhQ8aTvKOZBBZngjHHrD7A21CqfGrym/S5lCka
VSSoPHMYUSwU5qsWFh4qHMVfATwV2R++epk9o5GrmUKYS9MAAay+KPwnv+KpMeT+SFPzJiPV4xto
IcNj18XkLb9xd12msfoGk+vr4dF+4iWgDzuEJrukv0cwyPKW/Vk2YSJtU4j81dVRzYEHjM7u/K04
xXzBmXbOdThEftnP19GdpVr/aBlBEVxObcq9Vrl+F+xNTU8Ez+NsZ3iG2h0SqFgGiAtT9OeODnyB
WepQMh+EkQvSK9ejrGNgm+b9Mv5e8z6mYct7eILmcUINmIu3K0f6xVUokCNy6sKda19REJ5EjeNA
y7jQEvoE25/8xrwQxavHcB/CWPO1zLGC8Y2Rjl+VKi+mtevZjAxG2eUGx9e4FPXm9SAc21fjgOcB
e0tRPzEK0xr0Kz5/jMPRW5nPVbflDNbvckpbD2iyHG3p6hpTWMALi4rSejnXDUMaEi3heaaFow8b
0C0Av4xwbzIgQ+vY+UJJGZrlAydImxQ7IYqIUurOfparKHMwNGr752Tn2KK3gngEVQXzGQKpnsCS
geJEBqnvOoyVY4nq0lxE0IcxetQU059rwZ1n2RAEBV9Ob53NhBkr3a9UGujvUx+pQQe/V4ugzzDf
ZKO72zHU+P5hbWoYzxsb0RSv/8tMxMH8BOeyH4Lrdw7/tBH6MunsZNEackPOGHARulphatWu03oo
pyVs5Y9JcX5dvh8P4w0Uy4cnWcAzs49Gx0Zo7geavcYcPItgmrEdsBpfqGKXxDsf2RD8RN7qLWGN
7zVY41c6tMuTyvnhj/KIB57ralir7pbmGOUsYWe+EXCHxsVz8U99S/5xTqNMNYZ4OWauVbriT7lM
EzVb7AQGmN4hjA3Ou15mqdPl71wpqYsiqOHwEihiKtKIkStZ4tVwoc4nXYaXXRfC2eB/4PkTUjmZ
ptNzyI7+Ft84SMzEhZ3FwSjRl8W/M3hcyW4s9AdJhkeABKVZktzR1OxQ66RxgcEF/3jea4Y1qPLF
pXrDdCjEHDsBUN97sZLaG68VzTBZWNaASFVpLSykKBZ/ECrbh5poAchtSwPG5kaATUMjkanzYSBp
F+KDw8LEi6MJ/1UYqIAWvmxQCQsk9D1vij8lS87kyGqfK49Bqx5z0jgKom3j3hNmYALQ33ua4jHJ
Q4XNbrFeYk7cNuHkoJ7xI8eklQVhyJKfFBgj1ywN/jEk0wB+veZcrgN3CrQPdzquNjaHeTlq2J6K
cstMul6okJkszE++gWPLdgn4+BfPsRxWzQYkJO/0H7IFhPpIvRYL88RS10LsXd9JUpyFFJ7qnp0z
BgoI8MY2bJL4mlPAkFqRdVxG+tKZtUCALsCP+/IICfKQTUaqDSQNoD4W37+sKj62/tMJTgFQ/7bu
OVaPGV8QeEI4O+y5Q4D/xX8EIS95H/SxBzqucEj6FYuMctKdUIX9Ma5DRAGZwh3Dw0MdGjF+qBBI
fMZ702SP4dCih7WZxk7jETWJsz3XEPAHz8jMfqJbkbvzSNt6OqSmTi1KmoWGazMkDxEkd4ZdVwNY
TXljiKiSqjfGtKhLI0B0rZJUse1HD1qDOoPq5IXMo4qnbonu22+9GnA6gUmCz14nmnYV/9bgqxPp
+bF6pocULUSAo/+qxybLARlfmC76rmQvXuB/s8g6hWaFPKHP6U0Rdjr4cVocDguv0+HSmx23KsRR
WZT21JBVpdlUKEhqxk34wTOuw5mJgLYIjvtJ5Q/e3KTaI0PTk24hB6/x4r9SwLT0Rg1wqDBwmlSx
EuzfJvtI9EEb//WT2BP7Bjpzci5HpvWncHUsDwBOZEdkjhBRSvox3wy9vsZtcpJbwwuQ1vxa0e2U
9qb7v3VkTy2FRBAW/CMvNObpkvnvnjm1jrD5T3YWzFiSqRIO1gNhb5hNfJLNgQo+LglXmWJJKnXE
b5AN576MRiZpXT4N9EZ1RXFOrOXt6VfT62nzx9YmzRrfomcYW5/GyqschJNXqohmbSkYEkooJJhE
utN/tptcN8mRtBUweIACCqucN8EO8ETBJpmDGlniqXP6v1rdhTfTJodLf5ckGaNC2twk53hujFyA
Zhqd3UOYdlU9TRoV/nqlVoOUC8kLnIA5ZieM8LdqozSDKWLOdvY2XT0W/cRczsVMAOf3364dSxpi
qLcGu+rF5qHgGJ9LcMBoYYGBv3Vs0VXpjevDKQy7BsrbKp7HZ8AWALlhMDPyJBouf+hXDKcIaLbI
NTbTCFz0onU7Q3+WIadFhN2JUBinJrnWB/Dnc+II8NUQvveFfn0DdueEje14Xx0UpEba9lxrgRft
qbaJ9mp6eYWaW6dQj2EDP0F9XFnjr2HmKPogmf5SbCs4yZ00yi5/xAeLtKuoGbYtfQPGRHqvKLJO
8ABxyBrUSKyU6XkvsYkeSTKgbIUDXu1FqjMB34d+GXkAtHE9q0JwGBDl1GKIEHMqsgd9OLxcmQWt
LcAaXip4bxiXY2WvUXEgDVdGFqzqC0bEgg86Mg4oIQDZjc0kQzhe95fpu6FY0D4iBAbMMxOrjSs9
+EWdQ6+7bdmeu8qqgfCPBDSTpfKEmrOjqEcPVALH2DbNz5zfnfDj/Rqcz0WdQBMvP3VlcKOWFjuz
FGXppYHx44VRnR7Ys2QoeeeuSlhAfYpRYQ1vv8r2YK4euocUZsdieoOH/mKokzn8150mu8Os+qFq
6fE8BkTC4t2/yntZX9iIqyFQCQM7mmOK1fSFT7afu4pjQA/jkcaWuRd84Qr/GiOd66Gs/nGEZ1xx
tnssaQKRGrRHITpftGj0rhtwHroeAvWule5S9VzaqFS8KhogFQXxH5yveWDaJED651L0j+50bwTA
3oBe4yKUUi/Fh9brnIAgkLnFQDWHWvvR9BP8Gi9LAtdGGNMY1K3a0mjz6KDXeD6Szj266k4vXnQn
34t4Zdivg3EClzdtO/fA+e5Ki7SNIuJI233moL3Maza/vb9soocZZaz/BB+zlxXxx2U+km+74wNo
525OIw9a4QzCkbe+0zV1k3HctAcuUwnpf1giItvpTm5S5rwqv8FBeCfI36F6GS12ElbWVKpyn6fp
iTvsuUPa2as5tyFDzu71yJPUM/VJcx5jMrrSWy5TzSiTR6UmaH7IIVOJq247g+R6hmcdxYZ4gZrg
4qjTVPJigid5Q5S+d9OCiMbJIlc4AZu+LNKbltLi8TDSWei3sYFIf+7/ShMSNpZFBi74bkp8iIy7
v5JNAb6/ciFzMAJ2NAiotDxxNzdU1a2P4P3eHmrdEjTNdQdK/BvKSDK+kXEiOYIg/yRdMfU44e84
ohUiCnoF+oghEcAKSHGMniiQCmGHlTe7BwEYKCnqhzORJbu9m4gsXjzE38Az7e1Yldyd3QrRZw4z
vgvaDB3goRNAxk1E6omoXrmktjg+PeZ1hWWGvxQ7TnWnR0be6CCf26CqiKeTF7XwvMIQJ4x3df2R
qmU35jH/aPRvI808xm075S6oCm6Th2sHWbZPgnUET8KEDXcGlpkBS5pP72PflRQcEnVHuxvI+mt1
JzpRNxA8ELx/ilsWwixuhUdeFSr/IAcjjlitBNtKPnTQdw8uVGM5um7oYdX8zAOFuf2MAhao3lG1
yi8rM/rk4Qh2SdbbJ4tmhmbcNA7DAckuDT9K8UPj6kkIjXbGyRsHgwVCPswvBi2ZyD32MvClzX7j
K96/1MrRXrXPgQbCCXzEacid6S+zbqRpsMhfh1X8wEm6HLOX8aSdGoejLhJtCKCtUMPe263cMPJs
/s5H9T4azgCpYwOpieKSVL9E20VzHYqoMFUnY8tIwwg1cg8xT9rgxRd1TdYa4vo8NQrw6WQLM++P
21Zy3Fe6hyt7Wx9CJ8nc5ro+I/hYrwKPRJnUw8d5JF9ZVkQ/9I6tGABoxMYUAX32SfG1sDUmQGwZ
O3xyrNUfrYby33+L9NwC8NQ+y497YcElSXO5yPheej09z4B00fAhqOeD05XQ3ARXxJJ9C0pACd+l
W6neCXByMahzXrFL3IVEY+Msvn18+fmk+b/xS6HyIupsCxRL+RIxEzctJ8nsrHPGT6tuHOb4wfw6
z7cQjCNdlsYfIgvUcnmnld5Bk0yRLUWGlNscVNiVVCUNtOoOIOp9MZU4iFuYKb40uoMVPlGB41t5
ZkLav5LWMZv+h83S/5DiJYEJQFUP1t7PTKJHXYIQMhS4X1XDxR+brhRGBBffy1AOpnIxGB4Fs8f3
g0MCdjoYnwQV2/NTwrgeWaaqoQe0K6t9cnyJvYPbu+itGSg47s7hp8b8qFXGdV9fF/IdQ0AbFmed
YdhC6T+ldXgswAj3H6gAHrBy2QkToF1UwOr5hkv0Pj01dQSjWHqbzZvbz59Al/0FWhoMHsR+cCoF
w4kr847x8m9E23Z92UGf3oPhuwtt5tOv0cYQ5u9/p0fv4xW64j8OQGg6HqLQspOYBbp+d8dkX4As
1NfPvXUN3WlIw+quSVneAgi8q801c13EOP6am8cnHIZtWeLmrd1hgqwYZk+8XYw0SHqMzthXH4ML
eCBaqg0ROWcuVRTbTelQtVFY8UozOmeILjtDZweedUgtI3n05VVPbO7TmrYVHKzrDpu+wp3lpKiW
RcQwYKwK3qItFkj88J6AIorhz8LKajgmXG90P6euYRN9GHJNygD3hY4gjT89eVXg72Bz2DQkRuXF
zpYQz9mEFFcjD796Xv/vsH4zusgFvUCSrGu3/fBM6Fi2eOwtp4Xb3+Z8r1xFFNGFlJ+zXpTCh8rx
QMkmfbGyPnT1lNwoCfnDV2S5TwImwkU/mYhiztfJkymH9JV3Dme3hrDFpnV47QEd88C+zCXidAqu
xtvhvECd57VcZkGYlux+qvvS0jB0t11d0+d1xzPOlJQZcenn/Yp21MeKulh9wKGhg1RVtG/db91b
/w7xJQN6tuSmw0X019OatA93njnhpiYOMrOz1QSo/YK2Sg6jo7HzTmBPBMTLT0Rto2+zD99U/57y
6P2DbBEFXUCwjZS3NtIyUcUdI7th7cbf/FGr6Uruq4rE5hi9LMfPKB0O+D0yRC7le/frgM8hhsf6
BTfBSgKpVyajqtwycRccyYrwr3E/hgF75meZSngtUb32jTU9Xk68dtXaJs+dKf1x89B/r1IKDBy8
BlZWbomn5tWwrrG3vOrz+pjYKsw+HZX7SkkgsTDE1Z7vzah5QZw/Csh0lCZJZdP+iEimRuNUW5Xd
UHb/ZgYlKizA8tCmagAQb3e1wRDMb6BpoSZLarJcauMiLJrmiuOwUWsQ4ipuu3UfZVWl75ALFVhO
7gr2Jh48FZElFz+BdV1kVdSoaH9PbTIhvdsZIBtHGSiTCSeg1Qd//L66jScqv4JPcV0R8EPZa9Gj
vTfdiXlfHlBQdtX2zddryF8PeWgfeiR0woWOHUPtwcy8stoM1EW9eltjkhYIK1qFi+56OaPiyDND
0G8H64kkyvCSNYY0cge+Dq8rizrqRZhPv2vvHIkXSvwrUL26hrsSPAoUUo767wt0AXNXJgtOEuNX
Hg90s1Z9aiYleqo6BGR/bV7jJ3T+LAmHVomVeIC+Gmqmz0pT0kzANBzbyVf1FRFmu6MJno2AqbwH
/8wOGUL8dtUvbnETLhJD10o9z0jbW+lglXFhUDFr+xal7V/a4Kh9cakzlWPAvfl1uvkt2uvQNc6u
yFTR6Ac37qlMO0XR2Vi6QKTEn4b7O0Wo1FYCZ02DSwMzHrecjnRSa2HeRzWSPdWElzn4FvjqY1Rn
gufnHoDDVPSyWAaNdjAx1YTCvQMYcvKQQ7cadFvCKhF3paeF1WLdQ3UUl8Xc9o0gresejoJdPlf8
ZlcINk8v04LeEPHRGncVfdkCOhMRCWkz6vfMi5nmmiS5ss+Pqsyd2Jn1sGAzbsunnWCsGuxA+AQN
nDrIlisbudPQRt+5JTmwQjbsD8SdFgTv3QsxBSGE8nb98RODsp6sq39O0VvsP2vEAN1+pZZsMkLe
Wihf+UwKPkoo51e2p4p7UwuNCfXU7VqTJ+oPKXDzGkSrRCoXrTZtyjWRQt+ludMqXUQCZVZZQLeW
pJqLDhdis4xwAdMWjxyC9IXpHLPt4hoq+2M35bTr7cSGm0ILXLfOJefTxXXGQBIPEKAUHg+QMiqM
tF1zHvUjoOpubRFG255OvEp+BRjKyLOlkAj1XAh23aZp4A+GbG7xKuAWM7jBHTbnMckfUxw390bE
tvsnWnkeNRa6Hkjk8xw9HVbQYaALEiZ5rieI0P8aNCd1hZFy3lAXYH13lQnTdLQlIy1S693qomGp
f47mA7gVGeXHBEEIakJEqR1Nh5dGzs9l3lo+i/l2BgazDWx4SYecJz1U4hfIOBRXwCXwcvDMvybn
rA7WtTZYvkyrqwHXpHmw66f7BDWC5j1981vfxWipcOZgY/WfuXXMKo9Cff5HArRdBhDxe5nZex0S
NurvdHOaglw7vWs+thxB3AYDecLr/urR9eNiRv80iNMN2wL3hyJCdNZrZw7qPtpQzWUrwwvqevLv
dzILbaj1iN14kO4jFHnxMovooqKkXbuZglZD1iW2djrTU954O952q1s6+SwzJLNEpE6tjeByqYX2
TYwGRktFFFZlCyQD9gOGboiZxYq509jfk6DawvjSlSLMwMpB30k34Hz1MiDOLTX8Vs9YubyBwuvD
a1XwnuoyTisCFs+N2HqitENm4+0p3xy631Ru68BBtZ/aNaur06E5bi5/0llGIibssnlaoGTo1SN+
F1vZuemTC4i7oErSS3la1cL6Iov6a0hlVBKluyb/w0GUqXKHwDVN0arLlav/o4i2q+PN0zRMTv5Q
2mVizdRD2P6WzsIij0f6KJtcg8DRm15VLK0dgPGV5zaCaPdyxzhp8ypxxKCoVlXe5enHgbxd3KDU
lptGYgyxllM8LKXYNI6EDmJV3ll1LoH9pghMNlMKEzTKw/8JxWgy8vTNBA1TFrjoZ9XaumRvn1B2
rB87Y5GLQT6N5vfurrpuDfAjXdlDyBAw8dyEyi4sd6EMSlk75suvZRuWtmo3C3czusjzRtPsXZP8
sRlpyzz2jbY+EtZqsCLNSCSRMyDpXJhqSgfQ2JVKlpS7JlLM3SpMBKG/UmNXDuW+lzxxUk2F2XbV
T9vKO2TPNxItHYi4aojxaB4o/CS5HtoyclIXokr6vHDQiCqhOxSeuHeb/nnXEei4s2Fr9UOLrkhY
+rmZfqrQ7+eVBM4CEpF/rsX37EvaOHrTVmxs+d4WN3RwSblK8Unxsbe9tAHKHYpeQnN118xNgvMB
dh4UVwJMHcPZGpjRO+XWpFoNoxmDwdOpm0WbAIkV/ZX9PO1I859vJoV+wrIj/t4MvE01do2XMHgw
AhpvlyZ13MAvoerEcOWODt6TUYutlhbep/vrwfoHGgnSPxwUq2g9WlhS/PdZEN+nSRrIhLvyIy4h
4D+Zfx7LFURP2yA10L6T1ZqKLUZJRrq2iP84X21OjDAxfhdNXE5vXUxXEfXBPfktrjeS0EidZ5Zz
pcRLfXgIL0yAQziakHJjdzfhig942SYP2T0UOe7QDHgMswHVaFlVSH1QrjKeuhV87jjttWSIJa82
LVqLemXRytjYSS3162/XBCNiBTRRWguUpbvZdA7mFcAP3Me9rgsyV0HQ180CwePGjeTsT9mhRpPj
G6WF7e1RpxME4lFG4vjkni/ioTemvRLAVlEH8TMMFwyidAzR4DrWoNzLAvlOOhxEsJb3UxhNVWDY
tGHO/jjFzdXXlVIazFzJsetttS/knwgX7CHuK8U3UQjo81yJW/U9U2dkKa4NTKTcNiM/YmLJ0DnA
HMtFQP9Azj1LIeEBtx9tgodTipGDJtC4p+l4rYOt9yj3l2B8ZvnkpQgVGu8sm9x8g6JiVUxrGHg5
TnwfngIRTigwMohmK+EKSh1SWiTv0Gq3ihL7RNav9qZa9AoUFDkEUa40RZzkHWK6JvMznmIu5w4A
DYaSR3ze/OSMxHb8uSweLj50PzuDfrHFevPWqR1EhWCpJ9k9nrdiqxw091Fclh2k6WqDpLHWtL+7
j8La1c3QTXEyexOmvO3PJHt/uvWdZbVNMfJqVA6dk00SQwGLVbUDTPU+ymobPwNFkuYg9Qosogr+
binU9jThK2KScW8neEMlUkajMM2G6vi0gUwuUO/7Tc7WAc9USAeOQisSV28RYVGDJQXdRIdaNCwK
vdxqUR0temfv6ePnuVgXlGgoLBzj7x6whhYAXsLYGz60bqZHM3OplwTKaPTJCy/XR3p3FAwdpdNG
hmTD+xG3k9sWN1rdPvFmlSeIqlrqzRNjE7F9l6SQsnJldKPUwpQzKzrGzIdp9kgst82KJ4Ck+Xb+
tztUuVv25toorfXbMyUbDpag6Gq9OMnCsyXu8a5e1tE7obyHz5thQXdHwyIXPDkdDb6XCIxbA5XS
zfVEUlA8j49hXQ5wcxvlWUU9KWhCYgOLVGzbygpR2FOYOE22wo9pLxXuJdQU7GgOzxYRzd7+cbKZ
a4tODUyNscXn7h4BMBNPVZZNuqf2nRni5vLvj2XgJV1RwS7DrovM4tCYn6Sub3naaNBtDtRgI9o8
3nMkFSnF0DoD34QFRK47nxUaFoT2dHd7diSbzilpMoj8cdNGeQDi2+ZL7FJKD7KIvV7DEF31z3rP
GloXxNoN5OjjkzSGKS/QNEvWZgfKLtKWNEr+o6eid2PacXmS5BWIpP8J+NTnEVQFr40644PlA4KL
KA2HKQOSzRDsx2KkXIyjHWY//K0WBhIHReDlLqqEpY5oa9UlfkysqsHNcn3gygtvVXX8j70YVpRa
6GhaVyVSnBmBZ6UgkDUvKY4E1JEZfaK1qYX9xT4c5xdRxGctCC/tNRjNIEk01tPsouB7mWwAPDem
UtayJzEx0pomHJS2pX9EV1R1rih4G5HPX9oURFTIF+zIKWAO/QNO0pFpZ542kePr9JeY1pOzh3rN
hGaNDWPKoB3iLWd+6A8GZa4gsK6r7aAXcWiJP59fEHW/Mskumx3VtfbskKlYkt+B+KRinnEjUuvg
EA7uMOMwUicMhwhl3efHmuSfeGYzGLmFEllS1Vd40Md2KGQPeDrghmMaV2cOh62A8vwvm40ph9Wx
AXgxyfwoPlH/gPwW2uLxmVoQqp827g83rJGNR75rogkY77oIsIVbBlYDgjcfLLZ5wYWy5iBlvQKz
tltW3sQjlH0AzBOlwWTBkzDBEVDffJV2MbM9jlxe4jtmClRjC8jPa0VTRdnauuiswxVSj+58MIr9
W8tl6kSt+235ritUIjdPAfsbqZtGcGREI6yEi4tcRs/8rQi/eE9uIcWdp7FFBpUwMXXWh2gfEOSR
NFgzJbc04tl9Ivx8hyaCHQe74CMTBOGhw9n6rE/KCV7R5H05Y3EE4r/wUrvC5jZ1NFDzcTjd4LQp
xxlMV10Pon8gqThdEfR1oUcfU4kuel5SpC/Bowq7/IgDRUcMz1qwqEwOa06X3EIaGeyv7mqJVz0S
HAcVR2RH1dXdseln44KlfQBOd6iGUId0fOX0Q2FOlvzgHuF0Hu+TnfKxvKVyqHLhHAPIYICjk5dP
VXFSkovXtq/cYYW+fQMzA0NqY+7tlN6NAjl3XsfReqw8YxBxkMC6ZKmGpGo7XuuHdw50RGVR7+7M
MEc6MwLc0GPD4Wsx6ImKhzrz4KX517CnOosmq2Slfsi9WzPU3G5zIkW+2Z9ynTAZ6+FXIaJlBWpz
j5QQY0+AzXKTqWFcD5cdrbEJCh096ZiL3p8OuVxjmnDXKPar7hb9eTqyQNcSWrAk7NMWiRL3lyAQ
DYvi5QHOKagoVRfSMIm5zSZRcx9GARkZJx+E3kQJyX3oSk60SqveFtFykksITUb9r5VlGnn5c/7G
TYEnymSc7/lF0klIFy7H0r0DlC5ep+9DfKY7RL8IzHMlwX5Ra7Qo475d4Lt5HjQ7apgUZuoyynR5
VH5LmAFAxXhqoRp4CGIQTuQnkC7Jy5GC4gxmavbUKQpnYFpZ62SyWFsnWAx1/q11/yjQhEgxgjF6
OOj4+ft77U8fzSfkyu71Lw7kKNOHk7n3x1rajvhIMmuu7WmQREOtB0kf0FwsjDMZpf3rHrcWnynT
9uB8RF1rxizSavvsFvRFEb2amqHua0OVWBFhM90sn1VCVVOe8lsL6vShcz5ZWcMcdD+ARP7Nw3Gc
34vCEfeFL6Cay32Mdsq9sEhAKugvfjLTbKXScK2hoQNJL2QavaltVU9gMwPE3u6A0YJtYpxkyWI8
WBL8/OTFK14m6i0IhlNoZuUoX6Q8zYmBC+dHZbRrJwL7TFyxUBNzEe7CatajnSQfHPrj2t4/Sev4
WeAw53Ybkfx2P9sPEjyFjti0AqXXQnkzJyn6Nb0ZB4/G4kG7qscPF083z02+T3wXclj4rtV4Rsc6
GNfyYD8FvPrtTWx7Oh7E+1C3lBIomw0V+xAz0NpMqlutC1xNzyi3dMotDJGgYBILX/0DRX5l40aE
NLSj05vZ14JHwNKyP0oD+hdzOmR9eqqZad5tSxLko83pG+hymAR0eJtUVwGrFYfLsBw38ygw/b6x
3cScfH5AgdB0L0WOwDhW2USpri9SyWpJVIe7OqDtQQO5uQxU37QHASy11M5wkegN9FIaX4+RWFYG
utgP5A/i2iiYdTSkHrzxbDsErynzaGo62uJUUsVVfzW+K5hqW5uC6J9ZfskbqCQ038LKhkvKZbLn
jB8BEaI9YSe1J757/vJiePihCjDBHWacxuw/QLsDMGGd+1kXBdH6/4DIJymoRb9/MqCLgVwE3RFa
dr5SnDurDVAh1vO2BP34Xg1fv2f9vcldFNAcgGyYNDy+rmCGW4/L4vyuic+Pz5fwekOI7x0Hc8zu
RKjiTJmN/z6WkJjUPX62II7kgbrqSbdxIYUlPF5ktUBoXNDGXaytb7/QFgPbsTsfCILMG4aLBg/O
zoT3eMgpjl2yofgsnAqohXTY9toNvj3ZzqrOsvbPuU73IoLGkv19tUvmjRR4JWcLM2VAW6WgHt+N
lq9y+kLfMaKHzcvBirJyDgaczgFl5tPe2edt0KedU+nQHOVkPrivirtDq1QAJ27jeOSrNjWOAyuJ
3VbJfbIsSIH5UIk/8b6lhh+pygulFO6UVMrVbTkwotdc7NuouzG+IsbhiVeFaPIdBqRbreuDYRp4
CzCqNVq+B0+pkb/404TSa/v+nL/XFsZ8YV2MzIXC7b7R6ks+9UjM4C0ZhBGsA4qeeyr0PlIwLk+G
fgZYf0gb2ENABr+2gaL5ezKk81dQ+v2AU4LcROcSA1cS3DsGSu4qXnvwEIDkdamGcZNrh9UcgLKz
S8aSzr+nRw+uL+te3Y9YOxx6J4Z+vOwyK7mVkqiJr6/t8IlZUZ/OzOhuDlQ6NT3IVAxZlS4Ov67J
hXSI547SIpDuNe4EuJqEOzVGvgXU9v+vE6ZYAhU7dRqbls78mQhMgNDW+e7F3nJPGKe3uHyRhqmp
dnHuxhK8vvHdrMSVUpZOeoG/1Ra6JoEQpNiYl2GZhbIANYd0IR55e++RXlpICHAWyJVpdmzTzmrG
KapyIygTzUqvTJH2BxN1jiwgIBvCReGmH6ugzUltkEjGj6JmwXaAdo1EOK/Lt4bWCuXg+Gt6/8ZJ
khPP3r2MMvkjNQNLf4sXXZy8jctALwYTwuxH6ySKO6p4V+Qc/8szg3BE0RTXOZE+tGp105bLp6Cu
fO2rD4uQ6IWwtbTyQxlEjvtoAIfbhtnVV+LhkzV1WNhkjO+hiTUYWydYxejRcDZGKgFuMdnBn8OT
LElTOOLW/XV7vsbrmA+OoJFcM9AsMpuP8ehVPmvUxzp/XU4p/+5UtsZKvdXR3nUvTWicbX8BKRXi
e3Tx05CWAz4qQWpTZX4UgHV5YKq4CNbA2NCc2j6W9l6AI1oY51DqGv5BjuvgsaepX55t1F5xwg9/
QI8pEqks8mTszg/5Avk3wkIKUAUIk5hanqnfGCEjTDw312iftn8zKrSA37/yd1+aIT3BVE/14tL3
xneqS/b+vkll+GnHB/GsK1ZRsxhjqw7JLUQ351/pv4act++Ab8E/Ti7b+PLCgn6+Tm3ZlgQUJtxZ
8eTV9OQgxXu4Ip9oDf39kCbKlrBz5pO+kFZNgMMJiGeaaTEHA4HKGYgrYV99NIHBq8ZjvlQOexB2
wBcjYFfEM88rMGC2LV4Ld4p6PRgiiBIYltQPDvhVmkQA0E7WWWsYLQ7KETqNGzCvthX0P398xWbq
DhL954lrQsvCoDlEuWjUsQD7LP6itjmp/CL8vg1zwUhD/LMOzNlKco7hn7WaILZIsXH43guHMhlB
aIBt3/onPmXbetO/2SfD2cEQmwxbXvg+A79aWmAzW2hQqeRmDUdxrVOL0iAFYs/F/U0XEsiEgKv/
NfXcylriaKIBzGSilVAppGy5nbX9t/T9R4bqzQaOaL9Nwlj2z/K2SEvMyegR1mEaWvLkPVgJSTIl
XxvXvUuTBVmTiMzMtyi4qDJZpYhPbB+BmqGyMMAB3lTzJRCiK0BNT70fCYZ6MbYDiO24l6bMlvk0
xgy0iR9bFwaa1ef5El3xgqOfdYPRXU4p8gGy6YBZxUVPvWPvBj8NcsWn3D1MPm7VEEoWBQGm4D7r
NSTIoup+bwpmUxfUf2wv2e6oVDKbanS554v/euzTwBsE0JH2nBoA8d4iQXjCKb7vdra2pW+rtY5Q
lvlVeXcEUz9irXEzixfwjR//wCDq1/lf7XhwpJds3cU9DIAmfeme7t2RAJrbsoizqBJ6dlcTkY8B
Rtc9nJnFyBcGjFvESMaArHYo96IwgH2F/pjNKTMN3UpVmkT1M4FDjhMsIPz8HncLZP6Sd6HXeWKX
6/4PaDzi4Sh27yWH7Co8rxKzpquIe/8XXzjfjaddeUStnIJ0tyOfz5K9itQQ843SsD1lQJkj602f
pALemWRzOOZtCAruaMJZGlHPBmeZR1iwODazgoCpfrG31Bf4pvbVO/VVUfQGabGwFoJedv2RKDEe
ehGrqjurzqyze0xP2wWR3ZUBVvcerycxjQ/xJg79dczhRX6rfidFJvWIr8Q8nwsr9QBEfW1Pcbe3
Bh6T6f65EwQRZ7PEplMCC8HH/j+b3LsKsnWxHwuDGUCsPnJs8ihjQyRVl5YTavBRDczXmNTz9iOi
T+JRpyeboS7O81MlB0nrR/gl7AWFFzEjUYaS3I2cJUyOuAyVcHdpP30FpBQ2w16LsYfqJ9onoCYN
DlY2WlCmTtEFPRyGdxKpEnKfpDOBpy5244a0iS0SqTUBTI3EN060GTz1lbc30D2YeNRUdBGXz76E
USnowdS3SmY39Oe7Z1D9hchGK+q74nPv7RR50EOFyCfyCkGPROlru/K17N3ciKisF3Xi2nxEXdO6
7cjHeqM7UeU34rer1QaHZLtx4ZILocyGGgrKKWUOOTX9aOwtOZq1VqO0c8ocYPwYHxE0IbjEzvw2
+CglNbATMEEfrS7HG/kdR07Kgs0btosXVjckrMsGEy9EFOOommrzCRsh8vprie9WWXBvy6jMopsv
ke/AnPMEe080i+kR+0xyUzXFOk2h+Ot0RiouAli9u56eYgel2Rt/hsdpPKAfjb6tM8qKfoEGeYPn
XjGVV8oH/wLdaq62QBklH++AM15V2YmY2vELInMYJ8IjPDMGDjdwQCkFVbLcWoCKBjRcyKU8/LG7
LjBM6yQjFJGleD6YIoIPXl6qbN6MT3pZHfYz8qaniuT6EupFsloXj5aHjBPhRwRX0YVJsJk2/bsw
Dw4WBKylrwrpFSveKxWCJGr+toXVnqu3irFKxA7N9FNoIj4VvsVsPJUoKesqO0FaHDwQiXAmH40S
IVbz7tAB6U6NkYovNzEuNWCTLpAL4TFoL026sbFi8c4cB0Rwvmc1/Gvw1kFJZ9JtHErzUfY3pZOl
7lj0SrijbmOHOwCuToONwCBd5dxlhspywZ9Qzi1+nHlb/4Osae8Zvo+V1zG0x0x2wJRKekx8GJ/6
W5u81iGi8f0cIyc4kKfIlPsbN15Fmh0IoAJPiAJbGqxexmnhz1bGcVXz2UxeIf1zj/yMAqiYuhqz
xeSzTMnkc3ld09bFwDIQ991JCQ0tXioy7KfzovnFXtPI41xBcEBWE/6oUPY9QHvsTyuUETppNS6M
AZqhwP17Z3AqXnT9iY9uCnCHTv/hzbZqnZvr8CMJePEUH6h3xb6TRgyGF9Skt+8b6Th424ctx25P
sJf2cV+0Hdpc1gpZNDYhyUzvbNZzMFtCU54xPpD5mAfNdIzcU1AfVYGochshq+iXDRAtiqbIAzWw
/noUqLL1jcc5K7F9+JY9Obdzknduu3Ias2OQGXnGySQoQDGdH4SKK+IrJqxhsNicHm369drZA2XF
2GREZQxbaPl5OaD+s1xENw++umb5ZActWztaYLPMvNDWtXZ1UVhnu+DRhj0yANxpdcB/xynbZj5+
7gjmMrPiC1WGWI0Kh7RMOUXFSqsdEVjhSSoK/6lKzRYMDLhhYSDfuakjpUc5pS2JS71rgI7UyZ9k
egX0aL0A/YGtnrig882ZUyBqC+CojPkaWxrVA4K9e1ox0fjLJg7Hp+RVI/fJyocGszOiAmt6vhSc
YPrrWYP55qRZQ9WHDDDLQm25fTPj3lGbLrblrSZiVVJmige83NtuuYZTAX9ilYQ87j5P+8DvDNXX
ieUlKnwPhpRr3P/iZz8iFLofTVyjACupLzW7UA6IHWgwHmNtm2N8X7sInmtfolbvI28IBLlR8B0a
i1HDqUkvPsauPuz760oGY+w6cKULSbZO/xGtlzzVdVGV+1+MUSiI8D7XAdd2zGK7EfyHCFp4YwKh
hb8sEVIo7YKrKfcgNEG4g6Eil7dvk7CYjtX6Z5x+2cr1XcELgSSIl3fDfUe0hV7ESP4a+Ho7Yogp
jpynyfSJuGUK33KF09h1M8icqVZgr/+CR/ND/WEKIIe01+69o0dufNx64kAxMLgMeVc+hFNq9gGR
foN4xbaZr2w75t1KqqUIzjaPkU/kPH2o6pwV5PHwisC90w6yJWJUqx/N+P3ss5w9ovkOKh/GCZwL
PdLnolEJa7nztRJiPTj6Syjcpu0iNNmnz1eOcAsLTZCTo4J+RBM28XdE5frveUWaxlDJvOTllikZ
zwD3MA2edrX9YrwILRa98VlRYIcLhvbZwEfARNe3SDajPCBFPQKUS2srxm6Leml6Hq/J5Q5y8OBV
457/eCqFZoAAhuZyDEelbIbak2Zc1c8Z9cL4hQasdKMR22be4Vy7VYP+U2xUzs9cOf6pXfosyRiS
6N3dkMbb4wTVnRN2p7ASREoTjoBDf+TSN6MFHDKXZ6ks8fEf5ac6p83yxlh4Jq+kLBUDwDeL/CIG
w4j3Dgtu48Vw5iC9BjOHS3cfox1Z2my19aQjiOC6WfCMc3goEKMaIcRQKfjYsGSlmVdtxz292xl4
PwLj/wnY6Q0zOGaAEis+4V1m9spt54GUPPozkA9YmrGshbpu0cBTRjacjc15tjp4X7Ros1AhRRQn
NRoyp9Kkb8txg4zTI/MzYqLccRbkdjdoUj6u8SPD1TXschyeOvbHqn/MI/Lmg48AmHVXrZoCBElj
NrpOl0Et7dq4VzuIydi6FojrFHZ9L7hiGGigsMPEVxcsPFZoherYt1L4I6Qydt3PapAAEHApgHVv
g4yvGQp539gmT2QOmPiHDW7NEJ5Lfqdon0Q9XXx4iFPGMfmVyxB/J3I07R6Zd/lVSrVDL+1/MGnE
LqyvvLXO0yP0AbkOz9JFHlNJxHxkLMWoidCGKbTR5wll3F1HeKwHUp2UA+hc9b4xSZ/mT/c8yijs
2Ys97yANb9C7USqNOIEFWBm4W+PB6Ge1CoD9bvmn7ENjq03nRrQbUARH9qWs3aCiBhD1QuGY7FGE
rLTeUGGk1bwcDKyMIB4qpD1Q97tyxiSElxINhxlPSjKfW/6KKG0YjVx8kD7YSbto+6AXODg3VINS
7AuuI0lyvseeFWyLAToLm/a9m67Vui2aEG8JaVy46dZqBY/9AZ/KVqjHJNHuCXr2eHLQoaAlxrGn
9EFQPz+xt7bFQtH4mMeGDP0MVhkaxdvE0WLbHDWBX35Fb8NFYAL+wzYf83+bcMkEgcIGTEyXCNxJ
7OeO6qMsNVcQXmi8xeXh/DOe8vPY84evZfNk9VmvWlIsNT4TXIYVknCk0Cvp2N8PZrffaTnjgsEL
b4V0hiGJkr6zCSmUULEaESiI9a4/ujo39RKraWzruei5DlhvLbzsWi5FZGj2q6PtuNc7ljHY+r7r
XgWcthxAVRA5mCFAGYDOnCEvz7oHZ5XI8CKv50QNTL9s6qjsO6whVDGUB1YW4kr85UWqefz9mnc5
8jDawqXuKm3YQWVoJzyumu9oCAc8BdC9ibAoqEsWvJY/fK9A4BRotvgOjz+S9j8rkdtajoGFyOr+
BPgPDcl87IoaFzGd45KmqhQ2VgdmY5f5Wf0Ccqhtt2Gm9k4DE4pm9BineJNncumAkUa1WE5GJNnx
iTVMuO9FkuXPA+U3zXCT8/1qScPHE48HtM6y2d/LupB5cOTOQ4P43bgX+B2gg6nQGUxmGJDVecuF
l+l2bfUbnaMlsvlE+lCMYpeIkKQ0SY57aLWaK71ZfupMTpGACiv45yjUHtLQi+suuARs35ITL9SN
mylTKS+72x3smwEHCq8mGbqwx1cxEMX3oS7kwfhWtUwArw8QTh8qJ47mzRBr0OGdF5KJySkirwth
32z4UIQfgbaHbK88NwPb0SxNDMOB/odhYdkf7/2OqhL1KEsheI4Rfkn0Ltqj6UJGfdlieSiPaQas
NAzohAfo6JTvsXVSz9vNkcWSxbnPQRYrZXwFqRPNuiCMLSEjIdQs2AXTas7iO+YQbfvfIP6YX79G
QBK8nWiEsVBuAenaIHYwpH0HHskeu8/pjkDoT56soXqcKbBs18N/cgyXeuAPtd5/xPikZ9DZGTep
3Q4LisVfbkyZZGJFNzbvl0J3pWzOshQAB0zLx/6KiUlPb4b3+Z19lRjZIeB1Y6ahBV8krOydV+B5
MFrOQbtSiHvW5Si9bnj17x2utzbogZ4ZYHDGNj/Boow2GWGwgsgAtNOeihhVoUstRriuSZ7LEHpK
pUorJ4dWm5PXShbMoqzk12334sDb8RufwAg5GdFeasMIeL9BBFF/A1fpkihXS8/30cHKK9t5mGNZ
EkxVX9Wal6CCTPl7tI00WDh1Ll9krtV8z815hEw1SgH+vDSjxbKEu7Yr5yC5WTy9QFpiYvUP0cN2
LorLcoZMxvCOApLhpU+QOaLi8sybXiwZQDRr/G7QQXShuKwYCtn+sdgdHRf1jkqDRyc9HyoL1fpy
g8BurStBhWcxLkxIB2T59O+ybUzh9IFkd3OES95AJwxtmmTi+dVQXwLeTR0oTnR9ryE7CcxlRXAJ
CVEUVjcodXvDix2JLe7fu4vUfa8PbWRxbXFoGChc+2ITX+PemS8iqKXKjp6NtiIbCzN1KVZE2qPa
GzuTgcPhZJPSWEk4fiDvfPXHZY5TlpXnCga9WCgE4I7U85XWPObHM8M3ueFnmhFyd7vZk3GD2P3J
xptrw8eaxRSEyaLkXUae29R0kG/n7gID5505HGGvXI7459b8g2NCGd2oN8yM9h4E5BfHN4eKbrxB
+uGpzK8cVzUf0GKCgG/nVkNQFtUIjgCntT8oxgf0cy4SLB5EejXhlxQhevzoedtDLMLcD3MeuDoj
KUQMIHY7Nf5PCH3UtHa2hibB2I45GEsm5dOpLZ/4HZWPcnlCD6V8UDvyEW4R4v7oVX1nyOVhpbup
7c80lJFf/j5jk/93r8Utdf0E0eDi/M2QQ3WGJyUjmcQdnizWTWAz8R30UaSLyg5zL52h+/CfGMIa
n3qSPcn9jcNTEYYbfnDrJ7Fu5nddD2Gu4I9StcF/OGeT9xlwcwuSkLA3MIbq3Oo5XXJE9Yw3Fs3f
IyadUBYKMud/rCF+B0XvsXyKrxMABq94kJJIUnCV9vZBwFMaEz+wK26CrtGAc8h3wNK8t7PGvXUC
IP6YdElGVH/rOZ0w9REIujqcxGXPYitoz/pxwlxREzu1ZRJ7Ak9JUCW3PKbVN5X62R6A6wb/zuEj
uYOC06bdbZnk1GhYjU4a4iVHH2mJ/O6BivoBBp9zl9OJ5AU5adx3eqYP365AgslUke9OXrvIuZaz
dgwJ8wT4ByDIQMRR7njBqJ/LefVN3tzUzPp8owrRwhMXxz7cZS1xzcHTshu/BcuRn95d1Y8shA0E
JpsulJkYoYeHXZ/WwojMbkaKhfoIwW6usdK2Q7N022IJjQjEofeK9ElZjoGYVSkt3eQyJuXybnIm
j7Ub6PzljPuxYF32AOPjuBDsOBRMFXEFtBDZhnvfzNzTXqSafcGmrSa3t8oKl4zLwbQZE0EtrnTS
QoG0t/1TpKh7IXMC8xO0vVfnHcpwWWZilb6CBdI+MhMRdIKgJnD8QD0cjuf6hGE3ZjlFRInFXPIH
0lOLOjNTe9X6dobwElr1bquwSXkpFgmO1ZWzhooSoQYeo8eMvNI5PgRlFeLSF8fsFc3TkGSygWuZ
yOkr2J1WEvAxP2ov56nKoeHMBjW+ZmpglKsnzJKuZQPUi3+tc+KWpiBMacsc/IiR4vCetbG8ROmY
XvOHWL1Hr3MxL8lreOs9pumWTyiPAI22EF0XygMMab+FmN7n/sKDuq33ubUx0MYQOW6DKdU5NmqR
ePuUinqtries9FuxuqqKnUxLXzXkgZ9sxwwEyaNecwFQ0M7v5NjdNGk8NzsUhkKNI4Brntjdl3um
2KuiL+0iht2jtyyFAkEQZ79byyGEmQ4oUjpSX5y+CQjWQKPMM7VR+2vcHFJHieu5XouuPuwFP7bi
uostPoV7U2vl26MNOxqa/ZBC3ohS/OvL1eyT6EXYYkWWbNs+gC3UAMyfv2DzIMj5S/QnvTdj585S
frk9KcZcH/GglcHhVelBLbrKU/Qmbsx+R1RVNWXLu8LJmb5P/wF3uN1+DbbC824tjRWH2biTVqM8
w9p7LU86IuBPbqS2/r+ORLJwbxRIt5pCX5Zrdi6DGvLb8YaFsS+jaH44VKOY4VEfr6EDdNYRMoLp
CFyZH0nK6AmGaQ66RWqfj1ZKBuoVZOP6KxguX6dwCWA8055XIzzz7gKsUYNziYgzql/5fGmLw+yl
sbHT46RoDCAK+zJR0tc6GNyJ2LV1nyGf14ydfnrM162bDWd/RlkqkMjoO7EC4UB0Ut6vOG/UMaSE
0SSxMH1oQJSaCZ57zwLQ/u0eowbMQEPCYCk4NPoLXa568vWv4WdjDh0u+VHhig/o92MuFREPmziy
6w2DtZt9jH2iBoMZGsaVPUGKIXhr7aJNFle7WTAbTWwGOnj2jUsPNqIZTmZMHJRhp8rcBrZkk326
cwIGcf83jG4h8c5MnGaAz3TCYhEGm6Fj8kOezt6BH3pc6cV0UNvYTzUSOhdO9bFyT39dgp4JP5/7
MTbyliolIHv6a2iq1Pz3thx2Pb/l0e1seLr6ABT51iDkxH9PiAwISrH+7SFZl0qeYog1G8l9VPQK
2QjmsqQQb/+8G0RdsEkKPtnErbKiR5XiyGPEsQRxVrZzoXxUbP7rRDeTQb8ix1/CzKw8D8sgXdC9
9ppmS77j3THk+N7pIeieqQ+fyFCrckAriNYWiVdg/HjskkSZ5noa7Mcfp5je+AQ9SdSBK719aLQm
QqFlmXvjKBwv0KY4G7f0khcHngNQpGXirC0b8djiME4cRefuPhKYnuqZWaCWjxo4tCGUKWfxCTU+
LUQVqTsqpyf++km9MlMOLHlK7AwRT2q7M9SBmnrZiu5zlTdPZF7YDKtTWMdTfxB2QlnK2V/Mk12t
ZWljnDTwXJH012CGYi7DcKyUf8+Hh5vp+Ahu4cZuylTvzxf8k6PPuHbAaze5DDBTJC3ZREGCPAWl
qzakPWCnIJgFeKGQtZrITXfXERLYDoqp7g8AXdQrXCQ+msFQZxNkJwccLhGChCDovvApwGaqRqRR
+XsQgOnLVOpxBnb/u3wn8wiWvNx0YjpLChyvCUEBAIedKm40YR/bwkXvM/EYCW9QuAlZWmBvqHUu
EJfW9D53/CPcgelBGyJwXyOHGZVonEg+9lJm+q9Hy77tKWax7bMbHicQ2IPyIBf9Qjt9W6ya/RwM
HGfkqOQJn2kh/O21NRE4WJiT6Ov+JtiQ9IcrVagNnjqilSZiYhDRYCms9C+YUMcqAAI4I3XeAQCL
D5icQS+kvmCabwPsFA24FgGDmzUhMeG5ok/kZV3WZ07a93SGxWS9X4Cx3I+SfKwFR+8GsIVwmXY/
w1gzDVc9lUFam7nUCeBzbakgHB5MgHdGo1NNyX8tU4H0ZRsSwRGYQ//LzLf4aHYci5OKQ2Hx8BEv
8No89Q9rOFHSD5OQL3PEfwd2gnnYXQtWtrLV+AY9OC0CrwALPZsYVRAMB2WEYSV1/IhbRzAYd237
1DNPbPTeKZZL08WYaghKrliQvEF25joyhUpZUMJ3VJyDztaYedsexXO3UsyY7aHyzdUEQtkWmPjN
ImKb2njFymu4hqXw++GN+q+LOErdjlyw1mqXDlWOoxLJ/egoCnWxi1oC6pKMIZ3iAvvwRl372R1X
ZLj+rmjhzXfxylls/GVUyNqGvi3AKIysyByVyx/78j9UC/lic6sO9xjgFYfFFiPLvtULq2a2Eixd
sLA83C3DDhUlmhDQWq9EVUvaZtc8FHxVSwMZEsSsrZA3Xcs+2qp+BNk4lHQ/Ek/2bkaXgInGUCWY
++sOtTcVn/pNBiEyZ0xp78Y8I/J6DRja4ow9onoG+kID6v7m/ii8PtnlqK9k62wZYDvaNSZWlVXf
Q47Eto1Lnn7FaIAA2THlFNUsgd4d3ph3rPbW3d1ueN8Bv2P76Tr1KTDNrwxIJbRCW1b/mZcyMZYW
MVz8X6jiRoQpDb7q5uSVM7ttVw1QKIpPjbf1jyaT+4nzE3LODGD96JgNOh40Pu79MN54Hrm81OFZ
xlOVHXgxwX8gZ8LUAPO7tWONx4yucYS02vjA+VmQM/XnC+hlBx3emBj636NKvCpC2v1ggdYiFg8a
yR2HvwKT7dugQqu1xNcf/4HV45Ugz/c11VP2JKOIbt51yWhB5BOHSOqSxk+Vr0945rIhNGMMUFfm
9xVYAsYfhokpZ2P/UJU64CzDtrDzps9eOrFk+Oh4O8vhNTwZfuFJbWiIN/l+gnKde03oBF0UKsU+
aZXYExBND/zEsSy+rmd7HXCRR48ujbxof79aVUv4OVKpH6e4hBzfWh2+OL3gf7ye1XcQHmXbdLyh
+WgYEPPIoZ6pGfi8uQ+V1lIOBAuAnBEVHIDF/wzdUabpx17n8MfLnVc5Cq+X/QURYgtxMitoQrVB
QXMho6YXSH23tv3OPjzXqyFlQHKB7jGDr2ii4TS+Nj6e/e2UYNuOpgQkgOvnUzC7v6qNBq0IfLqe
YaX/UphjUhrbCipGMRYl719gXU1N6jNwJ35Tm1KVHFxSy8WvsTGDqcB6ql4XWOS1Rq2Piewxo58p
RTMF47rgdR7WhAJ274vcoK9eF2XIL6A1269m0sE1akM8xaFDePvTveN03C2RW7g1PJ4mg+3G2dqs
dWHLidssJb4WhK/r2uhbBUWT3BHUb68sSpuNSgKEvG9IRazqfrL3S/FUcLepFQLJy9uej3KnNpgf
sh8J/tAEbsQpoSpBNt6lXl8L7+EVfUDk6jxcKR35u0GDF42geYiVLZ/3CZjGIV+/5RDTI+LbW2tJ
xreOTYckl6C0RXKclup9Inj8zpvthmjJ0bSD6fKGQ3ydkh1ULsxZNml2OoNWW4+q0A2OKl6vSWmE
mktpwh8g49dn+fbf+pD4Pfop63/I4m/smle/dP3RlyBPeMTHYrgJPoKcp1BDX7XLXN8jjhdL+nEQ
m2wtMfetrK4SsUEcmTVc07DRMSpFw3kR+YAnGtbT474c6q9+2/e7gnUuonEXVrKdq4sLJoBkxPn4
vXUqD1k672oPhyFuVMI3v3yu3Y1/5rXWA1eBvtjT8dO4z/8LQVyCfbPXnDvMyNOCsz2a2Ltd9L+L
R9kaTsukpjNtSsxFhqO4wWW0H52Pc/XiKuU8opiPoGkQwqwAjspgCnH67Kw6HHkcQ3XxIGQK3dsC
ji4c+6hVujhPOhQGSwK4pEzRg2lQ2xvHPvdb2U2n+ysItZvT8GRfTCXiesrcf46q7oxJ+gjsqL/6
OhcjBFqYbcVWLybTkIA+Rghc/Y/R/1BATfClV1gEjdOo2DnzVhM7dJgFLqnVbzwSUaN3hbJHwxE8
JhkJoloeDNEnaPzk6KOa3vXeyL+mxPGmy5pF8QzVJruqg9LpSHb0lbiql5FHix/cvXqi3cxu0g13
w3RbVHXqF+iv/ElxrOnq5XZcRlGoeTZ92pM8tLVv1YbSlbR7GYp4q8mkq6V8VCG80VdAcvsgaRX/
T7j9pUfwAfYHXZvTyUjbqDtAmyj+w0xhLPgc+O+YcBg+5IhwQ01vo5+JW8TUmO2LYgJaIa8zBR8x
YBwf8pyFjmt3vZDZLDTXaEK/bWXGrKKD8IXwKTMZXcczUEb9zqHScowJJJS2nUR4xmkNKi1ScqfK
UBH+NoYapzlOwPuXLPXci57ILV1OicOW6BTkvPDYYGlmvY4kKcDlprKu9oenlVQaeH1bi3q/ceFc
u/M+9vm2skKbYmKrqCXQmmMsWyOJZXxdEhoYYoSn+LrH+ID7oNtiDphepIgSvSt29FQf3gMk8HOM
RvTAkrsdCZZHSKP+MeMlBlI1HYiHwsj1VlV6f71tmH8wfHYf21PmMkhD4/Qcn4VCVp7eO77NdISL
ipkEIPktRDY3KF+9BUUkgCPJP80FwV++Lg72KI40mbJOtWZiYmYfFZwyQ5NvBxVYxhLfzRsPbFxU
pASQmi5sQKJDAt3C4KFrJwxBmtPthcYWAV/fa7Z++qD06rzze5VJtmHg4NFerHKY24HDn7fUMErE
uVi0nRsIaiYZjWuFiKNrnAU5unjJ1rQye5z64ANAo9o3LDNWr8Bsl+iWTU5YgEhhOIEjiiYPJJa8
PbRNhW7AqKncDl5llsxsYNCjKyOgswR+cfjJokZfdGMFNv23pNV+AwdkqMn/wTB8PeGbuy3I5TE2
57xa2SWc4AJALC0ZiJpJxGKaDrdMubse0znkAZEOvby3yU1+stnCTCPhX9T9+cnu9DAhi2dFIcDV
/JCEFXP//OruA2Ep0CBYODL8JmqhWjLEwLrs8B7l6M8fBc44MWDCRCdZFscV2Pe4FyqNxt87HACh
ustegMNOhILk2fiXsjiWt8LD6mNpvJsDGfbD6nD7znlzAaC7zBrlX+8YLpgrvw+dKrjnUu6JKDHY
DY1kTK3XeyhEshYDmHGyBaKEP8DKe65+n7zPRFmzyGHIGdjQjYIjzgGTcb7KuDn/dFRGxnmGDzcD
khsON59Si/ZRR6H51eGBLYQDaCGABecSBbr03TyTk618igNKLKS5HyafzgIRQLG3tRbVoxXlFyBf
jraZQkuwN6VPJNA6T1+2YyrMmdpdjTYlqMd87h0Y2j+lc0Af9reDwUQhX6RS2PHY27rBSkO6p+Y/
eKtZo1+PyLEeJEvXPQKzgo05Xe+r97UN3xKtHh/ClpEl2nemh5JFPLM/NJEvdM3YEb3bmlHw2f1i
TBpgErwQHJTQ68EqRt65tKTiH5K8rbK4TkM3jvAEuYgGJ1lsCPBoeRq9cGZlS4PYsEujGIl2nwaA
78Ab1xJ1CNVl+O8vLB4ZLBAdgaorZ4WnOzx3SFIEIj3i/Px9kgl7b7OBRyFqypknHWS/M4HO/Duw
iynCZHnwZ4qz+PvgJpmfluPkyqA4kDYaxBm4ZtmpL4dT11leYToBTVLBV0PLo4UJZ5EjaaH7M0qg
/99mjLFxOXY0GBW7aB/OIRjnEUleH3m+5RE5C+/iSduNzcR4lNk04leR34QWFVbt1ld7SziPpx8U
dqmpnsTgEHXLe/tmnFgrpVyy9jj6sx5vmkd9fZBvhq7iVsj3FGgAH/BQAhjIi6PJSZDywdXtsh8K
8H2Uy+s0vOW+L/FJGRkL/xQXjvwNfFCW6k+V6mKwuKHqiuhBLIezmkPVscpFf+ATZa8VFiAi+9+K
Xl8UqU7AuYZNWrUCy1493JP3zKcTHFO0KcR0tmxQustEYKiVN3k0qsnPdugjp7Sq3tDgR/npjPs4
njxOFScM72E6RAaUogRipuY4MsCIQ+NhRtyD9I9CiOJopW47RQkU2cYxqOZFnRFO6t8Up9q6MIgE
Zlp3BmVqNx01m3Qo4dQmCmlL4CUq+qxiyg7ljP4AXOYsdZ9Rh7+VoR1BHAK20aXypCxAp3KPUr1L
5D1poNOa7U3DNxtpq0ugGrab54O4mDpQoiXA3ZRiKJtYCmFpIXzCJwgU7YkZX5aRK8CRZTSRhUdI
8hb0NJoN5GZ+WHX0Y8wfrVeK69QHYvhBUu2QCpwJj0OeAYD35PKCnWDQ2nWzCoyTYYq6Lg1mZ4rU
PPpL3r9rZlb14rVAlzGHSMbysi8qVoBkzydYXFqNHYDSo6EZy4RUtElblR+euAyRtkgjRbxOZL7I
3MrgJ3h4xLISXZdvoFIF87VyucQsQgGG+QPrwytJD1t3BLxM1aG1PkJYrFxeuGm4273DoFcSrL+C
UPLbpKEawUsTHCWZQ/d6RnsECSBeSiDV/++o1XclB7AKPTxRnLbVmVGMppgK53a2t5WChgVRHriW
tCbYsllbrDk6OiejzLN4Udpy0VnSYiLmMLCmP4qyDdhATrlMUtF1eq2wlNeZaqccqtI1g0axsviu
53CewIJOET1yJrGutgy0Ypv/J8MDl5DnmZbchx0HXcyPNDrXt3gzZheciHtP14TWbVTO60uQNeBL
XY3oU1xwDY850y6eNkdzrwpOF949UoL9wtx5oDB4qsy0sOzL7pvAAYy0pddHLdxO+tIaTADqjCcj
Ia1KAe+2mq9rTMi66HJz2SbPBzaWTV7gr3AF7hC75jzapo2YrzfAoL2aDX1ATYvZGE4kjXO5eAmm
3Zfug/05Z2NW9ZxbMa0+swKl4v8Mc1XOYauqJ4LdWigxxZ0JF2i9S+hdnU+TeL8j3TQXxXvCC4bM
VRze4IcHWLDs1pYQkMFz/aLB76QFiQJg8KpICOVqGLdGsEUKrlTLggqBCa4qhQiZ1XXFW/XYJJHw
oIK6+aIKwxRQSrPBTiQvc1a800QO+DtTU1GSiOFeVRAOCO6gnVASettWNj2eAKO+dJKEbw84K94o
SAiL5C3Xk0UOsvBLVfaEUKkrYL6FazFo+BGyVBoLqIdE7u96xVYiYqcnRAja7J2KDc5DJ7VVkdio
k8NAy7APeocq6CrDOoDYva5aI8EbMhUxESzsEjwJSepY83NCU0vXyFWaG1TVY0nPqbKrDJR8RAtd
rfrP1bK8/o58rJ68HTbYWpZj6RylhoqnW1+1cmAjUB6jlOUu/pOl0xyd9lGgOGk9RZ/EjKLFUbxS
p8KjjmVq33sSDxYZkcygy5UYsPZAFiw2a/C4EMVcJ/GpbJp/WKwqL1TJshE/T62PDLsqiwniMlLF
PEGKY0t0XYdvjjY6Fx5hGoFpg9upzdFBAVp3h6nNaXh7b1sCnDdm9iZCloTBLpihxCqyYVG0XK37
QVfx5oMvb4xagQktegsVxpIKB30Eh8P2nV3S1AN8G12/JyVmHyPZkt8PuCITBQ47+CDUhWpzJ17A
aR7djOFt8OvSZxYkllGQj/sTFHJUkvG84tLt2DEdtjQx2Y+wCxBvGnegaoHmfmrNvwmSHa8xd0sd
kh9LIY0PzYUP1xiSBnK07J+SxyJSx8MMkzdL8vuu74hehPyzaFEo46iQ1CAlC7zzv/jcERHV4F6H
5/6Is2cbWsv1bteKh5KcidwThe2+Bxa8rwVAAn1iugBzR6ZhBqFlT1raWhIAenWp1PC1EtibLTO7
acH+/yPSW67Dbn/SFFPST1CuFx6zR5hDQXsE3GercszR9jLy4AAYmJFJ4iIg8tjoUF6Qa5WvpLX0
jRJo17b78+f73wUpTcaSjLBtkiShIlm/ykNmQ+JxRHLMPQ5VWL/xMYP9xs7lZORkRMg4c2gSsCKZ
60NFOlQw+RapIwhveXv1Y9qQyoziwOya/8RTvDqXspzV+K+X3urZL0qx1NQjQ8l9CaNli1mKQVKh
QK8xk7n1+xrncJ6YoYq3XOACo/Uhzol6hTh0zinEnV7H4x1XnngWphzOyHOGkPZg8jwQGvKvjF3b
b1jkwWoKCZ8SEPCpiXUR96qopCLEPyJeqGyyPp40OCVHd6yVVcJR9qU8iL12XjDb/Pv1vufH4AMw
buoeONFhQf6WcXsjqQG5oKp5R79dZt9xCpObded626h/9NFnS0n0nBePJWvagjC4haWXmeQOdlIt
/d0D1agFajByMDH69yHviVJKWtje/d1lMW5zTl5+JbowgVsuFUGdiqk03sDNhDcZpy6dABuY8xy6
OixrGkYTzqqV3hTU7VG+lMAZ9Im1uSx+er1Rsnu1PbJeIsICyeeoUTIs3SzWnYzdI3U0sbLWRweF
ihMsQqrx5uGCGVVFUUjA/B7tPH10gHHn0YleBZmSCTGdj8FM2eUc8Gk6fZJU0yQ1jJEebtXLS+SK
7mEApU9hQdjbOdoJMu2oEG7SQ6f2ZOPilRjQEOXrGZV8phWb30baDCoPfBtolkh/A2yTCEXObpk6
7OENeMcS8GRYjb25leBwQ1JkFB1HxA+hdN5Fmaaw37TWI17hVcjxJerhkyPacIRSHfgZ9/6ZXd69
ZbiJxJZ9qcX6YpSyfIM7ocRl7vBbolDbpzjtpF50jAokYepZmM5uCseEnO/R2lQBluj2H/VRIxq1
3ZMfB20Z9yGil06+IADE8uojPJEDB+pPYVaMeHNIq8wA4gpUDmcN2GqBxzhJz8l5FsSbaMn/K/lX
Ed0iccGanHBSB+x244iiy16RhecobIRiQ1UX9qaJJvmLAdmAkaDGYg5gOiDW+SXQvFkdxxBB4HT7
bqSAlkc+2f+6AizeTb132kmdszOzLZ8NLIsKMVWwaJS1P6dhIQayuQgjHmcpMwWhlezgZpGHwqu5
sxaPmsDmSDN2kcmE5aAJXY1FioTju3cTdoeZO172gBiuJeqxhxvMjPI3FA3Q9C29Adtyj93WlhUh
M1KwnXlp73iYZ3uE5pYT9p8L89MUU+DQYzPtkSS70y/BXxa/zFrYDjm0ZBSpz6DZZTJB3/VPRLMu
/fjXB/NYcWebGNdd3GdrTPqERFNqoUZzLYAphlUBMn/VugNzYS1ZG1qLdakkJCEHXzNyX82Tr5QH
+uKGZ3pZcKxgGgLfOzqmMoC0m0pj6n9RKv2Y99/9uVMtPJAHTUCz8f3o99KND7artL44N+HF5DdV
4oqggqm0egPcV8QPfMAJXSREam/0J/RVeQmg7vzShtqQHNescSnP6Dkp1djRhLd3wrTVRfTdMbJH
U3ELw/0lmQGHKyRXKRoTEdh/TkLHK6xqbDUNB8k/TVtJQyfK0AgzDlpscym3f7rT9PSynRUSAZfR
iKu1ZyyiALKBOX501igkfJGL8wRFATg/xJmiAS6oCeh7MqriT9LDoWyQlYW7dx8ob6gjINhAI3TZ
GtWI2iTegttTCg7Qs4DrqnBN3l7KP7SxjXNnOGNaMrOTiIQhVSsx4AgO+qpnOTbVphzL9HT2pcST
85kANADwtUFqQNUbOWPGZVpatzH4o/IRSDyKi+Qb0oys4EVPI5zlHdoTqnhPH0c/fKj4QisYOkC2
jxoF7wA6tAQMy1JDWEBh6A5c5xfdRvFONdVAwkTZZb8GOxtDt5VKITNPoDIqm5dJV7KW6vg2NpzH
WvSHaDXs7MRVqksx6dvwUBvcSMdzRcmwl7j1vkdn86SunLdBj3jRWKLBhuXwF85lI+fsKuLehztb
FOhqkDTVpOS3IZeNEGf8mMgeyNQuMaPfSeyFb3eyQkwiNAiOlhxfsRXnnMBULLUDzIm6h73tSzzi
EgU9FaCc0pCbp2GNcBn42S/5orrviS/MStfQEKO0wdEfHEx8zkAoQWyqLHhWdqQAvyzGL3a7nnk2
vi067HDGHDK2X8OYzCFkBKoBhlVSgi0o2Me3JZFdRs/GTju0sPn/aUHpCUQH/tia8lCRuLaQSUxy
7TElQvmzyXRPGNA/sNWbcv7I+0X6Ndwg2LdPdOSzAzjzv/w3jMXf00+qvO2hPRfpmoOmV8kOCqQx
ECpVq4cbN9VhaU6AqI/oMye2PLfQz/LAU5xhmTdG5HJYjQshPcRNF+BnqnMAr1/qVBQ3nTnTW8j5
VXAPHTl/vYALwXXwExY89fp/+dBO9OLlbvWHpFe7GCS3bl4OrKQ25pid3Nbsm+0hpGm8XTE3haK+
lnJ3iQEPloE5wm2qwkBfoRvgi4Zlbt+B9mhz5JiPLhL4/HnklwRUN3UyRA64LmULm+OvP3n9IaHi
uHXzLtAGhHbBFC9Em2Yi9jM8Bh9CrTFVguc3vkXjZLhZnTDacXye+dk30jD7j3bU1cCvgagkEyhP
a/SVV6QtE1eTNunWH/C84X1uCRaUsOkOMFH1kk4JSA8Nx9r+fVdyVejtjtZY6hl1X6oAwLkyY/B3
XFsLvilNPvX+JvwcI7H7GyjbXC3bTvbKv7sAVmBAxCZX0I9d+6VanLLKo6NrrbtcmHBIyGVZRR92
18274LQ4MXDbxdnpMpploQk76NtigU26E+LJ5Ej2lasfEwIotu5ZjlX/wbBwbOUWSAWZowC0SlHv
GQfBCMK0BGkPgxokTD+fl9gl+JlNBOnkN7KXD6E6K//96WJrBqAnUceCyCAuzyic2L4eIUiZfEjx
zbKpZP6MivWdEG8A3xcdh9KPFfqdxUJ8C4kf7yChoqMo4pyZ8/c7WTUdIB6ynZV7Pr7K7TxXOss3
BWvjKWYWNAXRBMPyLXPUwbTK5RgWv5aGqZGcGU1mGTt2C5dIKAsgXdqsL4SArZiJT8n6ZQjV1nV1
AXmqUrT4Sda1HmwCA11wDrTSSufsWeMFekWqHH+ISA7g+yqOrEbfPnUf8XuTBKijnXRvlSu6cyyR
pdz14jKQYY/iCELO0IjkobAsd1FMCBgzkHY3ycLmdvhVR2rWOl4My+LKdGEtxxVoyUKXye+48E8Y
jSXPFD5B5BR5dI5xvLVdC158ivZVCpI1ZYvwn6a4ForRqgjf+8KUd5l7CFI8GVnZ7pOYmweYBcqX
QjraLOwnQWIrC/7W5+rxZEtZw8pC6ev2NzMWsLBIYDbTTY2T89/mLakXmzxyeg9yo5ZD+OU7RKfE
14Tsx525T93f/JtYC1x6B5q+kFtvY+EwhRdZJKQY+EW8hKHdfrEt6NUjUo30hZzTMj2f4Xd2oULh
P2k+NWTt8XjydpEQCxpj12y5cRpZigs/z6TaPFh11P9FB+fGIOuL5Yej0l/+kqNk3G7WmSWz92oO
HEML34any4N8ykkGmoe2VxsV22QUTF/U7tymh8XPW091lFXyUSbCr+tGU3hLp1NREOW6Id7ieK3L
xFcJa5O7BNJsKLaT3B/AJtSL6R1juphK1vl3ZK4IK0U0gcYFmkAziw0J2Bmy78bG6pWTDXfBYrYY
nElHIemu2sa9BOn9XEbTJp+mgEvWzYJ0QomLGse/Pl40yGmnSRCjiC+35DWjVn92fcGGTjzPGDsi
iYUjmMM2/dIBWPV7/lxFr+TsZo0JI90cOLFKAlc541/D+YtZ89YGOvsBPUmeVMMXLLAHk3X5T4u5
ecH8PNKyh5OCLj6duZrzsewa3aDVFUODQjqAZSsxbvKXe7rl6wQ0w0fynARUtNrwJsGtNMAO7Gq7
+aDPXwTUj4URyV8jI/4tvBVzWQhGpSuP00ZCzQfkyq20osRYjvcyd8lKIpZ62fkLzDKp42a4+8RO
TG9+MHGI0qh/G+gcf60EU/IJkeNM2QZ5RuOoxXnSo/RstApJsmMGdsjHR51YjO3gnDS7Kr8fq6tC
AB/snmCUeG8AztWB3u/Zb8KkuoyVT6RNNmGhfzMN9jjYT8dcaZeE/Je/hiv2LhKQaVotNfCfkbYU
9GSacDgedrzWhutNbuW1/o1KOa0OWuF7bNJWw9SotgjU41hgOIFhwR8LQGJHJhc/avmmRo4GMGgQ
or/hUKtvQ2n0ius2xPTtTAswBi0lzD925JLT+BVMr9ZHzTZmDGnhEnVHmblymlG6dSf7X14b3VG8
qTRk4KgN/8z7ElAlo/SFSRQxHFGmzMfowORU/rxafJYNJ8pINK4NTdkh/vh8I4L6j54yDyZ7biXs
iz9Jc3lZvm39U8orWtrP13tI4Px6QuNsynsse/ErW0Gk5M1AIg9lq+XmvL2LzyZdQ9mtmd/HYklX
LxciCvf/lMytF3ts9qTKBHJzcQq53GIsdM5kV6F0NvcNDTisgIWt/deaSrBF4GhEhYwtnzpaR+sq
StALr2dnxhgbml2FHnza45ayb7DosQWXrl2KLL9a32hLO0ojfOSc3oYbgr5d/Y2nBgpr28UWA7zi
L6FzQ4gT8VEr3JE+wQl1aJDXYoL07YoKmOK7WICEyp+2sQBTCBgrkgD+Y+SA8lA/dqKCc+NHK7uA
cppYCSTAWBjDX62CIGbKUs0OkJDuVyYjbe3p27p48ZpUrNf+BD81J/EH5zMLZWBAzoriPnghoIlh
D4/HbNxn9QuX4YFx4N5TbK1qIsPEDbS+Q8ikiBIptF87GhcTMmnI2hPJTB2jG5PFG6lPJ9yCLF8H
Neuuxs6rmfzQrG8rHOFPhnUIEepCySWEb2rc0PswVHMMWNHE0+trSFN5csdrl0A89RsGfTTLN8Si
iNrAK4LDCI8NpIVlunTj2SJP8wyP6iHGmZl1WuH0vFZVWcjtdFqTVSm0dVUWlDsMaalW5X7CF2nZ
U9dv7DuJ9yBx/DWhvX2yqK9ey2NiqwgD6g+06TtVHFWbfmISpJrRQIXT8/sHL6LbJfCsO/2Nxjv7
ZWf4xFl/XLHSu95SfBnIbsjqt8YiJFZkn4Kasb7tSfgnhTOIF1LFl3FLGev60lOZBlBE2acbTk+u
Y+BgxjGejWmNtUg0dKYuywEdl4YMkvP88t/bkN6yq9ftIvIDmDjfxRmfTXBmv5MBnVN6UrrRho8l
kJDvr/WwzbON7gILZNBwVou3mfh+h2EoSmdyBsKtCB+SeQ2ObHvOvzmnzcrI4+4uMP8jByQ8w3UJ
Uu6ah8sif99yqaTAZJvvtLDFKfGTVtfWvgzPuEIy3TmXEkK355z9kGouTDZog0zhowk3TepEdjkM
9kLAC8JmUZIob3pzIdiDg1d+JZs9ILtTdJeIzXck6wmJ/qLTBpd5bWFFznUJHSFtg/dEXgfUKbNm
kyU/mjPi+Gv4HZoa0yBZfB4asUjKSRcFirf2M9W/EfxO4xf+8QUozef93QfdsiSBFs/c2+41b6oG
MnzC+Te8cIebZsMkt/dZfz07juc9n/8NiCdipTIY5vn5IQrX++Uqhc9XW7cmxzK8yiwz4NJAdi/D
DJfz9S75k3Jrfp4oa2hs4jfrjDpm0K1B3TyMNz/Rv9Kl1b2cx4QKhjkEyBq05gqkUAKoUfBXglcT
8WxGMfJf6KuwFLzbRyz4Pb9PLD4lM0rm1iJ7EzH8k18oSx7ZZOYVttKn9uSsOqOC+wkzEgrAfPPO
Tueb7PXpjNNNTmnsRZhTqmKBjrAEn19llMAuC+BBwFI/+5o1RWPQ08SIUgAuD1FWytyQ3YOpZm4I
VqofUd2BtRLRfNlA5nNyL0jfBU9+e7I/u1KNlTEPmHuqM2vAyyFfJHpwXmFHjVdeLlN7kcsTjbjo
0aOHxmolM7ZIwCYhU5hIw1XvR709uKzs/0XUYeuoKMpywq4GoCYFjnDhVF3SystL3+0BHG34JcNU
Q5bE+v7j/ijhGpKR+CsN/qO62jKeQXDzTYA6qsaumUAeTHJKGTTOm/XRg9w67ot/iXtU1yDQ1IQF
BXn2D7LgA02jW9sfDkRVz7c/T728OY5liYzhYGAaCg836DVakEsna45gFjYF9DR4XgQdLxUA3vGE
VvTRDeKvzNpES5uVN9Rq+UqddUnk0CL2W4Q1cVtQaO7L7x/CXLBoq2iGzhsQV8R5FJhhqZCl7hDF
o8ECLVZQXOYyb4tKmKvkVjF0uMrY5qOV7BJAIdprEMXkhwNfZ68co5ezIHR0fV8hwbCGo9y+mpqu
ENyan4snsmdrIh9ep5i4J1rmE2Y5nOB6VAD5rP2NHf7z7S1Nz6tDr6iprnHQ8t8PgDxt0K+3B0Eg
ds9ObMko/FtfXzQ+cR9hMpYtQKT4ilR56mS439y5XOdJXUJaj0Ed2wi+tmD3T5zn4RWNWuYPhvSc
3aGljzKRyJjsv14Ikhn3Xvybq1dXkzOj6SyMpwBsuyTV184qz6T6NKI8B0ZjHiY7e4nSHfEckT/9
LjaE2YFNwBoM6gRhFBsKOfVtt1Ww0NemELuun4w/YyXGMgDdhgr52QV1YuLJrGVQqaYU9uzW7bK6
tOy/pd1m0XSZ1koBa78y+DRXHlYnm7yJRVOGYCcfO+arvoXMLbJe1GD9NzVClW3hshdem+rvEqsH
sE/rYxA6kqEPDId+n7QkJawO+6Dtr1LVrSnNZncJ4cf8StMgbDSoQnidfDov8PofbijTmp54Kf0Q
r14OzrhtibSFZbnJUQ5AVojGjMSIfYtLEXd+7zhw4/Ve+5ukAZu8IMEldpvz0NaS5dHFYFtURriQ
vN8zQUhgOlPb9BNMYBDOWH5DqkavWrWsKG5gPiIys1/KWKcLPqdcwenX47sdQcFDN8fRXB4pxko1
qj7VjfBE/n5OsDVbYqCE6IJwbRZK/W7LlsaMvUz0KlJWEZCuPu/IxVPqjfDYsMiujzvCjaQKl8u5
l263w6CQal5Rpyv1g19SjKh2tT17X0D/EXcA6yfkXbajoE7/AVhnck0aiyWunLqCJM58+97Ueu9C
uXgnvBwgGMoCeeBsRqjon/ago37i20DX8k6muCS1oOm/LvQVwmo9jFKwkI78fY1TefGn5+gn0r5T
iuS924RJfPKgTo0uROKZz6bYcs4dJ6IanHQCKjPvM/yea8685wRg/sTUAoGwQNoF++fcbUmbRncd
rkeKdgCOSaFNpLBF8xq2EJj3CYTGcIaiskY1t7H6btFomlkHV64KVVCXBq6eLFLWzU1oRoJ/w0ri
EmVEoO0NpogWQmHCvY+83q8zfcsBooChUkqoyk2r3411b7TFq8B0Z5imZpzRudwTYvHSbVxpqoXH
wzqlq4rYpDmSNus6xyPplF483FwFMuFXKzhCAkG4U6pYIxL22PT6WzzkKDc5glbzuUexa/PsLuYn
fELq5kUv2KmdafNA+i26b4xFboNigNOjkBFQUtTNvxLjk6AVdScdt6S+FLLoQoNqWRfEldaYkC0h
lvvW8xfCLiiig4oZfyz6LsHdSSP82ZpV1jNx2hyeNQZm8jDj0D8AtAgn/etnceV9gPmSbeTNBoyh
b/udwV25aftqZlMbS2I0v7IR0dEeTE9UgfPUsFQnTqaS+bcUdSItAucr7dMf3MB/MSGe1XLrs9sZ
QdpTr/z7JZb5i5mDIYgoevZxtnIFAxOSjPyLzb3M9DSIdfC6b868APDk+Tu1yMF0CQOiEHgnxaGq
9YMD4wVbS1+E/oBsLhFnU5Vjm4fzWfZ0p2TBR+oGCWVFA5eo92vjUl0LXQUICfNwfoS4IrOE2b6B
kZUJrzxFXP7wzf/dAN6Yp1U2cVZ2Dn6L5tjy3mw5Sc1qFdVGv6uh7jUiWBK0z5Fwuwnybo9sBUDK
5GfUi4Lrvr5vKx26zZsVR+K6OCG5U9YDwiuJUkHpWHthnmYRpdVwRN+GwbAc1macJDvP7gJJDATW
r1FppOanj1hEHq8Mggc8Wu3Y+IyqXEEVe1n93vJuRAWRB9AE1GsOSp10Ps+U5e0GkimA9FjUtTKY
U7DP7SDwtqImzzyT6IHYyyCYHKWgK62/SMcSA2rRA2CazoFGVDDQXWzNcMvzEHKaFDMg8KnI1xet
2z6rY2YcYFnffMMJJlAJwmcJga3UbHYRQvqGBtfBuBG+rzmwwqrMzNyLoPX/p+vaucL+cdDISD1w
zfWXFgc7oukjXqVsDSKmNTGFNL7e0HMda5uvfDmqcnqmjlBRiuEQ5VBOsI3h25E2sXXDpsLbP+PY
M0tgUnetL/bxjORhzu00B3VbBhE4rkb07q0Gyuk9emytJihFgReFdRte5165p1gvoN96OMazDqpP
yc8iJPAFmEnsWV37WWmEQji2btf/lSnlL9uk2UoyaeUH5G4PDCIHwLJEmAzNvko7yfoA/g3vB1qo
T4CPyNxl4PdAx75lLcjc7tlv/bB+0z1P+ZcHfXwpSSLbjQ0gQ5bahacYWLF+2QGbmKDhf+Gzmtvk
8UCjJOH/bVpdj+7UGSw/GSi1Ub5z2BUrKenzKqNDR7X9sW/u7L+mdOhoLhuE2YZDfpS3jr/aPJv6
YnwK5opIq/PCrTjJrzHOwLhI2EozTzjp7qGT86IlxKGtCFSd3GRLZEmkxcGLp/OPJxt1NSQ4b9FU
dv2qnerBjKCt53C0J50ksYoOvDavTCz755WxXLQFGPtmOSdFg0JoM6CmFUgsVusUczFMwYUqlK3a
5r/L8oGddCu9xj3bG68c4C4TdD5YLDiCOtDy5KiBplc2cdl8JjpQgL6WTo/di7dES/6kCL27JZs8
6ltxuKG8481kbWYsIfJWlLHmN+ghppTS54twL6daRYXkGPrKmrrw8saRs1d9oKj2pnNocF/PghOG
clCPYdASRtMBqXzHcj47y+Z6VyTda1EoUe/D+L5eUKdeF8kpuYyeJcSSxfFqO41DL1zAzbxGa0mn
RtWmzQW9f0W80gsOTpbBuGmfUdZKCaX3/n4KHkkNedSrDRpYZL0anePElULeKd2AHphEyAuQMt69
qSet4GMM7VRQuuUVqCdDfWmAIZ9W9zU+/Bfn2kI8AmjaHMg8Qeuekqo5k6E1TontNklQQjR4Fy9k
EelYsybbw+2ewtPhDSnrsfL8yTqAhVOpQfDzmRBEBekeQBuwCd+KEORe/GbjZV5W+vIxowO9rSbw
AeqneN0Hi2d/aq7A40GPV1mjkbhlH/D1G3ppdWXlAwlNnnUL9dpwiy7yP+4Dfn2P8QWq1Zms/gvp
s+Kl/2aWblBnWD5xHwCBtH6Nk+ymJGX8G31f73Qb6KyzOd8+b/o0CXaQcvT2KVNRtUeSLkuEWY1+
RXvf4UWQY5iUKJhX3Bjateo3O2WnY795vEl12w1dRvC2ki2Uoez+ANqA0I1R9fXo+G9ZReYyEIKp
kKKxssA2ims3/CcADcmPmuDgYaNeb66Wr25sH//Xss92bypb2z3pWzBERXX0ts1jMlXQMpgreNbU
UqkXCwb3Vrn0+ZrmaYCMfiGbO9I8Drc7nvF2OyLFsM+Q4HNvPupEU3U2k40yMu+B0BDQyD+kGKp5
LDSKniPmclq0p4o6eyYmvBMpuQ21Gx1Vo6SfIehJN9U5B9D834LZQNsIi2TRJ03ThHuWR+g3ZvPY
e7Ys8xkOLZ669wnRy1lHAtNbcucvfFadFhM/JAIm+9Z9OfBvVlYMsW/Up5t9Vm72s6szGohSaeV0
SEl5AP7/pDiFacmg18ivEbOV8S6Inln4TpkmbTKKzS5V1lVlDlK8CWXXpBPEVYG8MF/3giMJLh+e
JT1bFYL+ZHJToZkVCFMKo8qBWMNpEJMi0hwoyPAmezeM+gqPdik1DmjIT8GbiINGNRkehUkk87XL
ufYOexV/3JPZcbq3v2Fh/NtvNtX6uz/ZTs25HHhBDtMZTOehHfot3XuCXXiB4Q06uZOU4LOjegVh
dm15AVcEq0zOBrqJjxjVvflGv1YHBL+5rOxgY5/zzzWLfvu33Wz6dYrnZ5mxn5bLmFSKAYpGcDVZ
kwgwA/LxXbHEFbKDEn9XnWXx4c2xL77fSN4a6KodrxFjaXxsrONYtTstwkEUiDVryG5G35RFNmfh
YxWlu0/CbvNSNdkcr/zDoTdSAfynOV0HacUBNufij34pBfyRdR/0nvxKpXgKJbj2o26KqB2WS493
7HNQ3rpWPyd2d5qK5azRtHiiJu8cHmbhIplgFL/dMYMMzGckUh3TTO30MYmauOY+SjSfeMDLwcTu
l6RgksrvsVPKH2AUZC6bwfgYX48NuNzB/lEjaAZg2Xe2hPM+tyEj/0a25K5+SREhmklAaTACNFPD
pUmvi8PMC3ekPTb68VGQ1ta8U0yY/NUGgYvG8D2kRbh6b9srjvPKWvWgCx0/HR2FFof6jBqOVNpp
N+8+xstdeiFRE4WYlLo/wQtvGmKZgSgnXeD50BjoBuKorQpa76pB8t4o7axLUEzS6YTU+afMOxb4
GLn1Pr8xTwkibE7p7MxSryjbH3ZLwCdx5o37niQL5Wt7NnVurzqnyISLkK0sxs8cslD0YulZ3Gj2
XhswuNmlFGgQ4Cw6C1snWmZdV1Gk/oLR/ne6KaysjGT7hQo3YHLya/sHg2SZMFwAPkvrBTi8IjbT
XV49izq/T9SyIi8rcue/FwaWwmRH5Hf/hYYnq2yc8tmvBF+2KDVX9IMTKp7qc8VQQx+xXC6gk7z/
juqpjiPYhUZnhlbxGPE6/LRQrgoslsaEV//PjaH6MOyXk57P9RpPHNL7onPjSEUccTVaQDT5GyEj
jrX7+jBWcVG/jBRx9QlUnaUHjPhgRVtSP+WnXkLhR1TougCiTnI85vYLqEIGODlHr8+yo/x1mV9M
4Irltzte+D9nORzmvB4rmhHys65vaXpDJF/5x9KoOWo4uQj6IVLPh7nH/gC+Xqr7YZfMX6yBO+cO
ZmiKGZkQBhqy3BhtuI1NjyvKiJEUflJnEGCaLE9eTIt2kNw2yqU2ofE3omkOoW0CWXI3+Az2hmCE
jyPHwOB/Hb1Rdq0Hlu2KS8F+xNFc8A4kdhxfqb/s8qE0wbMmGJUJekqIsCw/YG/p+7EdYFr66yn/
hL6wKwLes29KEc9mbxcR/sHGyE8YuXS1pyfCEPCfeipD3k3fLuXjAnKIWCv8YSH6j8TcG3Xn7T1A
4wDrP1bHcs0W996TAx14hCO2C3mAI/9avkNe41st2joGRTJpgnHJ2+XwFw+k40GafAAdoKZr2nmI
Z/nWxDE+6oCLlzBvWMXl10iBUbkqII571KfWs4YCG+8Qi/yB6RIdpKKhDB8cvvXwCQUzhc9QhA03
5xwMRwP1fAlScb9lAexr8EPRRKopTmCnJ+nnkfclfuNOMMhiRo4oxrRaOL1DGU+qKh5hnrr6R3E3
mVIKaIyzLh56/E2xUvI9QhNCX1tZmgiA51F/M6zZhPuLnLjdIY+dxg3faNqe5CRIhNks4mfkp8lz
Y5Z4YE+WE3ZvE1BkjE7nNQ4dCiuypPpJWWaCc5ODk137bvOhylQkq+C2JQ3toupXt3z/EEnBEdXU
OtzuCoRMT3FKBWOCyTSpAT1++BDHRXy+puDFAtF2YBQGgCKi9uCYhEMY1yhTj3FNDL3Euhsp+HJS
abQkSYjjNiDnJu88y0TJnSO97C4KAWDvoc67vGBWe0E3h8gLXpWbqRG5wszZYWbZlSFpEokdZzXD
eUCCrq7aUA5cRawWD8ColvFHPk4xcQnPOc8EDI6TCN90UaHWq52XdjTjbPQLE3wURZ0H/k/vi4b/
pYj+IRkzs6XjtPGLgmqUw8nJAVloKDeCjXSYAr0fPg1LjB6jm3ljoa+T2REqzwRi0p3iyTy9Zltg
KKh/PVMIfWfeWUDt0FEIp2kiffvVHf646+b5HnG7XNZtoCNM53o0n3gu2YmsvT9uFxVf7rLzeiPU
KzoiEMjYBLo0eziD1cHMJ2I/MDtedG/k9JU3HQjVqqwD2BU0mKAa3aaKGw9PGw9QLmuR6aWPb4oK
UyIsBknGdRg8WqN5B1ysYU7AXwVUSqGoYggBabkJcnxXY79yN8VU6nMpOhycuaX59w610T2aAKs0
nfujYjGSuwdIe31CQs6BMIfxEmRdbd4/gsH5ozeeit3Bnq74Wo6+bMLwRL04d0RP2e8APu09c9gh
aDSaxU8d3xs5CO+QZ0R3wHwZzp3ljMxDGjl6Z/H4Z31EzwnCVUgyOiHqUVtspx2PMaA9Pr1hXmMW
Xi0UKIn5RDpZCAsWksB9zIdwyn8wJqHop+n3CBQXpNvs/yEDXe4t+brmnZ9E8gdd62CMOxH6u5M9
STokQksGDNbopr67dele8YUPOk7/MtuzrcexKyzqZOnLw+tq12Lee1vf3OJQ18d+e53Vtm6aDPue
Zp0r4Lxaah/W860i9hbPAw+fu+0yjzGLmwUVinZvUW5pDu95Zm6H+1Cb5Jz/MrBavnwqsNLr7ovl
j0VFOa8o5kXow9WeqHdx8wq0c1prYC9y+RI2DSwpiYjG6NZDAYmpToVz3oqJfj+HGdShWQRKk0yh
KHDtQTjgUuw62gkqv8ZgXzwqHpQpV3YWqubAaRx0NqVCVl6joSy6+GT6mkGnsMoON2dKSRc8lfv5
zsxv5uFzugHSXliWEQDDgcsG34E2gaztnYTjzkxffN1qO+dukaKoj2kFgdUEfH7NAwsuHA0agEAI
gxMrp6J2FwmIqVu6FA49bNqFndrlTPnirkvt7L2LFUHJoY9g9Ii0gCihc5lNGyso7FUaYQYagyKk
yQANeJ8KKhvKEacZSdAQZLrH1Y/LyI04qQyWZmTOBtIo6H1SzOKyTudjsVmt7mgWeAuow3i6pGS2
QDOjY/e3c5LE5iAtSxTUhZm5AdNNjk3jpC71mNaV73dPl/3vkg7MWDj/PcqNiYMXiYr/xqIMk9e2
Mg0FUNBmF7dobVDYKMRzk/RM+GPwJPu5bOhKCqjHjl1TVIjP0ndAZ/Xsu1e4nVVyDXxxNKTSfPuh
Fs5W4UU9uapTTSdASjq3C9axs7pAvFmYY6NM1jZGxlGst1V+PqvK+SI47jn4vz3Na93uFWu+VOAr
+84n8kJx4b85yWK8duPIZfVlven5bkT9ts3tF7NHqtmAb486hf4IDUXU+ND44CJx1u43LU/ocN9B
LoLt1PYsECliOgvH68oaPAckysOUd6n1dyNFIo/xJqnXDOVSkOmSzxsLNZufAhy9FM0wbq0EQ15g
VA7qitDY0Rc9Stx8c+WdZnfW0zQfLFDAwpNZKoc7YLYVKJLnixEyw/ACVQoMy4ZSd6S2KC/68qhC
wQJk6krWiDFF6A5nwbmdqUvrMutNuRuxyUursOXF9RCeVuPWcMNniPULy2oV9W8MQBQWRfb4/12t
qgAQY9zGUssQq/lAmr0C8RVfPxfIcy2sHzuHTkoQdGFIjMkqrShvBw97VV0sHrzwUzlHCV/toWgc
VUhl8ChygAwfy5esJeon+msfaZGHBXVQ2W87hnldBpeXXHAU4+dHVbB/zjMgM8QRnGiDXvXhyRzF
MQUzyfuFXYtaAHv0BkG58tToqoP5oWwwCwiXSWd0YRca7zbLlP/aaGwmxiA0CJKQlNB4ZNzwKu9g
KQnT+5tq0cJBI8YTJ0MY2mNkhU+S5KHLFjA1qH4BnvhDC55cPnlhA2tteKLa+kn8rUsuYoSTxFJ3
t9tP5JUR2WXoU+bB6mC4qxJr8zvYRyhJ5JI/dDiOO+MjrWDxU/g7iJB4eB5OX87QEa+2vKsvA8SQ
lpiRy2iq4wJ8nunx3pJez6MEQ7T5KJM8C6bm9v9SE8u96bdZFCQzfeVw+WRm12LLxp6kpnOFch99
4Rq3K10zdrq3FqzerJPcXAT1JMPRy/Dif0IMeRHPrjlzJ3xPWVDxd/8r2N9cQEnxo4iJ/7qLa0DD
CY2aLKTGbig498zzZNIpxquyK1Wilg4ofvbrw0cmU74+5cg2NDa5qhPAZiUdJSYq8ztMnurO3yoP
w+c1gl1vcnXHcBs+rqLJmZdxvHqyWn+VT7+FyAjhbW0ipa1ytMGhKSnw2PprmPnqkZNVUjDgZWb3
awjYhwV8/tlQHolyoJhnrZ71QKLPdSUdTnkS2rQi+eOrPvEu+U3CiB6OMq0a+rsc9jfVVmpBmNaQ
u2Ghhjud4Sm6gZ1wcjXbUX/S8N2AibPlUFZ/AIpOeP3Msdsg9HvWl9s3Hee2KMmGLZafv6hEOd5B
SYP0IXK8QA90AEBp6+Rx81QEAJUg7sMCUwuI1nzQJBGkdqG5oe5E70NoubFBG0doTQQGtQJQSAUW
8dorwB84yKY+bg1K5PDhN9FBcBCwOb9nERCW46ht7xczqOOaZ9Eo/orWRF0lIpAyhXhVWRAf4As1
qw7ITfCZsotRHH8MiudtF4s70M/ULYAK3UzYvlUrQXqodm3iRZw2CPHeh+rZhEyDe4qSbPoLCNjW
IKWNOzqmA0suWf15IVWMFeJJYGXZANyAk3JY4mqzNr+g53aT1YAdrmjsvLJCvfwzMLbi0XnFx4NW
VfX5IlekrmXcxaoJLAiWW7zuONNHBfZNQdLuf8mZtX3HZixakThW2YPSuvtpSwBb2RnG8/JHaxPv
yPRof0/Q5eHVKWZOIN3+AE1T4udsXj+FO7UbX6tJfn82KFa0Id5aEbUrigPWR0Wn4S15obJq5y9B
YMlNeWnbGpXKTNUiZc8lqn0QbgfF8pRd9VlEwLonfoTFPILPi0sNbX0SpP31/h0QONnNifgz53aF
jd7bA7NKu/oqI5H9WW6HwZG4ZKak99hxLY9wjzLzJnnb5hLsOwae4uhDVBAuilstx3QVKjRmQ/ld
GNqNsQdxIktBjseTIo8dvZwPWwpK5aTP2vKP3rKPBL/q7YKuTWqhNgoYvswcn9cW+u8atER11qUM
RIXcpAmy1ghiP1IDOPINtmp5Tg2/ql6s7DKHjgsCiP/L5ydJ8XyGTjR69hBK1AQxHfbzSAiA53ZB
hiQ+1OK+CX6KEZh+mgJF5GHannHCXuSBwktds18Vvmf+hw0TvA/pccAPPh3C9MpmPS48Aa92e2s8
3thSKl+a1HIVMbPfxgVn/vEdKgSeksVLZ8+DZEdXB82dEROtE82bJFKpxHUtbuIa8Tp/HtBgLf9q
PT6T5KGBN2Tu+je5zdIhHWzCd6mAtLrRgjq2UBxewTh0CXCXCa/ESTpCMkQ/QWjTZCxPbfWjWA+k
EmGpvEbz9SC3ss3H6otCLpQwWmsOtqHkfwnYsq6K+HohkiTr3aZ2/Xmnm7SvrESEEIaj9slJecRQ
7Zdv95KVyOugvlCtyZAtkb15mgQXYed7BCwrRwAFGwyFX8ypUUM8Tfg5IHI8LvHNWbu83hzeF2je
7hJvnRWxOkIa+CtAsyUO5YAbMLTlf1cSyggOvcuOLjuwzMADtePNRfu1Ea3ECTZ12Bbwc/VIkvp3
u1bXXOFq2YLoJUdCYf4g7v/QT2HMIqeVrs3K6Q66f2HHvVWNKjNDF00fEbkmCF67svwQdPPzju0Q
l22rFVLe4fGBuH7RNZAZKyHQm5sv/qlU7pbGioA71t5Y1Vna+FBq0LomfObnBevv1kd9lV3FASeI
1BIZXugqyBDpjw2fGyV05OYCVfqxcLfmMIQDYmCfrZ65ll//fMynmDtnov4y2bB1csD42gulDYN5
5wZcN7NJ0Xb+9LjDjT+PkanBC9z+6dIUH6h6SWfzFf8jwAJfzLwsk+xIYp/RKJ24+IjJLQ7ElryK
4rWoSeQHotm9ic14KCUa1h/GfUjLhL3dPEBF26boopALejw2u93mGPTcmv5X7wdbG0zKSuHloCqD
J+iM0z4DmmXHTf5UMYbrDoYtvb9nTxjXtz9pRXNDJb2CnmqG86pLp9F8rdJPJLl7kXyRMtnE6JBP
jwXT7556PwklVSFCURqYDhHDYDNjW+8RewslWzw/I01g+9tl/JIOHmu5FdJY6lsw+6vgfWMstxd/
5ErkNJp+5HqYYuP+NBS+nI8TYuGWPynpOvTzAfskXQDsKUpoaHopKLiJhIKciZRmYclxtNDQUJBG
I6mVqDAvAaBpVOhwRVfbN+B2vZMzNzvsMutqCSHvIhLRLt9WtYjm4aBEjgcb41y96Nc3lVP5GNRq
LxhctSFVxOwBaL29sGBV3uQfc5XZmAs/ydVzdaNVfvU+Z4E1mkt27ocPH+fw0+HXBOmwNGY3Btet
bAraiIMxsLnsTX6Jvm542sywFztf69GH0ADndjYhGMF6Cdb637FNOXAQmKbPQhYNQ1BnqzLxI2wJ
EmCUSwFvUkTkXvscgemn9vg4FJsQb9zG0LCds+FKAnMLlYFE2dFxqv16MtOpmxCd7Rc7CDq9Cy+b
a6h0/BafYnMscPyoJA6F5Osa54ZyH0cUSj4wvL2aU7NGRDLlSAqb7RkdgzAig3iZpS+kEj+Mm/A5
swZ+lJ9JfvDEc12HadPvBwm41I0kj2SJ5jp08xlrrsrowZutDlzgZu17DQjioGmNL28pF32IcBbk
IcMaDgxMgHDFhy1c0qtARe/zS3Zyjnct/xmeSCC3lRjW6MgUamNg1msyJVEsyZn+skr0CtdkrIA8
hZy7Aznb8gAnXO0/gTuJ0FN0BGikkN7EIbcjku37t7KdGDqohu3+tWzatuDzQV7SSleqJ44XuIVO
FD9YqzlTXzXDJQZEkxnVEA3f4PDmrBl+ueIP/iiHSwZ+Mt0/3c+rIsigWZGLK2MFAzV5FSHQfV4n
GMgJW8YcDNjCyCi/ND5GyOOMurDn9xJJXtVzHsW5pOMKIh6uGYpGap2iRDMAcDRRuI/BEap8jihz
QJHoyj2jhdgsdacnVHi3cDqVDnbQA/lkfGtnsSiaIVPgdfjk+e65Vdzkx3UNPCWcc8hBPT/IltRO
Jxq0hqZZ1jfnOpln2MUbMz61f2HtLvWklWHRTWMcgOFdxM5rPjQChxPgivdOTu+kOlTdqBHwUWOt
0100TmUolXS6E6TKudKpRceWT07EKlX8dqKCJwr/tmBPyRtDkvvoz2DsQYoGbz954xx/U8Q15S/H
6/sGMyDALm4VDzz3hVYd3QSZovKh/sg4UBd8u9OPcN2I7DRJ1UTfMR438WNNpHAS04m0eAneuEjE
k0OFYvlgPqkfE7ecPXEyUcX805hcjjnukVtoo/D67lEBHMDfChvkI2KEY/nkRzZC3CAXRJRINBt4
1fm8nJs424SDtp5iPexd7y5em9w24gxYlIY4AHUx7eEtuxZ1wXPYqlw06M4DrvyC3Zz4Gpc36byh
2NWJ94cKy9bAXmTtEOk1q7LCmIaQXVqjacwENndE0kIXxHVoRuwp1ovqF2r4cK2aUgiF8NbduaZw
4eZwiBXj9gFarhTrTz4uNByIQoCgFAXkhHHVjM5ANveZZVSdZY/Zq8GLS8RjpFoB2zmSQ0Ud7inI
UHsNT2ryHSAJnjacOA0RoMMpSYF1jZgUka0ndBNrRTSRVzwOO6kT1E1JOUlNZB+Qayni0dgo/Mty
yymVmBxBWEh9vaGj6R8QlV0saBgfKVxHG/8hzQB8+2lqXQIKViI9NZ85xOe8aZdi8NLXvvLCbpLO
i3Od6/q3AuegUYvx9NJkeW3gGHB+oUxtQoJHzDF3mvCREVPGJBKQteWx6uii6JNdaSszt2nNYTz5
p8FXyABBNQAMt4Y7SnXCrJV39NJ9TIEm5BYTBiRnSUODgBbFJVbKbLTxH/KEilwI6HIx/58Si5Yj
xa5MGwsY03rntVWbss8AuxrGBL58uaWdKhtOMFSrDmaWEuIhsqJDuDc623iJL1MNWOfKJXvEVv27
Z4vGm1zFxrqtS/3D82xA2qaRQK0GhmFdNy65tnJMz6kEFvK4jffVW9MdMdmbNHkwGVweaFH+CLSc
JWN7Wl/v5QT4grwzvYLGjpC30OWqn7PMW4LUiGBwL2Gt/hQB6S4psNrD/m28L/CPiXlh8sT1iho+
sd3FIFUYbl8pyS9MO9QdhwoA+gEzYGWEXVoVpLnY+ayjOQy/z9zaaFDw4uDNQELacxhFUV07dpDl
u5LuH2YUfLUvkUR8XGGnrW6s3mYL3QDB/8j+dXrby4eyc5wxi1aEzrpeHBrFSTQlwbooyKbaUdNe
maNFMaKRrctSvSrT63PD+dPZvEDeFh8aDgUf8DgJKxCriq8OesheYmjNAC6gTdzRF/yrdlENC1mD
5AoYFlvu05Tnc/4wEh0lW1dn9wKL74o+ovL59D/3uhSClURRNnCR5Zz5v1XwgxCaWUi9+5GOck/C
wfJduH8/vOIbzd3oo4W7ZnOr572KtlLfH81WTTyEHy4f8IIqg4EhxegKMZD+47It4g0AzkZwA7T+
SU+Vv387OYpdZUjDmMM8XUEDlREzf87MorxrpLByXdYYn2BtZze8oKPPW9vYvQgL2Cw6E16cTn/f
bnyrS/4uxExxg6ciTqDencLQExQZ/7JpUr8P14BjvyD3LOugj6rf0w3YQZpn+JOHUQ0GhqxnxwPx
tNIdAviiqqp50nY7xQB/WPpohP1GkZbNZJGjEynDDHTFgCIB90xbGkEPo0b+4oQuUQCVexQ7zQWn
xCTgdSNcPYE4HHxOgO8SKUkVFP1+Eb+zGUbxo4nsC5yNHNnparEgrPHpLdybkUR34hXNbUKJD7yx
MIRcOh9j2ZRBGANGInHPhoNtD8y4wCZBKqDc1GgFo7XN/o6RuKrAG6eaKHYMTi1ghGFFBii8NkEM
RfdUY3C9WeU+VQWymV87P2gXmOrfLhhIRZspLgPg3Oji3qPtDruH50g/puwhgy2B495/pLjwDqus
wK5GVBjtSX+eIS++WZq2m9/WmE96CsB1VXdMI9A7ABa48Mwl3dFruoe4Epuxtz4Rr1oUSukYdzU1
9pSl7zrzyr0RxnwlFV47zLQ0kQoPQwVmBXbwkgIRnEBocrl/8An6FmEeN5D4EVY7WUlosRSpxbkj
jhMeTe+ieRJubQ77E5uAyuAhA4epWwsqzFs7PdqoCPeiIR4zIu8gM2Namo07zsIvy3TnYSMsjOOX
kwNvhQd1UqmTuLCqMctEm1sQY1WDFR0//Q0FkK6CV+m8/DKD+fcKf6GxljgS95IYcKbDm5Vs6Nba
wPYE1MTjOMV7/DW53diFonrPCH3BzSexsggF5IhU9c57mmrcilXS47PZMcNiAPEbiVeDUAmVEYmT
L7pQQIIRlwDT7j/GYWjNbg4WKQfIxoo9zHDzqM9aDdvAXXgnK2DQCoYhUfq8rAJI0jfKT4hr3TwQ
FqfqlsIIevAIT2kFad+JIxQnLTTwhHEgLqF+5zgv8eahMEfQ2xPzzc/oMyhxTVLF9aQf4pL61nP4
EMRDTVx6PhOr6wGgMmEOiQcs2AI7G5OkIPi3QLTZVjMEuJkZjh9VAtIQHWqM1bEuVlEsjJdS0cLf
tvHz9tEzwQdAQhwjxiPUE7Qe/cjgvsZs+1a5kjH1sLiK5XM+M6OSV1xE82HhOeUL/TsRdPjLqirX
CoPb/AjscNCQpWky/TRBvIxvHXIULPHAc22ovbQsiGNQUEQjn2IkvSct9CBPvAWSMr535jm49u/Q
FfsBGMyxg7FsDKvkboSSGgAqmFAtV1OmYdVs4Lrm3FAJH5/Q2irdcK17+SlvghOGOE7qDvjlBvJ1
DM+B66nGDYcJEMowwqvWiVXpQTlRSGPxhopJhLOVL5iRMOLfQLT3nIgwqpitLhNVOYMH5DtH6IFh
ZqH1MxYJVJEBs0S5mCSKXuUCZaPqFgAzbhM2B8Yb/QO+/dPM0bMxUtKVTVyKpXrRu+qd7ywZD/qG
N9s9+JNmtPY1v0TQEQ/VdeSe6UWPw0+6rwes7ieeIL0TAEZ/2EP9dEqQUcpt0xYcM3aP2vJ4y2LL
sTTe+pslbtHJ0C37lewW6zwpRUWypIbhIlaNLk0rzEPTrnipuatlkxumni4yFRCjlmGfZT3Rdp9H
3DKVRPSnOxJlonj7jX8ewyWZ2asfmC/tGXERlE3iO4CnExaH3czvnuzkfwjpGdn5X+C6Vqvud79E
ufU7MZ36KEhqssjmFRvahrc4Ta0GliW9p+8k62PQJle9HU9asUUw6/tJYLrqaW+IF/OCovgp0Qrk
OY0hycOS51ISDHvp9SnFK3WDFz3ty5WoB+i6rK4xnLNecvR6BIrMPpOIRMfF+Jy0eJRkQujtV5GR
0aYE4jsys7sVDs9g1rPOjuHgEr06OUORtIF3Ioba5B646I/CkEIBgTT2LZFxk9m+9YNM5XzvhkOa
Xc3FyRwlCqXKrewFuB/2yHfWuG71nIRDJRd84vzfsS8dfQXrdbF7LDb1/xA6/GLlQo93co28o+RT
sD+mYVlWSmFq2fFAPCLkLG5tu8CV01Me0y8J75i8otDBgGYUYuM3WiF+lA0fbwqRLtK+6lco8ooD
iBP04fcO4FNdBAfe2xvE54I/vVeHAsKXCAtjf+MVUBUt6r07wOQKSTB+ldeZhd/zRKbL6kI0IlAm
sHLnQH6YuLE1aKDgnR826ERkhYCLyolHpUm8DUv+PDYossw+P+CniRCXhYxI5bm/LihrNz94uZoh
nX2zrdprhWTfgZCuHGPlxUO55Lt5bLzQzidZqLztDgE73cOGKlsw9q6gWmViZvR6JNdhN2fVB5jF
LtEMEivEuOp5DXKGGqzZKfBi742ZnGs9NsRzDV+lUFJVT3bYzpYOM5uvz894lJBXgn9JvrjhPZBv
QQsvKW/BtHyXxBREp8wqXIWZgNpQkZ83Hcp/WJS0iT6WxEo3usCXMPmpAfNR7KNdwAxIFHPTIj/E
liM8EpE/c0SvTJp1ynN+YjptL7x46LTnuKmF80Vx4gtvmW91sVCyI5yZVJQCR/nEx8dSXn7/5EbH
XJUvnTHXYJMe225yiPIumzzg+fkvC44nw0SJ3wRIOB2qVf2aN4rrH5FY/uqesxW/AWetOzDraL1D
KUaBAjUh8RGmpidNphMlETfHpEWL9u5XoXIKXCx102zHdyz+EAelbDSIzEzEwTpP+PL7OjLAMziQ
tfVGpW3wwzXAIT6Y6dbq0Ym1/ZJeOr/DXMWGKhgS+lwXJlkqekQ6mXKlLiykplhNvPn1eKJNwkZp
OZ7qV95P9yTtm6jU1J8OrLYHx3QWeSjnNP2vNVw22hbJQ77JqL8MatJcl+6twu6CJ4QVgLtbNQaZ
aZlVdJqGw+fk+ZmoRzE5GLlk4zFA8piDjts7rTuQiicQI21v2KI3heDZO3R5rlZTWeDCnRG/OOUv
EEL1cfJbnOjh2hyqzi0gNBbg8v4vxLdT0rI+rsgG9Th9rV91ej2b8MLLs+a0md2RACV7509C6Aij
aJxIa8L2QVlf0L8Qm+Z/7N+S5WPh//xzZNWIDX/dp4aBodGjvx3c9U2nbuHzR4uU1vwTGjod8I8D
LU4LVLlfvivr3OH4M8KKgESphi4d6vYtI1nusPeZIva+eKpwOO1fVlsduDGR94g0dwjaMM+uzQCP
MjaX3bJ6KeihmxnX72PKwVFlS4NqYIoJemktvcXnPGTD6tq1tWKePEJ/fbz0g4bnQo4t+U0DAAar
J5m6wfGYUgccoM9/zYi64MfUntfuIrIfTEgIRdhQMDYgO6QQC5LiBui9JxXivjR1PfVe0eBQ3lt7
2m3+JCB6yxe/nsqsH7PNElNVVNfovJk2JaitS2MRsX9I4jtvROM4ZnckmdAZwxZrFvA8pv9aUT0F
MQL8FrnaeAaytOlZx4LTnXoTt1ct8uLlrswPey2Kff8y6CQTTh0iFIbrCWczrrSzsUmRa+CPM3uM
4nVJkCjVo2GPNi/wZD5k4qr9KiP/cdW1uAWB2/hGQqT+OyTrVvjNkHS5dXEh/HXipzRNzM/BeGy1
pMQe4wUkZKA/gslPuAcw9MHKqbLgeogeN90cBIKJKtLOIDAtg2W8iRhdMT+e7cafC4GVqvy1/l3w
ccZBEi8MKLrpo06EF7gHXQULorm9qqwIwTILUHivlRp9AXoMjfkp2Wr1I4nUMivr6MIstbCNfE32
z+RmmRMfm0stRyXJif3F55vU1MAtbPUhOc6eVMjQWxC9hyhuj1VsQMA2qkn5JzIGRGYUj3WJoYwc
WNkrXOXxFEGIFEQXodW6h3r6fSwT0rDVCbISdZ4kG3/4ol5vEFgXmOp62K6ZuhOn0TrrGc22Md1L
CpI0OSDAu+RuSRiuF65U7QBto1CWgMivwz4DFx82Ad2UKIVgfOujddJVUAYSeeYRJm+p2oFnl+iW
cr9aC8luVjbQzOaHBvGi5BL2KPff0ItWaXddWMInDD51LPyK6usNguqAQ6wpkwKuAYOHiA05Usyv
yjJfA+7Z90vk7oNV5eI3yRK/QkYHvHVEJGDU0Ef7PuT70ntFBcYOu43dizvOm5UQnk3kj+FvY9AC
khFh6sI6TECV1ixZK7txx1dX/WREDe6b4hXzADS/RhmXCqBthWrFR7VPbsc7YjeTA+xnmOlfbtwB
QEanH3oiOte3clM0fvDZWf8PGO8v1onYBhodZx6fdlBdqLyGuUGXqbV71QSc4s8mkkcJVN/ucLBV
+eiVsc/6lDehFGAgPlPEOihCKOgGCgMftW4mi70NITbCPJ6jPNXnsKiUwviRIzrTv6CZLc29YDC7
Pp0ZIxlCq7ERtFxx8cgysCEQrMB73h54AfSloSYA8fD53wNc43cJN0Ds6LlqIy9dHtpCu9KqqCsW
qtELHknT01RA7F+GPCdJf1BCF+BmZOfPboZh3R2ybeyNsrbQI3rEP9vzd5XTqjUuWWAPSC7rX8+E
j9Gnzhgp5DLLuLKKhB6Q9agRIJOD9v4Vs8KoISj7EJqJvC3dkRJC3dPsSo/Hs2UxucE5BF5zIKwj
4Oinv3zhfuw1RLT1qk1dvThu3VSflEEHPq9Lz8wWO9orOClInOAHUt4swRA+DJYjxw8i/awlJnsY
qDGO9o1VaB+2MLc8MThFwd6L4MQrgXr/MyK/j5CkDAVcKbCEyon7B0VxsR0Yn+5XD+qEO/ojVFB5
vVGmswlEa2gtLP/rlXqjQdDy8HNQg3p5EqFL17hbD/+msKKju1HFtqZfRA088GmR5N0yv+nAPLlH
nPzCvFBNlJi/kftDbxCKWxVTaKpKZhGaQociUfSMdE9QSkDccVhGcltLJuU3g8P5AT/gN78/Capo
MXPGvGlyP2elCLBvTq04QrjUuc1F3mTbGmmWXct5u2Zw1g2lqFv91XEFHQWPaRy8HOM6OqGgU36V
2kSPsWcbfvEw/pO53Hjct2NwDLSFARHCNaskCFG+6jsa6OOAXerCt+y64G22Z/89BFhE7c5panAZ
x2FeW9taYkclxgYBdFJnZGfF112LPBl+d5o7d1RbOA1WBqRmDE02+Bu1+A+Y+laTXF0S57/AHQiZ
KX4SHJjmrQCDJp9llt9iQA/Vrcl+PZTK40+jZkWPLW7FmtwXFZoAoGQp0iZy6BmobH0O5dhRqdna
sTC6ACWgJN/nkBHWGZS7A5170NsnPQXv24xvPWsspjw5+dEofN948CY1cnhFeg/vx8OwT/HC729r
lfq0024h8R+vSpu/r9S/fyok14eEn/wiOaZ8s0NrF8jQLWFF9Hyz5Eol4GZ2GO6uPwVw9wCENqsD
iHE0NEdQuEINMHz8LB8ChQqNPVbf+6TJ301Ah+ynoY9ZovfauXZoTNowIDjVak9jMIyxG030oa5Y
VHDBO0TEQKYOPvrfeFJB0Koplb/vPzUqZq62IiHvNclfULPXBJJwoNPrwM4lBgbXguICuYRD0Uwa
luL566wtA0n8Cjv17lIy2NZfQnhgOfklE/EY//0Y0MT0fyEhlmLTxFcOV14g0Z9LXXiaM8W5WYqd
2W2InGH5nze4y49/9ZxzYcpdI6urS0cxUq4ODBlcPWTWrBJD8Ks+j34C5RzEW4x9k/Zyw+Eg9TUt
RhdOgYt3ElgLDvUZrGDaHI/d4tXFxy3lE0TrneAsHfQm5k+tdInxyW4iKizPVyuobdRj/1dXL6zl
dGogwoXnPlwSYyUAUwnpiw8j009DHtQsrzmFPgzhENo0uVlaC+EwVHVcAZfeUMgtMX6JMRIWk9Ya
rwLQFZ5h1+X3wAAFp4pD1i0E4+Ml+JtXe/zGIj0PzgrMsBOc1q4o4FRJNck2LHjWmqP610O3qQU0
5WhZtyb8BzqfhQqtipY3mrYmFVGUgm/20+p9jugjlDqgmxmC/PYWryWs7XQ5lka5K3+u5/uaeHMu
u6998PX3XP0x1LBzZAGb10Ly53IzS+ecJ8RAupC6zATrKALPHBaL4m0LpmbFLvIlLTGFo/EKIyDo
I/uyfP7dcT/wfjTaoCOS4FqoDqYUDqWacvay3KXVdnNjP2hOH8o0kgBjC7+V2GRKysGu1E6f/QLq
qUKs9sk1yv1bC9ktYElDzyDxPP7ZHXK9e6SlibzP8+wY1AYo3Z90YvbTw5QzA40NXOeccPq9TvqW
ur678bulnqVOSUYYYB7xYv+j1f3L1beTkwsHOXB7qHcE6FHMDVZ+J7qlkmgKPKKM47xaMXInuvpo
jbRu6ShkhKC77qpVXJNErLT4C/B3vMQ7Xqo4ETnFQIFst0mf0mDVjTWNFhRXBxXyDQ8jqswAzCo9
dC+Ftn5XNgjtd3xR5YR4f24OadnOHkIsnAnvKQDATB2MRY40qWkFfcRPxYyoxOPrDC45h3UPBO6z
ZUSGx2z+Moy8y5fsHk9uB6gNDsSo3qubzLKL6Ym09w6faqaDAsUG/g/6aYOoVFmIe7kLV/tSw8gE
5qCEeRVRGn4xqljl4O/7m0fmKhgPdO3uLCUNR/HrflqLFRWY3p5Jbpsn5LCYvOKyXGcm8vuPRmOH
qmOBuefg84KrsXsYiuRTFypR+y7COk2FfVCnZ6KWIErSurCRB5hAPbTTLjXqj4PsUcdzCrDqNg8v
eWUM00o1jlSm/ZWjFbbvVO3Go0YLlPHPnNYeQD6MyQCn5IZC8DfbbPK4Jj+4rcdjjqNuffj1sSus
Co34pqrw94MwsVXPQuKbC8OWnScjn5j/ePww3hRY5pthuU3eZ+OXcEsRTeleDlwYZRkuWEtgEPmt
CYlSYvDoADE0KyeDYviEY6yvmJEmGPxc2+Zg/aTzsX78Wi/ZVGWQ/SjxxjDu3CW2A2BGYc4cd6Fm
Wr7gNo/yleHxAprQwbBY36wM1MeL1XUvyT1GexztlZ+iedGyPp2nWQAAVli9oUGCG3Sn7Bhh3wm+
jqY3CmwgcwcTex3g5Z+rkf5XyoQRskL3D/Jn6gUi5ClWV3LSP5Nkm+3655l1drQBA8FnBI9r/euY
IbHbDgCJvnAJSWpcXSu6sf5XgJcDXO2MM5NFa3s/vZ+w+ltR5ySjTx0Qif9YTH7DJgMgwsSx3WM8
NQKy8Xq4gp762PRzAAwcjhWAslBW66gEvhnOGL3X3Y08uLnSs/CZFtOkhXv9QGdictDQCJ3gFKf/
MzvL6h2smaQ+B/qtYhr959KpQ5OvWREfpQ6TOYn1PLE419jKM+IFofMlJS3Kh+EmXTkOdJCokOix
6oCrpVKHoJOVt/8RlLFokUH6CEufJF6iI9oj7Ek41fplDih+YujDVTBoj2Ae4orHWZv8tevIJ0Ho
d7TrISUgjl43NAvmPVXwo2Y7jRlxmOkEqMbkd15h5WPH48tFkg2iWmj8nG7UVEEAygMweWhLBvUA
a2HpzlLzQ8Ikvqk5Yr1tGUT8w9dFMakDlYe7U9KqExTXxd/uGF427cwaaNboPWi22f/f4HTak8Gv
tXi6EP5PaaDpjbYKJ4DjQ5WH1cWGrVGTnmP93B4Ea1n9lJtc2Vv+iwVgmHlLhHuXju0XCFGxB3zZ
TzPd3d989c5PUnfhDHU/4XYxF9voSdtiQmpvMpURYeDu+o0XnAbSxew5uvE+8GseP6XjOlYu2UBV
pyjq9p80ABO/lOcANFP8yjB4bMFdylN2rV/hAnnVX5pYEVMm5p8uvh20I+B2ihoXRvXIaKWjqgNL
xrk0ZIGUe944b2rrEK9DloEd87gQ1L7K/d+JM+tdP122Fs8xx2M0yv0i1O6OJA0n/deExsblPtmt
Qbj4b2YprfK2c2snp7rmmi/gWTdpW8O/tngmMMI6Qeed3+GA7H3Y9ATDJZByNsoHDMdSLTYA/uT/
b7uF7/eFXwaGbUHb5wdXXh4iEt5h+IvPa6gkxIKffTkqIkiypQxYgHDzpS9CyFaeOrZqBDt925R8
eeHtziUGvFEGnUEO5zBzwIN8O3Awga/5NhogVMMlP7vnhus/NLsqB/lX516JANpNkEyCoc72VuPl
x27KIdiaDR6voBMPQtocXX3Aw578sJS7At/bz41KrOiRkgGPbt+j1du1Lrwx/II5wEf/plSOXRxn
4jCBIDe/1cp+kzmXKQhARgXdkm+98/e9gNxr46Jg1+O00oCd818cpj9caaKbw9JqnCpdZ25kGKFD
XufATW+AjBzoEoQJ5YN+nwcui5FIsX0ru1iND+Ke/RyZVmucNO+3smc/HKvss2xndHDSAXk/sfhZ
D5KJgNENYJd7HYCLNHJwoi4vZYkEuCkK0aMaG8JpN1bBUzNsNyx7MAqCRJzcXVowL5q7GbvCa5dX
3dtSv39Aadw4f6Pl+y6nrFTpDI+rqTjw1g0MJMI4uvN3mmEas0ixAQCyVCBGTnWJ1+k6mrpcCZ8+
Xnpbnv2vohUMdHFb/lr3803Q542at3KW4RYk06zp948skYYyTtuTQLf7kPl9XGLQnUMre4CQTmzs
WuX+VRKDLbGuJuSLTpixGkmvwxXnMKWDIelhYLb6D0eAWM2Ss1eKCtsIQYP8LniWHOvELQMx3zWj
QL4lNA5rbgwUMIOhkQGavx/qnGv2y3VnkSauRaR8P/FYibZ3HUhx7TlvjImsCbSKTS5MG0X6rM6g
b+Oui/9j1AmFPSWFaCtAWLAPeEGO2OCpwb6rWPFGXETqwCaqqr9gp8Z668zeIHGYb+75TPK/cFO1
VKrluT5QJvYBWR9gMsnzC6aZWKIEKtyAoaJcSV02ZIVi3xeI2UbCE3B2BHQVpclNfnyRtYrRBd2j
rtD3lvk3E+1LDJ8D3ZZ7sB0fVRjhh2ZVwSfHQfUHEzs+Hf6xHS61IOqbmtkGxM26Lt8E2sUqc8k/
cMPTp0WQcZ32MR4RPpI5CHim/xnAZI0jrhE8Y8N9C73/rQpAWKt+5QUVF6JBQWfEdNSmtl6iG70t
NSmqluNjoR4akpcUaWUW02z3LE8/W6DnFmP6T3pJ5D6wwcC5zfnrLP3A73eJSF3FHTyXWMvbtAch
wA7IN+XCBlztNEvRaT0sfFs3Gf5yYfOeaKvb3cNq0Du2IZ87pOnRP+r7Vo9YJ7qfvST8NqllFrmZ
7Li42ZZpOgNgcExvBkxOUVzHPGAojzv6rogVntAopz311VMDl9MJhBBx1Fe6TmUf0yr92ssGImfK
efuFG35KfLIUlnTYHQPDjl2wLx1JPQXGYa6/UR+kITn2fAsuegekTLe4DAa6GyIKLvt6ljK8y9+H
4aGL8YGMqe3U5XojuKP3/i6sLLCQLPoYSl/oI+hSPh0e1HCFLrR10W8QGC/jYqZxMIA1x+OttMoT
I424Z4I6lE+XuPK9fujuADH10YVp8uJDyQoCQk9XVg5Lavp69fbG+Q6KshbVTkaF1lZPeEpD0/4S
CrQ+VLvoekfXkWG9prjKPXhlNfSKHoMnd10FloBiPHm8mTWpCkLo8MzgAh0RFJAZZh5aSxOSsRUF
AkUNtNJzbDqmNCLKIoLO83YnXqZVTsxThHwmlqscBWxapN3CEfrEwd0MmbElRUWHNkrHLGj7d5ZD
clfKgO0amZHbEdF0IsyLjMnpPaEkMPTJhe8E3BwAY/c38JjCvViK71WP8zx0OAhaboYAZNB2qEus
DHsRlWbyf19ES3SwaPCwE7IpZ7QAir008fQpqlnWbWHEaJgmY6bnrYC/nQ2l/K5h9q0U7dQxf20k
ZY9EQzIemb9y+3aJ5KoXwA8u1dxhOYGTYnWyLZuXoAXRBDcmiAkgwYcSkJxSlOtu3arLZXV5QZP5
ZpNc2yq5cDNMVa3LWP1i9ipBkdrHXfVMgiJzJGvJ/fQ173EM64G3G3b+LFaMWhYC6cMu3trnzOdQ
POTbJnDjun0FQVIVoy3kn3kOhYVySX7f8eIlbvDs9WYnZ0lYA9PW/qX4NyIsNfGSvCk9txRyoVP/
iU+smAe+rRjqv/I5qS1/Md1iJv9QUeHTZWkxjpmrEpN1uw1Y17cVM91dvtiprlKMPKc10SBp+Itw
W4cBKIn+Vj75q3Vs/eyBE3A8Nok/zlMNn9DTSc/4i+/vj50ILGtNk1TMpiu+BbiT5shBCgSjgxIv
aAQY7g7YzBzjBP4w9Lbuh7Z28NQsFolekfW3UUQh2zWIHuqOSCW9eX1Hfy2RjfXXXkXUe8aymWE+
BCL+iKiui3FG25BKhR9YhCWy/7YzunMWfxepInD5IjiP3U97qfHKxvwoK7li68PrZUHd+QBzWyBp
u45vlfpAToNLqNsARug950RClx71yVdbsUxzeimKeNMiUt5vszluqfcvAF+7GEllRKbgCsGUFIza
j+uLJd0U+K5EPlkY/1pFX+5dGlu+NiU9Z84+d3tKOR2dUqEXg9mlClfRc0oSEl3mCm/1Adta9goM
k8W+rwrCdJ1+B1wvnMiu06OOhvZ81GWPbjqvphEVOtrwSOmBLm0ZdPPi1tyxQOJ7r0u6ar6AivgF
bbqaLL/rRlNXyAqPEw5/PCoD4BGNuqMPbUydg/uQs8IFCY5xuOvbsTbWf/ZiaE6lAB2JdwdGF1Wh
+cWpZEtYtZ4X2pxlN7N51+MswewafhSBJ9ZRGMouMlM1hYBv2UNvsq0+XtUDUAe98kzufSciAObi
EPJKWlWiKFro3Rr6DAkaoiJGAEiK4bzSfGrVjPr13wkOpUBPR+RLUVSUIohNKrkvp0xAQeR58ypa
utsphrq46DvNT7n2k6FTctabzqh2uCDjBB+D1IESed3uXBwDJ+PnxVm2Ja5B2mto0xstGvfDcPrG
tX3QfG+zkpwX2KrYVaEna5Eh2LYLj6sUSmqYvPkmib6+ZmE4wKK0Zgwsxlh5yFqqymYTQFC7zTOT
E9AzUlMPFT4wCGuW9w5Xx154iyne2WyML/C0z9I1/cg3v36NC6anZcztcLATc2zZI8PNVcbRfNVn
VDRYSpGIjH58RW9Wsl/qSAIygjY/k4ly7/Q+dIV1Ndpu/RAmqOguvcOrhVMsg75SMjw55HtwjMew
5tUB6/Am+AVDPMxD7ZdCFW0nWk4p0QNc4w5bjtFMROsglzwWAVWT5w7r/02diW6RGkNEywGjBi0z
ydx1KQb9pWRiETFsE/zF6cW63DVMEMVazw02XFQIrg/TlGhnmXU0QyRkdjY0Jk8BeGvYtrjSTzZo
GRoggCM7Owbe0sMXmdy6TB1wvKEQS510d260fHEDq7IEBfMxazHY3F58fvrP834wG6z7+skqwzRB
DCAa9l1KOstXXRCZckOpQhue17GR5tg0bUjsKshXlzbDik/Ivwl655OZVqHeRhfaSTF3Zi7vmSSO
vlEjgqKVq2rkpNxJkR8h7SoHwScdgc3L6XTnQSzJ6xTh8n1+c3Q7VoEaBjcwKQMnjhrt/PEFwSPR
LiyDd6rCuSdOPFXn8s+h7AZrUYvM3IRV8ambnxb9Vpdd5lX6nBrnNirXa+ON9pnUjX2IKhzLNQf7
KsaHZv6vY9KPlq7jHU3ZLnva59Jx5H/ShLkxFAqyMALyBATpAT7bbMzKBj9J3h/Ov3G0QibzwYaJ
3YsEFsNm+n8MEz66MGn/AatLSES2OKX2cfBXyYZLOxzO9/e0orwFn5Y4/TeBkKGhkXXZlOYnyxVL
dbfCxWh2Il88TRZOd67iyBxoGAYQMAvGHjJ1ukpUIwisZB4s6IIcG4DbO5PT86yu9taTccfFfdQW
wJhJP4ZPdKG+gWjg3Pfc1db5nS+xO2Wi6yJYsBDYQzFrDpxNTnB2kzYywsJnuNzf4ApuF6bu6dv/
jb3msGC48k6tYDIaFsXs6hd5MY7Th7CRE/mqgmh3FbLwNCnYb5tmNkqwhCFRgdqJLdMzsPkb6EGQ
lBa3AZT3MroCAD22CeoXJKizmUgdJxEfcF/0Co+4/fSJi65ste/BHy8k7rfL8F3NQkzjWHhkuKuH
R7pgoBwjaerqAVcJugM+NcxD18PoAr0HDxHZFysQ8BhnVEEDUNCU8tWoUYiVoyVPjmIUJ3or1xjV
J1Jpds0Yd0V1jnbSdVow/bOUg5UA3loy4g73LpqNNWzuabQ7PsxbfLjPBiIK5e7Uo+/u+NJQ8rn2
w+ih350ug852cjqnqIf5twNNpiIhiSM3Nqse4pkVLVk27DMZGrfUGb71HkTVyw42y5Is+nfcBIjF
yyx8F7uFuNJ25aO41zoMqspWDEj3nA1keS4YpBovXPAbFwdePYaIpqTxJgFqVijUvb+8wQaDZze4
/ZZeMHLjJUxUAPllpr+86HITvSmJ5+IVafbwY91NaCMhQxGhYwXBYRsNdV12a2RRaJoq0ddDZ6GR
2HQPOJPISwnlIHfaSBkU363NvoOudg69au6q7hcxTmPGTkYTbB3anzu68O53/N87oJn8f07BXMJ4
9/WPo2fWRiF5xdM+GkzFqvSryUPxR2AyM3iRC0XfJp6RRC/cDtkukeVj6dMpaMHv3fnEb52sH5UV
r0CFKTqH+3yYPdHZpyVbR7hxVkrmITa0A5OrmCaGj1Gw8BFkF3bSK8rbAidKSlFatwl1hY20L1YW
QsHhh/15+SN3FYGs8mCTbkjkVeuTIoda/rp+CLru0rmz3aLW+a9VT9qzU1790yPLzazhBB5Ac54r
BLB731rWcsj66BWXuZzzomzIWipW1LXmAmmp4auBAZUZTx9WeVSl3kqUgoAo/Wo4DECGugsZZ+kw
+IVC7hmaqvd6xu7Uq/xHRQ9AoTvsJfMwsz/TjFQRytkV74zYzeCTZ6b43hKQnJ6qNtT+295jqXwb
fj5DlyImmPNOwT7ExcWp0l3yASf7fwB6hwnrcRL3vFpp6suCxuFtr2dnSbs076mwAmZgyzJd1h3i
/XvqKb76MT4ebcu4FgpLt7Jy18j08hMCdm1D8w4JxJc0IS3lI9CAfIMVa8A4qxYw1xceQXAGF4Tl
1DO8g+XCdx2IUQ/qFDB13eCXbZ1hI5RUYvNZNWjvWJKCzBBPvBPN+e4idauEPgJITQcjYBes0aP3
u4RNpCnxS6VPrSSI0GaWTybvxTQfDyOJDB86r8Fep3c0rzIUExy/ToIGSUGMdcn4dRnn/Jp0rrSS
p7f8gA8g+piaS+mmhyiZYtRU2fK2jAUS1j/KLVcv/6MFcnXwHtWHVkbAJLvIocs9l6rjw5rWzW8X
pXZAS4DmOY1QqhdLleuimNMQIPBLnfGUCjO/TiBdw+iKwpT6+iBtQYyZ5dNuvsLwB+oM1tF59lJl
/SPSB2PumPoJlqwW+7lPU/2gG6CxCEynGyx9ozXPN/ULx/d0lQ8il1eASe9mTb3X2MV3jpZkeoy+
yYzB7LuS0AIzGAK4Ell12uNkfbFxz/ydWtiIdJTAfub2A07s+VuTFPo3sYXphjZEODxBINJxzya1
6x/8c0aInVhzAOq95rxXmeb7u92x2Z8JRlX/7Mdfx1PXcx5qqeb6CCat8qB8RvXMY+xp02r+/4oa
d00vvF+5OXI2zJLmSpBJr+tTHuBgZ0k+cyUbVX0BlXKB5bCyQo1zavFa9NOS9nAv36OHh5oE64uW
mvCI5t+IyWrs5U3KVM61Sa9cbxaNy9yXCFJrkxwAJdANHXnGDSYCiEkWnJxCzgDRNtsIIYFf2OtP
tLfpkfPaQlBC4HCrCGkIx6HYm9taPuHaQDRYC1oUm0kG4mMfz+4qH1Fbw1H7ki9eKHeWPH/tuEc8
+PA+y2ohmNuL95AGJ4FbPpdzRDDYdUH+P9vSwNDqY03oR2vSaHBq8pYUT75vrCeLvxJlWTFtpqIe
ScLZoeWNUn3T1VM60yvG+3BohKf/llhSEiQaDpwITyVWj+kOd9fguB2mq8yBfT3VyrX4L8Ce9Inv
1Gfcd4XKCsUnEF9LVW0f7sTUjz18/3ulPYDchUXlMS2/7lYO1dr5H50vVzg+KZ5I2ARch6HsrLy6
ZGPbgpQROAJVsG5v3d2oYKLDW1hbnGeZOZJF2RmfdK0guM9+4Pmd6HsdVl9lLk9lLZxvTO/ktIan
fhOeyzaxMiNcQM8XlSzK70M4OBvSIWm/PeqGkRIHX9kmVjHto2B3zWe7aGO2jXIVP4S1NS42W/cl
8CihOEWIKcBqm+jeJdN1uu2OVv/iNop5mMu5WDh7xbruRpK8MtHpwTUKkn/JMIcOXhwLQ+RboNT/
25/l1dMoaKdHia4pIg2z4V7dvRxyLQu0iZ0fva/NPDKTTz2AOadw/l4Nd5zQNI+fwICyhiFDSJHO
iG+nITf7hhNbed4duzaAvvxxCSiWEo794Vd/t1X1r8wat1W8K5r1JZYaGye5JictcnDy4Dw7UMkw
r9jU+wS1hh6K7g7CrCbSS7QFCdScfHFB/CHg6poDfg/UqAojzBZMMzf0iJWzaE66R/X2UnvxyO8c
bM5jpJWrK+ZRHlIHJUj/nJWaiLiYyaL3VnH8+XdngxpzvtvXqcJiORm/Y56QhJU0DBlShEO987KY
lWCIUjiOgfJXkqaL/9p69KTBYXmFtdKMVxWEsa3wWYsECOV8SeXU4gioMY77p5Rd8stZio1eiLzx
zXmgbIge6Uj3U2EPLkjImaGuLdVfFuT42/AVhdoiKnxdpm8hvQculGTw//qfqaSMbU3T2dGcyy5f
k4dhBm7ChDxZ27dlx4F35BdfXznTwGVlPP6OkzixN0juwEvJqJZJPcTLZx9jotTp25xUmTWrUm7V
jhOrMrOa0BcDyLhBluy4i1qdF6oDxlEx7MitHI38x9s9Rjmu86TDphHkJCGnGgKFhTERXLWUEhMc
xOC8SVQRZw1BYixqwzHkTun9bnkFUUC+MjtKIPg8Fin4RrRMaXIGDP0HpF/BHWliA3S5F39bHAlM
DVH8dOmF45200X69PxvaRbNVfzxJhDvot11ivIEur2wGq92vHKlyOrDecYW4lIlf9DK8+Z1dL9ea
jFz2T7+ZQ9iptupB4IgSeigCLMnPQ+Jp6v679SIEukHYrvqDnzCLWxxzWW/PrcExjAaMHNrTgbfV
W1pxrk1opIEYaGbEUhJUhhaiETbqcMDLkjVITq+kXpy1kByC1VbvkwLO6hek3H5/IQ1yRiSfJEnW
pBWL+gm0iVJYKN4itIfahVVUaV+ZcrzkWpRm/uy83t8M5NpeuoD4ezSYklYTw6TfGikzxicNElc6
iWo9I2SnRiwDD4+7I4W4r0D9mm0F/1d+NANIKPM+9jSO3MqNLj8SCNGIBi2WEy3obnmqIKlNVc2o
b7WV1mHqbPeFSHqovM26z7ktlW+r1fkgS1cBq8HaeZ8GSbfF7QNhrBHZGsbJ+ai9oFwMm+xQWsDS
dkrdcP0WiUiAwx8Oul/AgPjR4eqYHy6wM5i80Zsf/mkn0yvqdGLUB6sR+lM/FcdJf1jUxtySu5up
yxWJKdDLDB4pyiViN5uj85P37h4GZM5tbxjGze12DVApQod0rEZvirzJs9pDogeyoKSv2iVoL2vG
DJle1OL/vtia/2IncMECinLudwfw65JMIk+fyg1GCSz+ONm/TxTf7PhJw+ZaFGceMuT2KZec8086
I/pxzBdG1vTOWl9zGELeR7WmPvzMheyQCDGQc9nrnhoFR+o4JfkJAs4pddRsEREl+m9HVnIFoljE
kCqgBd872oubWvVYhZpzpv/4zuRH+sO913M08THDduakk477YNbfIYYSyKSqdXdLt1pFXtK9WOgX
12pT0fhBMSxzasopzTHTcT+m5puutFARcC9n6WU17x997aUrL1gJuYD5bTd2MvvLw9f9LQtCG7ro
bfmIphO3gbQnA1EdSazcWsrL3f13I4tBgYOaAOtWHXRvktXxbU0V8c8J0BhuWEgGng6JIOaqcPB/
z5eZNdVeLbu49Cv/W1d6lDm2qOqsvGg2/FzWmPWw1upBSsUrErQgUbmBLOLVifsnSaN3rGKEQWbQ
PEJrc7oKax4Pi0cHZFZVjyXw6rstpIIa7XDBKa0RmqQuxRPuqZz0/tmbVB2dWLmDQbBHYmKok/a5
9X4/dSKTmEF/5XvLRXanYUA7gK+Oc6FB99JqlPBx9/Eg302z0lded5CkbNLJmFG8CS7C4oBb+GNT
b+7DS+rPgspAw0e1TyJBFPqx9yduXwN+6PBujBBKFkZCX0gL6dR2zTQBT40KQh1EIWA8VMce4l8L
yfdT0VwboQwGnXjGHPON8tLquC74kWANC0TDT5u0necHZkkYIXobD5bd3o/iJHDpX1hc8OC2zd/C
GlcK36I2xw7hGDkp8f2E3sLziAkdL8xAWRPFH6U4W7DuR2yx1vxQ7JPyXxCw2uh6VuTT0f6c8HkH
9bZujmpHkJ2vOrMdvEhGh1rQ6zXiCtRoa+d39RdopfmCUwAMoD5bvOTorj5iCZPexHciWltTiiHx
D3EgtD8D0uTNB1F3qSkrSLRRDhaxpH77rYAG0t3MDaMc4RArKyQeFKiNwA0IJe96PSCBJ7Qfj3B2
bfb0vVj3hRCHMp39tBKKGZkIdYoCBWLsWVo/LKUXes755EGxU5HdRLbQ2OMCXtS3XyE2K+NbssKo
6uAwbalogT1vaREksThrQzX+i/jhY2oah/OQRbyUD4EOrxlaHwyRm59Y5m2dbOG1EuAF5ZH8t3lv
OGGyRkcNBoqvnr5YOCxBEjatCsYlNucYGmO4/6v5Ap/3FLucRpoUY/by1nqdAmOtIDLzXnCWckho
6+pQY8ZeZgUV2gDRoSrQW8A8LMcIVia+0y9sa+N7Q8RuuZslAGMhJQVtFbaSRIZyTKJcLba3WeSP
Ye89OpSFGzICvYI9drMWrVwIFjWqJXdapO1rVuV+vaB7fPh402teRUc17inhKjqG+jvWgJXOoYpQ
ZLXyy9LLwGfZ6J5ZIB2ChlYNR3scYE320HQWQko6QbeLufOwJY5I33n0F/1vfd81J3Is1p/HzPP9
mMtG8rz55zmfNlUkjKBkIJsGAGLP6svEJxvstCHvX4xFvV/ZFdM1ms63GTlvg8NXykBcDyQ+upAK
zurWLz8nAG1SDdNOXttGqpWD8RhebFH95h+wi9Jhqc5KGl80JZ900cc1EHgSL0+cLgnoyKlsqQBo
NPeokWMiOUuECEzXiT9/jX24J+CBUkjYZUvr1P9l6O7qTpxsjavW0jCnQkWUvVsy0/yD2kA/NVC8
ENTEPcH6jggG+g6A129rOp4X5JS/oJ1yabILqhpcn3WkKP1AXKuVJEvNDbTvylA/y6XT0JekU5lZ
QyFTZz2IJr6QVh9kB+PY0UklI9vIMBWRK8k8VcRTiCTW9/uc3/UCrkOCOObWGXO4bWnRvIOU5dj0
E6w00WAWqUxzOQkXMXRNTkuQaYNmU/Cw2891s2bm2GupXuLymwAlxDuvlsAzslBZqwUjFC6PgOJT
Hi0gjB+0HYcRwiSezCRMRf9n1QxZ88zl7EfgMp2WPLkVm4QPTo6XJZ+T7aQoyR+fiexebmDE8Glb
MBvONyLlq80vzMKVi2S2AT5kWwk55AWWugCxZj5kFdJc/bE/722HcDLigH2HgHiRAPZTEeHCILX6
EprRI7zcZEqhc43GGLRXtzIq9PJki8dFr4Pf3gSXi3LrZ/5NHsRSQ5J+uN4Fh8rpVYQKJUHjRbT5
8gHUixKuwN2IdYqDsxnbVxdhX0DdyJNcVEaNLUxDCVNm10W+IPjeF6/ZLg6iiSURqugZGXZQehQD
C/pf0TW0C7RudaaWennfbGYGTHRRsJ5Hv4wi6DJ+gaRLs2niivfrCD9H1gAIQpwJ77SsQaWZyXVL
Dv10MIPahxw8kYnVqLBgMb5FJp+c/f8mHqpJNnkTouZdCwZtP/y+utusV9wCaBpNKQdsChA9D+Uk
y/jn48K2cVVLwbM1x4bjMu2ZDcWSxdtnUHy0OrbcPZm4xMnZlCboc++7hJb9eQvxahvvgqckd6al
oIZxgYJqn8D4K5omixg+wf3Z8vZRNqhnBdakqjnrHPmyqpiZslVMK+Wm+tI8xJ/rWQEOO8XPYTO8
zo8mE6P9IZMCJHlWHuFQ8nicVs9n9dR9bNBSmT+nt5GwC57WVKqZjALqG31ZLs3DNvMyij1EGi4r
RTzTbEgjEtspEOMXatdWHzTx29MgDxB++J+tnJPOz5/tqjPftsKpto9fnTZLzw5YOFf0FxCS6KaA
+Nnn90Gie+gAMhT/pcR2kQGgi16I6PuGrNTvisUqUgNdOk9CvTl3/O67ZursDEPCI6EdN5+ZJUO1
U9rBKj9Y45PsjSjU7pex2kspuVdAbYjkkUy0jLx6uUrz3RM82QQt1rvclyUi10FwIvxwqfkcmgp1
opIJOjBOQOxU937thL1VKZaxIl2e05t/wKDo0x7Ac8FpYA0ETTnCzTMycRqaMjBuqKt69+S3wxJd
5SM86cWc0BhjxLr/LWoyz/jWUOQIUcAiS2HZyCwHjkiMeDWJ777/N0heR/OMAXShRQPNr+hcHhxJ
RbkuAJzgyMIYLj0vEPFhXJAwuW+KWDOEMLUN0XrzxkmRLHglxmGXwls1l1Vd8KNJNV+142BmB9u/
tyIJUH0CNJVgJi2CCE2YzomU+qU300eFgynSRFpCDqveSKaNnurA6tDb8TymZRssovZ2GFuHcM24
EPy7jyb1G4HTZsN0ottSabyMUbOSEgukFjgFxsXlEhs6MvcwxUZ1n+PxAuyfNguHtK+oHDrnGpBX
38kLt2Rkf7e2+I75nWhdm7imfKKTxcjoFPzSGFZpjgllTlVMVUC+ZFkaAIiroy1OGRcARic/nmxn
Vf8U6cQCQx3Sj9JUH5WN7qu2qXp+7LAySWF2a2kKiCuNaKiqIT5v1t5choyrYSEObtPCP5Pf0b60
N5WfHqC6LR8Tb1kMTyiG8jJEfXyqYzCyCCTX6ymXHIJvo4fOPRZzT2Gd94yi22LeBEBeNP+Fzkum
bgWY8HBR5N6A9xfe6xY/mohyEv/Fzl5+0UDtesU8cTHNGfUTN5f4kZayOEDwtfZ3QHYH9ci9aWWP
f1O+bEFcXWWcPhp6CZDIIMCwMdHT4AToi4FQMWRfuXt0xn+qk3gA6xH0S/kQD6O2aVSAvvd6MLjp
vWwlgMh1MAmsVvy8rj00CvLXSV4WjshjWeq0BhfwnwCmaGFsCmnWuxamokAwM1wzzhISNqyjYxJv
mcMVDMk+F6NXy4yL/GzNSm729xhgqhPD7WgJMDew+8exM2JWakyE2CSXzHjyMGd/pSdftp/DFOQB
Pob2bFFo5MuHHQIzMlMeuYkxWuFu6c1tgsnklitetXv+SJlgWywhqypR2wOA7QlHfJNCel2DbR7q
6HpMxEarMzGFAulOEsL9819aR8UUbiwJZzHPjOA2pFuJE3o9t10U8XDp41BeOuwSJee53F5AC0R4
ypuf6fXjUwzVEAHVEFxXR+30IBHM8YalcowZm6NqWhFiPfnyHsnTpLyvS0jAyRLgcokARyKnuiCt
8KdQQiV6azcuzoMbUM9GAFfySa8YVlIGl9UHWH0+sw22E3caa1xQWfsIBvXB6ZfiAL+YC1kTPy4J
tO0PXVTJCYeXBv40l67cAWiQsgGg0CM10NhL5QUOCESJY5h7uHDYmimzuEaU92Ppjmz42XgaS6sm
84kr/abSBQCNJ//pa6+UqVNuTwSQSBzs3DtxraQ8yDoSJQO2P+Lhf0wQLdXnMK/iWwecHb43ZPhr
ZNkkZmVnZu372xMnmD4OSXVV+A+Rxnh3PEyKHpSxKncFZYT+K3Wfo6CLfI6hSV/aO06t6a105pIw
r6cS1nsK/ubidoENPN65EOwl+YEpP8szw44q5HnN0e0AmvFXpp3WqN8dKWvzo2s5qtKFBzckQCoZ
1Ae7/t6oQAkcwo4S6lLSF11Bb/fFemYnxS2I0IkkzTcnbPrOc/VK3wJs6y4/xO4xQ2UIiPW3frJz
iFTRP2cyg91yRZ+yoplrE5lmYMwbEj5v083l0Ae79H+tEcMRWqRcePUk/oK8WQGncYNvbk3SJFyu
9ccOYRY2pb1efQHjCavg0nWzWC4J7JoNa71K8Hf7gCgJKW1vv63zjYgGHiWPUjKbC1AcUdvLyC2u
QqSjaSfFMDqxOdj/E4+NAMbNB2J8cIULwdCRioWkhNP6Uam5TXf+V/sbCI0eXugypoo+3ZxKrdGj
MxKE3an8eGKpJP1KzF2GqmmorZYsMBDt1GZHineI0ximAq1RWl4GsLcCz0/1nac8/fS0YHk2Juqg
zMKeUbx1OA7wnc1U1ma5kG2E22LToiqT+FCrXgi1P1+7otURBihe6crB2+E0BTc5dxWFHI7UqIjX
atCyWy6K8fxs12c7mSyoF1ExVwID7rYu4ONE9mfvIl6kQV836dUOR3CzDH+Yf5Lx/l+wx6aS708P
4lokaHus2ybAP34HYOyr6dDzeiBHwYhd8ZWpTOJAo0xrEhXrs7aAHiTRxPwp59l2Zp6PzUNcflDj
XIbUpglpt9j8FCyxbtHXc4BWLlveHR6zACROdr/DjJDA+r86eRHSDMxVXoF7h7aU+sHuDLd4sE5H
b7UCxXRKOafJL3PfYNDjebcJ2cMC+0iIeWFMFUL8b0o9GhdL5kW5B8OQBtdJeUSr/gv+FvYpIrOK
2ytK1RqDd9mbDsR0RDdQm0xSDkmN9Uk/V3AIXrmWkpWZqcUFklit6c9yd8zJ6EUJz8ucOlUWaX2L
l94osxCuqB+VFFNWOoSXKNcyaCTwmvf1e1sVo+s4qpkuwmPyRbzQtH2oMxAnHPeZKR4Ak+HWD7Ro
iqXM+nCPwGh+aR7RdrMGzfMS1SxlFfEah2R1XVpWar7Gb5AQYSjMyPYfVg3iRZWDc83uORSuiV6k
ZJNZxKdzk0yDc1WCHvrIZhjDxj/UcxzFMwr5nkaCn55y4yRPoabse4yyzg+5dhWU0HQRBzYjfqeh
wLObP/LWzucDaC4vVzQGeWtM3cr8nfAX8xYaCK9JLo1ytMaJ2EcQuj2mzJCxPuMPK0sNUYWk+9Yi
34Auog9IcIJ1x6K7hHpc6ve/jyerwZRwzvLQC3s3dOCjU3ypYFY+UsPmTJVpLUXwmQR3gC1o8B4G
ivRUnUJcNROoHhpv2HmYRRfrt1T/9ayWnsTRNxO6N/Dfu5PpF2FG1JwEmyzCi1w6RbJkGfLdHV0I
/jmbT/vgx3Mt+HzzjKoY29BMOmbfVgUvLntxDxoO26luSsjKn++dDDQ7sJZnBqHCPgtaSIiidged
j3YqszlHlvdt4tdQYsmANIuy0oNlzvgRrEASUqOSdgoBpsJ+QkHmcJ+7N0c6raHhjdaD0/RL+/5L
5SzhXTENJKXJcR+vMk43jUzrGx+Xoa3OaCpczvD0NZF+kcM2ZQcAjGhipVR5GM+DJgM5XNjGp/8k
lY5KYmiOCIHvMgzFrdJMPkkaRGsHF/MKr/Iyhno2Y7EDGjqkxHiyBqKhQiYNvkrmqzm4mNYUPa7T
b5WbKBHgUrLVH2aOEwnC6B4kYf4SfIxkEVJ1b64dQsLXrSOj3pErV4KdF28C3MyC0doz+8wVrXkj
PDXGTyTBy5VVXfiewIDpBe4zmSJ6ZtE05QhdhzpFC3RWVRH21oCCT0ZfGkJHIIuvzPdqFUfewU/M
vxoFlmN+owcWR0PmFlaZen1i9ARpds9kJxWRAU8giZhGpvGqwfVlid/UGfQy3TW1WWONUj6D3Kni
YzOEYw8vQxUTJYNi9fA1SiufQC/UAQS8r5U62NhidjVyGjDPat6G8fedcAZXmkSMRPvkBKToSXMN
TdowA33G1ONwB+0y+c17ScQw9PUa8GfLepua1mOMeMKCClNa2R8UHKUXBQ0H7HuAE9qORw7WdkSK
Zw89gSZV0X2n9LDS+5hfmPJxvkXWHZ6IJD9D5xoO0w38Z9CgzBBkXKaFRUz+/fFYd5r9553ZmBWy
3FAYMW+EgHA1bS+5cWTlGLS9KUoV7APRfa0pGvn1ubvPPzadDFH9YVukc7oeBipE3ZK8ic0nxEc8
fUZqynZ2wTRIHGJeux3LZSbF5vny9oyNTtSBqwbgR3IxGzj1CryJ08kCrXypO7zkGG5CcdCHvoEP
8H8wlyIkuX9Wjds6EDe1KaabfUR7iWZdBFlt737W+GPJ8YhBPGvBD8VTvP1tBOEBMikfy7KxzXuJ
FbyX2ed9ejCrfB8EvhkHozntNDPizgkBgn9bA0nvbXm8CTGm5lzp35itnLiV+g8qNah9ImDKeeaV
+CTyjb2/zmjHvI+HhcAxACwBDS3sry0W/3jkqwqVWHozxqzQwRASvninINhcAdqwj2oaK9J/ktcW
qpywmlwNZw9aLrJHYBbc1C0oKqpz7r3PbKpZsKVZBvjTCSr8zC+LGu7gY9V3mOh+clJvbPtZf7iD
K8OZ9u0xNDUbSmfvt2v5wV7InsDR6yGRPyGl0+NvZwPirRXB7nvOooNSYjF6K1oUiaaCGBUsYLu+
P9aJd+b5iph+O0iL0VFpU1qxc35NKX69Zg3CVyK1RE9/UnkhqK+XPW9yFuzjQ7t+l+zH5UgzmRVg
5btHKWvcPeQNmfGxpq5mpD7C2za8ZCj9evsnW/Wk0Buv6mFLbcQ5K37vOl2t/zD7yJaHB++PCnNt
Dj3pcK0Wj4v+sM/7KR5brdm4DTiOrxEE4rDke5A+Qif7wxso8AZpUiOxwWtmccPLDeBEv2QCgb9n
XFBkOvGEgHfasjRlw3Nj7WMvQIVlnlA2lNclDHUWHheV6MmVBpNT54oQjLLR6GRzCjjP4O0ve4LI
EecpP7PQXPDowsAcvbpaFPyu0Bnmm+1CmlIjFEABjGhpSq6BPSPzjPXPb1L/syINvDu8ihtE+3p5
64A8cxzOCd/dyQTs+jOF/hq+bA4P2xGPn7KVUMH4e1KjqbmzJsqT8mWOadY9MALipdx3F5gNY46G
tAfA1euv9VM9+Khl7q2t9VYynhLDewxBUQw2qQRgFD5dKgcdjGOCmbjw73ldy5ODXrtYfuvx3wSt
jqChZWW6Sd/f+yV/uluxyqFQz37o5pvmPUQk4s6+EngsyJ+rjF5HJIOMuSpvUTlh31FBZl+49J8W
CrTyaIfugQeD276kT9TXSjr70kpJk+a90kIA6/BqiGxCW4Az7iO7/IcBXLfhwHPjCzLPD3IfJolY
AC9o8PejmXiMsc2w28S02h06Nll/x5JvumCEjp8983eNbKidtCFQV/vVMe+nhwAUYSmuZHZDJ5TS
YNZVM2sFVdMJgTJ7fMBuz5SsMSgPasfY2lsG9B+FLHFqv5C6z0dV59Pi0yIpnWJBdP9K5uZKDeOV
rZVCyyF8r/Dh6ZHmvPhK5BAZwNRNZ1Th/SU/0l6b7zdln2KH0I11NH8IAo3kqKm26dmagmR69Rxx
bRdWEMOru23UmiRh0MMqZ74qGepsAGnUM72R0qfdTojEqwJEDw7BWQu/Wm5PuYVxdlH9yUbGdG3X
ccwOez6LsOiezWu6Xa8+lSarrFvcQnFJIp6rSydGaaQCS5NjCWF6LlfQGPxffuB77ftpH+3iYd+v
a637ZkaQu7BZq+XRjLNl+jo8iEZ2DAZTeFltmskfwhYj9dQC5B4LiqfmuAOqgF41k8nbL7j8WyAq
PYXXmBR9ysG+lou/FeUCw0A0N1fcYyYWNSZMOPEMZGggxv5t4x1iPVft/MCoI7eVoQPHblSyf4bW
cRQ646Sjogd3zjI8d/dyGZ6sVZ6xgaWU7A/0ZxllMmD3PNpGN1Is7Gfyy5QZoqApIhd0HU5g5F21
4F2ekT/sVK71j0kAZNZELBWwn+MFGnbr2NML86r884rYK7K7xNdhDJc6yyJ+OjEbvPR7rR2UuB2i
34XkHn/MFtd2AnkdHUNP9dtj83t+NtYin0VkHbzTuba+RET+xvp/nKfKBuzcebvhlXwJE5fPHrdG
vjvYFuLG6Q+scqqcPuehYLDw+WT9cNMlIeqep2G1VrR6icF0gLGMwwA5AG841UK7J0sYknR6mZ0M
TfGB4SOxFs0tVjxL/E+10SS7wVzFe5RC+gOQsoiM5U65+mSXRfJ/H59frq+c8CYb+nw5hQTP69iy
Vm8ITG/JHHnRQKaB0tco6XINR4dx3+1S2bFcr3hcgMGrBSRHIaJmFDq0qQ4f+GwzNttm7zeWE2o/
ktTt/jnwr7ZbOLmiq3KjpKZKvm2WPXZdFhnUQRVTCFWf2qG+gteiTBSUHsak2X556RD569DJGzOf
D4pDucqy1ypBIX9WmFm+0O2EYpdZaVGURd1qDa480NWltPB+2YDvMdtOwlGpTL23k+UdJidn7DOb
zi99vsGYjTP7KIlUKjKnoUgAn9L43ps68+gRbCkut61ZhWrqAa9HbRNG4ZZOv3OuXNHR4D3vtrMh
zzPul6+9kqK+SJ7Usv2Yhw7trPtbnwkwarkjRCNbIpe5iSD6tFC5OweI3IsP3hmpXyYOFSuQ8d6s
OjpcOEoM18tiApReUGanlcOFnl/ZUftDhnt8ptsMublZ0C4PZPiZe4Qjo1Jz2O9NIpM1GsdP+F9H
UFUtcJ+bkbHDaxp3RKfLhN9GCCdSuP9zMAX1qvOPGSuJ3jOWidtS8mQh8sXQJhiSF2KLN1rXbjU5
OUMV3+hLcR4c4AcupJCofaX95PrAu1tjGM/hrZ/rEBd2k+QfQwxmDYGDHjjqoE599dce74nmp8JT
8uC/KwFuvtvgRPLMz/36+D/H5ASfw4HKvWrMl4PElOrtj3IchSo0pjNtn+P6pFTRvYEfghnVPPCc
oOj81BhmBLWhhem8KyzIHVERgUSvkNH8ZcdL/Mw7lbu9wW54V7yooc1bahYZ9YF24VJEaqhR3X0g
sJKYH4hfw69FsAeFndNMYyCqTVp7NvmaUUysgLGoA8X0LPaxEwjvvZBsbaTr64BugkIMfpN2qS/P
ZNaJkd9cc1aHp9gSE1r8L7Em+zv3LTMkHurEDXn9+7IxuHmthICdL18Xhi3h9TLeW5K7VBUlwQ8F
0IQHpjHiYbxqp5/il4ReOE8qFuOR81fssXMtHVtvAL3ZDFe4IR6zUT38bJlgTtE+odqRnsC1rdnF
804SThgAvNUjzlHxG4PjvPOIWNxJWICskUFvocng4Pqx0/Yg+MkHuOC8Xqn9hNTXx0nJ7xEVojui
8nI2Pt3Wc1JwT4VSf55ypHAQbDWgVMt/AG2Rx2KBGchjsYCtGR5cjW65YEsjTALSgBECuZOMW5uQ
ilUl7kMhS3bgSpeSCGzo0sdXEMM+PDYKHbvmITJCrLQU/84mdEceX+MumTVp7JkWi7lAHwqJbVZ9
uGz+6PJ/yPXzU0K3G+NaQ6SCpQjiIwY3CYyG6B3TIZ/xrs86y4E8Wue2uHHnGcYE0AA3T9xVIlOt
stFo2S82ZPrNfcv3eNYWX9iUsKxmBXa92AY3S4qCUEiVyh7iqWpzYT8vqh5LDVuMrWP99ZK/7vgj
Ja7sgYIGtdKedU0prvB7QyrvMTOYb1jbmgXT7nlUp7JUTH+wOhcGLB4G6lKpp5x6RAGK2nGAxSSn
rZ+q2dHbStWi6Df+LccSDG4yPeR/jFD0qAxr9h34ekN9t3iKYiTd5z82LKjB4D8IMBTagImX88Tg
qPnqaWJAJqexJYz2pnVo4M+hveyuurIRDKHtyhKvaAugURSUNd/rYca9EYJ+bDUsyB7c4HyMXVyx
EWPEheX2yzplUM4+egqszN+Ti36cMIjgu1BmSdhtRPFoZ5SskJ3XzRn7iN+OnPzm6kpPRq6nCazO
AWGTE9fh/k7vbxAuDKnIr/nW8epou5Lin5XIRM9ha3u52AgB8ulqxpXVa7KD34On2pCkKYdzKaK8
xiNJE2/F8Bz+/EKbf5Y9rCWU3iyL5L8qg9nCDr1WKh9vu3IMTgcbMh9OaCxy4wRrEA07LtxEqyxs
7hXKMQrOhKu81r7O+yH+g8qICZY8+TxdSsXARKKqgMxlGlo2jqBvuhqhIIeP7DvdbIDBwGJ3K1gM
FjCNzINV2XS9jokAMrcHR/uT0xDVQlRbssB/qXir82iADjoupvVQbcZQL+0AcFPOUKmw/oiUbyp7
wSAgAjtaewr44NsiiIBT0mltk40CINtZpfwYkv61bwhHa/t72Qyq3c1jw8ssECEk4Ew7U6Y6zx0i
MQ/gGfeEtU/zw397iPz5h1jJqtgUmcBpXw9xVYJRbVxdidm4ZIgbbnsJPPgTodf7HftI8Z7rn1fC
tYDhwEJ+b13/MSMbuR9rszSdIx0KNLRtjlSv3JlMaktqbcr9oR4x1vPIvrCjMLjIsjjkiTRr+l67
8I+ZhjHT0imXDSYwb+q688zZ+cVUxGfCX+4Rx91prj46Trh1wjMqM0IoqwjiBltCji6WSVTfU4F+
/Fmh4SC42rQwEWCyEAtPVeWh+PU5KwmoCX/U3b/t5sZ4MFAaUSEBBOw6yqSloaQz6IwsiXLoFoWB
l05VYO6xHlKwhEGi6diKnGvInROYFdm2j/2hefBeNkWMJhAePpJOf48TumL5wxAgncJdSdzebMdT
PtVHEkw+h0K9/fIozFiCmamsa3QtSq2ESpuhRXLFA4BtX05fAI3BmLTVxe5i7ScTvBnyN7Zeb5Ja
x864VDW6oaXgrroOa13gRaeNKnNPNII3ksDJbsoMP+EYeyELX6G9fKyMjpbTBoUyNL3mJ52vbrTk
F7Ull8a2XyTw+k7gHmlimPP3vyGrF9J17bg5/H0nQS9uVTIFrCW2mGTFY+PdMa+OogAmUdpXbSQf
HRScdPciNn0oyWwDf/gtiz0hLTIwkhrxB03v/bfis8dTpRQQRPK2MbbWdysIs2XnQdQdwS2LaT2E
vPAPi6RxmIEBoE6mXBzJU8pBGgdgOae34hu4mOfPi0TSgRSkb8YNuaG079Rp7UwKzpUu3p1Ogz0m
/aa+AIUmtHSadlxQTELsXx/lwl8xzw+e9OgqPPL11MH9XXhtL+XHcxyoQIRPpWqpmCSvk4FOw/lm
wcpOw4c4EX+cduJPMeevwvlX5Vb1k/w6+EHKa9BuXMw2jFIrm4Ahl+WzBJltO7aUGLyGufU4UrIF
fYXkrxZyzZDgYvNgGH74wzjUa64bjtNxgVJjcxHb/I1QsnMgZjpIlAnoUFCNhgX6uOwwZwqFt5R/
ZYOr+KhLnbmMfcPRpywQYEiZCvlg7Zvz/Z5oGg3Ysku60orhLFhKnOutSrMyLq0mr4Pa9J1LJTyl
a8+fkClpMzvEh0e94dxZ1P8lDRjHR4WQMccq3M54QCNkYB4EsFLDkiVOeiOfyXbdvjVTVfyCAn7S
LI2w+ggSu4JY+gZLSHq8WwASFstldWnFcEFS53tNjmhD/tJFuC0vaUhLfL1FznNg6CLXLcPdDdmU
iweVUu0laE51T+OTTMTOCP+RvC2rbRsrgnpWr06fZBChtYNAYY0metOuykcjDLGm6F8ahYZ+k0s2
Zrim5nG01X84eAI8Y8j9JAiPBgswkmMHm8XlG2bw8LfIHkxAkJ9JBqHEziy61zfSxw6MLqNVb5uu
QZyeEEhsGqKqn0l59HamtFUQ7NBNnH5BvVYXyaAucKh+PH6bDz5b73oAwwAqBkjIm76aPDYNsQpo
C8q7eZ6Wlg8oPgSKtJTWjY7/1PWg3rdMtgEGAbUf8DEitoE+IieZLwZXW3+xOzRZ2GUCwscOQaH5
caIlIYznzPtnuD8FvBJbrIB8l0UZe+fpy2IwsVbDAl0w+moW1MwExkhBugeC23Rf+esSm7Lq5gIc
WlHHv+kFVVkapmvKP3TCJzXyUVSUDgro6QS6DxElEFqMsmksbVLqtASRP+lWIBRWLMeFHWu6C6Ny
u8bi9ZpBcBHjxTiCd4ry6ry9jeMtI8tDbdvbYIntV7YBEc29LEc/r9vWaM3e6UrtVOB7OiaP7vhZ
gxhUQopchfdwRI3eh8YEDumkU++7eYDyQA/GyAe6GKVkB9t/9ua+pLN1egoVCqQpYuDOgEjDgi9+
xRlUxK6I9aVpnU+9FHF3EzqNyKQRSPOBvZVTu3E6y9NjHTVqa+/6iTia4k3PxYC8ff3emOJUnLZa
63MH8ZuKeHU/DpaGllQWY0tEt9ygcD721xO1xnefbLzL33FSkKpF9cG4JVDciNPmAhhSK0GDlEYf
uwIFeiCjKjqZIQ/NYZ5HT6UqSuce0AZpinJ+46ngpAoxJ8//HXwmfHB/2mK+o9p335yPouzLqLO9
SN7ORYZL85wCnUL99yQg6Pzf1W3cKMKHF6lXnED8+6rqAQYi5QFg2eUaVlzVLi3bMdtio0juemBb
V65Jcn3fRIWf6rtoKTlg018T0HhWbDWfI4sO6GnBIeeEUnA1J0ygs0A5dPAXZG4qieZU7yG0QS51
2sHXpQU/aQd8Sr41VS6eAwMhGvmuMdrTogP8vEpkFPcQiH+m8Vf5SLu0mxmkLvem98q8PNkl1em0
clf1t+iJO73an7ipb0iYZu/jBOXOb0t49l7djjCg4qpSbBSK7fQ6uBOePdnoeIbtu3QcJuNuFsi0
EWow2fTgwounQxOGfbXSDvSFF44xhTI24VFHHcTIOYRr5Cea0Pg2FPDpOeV6QV3DPZ3lvow2V5+/
w4FpRuw4mXr2tuUrAum9JpNESrIRBvRdYNy86aeG62jTgqZCQj2OMP5ohL4RQM8GgiB1fzRmMxuE
DhEU/1UhhU4k2mi5YF3kw1g4mKl8Yvfkn4aOVSHAVLAFU0PdcNTEWlaCQX20q82B9uyVhHWbmpWM
X6AW7ER+KJVGZAmYh7w2OHhDvvBEuSr6tIX3asE1S6TgeDb3lIAo/wynWDTGExhrFGy8mtS9Cca1
mSfja7dgbA8IzKcsOZMYplbYVJ0agvDocSnpVqZp3AvOV4XS7LMHRnjo49sjAgDB19roVhWbMJbl
SincF0FKBwRaDm5VbduceolB3I/O+0jBJosk+H1o8EEWnkg45HPU5eFQ+xz4OMopP+dBTg0r7PC8
yA7ynrsFKCbXtuH/Q7WtnK1YdxrSy09mC85aq6fKguBmR7CqRgnZP/3ccdR9ipHcLQ40Cnp7TgmY
G7Fyc3kVCBGgBJcWpx5dTdQwNzDXZBrhjvs0Ur/5sUs7WL64Yd+bZKjT0BYb7eTWFrMmcS5DcATv
c3SOCVrXksaRFgO2SUVQh04fOJRPDa79lmysNIZwXpTTvz2JEkurmdkjUKfKYCl+sBIkeFciWA/F
8CrW9GjxWyzqrPIwvzHuBmhu+dHHk/aVfP5UIPgcZ+IjHsfwapxITq0h/RNXHknk9uqTW6EMC/n0
U1ZQpBzveReH8uNWIJcMpXlkC+0JZFfrr9qDQimht2LyfDJguCe3yGYam9/XufMv0GyMTTmd7U5g
YA/0vO2aj4R2jKfoele+28cnubvCNds1OD5pXriAK2+mIvK643npQ3JTjG/b1xSmQzLp4SUEYJfs
a5Lw5/uL0LEfxgwgM5mV2eoZQFAnISJnrvvyx1fN+mPxYiKSBn3qqKRYuIr0emEpZKu1s7hbjwZC
J347xR6lq7ATbC3nWqpUm1Eab1ugrNBMdMjKwDJl115+2Lb8KoQKzfd+XY3gm3KuX5kZmfgIikqU
o/hY/XUNiZcAR6tKBLRtuAD2z7QY+rf3xWYWNoP+x9Sql2ZD37OS8+s1TXgGL9FFv6ijnVHe7msr
erHvFCNculyonkP/XTQXWc65/+/uBL14+PN4TRGX2EjnStSwb95Adlk84HG7K8M4KuGPPcNR6K7H
YOtlvrSqzz1sTl1dJoQHK2bupxIv7E+SIjLNfO6iqVpQH+jbCUCHcDeoVFVB8UpeuilZLXfxUEas
rTWHApAMuKxqVXVlAIj07Xu/j84J5UIppmXhxQ/F9U4WV5SQ2QOtvnKJQbBHX3AsGSGJlAQI6iqp
fH6Sj+cxcy8iCkFcO7gSzx6Zvvl+Tc4ERJgmJWtMKBw7nKa98TjujTdhCFg4jnUF3gkDG6q/M6Bi
xYHJNO3AF2lON4AK5GoREZF6duHrtS4VZveiciClUdYvjMYK5GlJ9ho3ZGvSmB3doRg11cVqZmWG
keERkWCjcJDT9Z9Xf9y8ypyJsEducyd3E2n2PD+rGCk0tt3bqP6Wy1SeAubDWIXXFWgaUFmL0rZU
8ho/rYaWfzmZGrhDavapgUlFmtFE2loMu5JF2FMWkIkt+Hkmh6MiZ5724mGK3STF4J9FU3qlS6aR
EeOiSmsaiELPJVQF4ZdJyE5eID9I45Msl22CcyfKAxygfgnxHT//ro6NgVRPdiNLjR5SckyEgBHK
Op9pM9AGdHTmKVGAl169C8WYeOkNXHbngJEYnCOp0jyGhtsV/xFf1M+YvCvQSzDERHCV0SkRlI9K
JzyqeHv+EKGSR6YVF3TSDtbAwEn3qf7uzkShI4tFtKpb1vIwHyCHeE319SfTT2rylUHNYUcE3qwV
62rT+5UZezTl6bVJyJqxzGtphB7pW/s1uX5/fZGENUW2niMRM15Ry+nuIOhF2dyzv3/O+XdOa5lW
2YUZimTruSTqdpGUErjkTfxiMuhPiO3cGxwmzL/h27cg7YT2+hi8x4XWn5fbw6rETHCWxRCLYHhL
RtZAGWzCOHEvplXbMsgKO8U7Beo8AWYG0iF2xeosT6Yo9RfZrXspdSuKclHv7GufVXi+7Fi1NVuf
F8bqUMku0l2wNr+4MaBlouaU5yityrCiVbZlpgkh9JfEQY39+NCKaVek4jkdVATN+RkeRJvHgcqJ
Swg0lF/nR/UPGLLtrtIYI/mMoLMzZSHjboigyrbgAjwFiKQxAB9JcQHWftHdxeiEscsJORylewkd
7W6Lx+3AduCoJh/2gscVi8G/OIpxPZ+o7nPcuZBN4BJfwOBiNKPiir6JtbfgZXFc/umn7N5bnjgI
EdZgAfVb7la16QqCuHAOu7smNhhu+x6C13zk4gjTwdu9g7eGBmjyufiFJ09CHlCq1ZrJUljsldCy
EwPqH4Hj/Q+mCzTOVTgDP8m2P0ti4okzAVY8cBoqCp1o2aAg1r0fuhWM5X02QbGKlREYt8G7q3tb
W4JCwwIoJFe/daoZQ/AD1q+P+O7S+79Y3CTWKbSBbXFKV0lKjZt+zwxFegFQXz0eYx+49XIzCj+h
6aGEscMP8YRdN68zJso5rTGfunqoZnB6Ns+PO00xs/1teDtxhEP5PP0VP918LbNSB/x/9MEYrlsZ
e7WCioLQGLcV6gmlFRaWzUn2cvJ4LJ9lTQ5+bhDnWCmYjr/s+AtnXdBy13hpN7c9QsdDNIhTn0CH
6mhrev0AaFS3UOg4Yd7iTcCd41ssk4N6tOGhFaoorbLwi+xUbfowomMCAULqeXFKLv2PsmYVKwNx
+wzY0JYy0H+QZ0fOO5wkvY7MPx14bIQYWoWRNFCAAtekgYwTy8NtbbmC5REaWyjYIT+yY1NWMWvb
NJwBAmegeSqL2QXpksyAuUqXfH5xQ9bsevZSs7zQXBjYiTdbLisB/l5pdOrCWKW2XZgVsP7ucIv+
KPeYxriSUrPyfhvqgf/wF7sbHX5S39AY+lX4tuySJb6AnhP1NsobTFsi2Oj7HVICIUCuCnyymtV6
IZ/DnlhhpJ3LZGPoIrl+jL/VmTGCLSJ4XG3cGftj7ttIg7rW2SIp6qCw81uU/i4cfcysJ8m1Js4e
2zoW9uSZL7TIh28CN7NpcviHyUTA0TXP1FfItXKu7TJjlOnTVjODQcJpVX8iajqlv68M12p2HkpT
rEo1ruElwQCDtWpPs0JK54D/apWGk5Eey04qsPtBaXBaojU6++f45DQ+4yGSzVSc+WANEPMRhUl7
6ccLpxLxvH8hRYc187f80bkjG1Hk6tpWhda7YpW/NHIuhLqh1bBQD6jdRyQoVXTeAEAiNGDVnRaq
N4qH2pk3+q0gLravjNuCFW/QyVThLiCiH3/u1TIjxSS2qFMNr9hNFMZhgLH11s9Roi7VGE4vgbYU
vueBTF3VipcpdaVgxeaH/qLHDmnSDx+NpQVBCJbk4il6XAZAIao61JhOUE4tr4/onevpOGJiogFb
GsZTa6VOL4xny3w8GFKDvVPRlRIt0ZSXhu0qotvGqGvWdyz2zg6zu+3byeS1idc39PA8hEQu+j03
V3063MHpiENrRCya3g1yEvhsI9hwhJGYPo2QVCEbuUaDV+XDCgMUYdkdymWwPGDEHyLH+MsrHotL
C8ESDqpFvKQ7Q21mcCuPQ/PM0fvIDO74Uj73kmDD3Up51MN82FSpky1LvBHHp2du1TQRUu9CSdqA
zoHOdlYlMcdwwiMZz7tOwMeBGa8DipJoZ/DBgUKf0Wp5kS4KZH5wLX7uBQ/qCa8ZaxAxdXvUk43h
KDgy6iRMGjGhhmdVIwgXzqldKgoCtSwaUuwgcQXGqfZSzF1GNb2h0EFe8+d7NpP9KoH4WKG81kQX
mmqERo2jkqrs3Wr0iIFeZPAD3+IId6an02KkHZwyVx/9DrFCLIdsReIKAR4d34vZFHJip88lHRnT
1PyiDbcD7QN6wc1+3i0F5Pe0PnEpe3b+YM2INw//OW2zEPUSR958Zmd1SCX3fcDuNcMEf5cvdjLk
+aJgpHlx9jqGi4cJQhAINJbSgPnHluDkLQRMR7QUKfqzYLfg4VC/wfc5zOJAk/QxEXhrk/pfdHE0
ZGp8FjokuIMZUzlw5W+Vp9u6ewMa6V2ixgsEl8expTPHkbNTlQaHrTRM/lKvCqBFqGMQt/Ows11/
yAzfIaMPEEgOBMcFE/D77uHsTD/3nPXIiyIfgDGfEUqbVWY0PUNT2q0Kw9OC8CU9g4xUBGnvjL/B
PzCxNRJpzZ7k2HqN1/iCZg126AOQF3mGDGnFf92MsEzGF/z2bg2B4++QgI4zzlmjUY0xxNJYZC+U
RoyDV36agJ64EyijwtkkBdA4ZPQukdCAfnWkI25zidb0VQK+MV/Bhx35AqGhOKgSVa1So1SbrOzO
9be/PdwXmHUx3sbucYyjSFxyCYGprIn7sy5NCBWzrk7xOugHKQTJfnTsE00JAYAnVi/bjOCjIowx
lLKAlxLmj5ce7b3Nl6uMbQDDeQ9vsD7AYRw/DV6Kngq7Qb21e61cq4z/4KBDjQGjOFyA4/5Gduoo
l5hQhK4soaSuHF0H4clcujsx0SlgfQEp7XEGRpnFcDGmnpx/MYdNwhfBUvlactozlyjd48A6mJcP
0EPgRk1revt6bkYlHtRSOVgzqijGRjIe1DdzXZoednVL1GgviVKgIpP3HJT0RovlbRXM8y5gaS9B
zDDFZFnzRD6iOzEwLD+8TO6hm2cedtVXEy4z2qEsXJkJ1T1EyKrpsh1YdPYoYroN+vOvPYHD1xbM
k40d+HXBIaK1sNsWNaEmSiJJfBPR8m8lgOxZoy7mlBtwa0b6JDoujEcmKSSCAR5ZIoj7cnHlRapt
zMoe3O8amN5uHTr5XwGA6JAi+zrCoOyIx1IqN5vgw1fvM9tMCB4vMtrXj1dm/cC9Aa29/GBpPrcQ
gzA/59T0yTRSFfqPtC9x7Tj+yPuXbk70xsrvRBLPNtKWt378GPluyOSEmYbeym6NJy68P8v2UllU
EXNpKng0KPadWfxP5wbCTKlcBcmG27NgLF7PYE4Tec6fdD2M1cSw5qhIaKfzk6rIeyu8QungoZeZ
yLx06cpKFnrPkMu8Vwt0kJC+F3F6c6m4MtrH7Ix6Ziv87dqySEOfSsmBW+HDMomvI3uf79OVrLqO
3G8i3mkX3ac7ntZ+0zc0DxZ8KDAeLXbCBhQYAlAnlNhYyp/8dvpdLd6bICJjR14hRq67F+rmPQWI
oULXuQkvpN3uVEz7aLMBWFywXJk0f2PoxqsWlVRx7RE8V4gu2Nr0LagF0SNbjCFPXStL83h5x7a3
pYaWplrlAyUsNGU7NVgzv8lqnXLHVnBR6xZmpT9IFxdgZzWnF9oWpjd0m+vD2nbyb4JFGTnDH4U1
n2gi7ACqVsbKDVdGlpO1/wLYIhhtiy3QIremwxna53QL9WHVa/sXG3+sZgaOyZEP5gRPbeALwMP4
YlUAO5t5ScagwuR2YV0gEl4qNPqrXNGAkHLVgjSB6CtcpiCWDr9g6YhcxlYUftxJKUFwxka0YWX+
sbl6jWT/iqPG90YynZvt/qdxg33Q32EFW9J9e9dk/FCsrjC4i8xSN/geq5sSbe4tzV8zjhc/I+Tl
SXGqSieQe5xjg5/W2C8VpNcfdoss4DKru1NoRYkHbYbo2QEgLTXDUvFZRHobR0oiJXpgo0Qyny0o
J9qkXj4cvSoO+8/Eir7z7DBJsZydFBPuy+cmGx6GzKGNHWE5qgIEU5kH8kBVsIMOZDytNba5DXbC
9OX8vMfmIfmaD6osYul7IbMo3Akn8q9nlb8G8SJnVromXWjl+i3dIXwWJpvMYQVhigK+zn6/ZSx4
eebASsJniY0P++1jwzEYGTU+aB2h+CLu60UKoCYsj0Fxy3JwznE64tqXT/bIWfbUygWf7v5WYeAY
rVhuamwU7iH2pw3fPTaFdDTEPkV03OYuWf7MgRwMYHUhGcm7zKeyMWT9pM7Jlrh9wQuzsLED7kMp
IRPZkooufQxKI0vsFXt7d6WVlEeiemPRYYoic3hj2z9Cf5hSUllmu0H90mkuY7Uvt6cE7ZYear2G
Jb1fvWL62Fj+5BslfAOTb1xifAY67zWvEvhkeyt9ZuS1jhs3RSRHExgU9R6zj2dQ5+5fAY499Oq8
r9IDPNbiUTDemgY5eQquZEi+d/9Ky+xGdgdp1o5JWHtyePOputy3nED5l0Hkj7Gl+23rHchco2EN
siHdtjZ5JHnkUZPazQBDhViXq9JdCebgydNPIOzLW1Ez8XD6/ZqnLtDLLM6JRNXsZLaX9H+Yh4Oc
WwpWVf/8+o+4jDS3AYWZ7qP1tZLAga31AlUAxDL1nm2jyOCXwKrnb2UaEs8q7PjHkjb3bJXKVA/J
YOcvB6w0nziojorIfrfywhCCBe004B94m/BvUKjw3w7EzK3TNhWMFhwzmswctqApbAi5fPwFx4Rt
cldrN9H6klsqzs7Jg912cj/z1I3wUW/26G2gnCmT28/P4l6qmH5swQ5Dsrdb4L3CXCnbuWqsWrnA
2QlJ3dYLKffKMmlKur6XqysvdZcUYCiXyXgGtU8Ed/a2AMZS/jGl51Eyj66HrvtLjjy55D95o56S
ROWEHh37UVL1Jyz734Y8s5i5oZblMyE5cZsDSsc/76Dj6s3ZD8qUMXBs49JUKCBq/sX9bFy3Q4BL
8GNdXxMkEB7lha1RJ8FDu+OKp5Cd+QdaCDzgsg/tNXdne4Ti4lHQ1adGyG5Wt3aKrYmM0lK7Foy0
SW5Tkk9sxG4Cz7Bgw7fAcqw4T1cnpkbd0jfWGhTyYlqjhgmKZN1INTRQJ3y30dnzX86hqi5q8Fdi
AbroGYrlY6718WN0wqFA5gs+AxAMOOKWjpOh+j/stHD7QKKHaZFXnVR980KDpddU3VG8oTj6YxJs
x2UNfluNXXcUwl5TsRiNHiMRQkEJvc1DQwEam+a7OmSjuDc7x3zFb2B8scNUt97g1YBc6Q2UnEol
r0kH+6iB1lhqoOCqFtNYePcE1g0XfgHxq1QTRG+v9HKjNjyrP4LsfK6Es111H1e+Q/Gh/KtOAs+E
VvHh52u98+mN00K1hkHgyvAW97RVGPm3roYAPKDxgDJMD55ivnkI4Cz9Xn0XMprWaExlJWSNQlSu
Y1Pjl0oMsoBFyuj9EkSO/Y14CIEkWH8mq8cYZAdAS94g5sP6FAA80NasBMs1OAejbhE/lQCb1xsg
m9xgQcGBEmcb3CG/NwBsbd8/04RVanMWUF2KLKgKPQR9k+w6+KOOuQTHaXRheU+t7kxJJm3yF4qn
VdRPwwNZj4K5YBf3Ots1tJk0YrUNCVJxfhzlSih4Y4cOcw6XBNUorBM9Bdiz8YwAdIMCJ/2JF6j2
UAdAyMAQkV3E9EtKKhrx1m82aGnqltg846ps+8fwF0NVpskdfvIXH15rWvUZM+F40onZdQiEbLUg
oIejwgB//CxZWsQFIAoRgWRHQgdkM3amRbTOlriV51aa6anZNHXWVPmPAGha/1aT3onA4l8kU6SQ
o78Yqi7NOZfUdYczzHJ0Vd9usP7qoWO2o1pygt/QXXkM4ToAFbWIQF2asnDPmXADEhCtgf/Y9Smz
trjcMtc//SL/CpszmJcb7+lkgtduKTsMay8UT6K33WSnqxTH695P7MO5jDfb6A8/zLR3iOaqTxYC
Lcdwqd9Zo5MtWUtNczrM+mZnOl2amysZnlG/abdlOg1jiG0cB9jHrFFphd6tYge2aKGRvzKKXPmJ
RXxWfkQ7kR3+RRVZEdwCOWIcqZbf2MZ8WM7P0P5lASJCgisvL8x91uv8//1lPKXM+btzbaXFd3kI
kBWiSwwTyxnEH8lTNpmyP639jecxIvtvjd8XNi4aL5Ap3gsnpzuiynmMD0upYuF3NHwpQB93Af9C
t13yp6TpVNcX/v46LfdWAX9ZmWKw5/cB2JOt+srMTHvr3RRrfYb7OBggEQ3w5Yf5QB8fXqgLmxcS
9mCfAgc/MeNqjsPQPddMdXKbFLSKBmGURCpHdQVx1zb1M+DHLukW47PAbqlak6CYukdp+Pyo3RE+
d9Z6ZsyT8zsCIXEbZXFQ+bp4YsmFl95oWkOs7RSyydf+YEN1QVtqLChurKb7ijjRan3BiRavlVut
+RsdJU79rTfJiLexcVW2ddLPkAkXM4xqABJOsZiuwJue5ZaC6cIMJSWL4x8fq7eNDKPf6rAuUPHu
Y9XZ6CermVnA+S+q9oe3z9s0bNh9RvoJGTQXOuhRN6ceoeDwZoBGZgVGAlW+EVZqPWPkxgcxJppd
idLDqlDizGfHfkqWCWLxCvZJuxv+lJpmbvbhnU3QnRbbgG8B671ylgUaODnQBFnRbSr2ogrU7pN5
781rvEtwnVJCX10Be0gQ9BN+jEDjcxvr5k24fN3kZm/GrrINz17MFv3a7t6zjtHBTBpMmsWWKPjl
HyKf3gcNQayv+suinJ7kdMyFexHoeGhCFsagBK4Wv1b+Fi4HGlrMpf4sRGRJbey69pVccuHr1uib
SPVWgRdRNBFG6BboV6z92ZiMdGGN6TvjrAvn+BWMy+MUtVsLvYaid0spAOfpwipF9uCDO+drNFHH
b/sWCm5IAyzgPYltatxqdTSJE8+qHiwZtjYCQeCRDGwfwgJZ9lhT3Er534qY+PSC+RA1gBFB2krO
ReUuqYriO8LEClWSGFShSJOjeJ9eovfaEBV7pRbdixAlett4bmCqOMbWGwpyoiPK1l55mpG/IHda
hFL6UXaVwNbzON961w981rWw2jzlxYpHQ+Cbo9oZgXRlWdEKD/xrN7yqqFCQFOrrcE85BJ3HZHya
FVnJmGjXG1ETWsxonKTD2G3JHfzFx3Ey0ocpU0wTWJTKN08RrqtZrIqbp/MrroF7IePk4G4Po7q+
fBpHAEKrvI66fanvPg+hQwpJNB+t+uHDjjLrr1SHTtYrwnDiyCvPHrKEG9NT2W9UduxAt+iIWBuN
2du9UOLqgwZPcKJCafTAGaqsvLWN7dE/FkraLtmPcDTwONHep9kHm3e4mr1oJPq2GJN7FDzqspES
i4l7GGyZCXBIrUXZjU4yVaCO7ktu5TWuUogaIB48YJClsnTpQT5aMWQo4Ii2g8r4kKmtnzbiLz0o
x3160lg/lDqqv88BVjp7siNrzCIG798zwIbNKH5XJIPbGAlVxrtdnT4azh8N2jfAis6um0fJwJ2T
iNsLis8ZF63m6fiaUxjqzst6NeB8+z5c8q8scffwn4lEAEKvqV60l4fba0aD7BgAjNUyWFD/ZD+j
9oe6ECLctWYBBCrGUcGvyIfCzQ/y1WKWfhUkNslEs50TYKturG0FTsk6lYz97JFXlBL28k3cGrX3
Aqks5vsJuJ1mORq7zH+s2X3k2xCwNGzoXuGN85RVS05nOr8VL+V61Ks2HAZxr7d6RRyCbOSA41ed
nLl/FHcDFI9+TiCgOkkntG5HJUkd6OgludZJgUQmXOHtTRdHMf2v11+qYsEsNsTHIueqv5b0JyaG
GO5ijBVSQJuJkbzdpre1vYMjuOwi9f09udHbA7eke4N5NJCwU6TLM29hM97XA4DZ3c8J7vQhXFKC
WpVoy4wpKBeG2steOcdUDkQdWyxWUktyiQcjc8NQWKvhBmnbrPZ+OthFWLIxsvYUmC4vQAg2wif0
ukujgwvBVrM4cjYHTI5Y1PDt4S5hYJ6j1uTlAs1qA3R1+aZCRcaW3G/YWr9zEAWAXptJi0BECTNx
EFzUJ/EW1zFqUyFHfEAG3h6lbApKcn114cxb14zyi+GroaCGm3vKR3J3aHnypV+HFID77s9SP9Lp
uau1uB5cL+r6cvEsijaDqnvIdDpUD3cxTrKpQYlSu6g9Oc8ZeIMX0gHe6h4gmmSzgJdQ4XpNer3f
FsTlww4uiFIDsu2LkMGiksVyFJZmHhVSph+LbC5Ex2ZTrJz+Ntwcl02T27YGArcc2pvVicunyX1X
+hEejNJz2k+WyEGHOLckH9Vf962irYYaY/vNPZ3OZPkAythronzorGvvcXrQFBiNilD+o0B3fwWI
Xao9MjFXgIkgbWkMyRLMmaSKR/+w1zcGXRiwNquDavP1YbX4q466pdzvlMe7MuK00hvE0hx7UsoO
Cfu9RTmAV+WHRseHVYGR4eFeRCDywnklEemUlWHwhBekXOpbvqUj76jEp92QJlf0U/K/8W0l2TsT
EKuAAMZ8jfjJvI2x9kkL2W8j3A03F4E728IGjffT1bcMnAqA1MOkV6k2Ksrt9bWWycKL5K9ZR3ds
wq+pvNCzMznGbYfIJWZOEcH0LDkhefL649jKdZGE1GyqgOvDgJIeWIrxpZ+j0NNBQVVu0Rw154KK
XqFi0kA+oIwQWJo5ACgmEBqrYzgQm5Aye8xa4gA5C6zdBznBjfOQJMTxGdGX4qRKuAFmgUY7h3jt
BP3lz5HuglEg2AHl4AFG8aS6S6swyvxNWlWz/hPIoY/jzoES620ON/tcsHazA2KlxFBG0jOpBEq/
D0DrjLze/koKdTm1R1f4m9UZoGfPVy9/iDHRAUmczd9nHbH/5losA3oV5NsZJKBQMfirCkPSULhD
JCKxhNmmkmo6WQywLxwpSZ+VCrwgnzCpuyghoShzo7nfl2O0Tp8vfX0dXOsjws67sVLKc3V35QR1
Zxw1/9AW46xeUnmB5bgHss0nmE94GO8uB9MTOWMmF+u+yXfETqzt0KTVH1ffPzS70HKQLzwjYAGJ
J/OcDF48mQizZugvo+kFoA2+4KyjUHMhQUVXDzANQTco+C7NxLldcb7tkeWfpl+DSaOtQeGegIIu
Z3IctxjPqgqc9Yb8kDwmbZfJDdlZSQEkgWHdcKVEtqTpoYQwQlJTVwJH4CrYhD5Ztqr/TACM3hxw
dyHBj8wzksKiCZvxC4Br8ZgM80KRa0aIm59uLG4WWaEkwLbLDwZvcEeqAHy5aQvH44qcQcnIc2o4
gKCz4dUU93bgSiWGahCAa4upehgxCb8NXVbzMBcdlz2h82tLAnrH6bVgpxir6DoSWdZ48tBvm6OX
yg5wQcJfh1y/AcBIb2mOLe6RfkmE+WARVvjNWG76AM9K0uTdATHpP6V24+3O8QDFz9LN2idN+C4G
9SreTcmg/sWw77DuOyFA4RBlldvdJgVoeRzkkRg+h/PWgOav9p9aUHahIJJ/n6mwBWaWROGyjNgz
w+dY2lmj+cZifourGL3VBBNCLq68OTWSZjYMevvcLttqw9zjt4pJdJwrJCcprvPohuaUd7mcAlo5
5tH6zBmq0y6V+N1C36Xm7W3oLCCwKN7wPH2llRmbcX0RDN87wrAfZTKdDddtuUhE44y10EojmKPA
DjdoL88nlSpBQFAkXwQpuzjjRgw8hg/hkPXjPW58yP+oxQTRHUj5/8RUQbHt3k2fPIiklbJHBuvW
ebAEW8lADda1yoFw9psKhi5252+b5gcWO4d7dpNVyUY0hNXq8yBathGFnwTOGxaRSroDWvJdtV5a
ApXOPYIkvSQQLY3If8E/o/S45lIgpDKKSf7F7C+xiLpOndd3tP4Kx/D1pTuS2OZirXhVPW1PZ3Uc
eSikrJV3k53pd23mtPQV+m+f64hIxijZL4nMnruCnau3SMXhurxGajq9w+FeeSrKhWl9/kyKeAKb
id1xUtfHvN/Snj/D/ydBPKROF3KNpt1biM7I1ys5de/u+sEjnN8N9PYoZATAmZA9uv5ukYY0pBeY
rsI5tZpvr49b4YrRy4iI5O9wpjRQfAqGVlWrhjdnsXvn/8hXdNpOvwgq6fLFHg/fHxnPpGKNe/5p
0JL1Bs1Vm+7j6q4QEBDYWTQQ3sXGaa8D+lr67JmvsnsmN2ldDK+WoKJYsuuoboPfFnZOIiL+KzUg
ymJWDwnc6Rz4xo9Ee6M9FYFOgc8Mkgl3+fvGS1tg7ZFeKXdmI68rk32IVOg8FH9Nrbt91VQIhJ35
dRGhebMpKwK9wohtWA161Lk+1WlWpWSOqD5bMzL36sKvGTSC8ocabrMdvl4p8MHiB3rNPsctlFN8
S/luJ5KMXYiEDGsZ7uc0Hs+V8nCT52UCywPQaASjuzH4As0sP1sk4LzqNHrgI/RiWrCbHcIWpaJn
+KzUV1FZMUut/SiPc4cOoMnv5I6U+ta9waGgyfCD/iUvsVjW+iSr1OzrkFjfFBVxCbiBa1QWhROR
BWcMUJ0+bnh1fnKZhCUttdaQ5UvmZMmKwDchuwfm0MFyn7sTS91EyPlbydl4Sk01aOgiDtKabS26
zkf2V8BGFZWDMTJW2vScI/CqWz2FWFFGM00tyr1YdcSQ9Ne92A/1PnAvHzyfRMr0wOILk96UgaRn
rXkIW25XSlTP+7JjG7OWykHNrIGilCt4KeP7nOiU3ieaXuNcKW3oZf4UCkco68FaMAGUxcn8XQxq
HM1N2BFsarlk3az2tVviVUY4Q6D41WV8P/8OvTtk/ziaidQYwCXpOhs+M5BE3ezXLzBy42FdCp6S
NiGoOcpNoTvjqQGxuMCa+VEtgKvcs53Fz381kutq/KsdZ4KMYyHe+vuDBj1ZybyGzX+y51CU54pI
XkBVJ6kTX8c0oYrKymFn1e/KsjVs3SZLPNl8NVIJfp2Q1LCYXYsEAM/HhbmDXL+2O8QFA+cBFV+i
M3yDpSEE6Mgj4nT4rpoOZiAW/pFNObVBvipNLNaO5+Qr+TBv5OA5GvKUWE5r2D2LIJsE4Oac+I2O
zTJoH4rBntUTjNiKTJf1zLh/1Sp/m/VvslNsQZmoDRx7OyDxdvXkyjDLC9f9mdwhwbEYOOPFg3rK
bnRhS05wQXuiPOhTx6dmCnEnqvUitNJmwZaZT+jPh/pZZdVXIWT1x9jafWI7UFBuPFUn8MNMSCN4
xWsZuTxx9dFp2g68Z0/NmxXuPzI5Tb48BJEpCoNn02+j1OX+Dg9F5L0EzI0wkCs7xFgxwJiVzv/X
RQaazqU6nJIt0oow/jj21QpIESOoBEl1qKPMqm55vY0Na7luN840BpEJxt0Xl/lqtrIKuqP4sABb
L1G3BNKjkOMUDsreoJZmE5jcUlVY7hdcayThmep7Gfcj7lRkqG1c8CoWIoc3kzWqwCrvXiQeDHIE
TuujG/fywNIHBdcSx/m+aIeoJMZhgOgxNJdAUkguUguyHBo/qwlN2vP299A7KSj1WBCpDjrH2nea
DVOlmKgLeW5qcJf/QDUFiOleUxV08/7jPeREmreMfhCyv5SaqSd8ug04QOiqDIf/0+RN194dv7h3
4RlxxI1VTSccBG972kOBrgmavd+OrOZ5VuSFq3UCXKhcLhHrFGC5PlPPq0Nw0qftc5fdAbF7ahAC
1O3/MoHPNRE0QcJJcKAA36IP8Ma2qKnHqLO7D9GRJJ+hb5jCFKoSsizbm7hja/nGQzx+hvx3Pkvl
4baDzsz0PcetuUghL4JoyKifurF3eU7knSrT91ZNCX0nOqrcbCtW9hKvjaEHsyQNxKp/BFDF2YXH
ZbxKL91oyarvsetcYvEQHjZWngyCTJc+UyG3OFCPqNyHQgHfkO8CGjeTX9XVB71eDLJy32QR3/pF
NH1V6uxPXz9KR/okavvjGcvXZalrAd7o7dBtY7OE+VA3VQ/P29Zg14wlbTIpWZ7ucsPMB2W7WTm7
71b3xIqS9fyF1WOuU+hZ0d+NJ28nd3iDr0LsDOfrEA0eoefDZQYYi14QM94fx4G16gdLy3IhYita
GKkRw9/RXKL8csdb+EV1N0gR1tlf8MHsyczm6cn3kQYe4IRgsray3CCjkrPBVSB74R71XahDANSA
sgc8AvzMMt5/tHuBSVlfoOEeCIwPYkdegI85Vs8dHJ8qVE+789y7IGa/Ih+IWAn9ulqm57o+AY5d
yIB6kV20bc8hOeCaPkbhk6kMqeKlib1CexiHTYZhQRakIZbNfwuPVnkiLEBMOuOaDxljU4EBs9kT
GbT8AmoPm+lLucHKgne6vXz6QR6IloeFbSMQZ1nP2a/JIeOGrH9+hIryMEyG85S1Ka7CPxyNxzik
/soI6scgivcPIhrMQSaMlAtxNPuJMOWwnZtBlLYAJu7zXS5/2vnKjt3T0WZdWa0OzetYh9WUglQs
CWO4AmtKQMmR0KLQ3qeDG4LJvL41sD3L4Ih5QAWud/rq28BmJMlhVa0XF3Gxmu1/tQnrKau5mLBn
/y+R9GfV0EXLLBbLO6ls8ZkriLYaMvM5u1J3ZJ3zaZfAz5xO17rkdrvhdhJQOaWc7Cx0RRSIXWwp
jRtzegxXwYOkZjqS0avnixA2BatQyi6IB3Qr0Tv3w7HvpTatG5/YSdYbWPtsNCim9sEG9T5LZkDl
HofM25+uGl6Wt5hRwrqoS4pebWJtKFX95OujlAcVdQgbHqbZUB/cdSWqiPe5qR1QVhEP46CLFyMl
yganzDwpRg2EWJU52O2h/zuLW147Xsbk8PJiUEa2OzQRkvphAJPkoN3BG4Ba+sxf4Zs0UBcO5ro+
MLgxOqQ87TTmyifjEXZca0BgnSowT177koZTNAwnDmRfl/sSkvV0zfBmS1KEx++krc19oWd2ibCF
piNBduZt/z8wK2vu+7xpThZmb0o5TPF2SFlN0dAKjTI6a1+CkJJjTR/xWLK7pET1mrk3E2HFIAz6
GBmMwG3QukfoL+F71Bk2J/f5rULaVVmPOrbIWe0lyRYOH7cbVDdDcZS6zjdm5Bqaor+mgFkzuVfu
kPal5rpJk5Z6Tz43ZFXVIH3BGLpXa3FMotLVqFp8s8JZbsXMKqaEKQDyt9LhZrrXeM5tuxEoKJgL
oGWEHaDfXifNi4qSbuQ64lCQXdAL5eFYMRyjNxri0SXi42yBxGeP9g8cOHFlrAU4ykeLAFlRCKeJ
lBIYKT9pdPzlask1k3A39uPbHH32IHVXexsEr0k6yU2oadeu87pNHSDYMAikZm85+Tr8u1HJdHF8
A+5ZDpTFKZTEZJxsyONekL7aURHczUjUWBZt8hliPvN9ZGDtHB04NMCDyZozu2UejT30LlAYptVy
Q6TNQnDkztIQmEJG9bWNV3uBhl/Tn/945ysDmvANUkdDtnye20KblpUGaVZgYsx5lKXUIUV3EQVe
i8UshDqhIyBi+mSWlWYRz4d0vOUbMGBC3rdSrEgLKM1ExCVfux/VbBWOecC2XgUodBOiNkjiR1Ya
3wZEA8PKd0tHmtp2b/DWDkjtpIfZttf2mhlr5wX9Wd396csENtGRUpf0BTmHv0sbo8r0teqZuWBX
vOd/gAD2p3K5XSjpG2IGjxwri1OyM748OxX6MfbBqtBKGQoi9s6m8NcH/G1rMhsK6gCyoEZ3hqGS
GVOIELOHAT0IVmY2p8j+fO7z3aObnl9XD2Wy6XMYucbLrgA0bm6Kzb25wvY2gI8VZjZHMhyFOGvx
iVQyICKROkMd6gUQUoiyidKYvT6mUYpjHIR3ngBem5RlJz8aA9cZ4OV5w1ABZK/cfX5JNv4Blzq5
SH3lyruepiU7aLErJmNUShQyDw7yvTei97Q8qiynKuFJbqFmIOxK6r3XUYtpxF15N8W9vNPSCm/c
cTIROjHBYWBESKJ1ZY5ctzAES4naE4P9e+I3i/M73ClVQIo7g/RY8bcxnvuevdemxJeXEU94vASH
6LebW5kZ8waP2FUK/KP3BPSzzJwUzzSjjmcIiG8kAbczXr+brvurLZ0hYvpHmqHUOj6ngd49Lxlc
JHy0px3FYa2TMo524zffi8eUSSWaqhDgMzfuQW2PH3J9fZR1ar18gdlj8DjLnnRpRQRNbro0aF7n
sN8Yrdm7vjpLaSfW/fxqpUwtTORH2kaQPU0RDeqNo8GUyQVAmLCsPM+jGRSO1RSkLewariKKZ2I8
EdAMvbYWevnv7JUJH4Tvgcp4bviD+A81+4Jvoi8d9KFMuuU/84vdkna3149rty2cMrleyxLPY+Vc
5vthicZri5A0AJYmoBnpr2T9MwuKdBPDjSnzAzHmIn/Aw63eJ0E8GsMSjZKzypbYfp90Tn26l0a4
KX6zcNtHfh07b2CR3fRFU7uROSVALqChK1O273ScQyJspuPRuwPhreJ2wlaeH+BhAmHPYzAwN/3+
wu6gELDmsOupFCTqKd+0bfoKtmOwp7M0URaBU4KxFgl/kTCDM9AZ4dDpp+K87t+BA8voxIoq37Wo
epMf9jBre8Q+3Bxmt8fS+E9AUypcoBgytT/RuSibdwVjBl8xktxjCqS8oNHYVMr/E7Obq9vz3fZQ
4Wi1obJNYqY5Wkfh1/i18b+cxaBuXyyy8NhHp3uhrLEYQNWCifRMCFhzMPJfUHCAGqOi/onIgLJh
k/uCtcPE/iz4W/BOr+3hZkDbhGUzo9PY7rkTrF8Qgdz92IrGgtQduO+xOnHtR7eRAWlP2ES0c37G
qVhhc8i8xVslpyznve8s3W/biIxGgxHkcQN2hi6nKvF68Oklpu44oK98WgnC+vupulzrVFIy9X6Y
+wt4IGpaor//Sl5SHyEoRys+kxYIfWkRjfP2Lj+u2XkjEPqgqdiCT9lQHAiVOxxpP3QSJjx6xxPm
nQleTAYhidW16p4OxWOrAi+LMMyt5N7a5CYXFbfX1sUS3oetrDoNFZIW1NFjQZ/Ddf6YiSlk+yv7
WWTIdeHdHzkkrtvNd7eGzwzC6hYSrJtUSSLJADwETkE8WuVVYmQZpj/M4rUGsYIEAJ1W4BicBkok
dbiTzf4jU8qx2DiKIxw+3dYJxOonS0aKS3cDltk+bmHzDovCL2+PDsWeSL7yyAra6cLl8GNlq/3G
kSLnPZfIxXrO8kIm4/gH0ER4O82/T5r9n1dnYqER3PcriNCETpwkRPj+dTcJciu99Xb46sQqd52a
iQ4VT/XYnR36VdyyrePRHPYKUH3iF2O37iboEPQxA0sdOqNr8Zr0gybjjSGfYzLQ1ft0Kh+2kcWN
9+mXyzFxycpmyN7FnhgB1NnI/L1Ikn5YefhpQLQimzS76jxNjk2z0LpTFqaX2SA2Lll1j/D5W9mO
dP/jGkzKrAKX5IgS8iMu6LXz2P4DDf8mE+RxVnDJUuvKs/AWCrpuGo1YocsCjdwBJTNcsQ2gAlB/
vfGR+vt467XicH5Egm55STZ/6zkVxilzuTt/7v7YBMGiZVbLSQB4FK1gXOLhgrRVGAVnauhu64SB
Z2vzneEPmJjI0/zK6bNOe1A8aPtGpB9mrdZpvTh1TCccBWZDuSF9MuQcTzRTf9oy4h2mOVMAVNNz
4DTy715Bas0nPgqUoPwUpf66XKgPj411NWtS2NHqo8TEhaqqyfe3UncMBfUJeHxf0ZS5viojp7Gg
Zua2K40AIerOB5EeHj2maqaUoLuqMNYFnRFynkqlyK9cawix0e0a46yEp7iFC/aYOB+rKv2hDYwV
igJKk8aRi0xs5u9vCoSGAgcia5x/PIIiObna9/IHN8H7a7xhg5G7lNXaR1Z2/5gtahTE5syq0pwJ
/YQdpEmPfcMxuYAMyEEqJ82dRgudIPXA9BYUCvf4mO9icMCGwCiKfPzuh7UXaT6YyU3eaFGGdGJX
48Nbg3XSS/dkg6ktbrb07/n2oZsu0Hi2ZR6BleM1ASFXhubBBj1dbXsrKM9vVrCE2vVP+jxzjYDc
G2/3jfV7GiYglPmQ+Ac8dtTez9DwuJS9x8Z53EpmAxENtZ/ollhWznPTWP5MLHOk7SXM79fMkHt5
XOAEfcIsnDXCjcvxyMciUMOmWwdINBRBLAz32URxnQrHZNhL/ARpMJn3kBBIEC56bBDE+2pve+UR
ASx7FHQbTMxGoLJSGaa4BuNXXal/OYz1CNv5KLnvdZG2l1U5Jw2fDg7/xp9NAYUDPQTC+CWJbCSc
JChcOgQrboUsHdB0Cvk+Ux1rwXaAeUhpo8OEk13Uyd0tZlevcDbUAtMkNm/p8YGPcz29reNfRRW/
sPfjpabbGG+rcovtMfWxUDOBWwPx3d+al7pOcrKHXh3rSTv15CXWF1aeeeWxbpVkG3RHTQRf/QM7
4t8x0qX3PnA1m/kSMjuUsy1gNMP5lHJyOGypPF3X29m0PWKrlax3SLIdzJ3UFoaqAd6lKW4s4zdl
DOW/usMz13KEmI/chKAHr7+KhzYtTVFqJldqQkkkzbQVdR39HteTP9UwtwWDEvm9/jOtLWUSB4b8
dWHM4zwFL5w+JeT+g49xDsubmwJT474ErPkTraYEdxblzyPKXIxJW0LSTCFW09Jmh93Us2k5dpWe
LsakVifq2i1dqQIRNz42HpIsutK8CmKxqx+n4FTakIqxrPx6s2f9CS6nq0LCpYN3f+yEW3Ob7/SX
jk4v5YaSym8KQKL2yKo21175c8SLGzNmdAAWmQh7NUnNSE2fcC+7Ttgvct/72TsvjhbccmMpP81N
3koCxYMIjuE3qWSk1It+2FqZntapa/DiZcXqVmz+6V27t0oGMXTGfeR4ok6cVpZgl3S4AXGhwju9
oGmkwDG5s1wwcuIlyUQ1Y57opxFUe3ZBMMdm5xrldmX+H/OIHvn+Mz3PK7aSs2sorF0h/0eP/Ld1
ivpBe0c7/aSXPT1uzU5iaC4Uihlee2HRbmdsmMi1iuYQ5CdAi5KHc8wI+MnRQYYbfHKzRruvG76j
7WR1HuCZeTwla3sZ+rnZq/z9QwI4v5WOBW2fIRvy2puiXCVAQBTQIa1tc/a+QPz4lks32XJSV8dM
PSK26C7N9M9DAE5XTV9Y1KXiOmrIzoR9GGUrulnkMa2JQLt3Kbr40JTKsQ6aE+bLfv9+VwG3sUVV
ibUMAkFawymnI5g6h+82xpx2DmfDmnEoEhKj6alIxJ4TwCZx6BBZdTIKv4DkBT8v/qhtUBM6+YN8
zSsozYNKRVa4FY6A245r+N9MvUCTgZ/uN8M8mw7QjprK2potGSNEzFdQk187xLFTgh1AIvqoVBfV
C5omR2qyvfBlgvMM7tB41he4XqbS1I/FSgS2hyKhLIxPYUH8cjXedyKqNPGRnYC9O5Zhd1k7ceiD
U/LpCGZRVqrXOn6qfL5qYFvGxfO8EloXb6Z1c1AxsyQVB/UI2sI68mhGXLS4pG+HjpnIcimorCCQ
hs4UYdTRP/53DOPbmDCMeua9VHnEgTXPnsoZavEAm6WKQDw22dv80LzyU6Vn/OrlWdLzRmKAOEgi
zKsLp2IZJtYX7buYsp3lUv9GnCmCEDghiK3uSUHGWFhaS8CUGoirv2K3lhPCQnFkY13BjFwSrfGT
Bh2rsakF6p6/Yop86Khx6qlcD5hb7VeJWxmMg4pEQ0RPVUxGqbP4Dm/F6oW0d+OlSKf6zymecum7
V4H9UFW2hyekbylxp4IcpADIcuMnW0eG5rbbYwGTK/LtWudTPkuX0utHtNZjuJE5yDN9EUU7QKqb
SxOx7t45dKBoEpde4Rv34DkAzu8h1T/nB2ZjW0CpOrFd4EFHRZSvMuIwm5nGuJ6GOdPn9hE77+t9
1JdQRdAXw+A5cuMPpdhpU1OkyNe9qx3oFfylkzymhj5pwseRI7gzk0HMqXePgnXs6hVMTYT8HmC0
31q7xu2Wks8SZtKSJZdtkLs3AzqB98k+eOkU2iE8qQZunElK2haF1/itVWWvRfitg1BCM5ObByUe
A3D5QuIDirgyI949yXNjODEAoJY2gMpOACJ6mv0GaCLti3ZFyUEjBehDWxAtmZAEGmgCDlmRbpm0
q7uKGPeT5qUJO2VAC1jWqg1iGNjH9vPpoFLI4sc0EaNe+ByHH4oug8PJc2QTwPBOSSUkHMnanovq
8EiypO31rgkfpAUAiW146gj1JL7iE8Hk01hlg6eCrs4JIWkzIAXfRm9DUsttPrPnmhvBAF8yGS/3
cWBN6olwtwqHsJCOUmtbc/INrXLZBO0dXhQBrN3jV4MZoKRqUiiUaZFWlMHzb0gZa2eXxAhTINL1
u1P1HGjWAiDa6pE3wnumCKgEH/B7D7jOOAu411DouV/NWeB2RuugIsbiyRCWXZCDIanF26fNDP7g
Zk7+gPV9nqrUIuXWW0nGYqsz1ViAVHs64NjCRlOT7qyDPIyv1jTyB5lK47Np4yfqqbnU4bSSMnF3
rBEBq8LzUI1uoKdC+GrpmOcnRoNC/FMzLdyKCed5A43feqy68p6NVfg0XygEybeUvpEEAkJQyyBp
7OP5cDQngoc0S+q66HvwM5kyoY24wDcc96iu2ISAISI0Stj1psGNTB1j04vvEE5YMCpaM42VhGLU
5f8gCidKMD6HtJEuK8w3QEQYZ9Xmo3UZNqu34EkcWzZFllUlckkSwAyZ+QcepDVOhMwtd++opACC
fmKi8cHL37xaQ9w13w7J46yFB6kBQHuVoRMu4KUVkRYmA0vUXUjrjnH8q+2ATPpvT6iSdzDkg048
0Z0F4ZnSOCxhZSEwdMKlq5DdmCXFToZQkKFkdQ3DH/VcBIIMcrnXyiZjRuuP5XbGroDxPxuTIsYn
7IN5BQEX0R8jq7rFJYGJmASNv1FmVCsoy24lnNl8KXdl5GF7yIQalSnq3a9z7TqSvvf4Hh7G9f6e
4KLdql5KHqWO9gFRLe1Sw/9Fh4BQ7S0G/84tI71r8jya6MGiZo7u5gRjch/ejpb+kJEDAvbt7boF
x3cpTmzseOZ/Qn+t0oGAXyQbsGFtobzQESTYBjJeLFY3G28M/JCB4BD+Ho98JtzWfNmY6jeXSOGO
EZ6Xp9s04vRJCWCie6QNqhIIQkgW1H2DTH4BYGXgB0gz3t1Hu5VkONyuXf1y/A+VHlqyXSUvfYSI
lJ6xKy6s6e0hDJSpld7Ru3LP3iZSVtAYEFU8/jIE26Hwm6ZFDh3nVmC1tmbpE7ZIG+2JEhB8Ja+T
c9OuOL00I09gHYeSIZd6Mz+F2IQeeomO717RDwIhqp6pMvo77Xxw9xSDTPkJ2TyX7hCzop6AKAsa
YcBDjNpDGNzqngNf2W/k7HQ4fbUSd7aVTtb2fz0LqVJe1dhVdDcBQHJbU75dSurAcH52orSQg1u2
zXVFLVmWOfSldRfikvcLUq6uR45yjMMiD7Q8ItekIspSB6Drd6SNssH/6J63PpL8xTALiwpYPn5e
X/x3q8JLuyJV0L2xz0i4+7zmh+u/LZrgWY3HYySAvgLsJCZBHsml2b/x7IfrK6j7X0vvGc0RIejU
A6nJ5a1UKeyg7F119RSUm425lRZJwMoHMu0E80DrYD1H4LlWZKrFqBU3Kh5AB7i0OZuB7ut/+Hkg
S2AYW/0dgRD0Tx0zn6vmrVEade1/pM66pUKP3Rp0J0Ok70gFaiZfFg2XcTfS1rVCm46eoiBn8LeU
bPVczauFHfWXKi54DaA9bqS3S9MBTZHMyCtgdnbC4NXIx1qzV+0oPLjlTHHta1uT1+MIce39KgBq
qiW+cgqj7IyTVY4MsN177/eg6/+dQwZ7Yw4OTzAQqJLwSv9sMWeD4hyy1SHrhVZdVnq6Zc0OOnjI
1/Y/W38lnATvQzh5kSGPDuGnxKvZD231Uv3wsfAfUnyS4TAMixgYgvs/mlg9rEqwwWP+0SwmeMie
l0ee3nLNZbvY3SXWOd0tGPqpvaEefY+WWOf2Jua7uiETSo/PDAGsiF8UbZA4HHbdpbvOqgalUrox
JDWJFsX018YhzsD9oFjYiYzVi+vtgiFiVuiF6dLaDJTWIkiiUFW7wm0sXKCIVSHNYJIBjbYrZJup
gLcPeo0guqj3b8AQnWuBNMT9s0Y4xQbRfewGdhmt0+HsAw6SznCoj1ACaR4rMzDaKCRy9Fv55D/R
Bn8fzBxu6nFB6IRH7QdjlGBn9dkSJjAeBdL6RaPFSlPbU3grTts6Awb6sWpMGLSrXv5SyOKvkZ2p
u9xkDjhpNsR2ChiFP5lD+6HC2KmGBhJfpC+hjIBw06QUw9QUpmE2WitMRIiTKmPATW6Bfs3V8tGI
uZ9LuDLB+c5Ctzsze5E1C0408ZxlbueRwbf4fB7yJyQO7lR6AEaxScQEicy/8WHF9SP3+tSszm+i
8CvM3Ma1So07vY0OJ6BpdXNd7cN1S3MD2Man0xmsN53EIXRqWe17OBX+nmoUhuGOAHFM53Q03QC3
UfxwmoG0OquklT+ZJ46+YKd0vN7chWikLnjkMTCce7wEnJCEQ1RWNaNfFHFWlQnc+Qfqv22beqhN
7QmxbZQpQdkJ7XpvJ9BY84kcxtjvORlrmZMdFZoDmmSPxIAKBLJfZJpjYz8zY8auMzLyNd+XtdFs
KcH11NcjTIWfica6LEeyY/Xi8YmTCrM8krXdr7Mkl3cS6deQAbVY1wByG01hrRaVvKpr03OOHs/q
YWjEXtuZPfr07uvZZn+yytiLbDJoOrnhlR7UDklUvPQbC1Q0/ii2S4m4kHgxEfi0ETMg0Igho7Ep
KdloqKwggu4yZAckfxwwNQRQamE3XQGQtIOOHYav0OjvxOaMmnY54XzzgkCcLNuYFS8aajedRVMN
nSXixMvWMMsrmwUjveAW1sMjTNeKCb6t+2J+DUj/1EwLSmfb8/E/6+Uxm1L4Kz8hIeFIyfzJl9lJ
YHz89EuTSxDg/9CkhoS+uSPY5zKVqmMvUcQwasikkQBNL5UhokQ3J6jN3OT1dI6XbZzXMF8hJHIF
PEsykjWRwjhiehI0rvdnFzaEHcctIGDyP2BiaYonTV1hyJYNKUV9bytDJUxBXPgTZplt60v7CTzP
OMzwQoYKr2ea1PEHwMVmuYxjrkXgTUkp72wawCArYkhgMbfAxZLzXTfTZRZIkb/RL/S8vfp6Ro0+
RRDxQWtCDGwBOuBh7yzFUZwjH//qFoXB2wR7mWPPUdq2VWZHNo09kDPNszEXoMhpcC5yQajJ6ZqJ
1aBJCfcqZgoj5vCxkEos4p4i2H3aVpZBwLonB+F+ZTt4A29qbbclBoD7ZyzN9BGcaLFGCR8h5Ehw
NGfrqNM1CY/3+geeJB21KwI59KJ8scuCSEcQapY5/8cc/J5gBk3fej4DM9xtdurcBjYt5/xRGing
+3yJ73MqJ6uhuO/JADtSybajsZeXGH4xg2FQtDSveMfy+kufZX/7YW21d4pYvZ/oNypdSd76weBk
6EqVATalIthrmdWdJgeHAi7mlBtwEo2JOWiEA9EWA5c1WAQhdUtn8W6jP0PfRvCnovU9ZyhprMv8
32xeqUyZhiAPEVhYO3lRNVZl7u40HAdr35grIUHZI2ARs7R9j5P91KCsLx6uzYoO1F+VDbhfKQHB
1gZtfPlL6uH0RPvRJiOD/YXuHVpSgKQmRxSJY2pdkMd2QnAHpTVcuxes4O5r+CvFc2W8d7nSDDS4
DbdCxqzedPSkY0OBlJISseSnEUiUgtz9Y3/RZE3qWQ/fbMr5BBj376lPy0TmY9ixVJBoqCuNXQRf
r55XgqBB6KbEwz+BfscQMBKD9g/XEOmsdNLxD/JPO7uSMtkPTsgYYHZ0BvEY0KqItDwJgowUxdyY
+wE65oQspww7wmVxnfSTGa4xScWKEHRRKGZFFM7xKo235JNU8C+x9zWiFpFIbW4qtOsCxCTUW5B3
Ni3Vog4sMBlUfszXWhk6T3gd9CsQldQ/BX6dt7H3P+QP+upFJ4aMqrzEuoCYCxAwlblB7ttOIaRb
VumMSEGba55FUk3+Ixb9h8IYSfydJPjWw94gjCDPX2lMPsZLmH2X3R9BWKYpT1nMRtJvmR3O/v8z
opUxvb/lGzYjWUOCo22qlqJ3dqgcRV9S1l9b3fvzwa/kUB+IIXvACkjRUlgMLHTtl2nuRnEru4z/
AYE0PTyOd/HmNDIl+x5s9ztm2kr5+lzAp5l86riXHdq3ZoJLMI5I9yt3ArsczMMFX/NK7I9IAKs1
4veK8ZDOVtP4hdUF+gM2nNImsRlCtxe+ahdULkq8EaGK1SViAxpd822dbw6r+l0o3R+bnvza7E5e
mL2d8JGB9/NrnZwBzvBho1Do5ZmDRDphN113eAgFzWwO9bsznHqU1W2byUMos2nWYn9Win9PXNxp
0qDkcEy0i4wCHS2sRG1mXQLMKYs0ITEhMC7L4W1hrCVYhRwBmJ6GnwrpGyD4BCtwEX4zLhf4gRGu
0Rz0wcJWg2HJjoDbeDCI5r7XHtli5377BnNvplINIgAw8nb0LcmdgqZ5Vkg6WSph+wGpSXDIR/N4
A0rzZ/zKM3k9fgCfMDiovah0BaOfwSm9CHgYODfYPc331yCVqAJSah0WI5b/V9eUx70T/1HfOe/G
yktQUEQmbptsTRS4/YOsuyCQ3VJUZK1NLA/hHKD/Ifm3AdevUTOvkH1z5McPxpgOFNIQn9Z4c3FE
9QTG1eALt4ijEw5qEMwdtq9oc85EhcriOtPaIeupqZYdHfTIKYcxJjW/wZmox+/3JPo+Ws0T9YR7
K8Q970OXrKU1DJbFgoBTQ6YUmLlT27O7MeEoCdB2sZ1lUeO6sq8dOBmmopX0pBeEzKP4Mhly47gm
Uy8Kri5HPhD7lwyMZRtWpdTLxBaaoqz24pPlZPlcLUeBjhF8t1YyyUIsSyQ+59ouOvBHqDhnBLjz
nsSlsP+IrTo3srv9ImpWS0u3BYpXCwWPcTG8VA2lXfQSr1rFZZmqu8Clx2kUH4Go63lbCRHox/ay
XTvFywO3FkSULWD/sxTXQj2TApZhrpdl7l0Ve5yU/LGVlm1HMiE1tkX6Udai7GnLXQyWgaxfNe5O
/3XTZkGkqx2OsX6UynL7XxTRiBGlNT9RS2UFDsp8bKhTWwN1RiBMPfj9Odpum1XqnqhwZPe030iM
9IDS8ZNQtbCtckpamdEwubT1jN131w8AIKTHKhk3ouDyeHEDVCtVOvZMAJTWH1Spdi0wU15qCvwl
PtNPEPFGp+njl2AK8RjKfy2rcReeDDKr5A8iunMl7zLYp5E3xG4k/bTwCfXVVCscw3+AOjsZN5w8
kDNyUqZsTweqSnGlGa5DhVERYUnW/acFZgzmVQoYx3ntPhXLumQGTvKOvqYlmxT8d6MlD/QAjw/+
MtofzJu6KDF3BPhsZH91RkJcf0QtSz4lzSzIM0pVeyibi9e1cME4NFbE01Um9Er4Ljl9VogEzu1A
V2xZNLU809wRBJB+b6ED+ZYVGWnw/b1OMZMZVJljtT5w0vqGP3H/DF94/okLXte8RnkeU+TnfTOp
hNBa1O+eyjByss5BpSnpKVH22vDMM+TIXMFnLjDtz1tAKDaD7Yrg0v5/l55epC2uviXPAfCnRbXi
aNkI6Qg9DDmEhGQr9ZPViYRNcAVl7O3aXgf9jaFNuPRQOe1y6Tnu4xpSH3NXnzEs/INQ4EjGDP6s
a9cXYKKHeQQ0J4sPsRou06BeJo77RPjQ4jGvHkZm9H0A3CbGWRPllak1JQArtw0fes/VoRPv4dOD
PHDJkNLW9BcXLMQyMTo0m5f/ZmnrrA4HLUZqf46HmyiZzGvhzAyuYiNDN6DfRInm3kiNoYLY1Pkt
xP9pfOK/UStg9FXlFr1oaX1gV80mWeQUS9VxeguA0L/KJztoY5FkUdcupkDvUmkS5zJn4teelufv
SHrQjhSMCgu+XbWTkJc12ZyoYu1wi/TsqH1RTvEw5ewHEX6BuNgFqShfGdqWzYOr+iT4S4fT5eJH
CGk0xE/Cb0gwhmLEtGRsj4wWfHopExBrubL7T0d/xs5w0JeIw0zPqDJWOpaF4o0w/IrM0f0ZJeSe
Q9VKs9YuwflRVdFQfsPKz1EvOujMXY2NOv5qHLMVhx0abYly8WmaHuqVVAsGJY4XkqM72NivOzKW
YU5yfjC3DXUOwnF/h8ihIz+Yf6RPQMSrFa1e4DI2KWlgqJWdrJB7QyUSpeV6rNvCjvq25uXzFXb5
NKDz9pxRawOjBsgFmskupvlDCrkOB+Q9PAv9+uGQD7bNdFpIHavdMg9DZe3yLYD+B5fFHHcKFgJx
KHfo1Egbnq5uh/0BPPvpTQF+8TkKBSrWN07BtYDFobcka4QskhOa0GR8N04EplrgJ5vJawd9DA4A
Nu+YZxhuC9wlnP4ynSow3aDpaqHge0lt+O2eG5ALnusvFPq0/NBLs4pvlujkd7EDRHBpzsxQASjm
MKC0g6jz8UBdfwy49/KWtNf/VQFHBnm89U3GzRlZ7e5M5TWGLVmDLjX7Y1RgES6MVKYl6mqh0hsU
5R3RCJQNKn4qWd6f4M0ahSgTtRhS9fEzi+iFvKLyFmJiQuft3ILwJ8YMPWMpUp/MObBxyHpGlZ/a
6/dXDA4RsHZQMwClh9RZj3yN9DoMZnQ3ZbH8LXLVfd2DOg/Zck3DMQoZTJLy+YSsbAJxrK6B7mdE
Z8mwbfijLSjeVnHo+gFRkPMdviD7cD6WqCgmrD4tsDY4aaofcuDl4Tvhej8yraX5Cxh8fpcd01fP
CrDmlc8qowftJi0vak/LGgaG4fTtqF4r/UIKPqQhljpOHYcb/V98z1aPf7CKZw9JEJsWlxzs3UPa
CNiZeel/Fa34Bt1zWc7fWymZf+AvKDOt3CQ66CHQafrPGX+hRMltO4qFXotl8zY91X9vFvzX69j4
hTrRxR4JyBPOodS+DDlD19ocgtlmSSUsCN845fYXcEsdl4CXr8+Er+9PcosexOyAGfjSMgEd4Fry
boTQQDmT1Rs29LgTvS2qhTplXNfNCRV+XlUFuVi0KOg6fTShNQmOgI8aMwu+UeZSIwJcQxvBfCM9
/mMrrOZ2AfRrKrnnNNW1IdBFixLRLvPFmsc+VSev6bn/E1beeWxCVeVGROqaxix28g8r3zjNu7Q9
AQWPZ58ORZ9FpW90rrZ8Nw1+2MpwyhN1OEpfDUqQHA0U7fCAtOUITw+zNkmoU/ZV7UnuR/0aGJUo
7wepHi/AlrocnRRM6HDz4BfYEGR/Zq50SFHVGkkuvmuA2jqpbz2rxjtpIGzfedPTms4Oco4yak4K
z6YGshjum0DObIMivK1GXzo7dhmB/bte33mx7/pC0756e9qSd11max42B/mXLLxB6t/BcAsIX/mF
26c8+EMIr6O8oJbPJjITXByF0TLG1nOsVjsNQIN1JQyEihly70LlUk28Eb8HVAI5YVjpdur1MZOH
zGccFG6goEfH2BWQTNfuIUSDfiJMThEm1UCXPAym3RqafkU7Tqbr88TVt4ap33cQfe7DpkOzr0/E
0q97yKB9f2RiP/1Zb9HYwlbwuJJG04fYRffloxZ0BlifTYLWRK4oTKSTorjKLGVcwFSfCHVUY+Dk
YU85UPDQRIr141SUQ5b4SBSU+17o9w7V2XuznPHiykkVM/wZtFXZoS+iDnrtMj8BGC//OjI+Eb6E
IozgKgfh8PUDNHgnqGFBQLh6+fo1olsJxHJ9QJOrZ+63uqG7BaqdsR/RyRHycRTpoGg4bfMvrUWw
Trttdo5zWnsCpJr7wSdEMc/RgunlzKVArkgGqXmksklU55tEagm2cDU17fv6Nj2W6MnJVPn5teNp
LHONz7RpTNQhvxnL0ga60uxERqVzAHjLFzkQtFrAowEzGI/1+Funv+zEr7wOOSMpN3VDuEww6Hx8
voU0K1hMiG8c7iHYXpfVQyLNJvQ1xqqrH4PlNc3/w1v/OaqVM1LvrBleMZqF3m5DW/LipV+DgXNh
CCi7mgW1jUlKKhJO+ETy2DvaYKbbX6D/qv9XC2H2zBqoR4hAWrH8egAlw6sKPn6g32te+O14zLrE
pU2jnSwks3nhffCB6F5kkxNU1PE2p+43LwuzB0fLKSpZLa4cPg+KOWCBNvs53+0QYWN6qsYq6udb
tDfTUwEdEJskTIXxpQAx0BouZCs05gPwvZdWzyBpzCEelzeIiBE+BrQyiLpoymfSPjAfpsG6cMQf
HFNxniS59H4osmnuDuLLsUIYUD/mzLFDk50gezEXKi+FuCNJ5CKOseNVd+0j1I039atPCcW7+hrD
N2FpdxxiYNDXoXWo7AcVgA2L7vyDYAQkT+FD7GwL0NIo/peXbJdy5HEE9u1kKWVVOak/04M3VzKL
qo8steNwkp/0j2tQrpO84ZpgvM85myeb+QqGu6/4PKxKoKEoCUmEiAi017IQYL8T5UDgvled3YiD
qTVIo76EbdtEdGt+DJYNgcFj6fdzC7OIXp7vnUoBpIXiRcYj5sZjN4PD+8h9aj5v5Cv2E0UPqhX/
o7gcUN8XSvLtmd65woRAFcpHDE9ZS3HeJ8eULVpO30vuAMCueHqcGRxg19l9DAzNyL5sYcyRHgz1
M54ZLqlxYj1KUKItHoZNfzigmSo3g62OGWXXW67gIHjNgYRMITZkgepgqYHU4Ys9yvDGKpZJJtcA
NKwgrC14SlAohNX0TK6AEbGiSyXddqtaAjQEucbdh1IJT2oZ6UeEyT+T6yM7nKZkdic5wbix/AUc
UkRhInDbTlvU7Kl8kN+N44whJJkixf+7iArV+/8IgZq+17HbSrcNGVnP0un7X5OfP9ppUIbsknek
sYkiMKWZyeQtyVHoHNfeOXf3R/21AKmZlCacFXEurmfJQRX+EnHLAZtd/oV4qmpcfkYyj4KHC7FR
IdGigLso6nZrdDm0LqfkmCaEkMhuyVZNdiKA+qA5pB9s+e7aPtZzyom30HcJDGqDEgyppmLjEf44
Mq/pWAWevJXNvt8ySnlDwOfT3HbKbLrAOYGJHu0C1T7Pyg1En7U522Y22Nh5LWwth8grj9c2L0wf
tF2a7IFQJwenvV0UtdeBtNv2w5hKKDuSVTHsdV4uo5FTx8zbGEcfYHZFpKtjeijsV0tFuos8btJ4
5AJLXsFTFOSNkrnV5+WBBAByMN/AHRrrUa61FrlaX2vGH0uq6j82BZVrF0fvgmxlc2vcYiVNrmp6
j5kE5RZLqWiN4JUCUTQiuRsmSzZ7rOBhYzTcEmf/+pFWoKTFgIscZmOIITzEGrlkJq+Y74ExrNIk
5OyUP4ql/L0cPzq5Rtqh/vjplXXJM7+lNljw0jBRAFDQUFgasdHe+0IpAUODsv/z9F+vfU7uZavz
xOggEhE9sSPuYK+t5WZrEdq7Kfqc6v8xY4xD3VG/2oShFiN3ilmz2d2A7sKq2+jVF2+PVvrnW/vK
uN6Gdm5wcB71HeGAXyDAPe3JamEvkzp0OpFWY67uuw9XY3i9y1wc+aXWPRo13efhFIMYdhmhObc0
rLcQJJgkMyHKIUuz72pXT85Ulap8b6UQ1Ib52YbvkXQVjrLRt9bTrYW/+fB2/4eTwTZo+0f7gH0m
LDqhBl58weR5vJkyGwD2eOjutBptfm18P0iVJR2Ev1xtw4wPFPIdIKgcGEb50YzhvM1KN3/f7Uqx
//lOy9cQ+ljzefs2EZ7EMR6WrmJn9A21NLxzY3kbX5uU6SQypzTUFVoLrXvAAJpIfzks6fZfa/Sx
8ZUXbJ2UdI65LB8S02dhb9if8Z1BpZfh1q2oVpghi3lneAZjMszhsSt0zgSDbYd9RvL1MxC1cmIw
s2ZxkHSIVpl4l0Ebuz+Ya8Ns00KMnhRXDvpgDS8SI5TZ/q/tyGiMfPLrCLXbkSEmo645FrQqrAnE
+R/xEmUW1dkYJxuOZgu0RqQZORIy6MA5zHK0WOaZU/fqDoEPrIAGCJIKBg83MsCfp0UKYIo6F2bc
b55gIle7l23C9FssYeDD39J6TCFa2YEDXfDcevGiCe72tGJGUqnK/OU9qlix612BIJDbpHe5qiB9
fA4aK3XVZRt5KgDleDZTSotqwPBNqoeCa+8AjujmXUjYM/HEJLb/OXN2xtrKVGmBsRfY4x7xEpHX
EztOu/My5+hXrBLnT66G+79ScKwESJ1h+vbgzsVoLVZwRa9oMYnCTnQZi+5YZ5DRP8RBTJW7gOs+
kCb+MMgBHyLFdqow+EzehQWMW6vo6NhdNAtRcfhWQHqIpW+FDhIhebcTO25Bg43C7AN299vp2NPN
do7pQB79C6uWcAIEtDbGBAMOo7rvTzP3cEZj8vJ8TlyZpurQ2XCpaM8ZuQSWTEm2VOEoJ+uu5lvw
GJFkzba71Vx1ojy9a/C+he5AP0ePWaRwDjQQVC6vZStwM5wXswv1ueLiLAE5bwgOB3D8GiLn75e8
0Vn/V+zRmkV1T/UOLXGgCOfIfsqlhQX6vjNJw1qRgDZQ6ZzYY2llyLZpjZhFHsBp8Fms5wQUvvLT
OXxg/Mf/IetIFBV8/wA/hA6YLOck2YG1Ppqw+KMsJifH9X/NSKd5O+k4zrj/Md9DK+TkIEqixINu
KVR2w1VBf7zkYnwMqZK/5SUyGwuHMg2OgX/ibh4EoblTbdn2iVMBrsZ8IKLX3ttA20yPFIH3K16N
D7ZgjGAr2hntkT5yA11pagVhdQ7szMxsQiKQypc64tXgGUkr6aN0az3Nv2KTEEySoxJ8EFWdh3CV
I1G+e/PwvjZSb0/bRTkoHqaOPhWD65UCHG2K5EV8zYSSUsrufHox2qVHI+B0O5eDXyBcv4+l6fWz
O98vR20RVf2ZLmP2PShIQp0FzBUvSsg5ZH0IfFtmxZk/0yhTKI05KKjjLRq/kFdbtl2SwzBwfjZD
1OTSYOdLGf4pZKgFDwMIOuHn5nsvrw/7tVQpKKFDSkH4UsR8Eivys3t4t09uItreNKstF5KXrzuH
hapEVvKq1jd/uYZaSPNeW6PrJ1ptWj4DWN0i2uWJah81tGaRJzKOwcTJ1LmtqaZeQdMK/z/twsuV
NjQ/3HRZAaFAb3zJ9SUqXtAR3dIdvxHQkKqL0dQd/RaYhRYJZbKqBsrF80f07mYz6MaH10NjOnS+
sqm0COKVZBQPOyStNu3n9xmYz2n3YZmOqxH2KxhPis98snMbKSxoGnG4cYzRhp5PE/QJ97iyq6cX
vjsuI0MzTZ9qlKCdBLYf0UtsH/zVDEpPrONpM1dfHxD+qqcvTDVgzD0Oc0BUd/BEE4LMvPORZ/GO
kZ+mJJ1Lz9UnGKcHtg36vkgnTCXSqnz23i9tsg4/6HXJLhwPRW2/pw1XE2fuBCKYfOXDDFdZVscb
IVNt4NjtrLc7rRTvoIgecgUJNFEdLDDjGF3UWOpEnQZeRAVYV3zhZFH9JSzzbPLwEB24st4aeN6t
RTOc0nQspPF6ch1sFAuGleqOoljdLtWHn8vKtyhVYpW5W+Ow/COL3PA5carKxgPsVLIYQU67Cv+u
j2P06IcZLvf86wYFiNX0dZQqXg+gF1H3Bh3jY7USvUJY0Dh90XoF5UEqxK/TgH9Dmb4mI9x+qGHg
2Czmkt3L/bgMoH++U1xOUWDDR2hGMQbLoM5/6x2MAyD7J0cDEU3X8bfnqecoOwxcikf6EEwrLFLp
+aoGHw1SocvBZTlom1luZIL5LLlm85JX6x07kE8oyFiPrufx8GT3h2J5smSuUGxWVgrJpe3GpJBI
ewgzDwiJYZvIJYNmHvowKeKdSABZiqmmcaYuEtijkpXH+KCDQsglNkP1Orrjsh8BsORps7Jcfi2N
/wdyA84mnLjYDWCcCwyRoRsk/Jb6zfAlzLZjsMvAtRLf32238YIcG94aW5u2c6Me5dKWsJdn4X2n
LRyD92cEEuoPO5yFyMZfsxbCMSm4gIUrK0r9qt8oGdoDbodu+xSL3mkO0hb3T3DzzQjMs5ha63lQ
njp5ELeXEF40yKaqRj7ZpxK9NMsxZyv3kgB8p2Q1b3aRNb9W0seOWlv8qhpwPlXJCjTXd+Roo3sV
ykOggStfGPZvz7pSRJ3dCUMPW0RvjvUH7WCXEEMkSEqOGdcHVx7nODxtpZTFQer3No55YrktqpXy
g111/iHuuslGp4Mk/bcu47DBQYETl0cbY8jjXlAGp+4nN7O0nx1Fx7YMeSS3OYVqEWQl7E74U+Dl
lwr6RdtQG4BDkVj9jHocAVb+7Zkq8HZubVLrlKNVnVMK/GXyxEBbEGu6KwNaeiC3p8T1jva4NxFh
BupFsvYvipvAn9MZv9R9nlDjiW/kcHfK58trk/iPMXsgR/bu4iiut5DKEeVo1e+nvZ7DJzu/F/AR
NUzZoE+9mfSHBo4yPnA8FR9F8njHNGnEATmraJjgN5++U8Odg6A2PZZyqM+QznSBz/bU1Lls1WsD
aYdbR6U19znEPa936QJ8H6xcdZAvYLY+jEXhy0QoxVWR7vWTb9dOQLD26edBnkIVwq34YOQDZojG
ysFh6y19dFIgcqfC8vAtjSuMyNLn5FL7O2j/qDYEpqQelTD/jf6NY+HyqAjcrRJfydQpXaLswZD4
7yieS8v1Bdi5EOPGE0e45U1/xsBLMuSjWb1jVdIF9F5taymCizVLu6Rcc04EXi5ufXF8D4uKFMXT
0DitW6cAh5ot0PMy1mYJbn+NthQwLlCjzQSos39HMtoZNdePw9dWBxndnFwtnAkXnQyeC7RhkRTz
c8QrOH06YCVZOKOOVxc5y+6BhKoQsO/iuERtm+ItAvnz2H6HA3T7K6BLqn1MY1B+UiWaF2+kz+UV
6FLG+5qA8Ae6rPIvt9n9z3bloheUhvsiTEjlSlEr4XOMOYfqi1uwJVptWetMjuVXLz+WaIORnLkS
gL+fCSfzKGGKsqp3joXpDKwyJFlKdsYRTLzaY+rT39A4p4YU+UGnCNktCCbsMzzNe2KBtVFBmA8n
DZPgM5pBzju0raMlHhwZfrUSS+PEpj58kuQtRN7l40BwU19syzPkW6uqcNTIk26AfvO7r8bFZvGo
w54hj2tjrYPSiE+f60XOFeY5NFXtQpKSLe07fxlQtziJy72V38MmZWrUFNOZvpwJxnm5t+Bb1NTR
PxvpfuWCRKyM95KC3fAbbNASFVSiTydH5uyKKQI9nKMuZweGZOHhcE64e4Hys8SBovmQamEneru2
ALk77hNJ6UuHimjJ2dRwjiEMceeCkEy2zHgEef3giGlPaYMBVri4HZC0e+8uHl33w+YWdl3NaCLJ
arnHS26IEqYxICiWrGfgHDtYVOEf0bm1FWLls6Y0COUZacd8kN6y5neX6NNozVvIX8x8RkKy+Ylh
7fCg3TjGEfosBvuJ1V6gdgfGeoM6fPIVBFzNYwZD5r03FynvtbYIQ8HcedHk6yr4T3sYnML18OcO
hY5xes+UqBEZluw/GG3Ye46ChtcKN5jJZCrmdY7yTh7/IjGKtfkT9bp6cAKlVu1dqrMOsbcEQKq3
YkspS1omrAX3MBGvOXzribii9ToFRXO1oTBeo3Mb+x5hLCNFbXZwsBfrY5tA5ZQUyKi2boHYT/gC
9Ztdh/2SHxp7IdMAYfhasSj9IoBLznr6OROQkz7p7SgT67omtZBy9QPwH+70dbyTkvTjB2wvA/wo
KfEltD/J6ed1ORZzzhUPmPFMNNXKLd/OIr3dhQhl0x/Wkx8HgaDN6lLTHPkDIvqGvgD7agg9Ql/h
vXOwLHd24PgCr9hJt3RTgvwtGSBOlkorRH7CJIHKZTl/yAVbqSYtgmtL/0p+s9Po+loSP83TJ6kb
6HFcwlGSOgIcx3e9lfpw3gj7zqgT2zcUgPWZcebyazWsaWLCMuPTnaxrT3qpm06jbxJPdUf9Pvgc
I1RDekdLEWjfAeKE91C3Wwh/k9ZhqBqOH7ktblE69iGMJHTexazz9W/ikU140yk5BN/1Xbk8QA1s
0JJbxlogJmnd5ExZhJNipjGpkEO5EnA6qbR4MXiruTgfi1ytFyru0kDS8bfn7xITRtROzU/YpV2b
m+N/WqQUf0cPiO00/qwQtnvZOtsBZEgR3c/YQjXiYde4L0Qma97L+lal2DjUHZTX2Ys57doeWE4+
3zUWId5t0tuJQYfgbUxFmAAbCViOJwdhEn333SwZyxpppbojwSsiKa9vd5aIsZZ5uei62wtlZ/dW
y+AMXSOBICdNs6W93oPA1LP4AxogVoGUstFDSx+z0r8/frGA5A8dyqtkNJQ/hYpoG1bNH75XR7zn
k43GkpnqqDI1rs5RpOtJRgGUF3DXmtiwapRaXg+VhC0Y8ZaTGHoW7hhXiWKw/AjwsO1q+YcV4biY
xZD0VgBE/SeYjHH9OkitQbr/QzThpvM96Q2OvTLF/gZAUEbykze3Is2OSHyym0fNITB4Lxm9GruE
oHM0XsDkC1izylHE2/B5KtW1DYd7pcXiX1/0axsJWQH0m5PYjPRMw8IkWKg1Bf3uhEpN0LrPS5DI
PqEUvMWGC5CKaNonrIeGLbM7mrFR8rsqjqsiNDDo3zSsrPKlXoyV9G+ACjyVj0IEw8r46ifV03Ch
4xuVKxS/+NzrMgTAVdKWmNoKtlMY6qBNLyPT6rHZoeC0sn73ZuQeb1slkGH0XqaBR658oKO+4ahj
Za68cwbbtyjQhbTbCzJpjIy/Bl13nGhSBYmvkPl5ymglxyY1W2q0aCzKfSY+s5DHHk/I1rI0ol1y
P4H1Y+e+aJyp/k3y+09CZwcWmNm1kH9YW1r5zx31kXImixTrBZHeCdvozx75wgpFYqqZX3V2jkSR
3mdlQ8h2S5Bz9fFeOZUPJ0N27VsIKCyKeEv8CgFAS55HI93QD9bfc/ozpja0UEDVmjojxEhYqknF
tmN9l4i77DBKBgpdT6d68pjC2ePMyIt+uF45aWu3x+Ik199zsSI6GLkksmnUb3jzxK5rQZtwOpb8
YSA6ZgTlhidTHR807D81stG2MlZCcgnCWJ4jQRsFI5h3rHJZ/GFoI2KHxzn0G8PHM1TbHP0BhO0r
HCFhFXKpL54IHhXXLFxE5SxSFsVIGbfQqof6W1vqtOAWuc9mRsTwvVEU++LFRYelis19F/Go/Xna
ATl+HqQF626HIrjwUKLzB3+Sgi0rqt4OZoPPym6IIMSvic20iRq6GX66VTIewxWvIPoz9+oJ9GeU
hvL7vk0A5DLC9qk0SYBfYmoZV96r7efUl7vXza/WRD+W2s9gYuymYt+uv4FuRC5VijxR6R+Z3l+2
t7KKXnAiHUiZuXsADX9EvtNzDJBFlDXbXH4MaLbZFifWOUwWgwy8wlRmzvn1gXLQnxl9HkRCnRmy
SNwGa0kPfYDquAL7R+hibRpj/db5NqmYMvqEWF+sJAq0+SCF8xmaabSg+lTkTmq5iSS67EX1Fmdc
f5j1lDuIfPPD+UBq+ETZzGDe/tZiQVdIKnkFf5b5cfOA3kNXuMcKlyono2hC35RHaJBAvaG8/49I
hx+MexszzCs4P2nbySGJ1OOZupiS36fm92arF8Ie3njlmRmChmRt0TO9yAnjgZOf37QEaBduHmv9
KZ28ScYy39vUTy+q68eJbQ+E0mOBT38G0VcryypQJL4scpUJqRATnOZDuxj5+/7RuRfzd/b3XD98
N9rrmNxxIzir75PI4VP6Y+ACcPG1kD0CBNbNDP3+mjZdBiyjz9QjgGrM/d0WvViMnubzMhwKJnQI
+iSutWpe1FRMysnKjZ2lkD/tP7Nj1qeTGq9oh9dl7ynF6HhqlL2pH6Rpqj7lsVRdNyvvp/Jjcyl2
tIP4YvuucNJB3WWb8LK7qsnT/TfkbCK4ri9+eThGjk8fvA9cONG42ros/GcWCJ3hiiMa0REpeXYe
z32hiPwFXEG14ZCiHSbdI/UjkdiTh1WA2ArWMQfN3Ooa861OQxxlhO5+1RTwLZlad9e357tqxdP4
85KawIiXHSyyXE1s6RwVduw5Y/3ftZWJJI9aWjCTpwCyti8Isv3RMWLL9XsKay050e3ZBNfEgx9s
at/7La0Y+8Nwwytx9Ea+iO//orKBeOailz/5yTzHNG4SHmfcKBVwwWxQ5YE+oz0p2Emv8lUCEtKq
60mN02+XJctPIROYC1jVmliTTGKHZaCSI0fenvexFCgAQQyt/re37fqzQV2OIbT9g49WQzrsCUBv
w3huOg668kf1PA7/grU+xRigC4aW1v0yAeQL1Siqmkjq+neFUgJylTnGS17Y8z24DZH9w5EfyN2E
rRC/cQEKQeDJH4HJKcS+0l5JmCqbozUdDGIAFWDfuLL0dio4XE+PHE9dy8zfparZgsLw6NqOKT+I
a+5hkhaH2l8ItSS2CUn3Sv+NocqIL+LVHgDhIcnycNfgQGmO3CVC4g0OY22Z6bWHWrUKHhfaAaHj
F3EyiucDIYHNjWZ1fovCi3duSL369XG1hy6bdA0Sz1QE+XmUOwNDNna66oJzIhC/zG1AGwp02Qny
eUtiZHUjQw09VXIBHEtylpTccJx0ifgatF0GgNFH1Hg043ZNR03ROeFiAXPopNofHmc9Rl0qXLIc
85+vI++dM77R2+E14n7V9TxyImt0g6eKwYixzVR6rRBo+CTB30I+OeHkNpC5ROi5Qrgfw82vbVx0
eqg6q7OfbYKVT7fq+jts/oIbEHA++yPWF/nYExDiWw+2y2Mcr5xWH5Dwpe3Wne+XlVZiHU3H9uSW
P6bB1NGFFesCeNsjhFJYn2WSuA1bPBwpSjWvaOwQJCmIl5kmuvNVoNnT8PGKdkWpYz+T6bVixbTN
dAICgbf1QvCB9513fIQ1w2uZ/WuZ6Le1+zh32p3GqSKZz8kQMLSLoShVkGj0Guy9Om4P1uGrk/Pm
0br7KA4tvRaAVjdmsWsO72T+K39RPSwCdXe1RkSnhlSvpWcBRqnXivYWMD0xrZz2nvnq8oBDCb3S
cbZs0ygDiKHncxslAPpVREcDH+6nGiiPjZzYMOrgITevHJ4nYQwDL5xMG08cBBmo2LfKDWIsl1Pr
JLHRdgsULW/JoIcWsWsIsSQTh0LAdAGKRqBi/N5L8UWlrkrSZzoWFA/U903oVd7cEMsd8B1CReju
eWx0odxCRn0kq12+chXpnGJKyuldhzIvCsnxuEsZTizwuj2d2Z7NVwZSVAfO1c4CQHKglo1vGkQ8
zU/cColYswh4bDR59Ndwx8lqMd/bI+loBVk0pOA5xxebJ8ZxaesaYh3mqjCGYUl5HKUA1qcceORg
q4REJfgcsdN+RKcRSAhu56qAy1JOBX1hVf9m/Wno80rPT/tRY6JmtZLbMUT8TL9CTv0MhyVEEnwv
Ri/amBPUltJqeBgAUr08USb1Tx7pQIPapyTAdFyccR97BIU53cYQy8QPVkaU01IyjSGD7M8dVRFZ
jkW3Sa3MqMhS15wsWnkuh2QkuNsbCjX45gNADy/hJEbdv7ChgSjae27YMgcCs9YRINOMS7CtH//i
rosw0Rs0n5nR/VST2KmhKcQX7jISc8sPFOhLCgJF6LRu/S2fj6yhD6t6FrJLEriKG8CjndqSJGKH
lWoLDiUKBdepf4u0MCYOGl6XvEG2jk7MJihh5ivCawmfRhWXw32kXsynNL057aHfu1mT7dNVG82D
t1nk91eeufPb0ZnuaXX8MUxHZrEmwpR9abMypP1znH2VeXhS9aSxkAuH6Fk8TOmn20TXAmTPAXjU
VOqLUYYrIffADvcvGhFprbHM1pFADF5J1g351YfCJYE6CkpXe0x39Y5IFusY6hISYjbLaM/DXt4r
ktEPuk+OeWGGSVTDAYQzTZRmsEvwbfxKkcvhQtr1PQ7JbSxJHIBBSE82zejk0oieTFAdOFQqsKIe
2gyNxdFJBY10K180BNxnvC3XkuktUmuyHq85iJ2kzQS3440hH3V6SpDzsMYSHk91mwEDJuWF98rd
0yDEUcVPrASbFsuzasdgPtRTYLvOLcWhSOCduTuvndsZStXBC0n/EqwhloOAYttUsuoPb30Ab9MS
bCQo2+ZEuXgyRLhcHXFpoa7s/jCZInIy2vS+Fa2bKdnPQXXgWu7zi0qwhtG+ew9tWPsm0UqY0Ry3
M/f+s48t5fwLfcsookHXbuTGTXYEeJb6PKJrwNOzZZBLvPdzR9TEekthYgTNchPi8dM2yh8U3Edo
2ucvDvDGxV6At5FUXsrLoAe85uk9+4oRkyf7Kxi62RsdtxZQcPx/UN/6aEdjm1U/+nPfyYC6b0rA
g+VFBUsisjbK+X9Dzrzb+VbLxbRxGjcKVqAmqZE0dXywClGGF+5F8MsZQTYQHr4luUggHSUv5f9v
Dpg3gd2UCX4/Itw5S0em2cQMaK+jUqPn4V09D0bucVCYDv0dDkO1CEAyKyRgbRewSo+9/BBdp6HG
OZ1eQJil07AhHKMfl36DI36BZtCawgTsv8amA+aNvq+gfbdupHMpCp4cXFeKVS/2a8tZt2D34rvO
ixF+AAjNdPFuLDpH9GsNMqHDWzBp14sJtk0ljaw8p+XWD5oKUlRMk/jnuACffdBfOwzDiCAsFW8e
QvpO+UCGRTCDQ2Br63owR24tMWGDeYX67R2HPXKXfMK0cSO3xXLq/Etxz+82dC7EflhHK6kwKMiK
lV9/3Jta8W07doiU7N0+E5RBRtBi+vmWr5ef4oAzR/1RmuQZOIFnl5JxFL5EOfQwNeAr5Kut+KNk
0im2S6ldx3n1954ADqi84269XKRoRa9kJrt2JO0R2fWPx6LOZk9PQAOrF5def7wsZMMeMhQFv0Hr
QU57yvyWbJBjGP+OhXqHZLL1D/AzWw02Dp/yRxg4JBb7q3ZIQ7Odb9tgD22Zc0S5GLjXjlN0qBjh
dtMyYRGkUw2Whe4lWGdIKC3SWjzgxYnhr6kqF8tTEomc9U8V7k8zVsWTl+dkiNbxYSoob2w7B+5+
+yxmFsk8yWY8jS9OPgG5yJN+ZaZYI9jeQA0z0q0bkdubcdJJXoPkyi7V8M4gb9WqTaSpL/4WRZbl
8tX5f1e6JWsxLm8aqTeeyDX2xgpQ441LUnMEOCkocQy3K5WQmzC5skglBrea4Fjka5LjJS2cvch3
fCe3G9HqZ4dzoGora5v3QXJDvWYSm0SqOVYYPn5bnqqB31TGdHmWsFLrCN7gkdIC2zEhfl+5Hqgh
J+q+A/bAZB2x7pvnbcBmXqQbC1dcZoi1oNd5cPLDdDUzxtiTgu5vWQ22rQbezbaDbTp+0UasUcAr
G7GoKbBFd5xODxTXX3qOr/zkOYInkzkG9ykLlZX170hOH+ecm74rvSjEKuRJiPZ0L4UMzrN1NQVI
IhvHbmVMBTtonWru0H7F/3K3N/x3fwT4MJAtMvmKiL3l681iQxCoPc4gH8j9IFsmwRnQB6ctjob5
AtBtQ2OVxCdPT/28A4DFQihwtYJcc1HTN3f4dceeFNe+htOFXfaiiwKdh5pK5iBnKRqE9iQXtDBx
at9V1LC1EfjT/b5GS0yhEQL7id3cQBNxvYKKJBuXMjkzrhgiLN2JBxT/weby86oG4YoUlsxiN50F
8NZyK4xGD3pmULXf29EMG6uRRhkuLSZmQWsn8XINZiQykkXFWejBOVa6zZmzTcxG9qq+lD+xxDIM
4HSiyA6Lskm79gfQMqkFZXS87HkYnGQRANEqDjAQVOVQd4ehgfU9RDq1EwyiqmAmU14hwcc7Kzpv
nqevyqOvyXqhfmFv5Qmlq/HDSbpCjX9YEzKk6ORXSC0r87l91lJNoWCjz68y/pdvisnFq9qcbWC2
yb6MT1V1tjvsrhVZMg8sxlLH1+GaGsMn/B1D1fsCXcsUV5nTKHumK4OyKTCH4thhkFoxAgI0/nN1
w7snuyGWbfW0xvebglbXoCq/gXWPnzD+jUiR9DmIxk6wsAxzUCsnnqopXMfP2w0ToXRbLf+jcXzF
9f4/5E+/f/+KZGVq/IQp1qHotCF3NxL/IuVcqzNlR0NqNTZqo67x/5RS4x+AVzlYQhbax6d8CYQv
FWW0g8KTdci32j3Py0tkY4/LwRuQlXrfRhWqS1qytHRudoSuecTWYiKMwjRZGr0A9sHwgPPntqvQ
Betr4JHd3S8gtH38UeWXVXwZOegOS+p+6nrK5IInvVwCpYPohNZoqWHNL5wJLFxoKQoEOVq2tPka
+kgWRrsnppsyDP4tzyTc3x8Xlw+6XM8yJWifrKHI5p1cT0M+PHOX3MVeTO9yRCOKRsSzWral5jzp
QTBkCKEzlOxvAQBtljXzd5WKdau0r8NVZSzoRvK+1FYDwxbY8q73NC+T6iReaBZeDym62LmucGAu
U6p2RIcgJ0CCjZ2sB7IKAe99SRkCnqZEliSl5jdx3kzcHg4Q2GqaIg/X6qY8TbCyYAJQonCzNDrg
Nhh1ZQn7FoeTe6r05W2GDlxqqSLg4WflZ8ShSTN9RcUgDc9+sxVM/LiPhJbNYABxTsmP15elwrlu
ThP6GSEE61VXO6A5tOM/rRafn0t7Ip/9SZ4vkM9WuDS+iykZjPVQEVdTLqovgeqPTUSO9ueY2XjB
oIC5w8J8D3hhzLMMbVN8p/O9/E+CMsIOAf9TiDYdvEBUyYJlCqaE7T8HFScP1mZd0kAyzcQttILw
O8s/he8r0I2YDf1GfWVaMI3QzwOoBaWQEtqkcTd7/L9la9e8t3RX79sji6iU2L7aPTvwfUR1F8Od
hhkiR/mfyrBalViqs/fH6BPoSyHHEwaSUGvdciQmSN9ibTozVr8VjAFHRfi1A885SrcdHGWXGfXB
O4I9uWYAVtMbHJJnAXJ0Cl4c4oPTorAOWQepO62Tmk66FtIps+E41HTvVut/Qhj+FZlZfpEGRJtE
o+XqvzYySOzj1bFA/oOCkzYTJriWWZnwXih9+HB7Txk9R72phn3hcJv5JKy2G26AU4/AnC2vZfQu
MHoY5cISx+e0hkrHNk1l1DMAOKWROI9WLAjThgKMbu4uJz76bccozb27T6Vz19jt5PBOYaBjyshg
fL8bA0J9Why6fzhZAdrC/7nx4UWbtB+MIqPRQtsUIBc4UtCt55tlmPS/GC842mL4QlWqft4fwWme
brPGuCX0LL+iVKH7tJwlaR5P1mLFpMwG8SNL/G3OyAhuZKrjQuweNmhnIl3I1Wf0llWDeBFZk8bt
Ai0XGRvEXQW31MXFJ3E2Qhdnlfal+05CIRl0av51xM/RsrNZ3PDCvJxTPRlDhMSSIG7yYPV4uLcT
lUoesCscGpyPCAiBJK7MQ5LNKzwtb+zgQIFxQv464PKrwpDYFecXPSORnBjXsSSYmNx4mE4zn5Nl
Spvm7B70ZtKJ3Cfkfs+FcytU9BOBje3FaUWYSOY9la9RKOvm0nsChpNz9NavOXLQDxiKe0gUUBkP
bb/9OuBeVYW3U10sQAbPFGASc1B4HSmz9jGG15+KRkY6mPH6qnDKGsbjrk7THGAED1FBTVmxnm/5
/6wMi02H0ENUzlGyEwnRGbUcTr0tlC4LIeMZQfa6uBX/dgE4LlEo8bAjf6UhvxkoYoVnieV47YZx
Zmyce1Q4FS0Z5e7TlDFucycTYeYJB8eGkDApvAEyLWaJvesAugxuCyJMtCe8NYD+XnrkHLxfBBxE
FihQvKpFJJNoGr6SSEXzsYv48Vpqf6+O+eGTbs+Z3FSR9F3oOLpX/A4Wuj1a+x7L237M3x0y1yDu
Ncujikf5Akby1t4A0adZnXQW/yfIyxdoFgcn01gK7vXbA2Y/mSbRQNggrli3LL4+MDevAtB5y2Ln
IPF/4dY8zcV9v3PCI8giF47qfzVXzCc1S+kMc5c+oQ/7zOF6KyAgVBcAr7UIS0APyZ61nPxhX7pj
YOV4LgGZzKWnBIjckpdfSkBWX2O9+C104f17aC1Wg0ECRUzRqmo40VK2JNgoKuYGZ8WOEbhExRfT
4OajAaMKNNj3C8XezlNqgpbljvudmtINKcVv/uPqDRdhMWKtAgEiCQFLBIfohQJ+r2ky/2ScPqba
J8gTxeX9+Q+TBs7Goritpx8Q2akAlHDIIbfB3TGHeqA6RqRX4nSRapFCPZAIRdP45W1fG/uhxdsi
tIKfjOX0YyuPUBOQCNdo4eoFcdhpXKnA9sNCha2aSAf/ETg7XRaChyQ48Vu2Ly8L3TTJG60wEBSD
OrcTq3EMRkE3Sahj7n49MJvBCVO01RcBaOFBsqNspylksUNW5YSsUyjgSzGDMHaztPEu3UU50w/5
Ut13PbcdPHM1bdnGffOBtRL9MhT9eeJTm9OaGcyMFg++pbT2Yup4DE7b95SaiwyPMcjYnL1kxUsO
qSShGLBVuwPqNivYoBJ0aVs0VS02wg63oIeiWJ07D6kg7Xy/VW11f3vlJevUjCzYgbD5xwSt0UUf
mQ3c4yeSMmEwv1WjEKrlEpzynwuv5cVIi9V0JBZ6agxeKqMiEqrwCSBW300RDkwoD/Dvxpc2WchF
HZgwz52LNc2Op7iuhBU6qUrNIiH9R6rnbQVFsnn7tWJu5XK9RpkNk5aam59ie4ePUawU9GtNK5lQ
CCVn5WDZCfkWlwtaLBSw+hOtfhEHWRcWKcxR0b2YrpxOzpVLYI+eq0ZfytCnX9pbj5MjU1Vdpfsu
CN/3EXJhPUU/hEkuPgAviPYx3jjzNAu5qZ5d3JLvHbOrPpvN0ih9iVdwtQM5ZIJv9T3hffDXVr/h
kRsBWCPkRQWGlWZSTnwo2FZRUwbNrolgOUppX3jbCWSnBYx+QtYxbbMnEcMZZZV9N6kD7AW7zLmG
vyGo/VahpwmF2K9aP8cPcbvRyshfiCFbc8NKorLH2h5tVVdfOVujyHAIw8YWe6zJ1ceWweMHNCNZ
rS6KFnRE5QiXpEoPmuR4jvhdVh1ZyXp74Tojp66USb6xPLLh6GBc7pn1Ia3rDm2Crhg8TNkaBgBq
CPdicpJU7X0MnjZq9E2C3x7Lwc9aYqsPQYMmqF3Ekq/oRmqFMM8jYhP2rVjwLlqtH6aA1pMFpd6C
y1hGAFR0BsjyhCXWmJDgUgdC0Tgd240dZakF3C7tGFp5oGtCvVDe5X4nbunaZPomWkrM3BxuOub7
Gedvrhgz9IktuMIzp6UUILKqthQJfhtZo46yDev9tZrNzp1/1gr+8SHwzDKtexz5zHcPt5+3YPP0
QyuKQbRXPtIR/df23WpVMsoxgyKnnbLg+hVuTCHJ5jYdt47bWkOOtVe6MwCjETKXs5qM4gTe1pHH
4hkOt5SnhmE1a9Ge8m8DlGs5Twlg11CPaaYXry4XyaHkjLXY8B7RrqCcxh8tcY1FxRo6Ro5X+fhY
TZMBFd9H1n/NX/ksYu6BYY8/WTA1rPprPBTZogh56RoBc3vpb4hmr488kVf3RUVmSvHqTpugWBHB
lYkI5z5I9fhRLxy6kB9aQIcoc//KjXQJ3I+FPgW1JJXb8mt0e53MqUskPG0kTBvbjssbw3AT78xS
8S0xO9/ohGq4G0FGe8mxThOhQync+FbbM2yQzPs04+Nhdmj/QUeRva7uxFHO2AN6WLvWZ8SFm5sa
ZrvDYCJ1cCQwlfgq85ATmfo7g4N4VF9whFWjh7BifTShBjkhG5ehGDI9UBdtmHDg016CEZpM6eGV
qcPIEU1iwmI9xE5c02U2/L6u1sD9mbgOuHvpGhfWXmxMiP6DgosjfhOnu/cCvWI+ytOUIGIgoFtE
n0TWeJqzGs4Q9KLRRNgLcakY6fAn6tCKxflcO2ZIA0f31b8TUZankmu5CVK7fDu467It0W28cltG
N2IW/oI2ih+YrsmIVaZt76xSSSK75g3xv7WtwqZpqtEIKvvjUh/dOPqxpUZ7UEgMXP4LxVhVx7UG
Bg4j1zZyKhNDN0OAk7PhFzcz11AzIhDOVvs7V1PCH2hM1WX2XHVfKHuWX+lAppJ5dAANgLqfo8PJ
s7ps9RzLdjFLYVHwH4ZKTI3LXrmXgWh9Ku2gAi28gfb3/FjIai2/iQQm05avmxk63DJMXlJMl499
Dn3M3wQhPMMPDKphVWlIA1zryrMxP56K1NUX8dfnaW3vh+ZQg5ac5Q8jClAzPkNUkqq4HxVqhXQL
+9/v6Zi9Th3hT2qpncF+jwfSesn6yHt2AXQ3CuGhv3yiuaKzcwEM4+GbhLhahMuKlT/zP7B2LXoJ
ORqmWnFXGTbllPjN8tL69hV+IMKKUppt46i9KvF0kVyHmiFDOODwtvL71Cs9a20WBj4pFoDDdjZW
9tuL/x4IIGW7DcHLQ0kfilZA64m/7x60A3qF9Qu2PA3KXYpH17toHcHYYkevd0XE85W9nYSTUotd
tx3gyreCO6rRfGV13HLz+RKmu5WnUMOM+F6Q5eRN6jVdgbBsC0EKkgg4yHex7VU5ZiqwAEDKry3O
C9RyHBwwRZ2K2UJCxc3AlLgheTlJgex0ksofNOV4hX03RW9MMXHL/xIE0zjbbnmQ7op/hKic4BhJ
psIjeLqWuVJWd0viEJVUvKCw0hFmKyPAvMRfGr+uHJ50pdqCwduexodI93zlZeDCWoo8FtlipFLO
YGydj5nA4BwWYgsHlUaBFOeHZKms28nyoV5gRSJpqdsRtS5SQbvZKc0eMzzNfIN6Sx7KoPcOmwmE
92BN3zuJZQ5iiAcEW6uRf4ucBBdLipWa18hI6H4bi+dFIwmITSctfU0X9MymAqMg3p5g6B6lSJ8Q
/KcBA4nwn1aNbGjJ0Bi0iOr8awfug4iBW7dNSLe7vn/y7D6vHPhPA8Jru7WK5bpCC8OxlR0EsB3k
FFrTg8S2lh9AyeveOoxVe/+lBkHyFzcL8+SYb2LNoDGa3tLB8A20Bs3timv+iGN23ZQucXhHkgtx
NGJXuICskheQnZGOzcq3bA+4YNcNPyr9vbm1je8NGoofFNlPYxFuapxnFIzrNhdXOvERw9KXvEl0
PquWN04PLsfDQOyZ+J6OiGe8XgMXEBkxc2tOhvc1MO9xlZ9wdHHNZmLCv5T+iWGInXexvhpnzMzH
N/uJFVx9Rd2M4EYIiKwGqA12JFHmkknZmZBTHdLeubl5jh6bCMez1hlxg0awrsvPC2thFhi7+drb
RbTbFr74Lxxq2lejxiA1hqQvXuUAWGyzptk0SW5Q3tcQ4E6W2yglV26lBuDO4Ja56oZfbyjgOwDh
qHpu7cQaDN499ChbX9SjYv/wwZ0llJmleFqV8AariF/l9GqZZE0svgZpy55XnH0aIkw42z40W98b
Qj12gi+chXEw8ui/kRH8P19H8EouiDzF8vCSMsHCYhDpJ9raAtkyZMbuz5eO9MCektJiIjlmOjZp
6hrn+rAz33ZjkdQc/dLt3uEeT3lDcHdo1qwEuPiVZ9sUX2X4gh5pfrNwBnNIMoCBy/iV59RW2wwk
KcCZMEtmsDMF2OPTqSteTiNjj7/MOw2oqec6XJwycjWqIticzv5EMp2yFDBZVRahHJ6l4S06hGlW
zlAu1sgwoPGoECV1B3apzt/kYcj1K3/5wRNT8fQ6cIADppYseAm8N9B0BrAhRzCdRI4fPYS5vkoo
Vw1TM+NiO3zGBY29q5v3qoHBQqS9MFzRdhV6o+K9e5lTl60HANC5xJXGFjKhgt3cuJS6bNp0Py/c
QR1BKU0WMJ/Dg2n0lgOfob1538F40fv9NhX63GAsdc4FXvdjqJAPrKjG275k8//FwfwWwWg/r508
89QMqPeke3EjIipCf1ZveIsRZeIrOWljVlCB2D9AZhadCi56VIU7z/L/5g6JzH7qFLaqkAVTNLb9
xDJAqEJufwRaOyDNPuEAdefhqBSGrbUvftK8XsHCwRxE+OK5IMjpcl1bshViyhEA0BXxxM7EiPEL
dFJyasDWLkCup51YaH/Pe731vBVT94yB2UIfSXEQuAoRi/jMhY7n7E5ciYOIOFP2cSJI3nYzK9XC
YreWBX2GStlANrU/dX0lsiofzCxiepG5mOEp0BJ0Qdk5zTmx/lbXTiVjQjbYyIMJOey+B8538czo
rfQWSJE5wAjplBovXV8E3/enpU9X6bOPZUG7O6uPNY8OLKoGo8ZB3O+zlxVbC058LMTB9O0AfQCC
vdvG3OponxcU0Zv/sgSryxRYyjH3B0TAf2xbSZo6MFsrfeuZtk9wqBVqXzaAbJvSVgSUozy+rLwC
CFGehq1YaHvCOlJ5af5bF0/wOf03ObE4aAxt00leZVLwzGPsQ7CyfOQtYiNH55c0VsaB5kX0KdWM
VoEQzMgAHEAUXga2Ty86GoeZd/txGIwqZVT5oOVATDfLmQtz9q4NmiEp8NHSdtkVGEPq/fwEQkgC
XtqeKJy0cehN2yzkJP6P7etoOq+efWuK1msD9Ukw+v/i2r4MhQyvF7LCELWvoVYbS4mKZqHUxU7r
q9dgqehdm8ubZDoruuvsmqmfMeyZHia3JJdC8XyXZJNygZTvaMeVE6TnMm3RGM0TFsvq7Xol/Cv7
AbAqBSM/Ljpufq2Ja2Y2qgv1tuesLtLpV1iHdDM9HRRbvCorj8lIU6brxDp1Z31QuF2+XdysxOsC
DnNJHmTtwUoRIdMCfvtgI3CB5cp5eI0e6Rni35P2mya3otdSUodSWtmjwL2qBN4biStzD5s6DgPu
TTWAyt9f0/jzXfBu58petGng60tgf+FZMmg6RvI3AuBy/PP/6oXv+PZrTxpJD7xEyPPpfSPoP3uB
E/qWklVqujgZbfb9iOLcU5T9Y8xYvWlJfV0qxSAiv1/eOIEPU4tWy0MokjR+AoSbsrDGbayFLJDq
kqFOl3paW1CuVgRP684f9g+J7MWKtA3ShGnV8m752nchxzPkV1VMvDu/ODh6+sv/EJbVkVdUch+W
229Ro95H4vv/DI+4HZxCPOoqLPD+FOe9N07NLTEw7Xis9AlXGRN4HJo9PP5sNKFPcEMYIo7TC8r6
iRTmf0R8W99TUyOOhSTnDquGKZS57lBrXOP7aJ5DL2m9HsS3uv9SXaDdCn0fqCqnP/UpMJMOdhox
XxYgJmciC2FTq5K0NB/I4ZAB177OTadz0Iy0K2PqakU7M4afIE7bcm9sR9XO3z4WvfFYXxPC95aw
/eQCobbBj+6jOwEIUuvohRsjpIXRSnNmOLwI1q+rQCS3fxhS9G92KWXYFgA9Xf2+MBhsV0/UMdDp
cK2Ehr+HcvlsWjuDleEgVCyf4fBinJNHrL3Lyr12UKJv9S/4UkwTauFs3vB/ljqh8rcD4iQrJeen
46ExxAxBBjuj5ZwFBGyV76xCIX8zuS3dHPrh1CEm2VVi9CClI7lEy+gbYdjGBKg7pR0Bt137zqCy
3zm1aT7YPFyRvRl62OtI+767zPDOpjroGYpmiBpAfZTKkKowzleGh5unIvHIg0uT0zLdHeAAc68U
HiFUdAgUFhZsTKt7ymxRX3OTOyFavWap3PhmlaDOhLtVySjAh8n1MN6Nx16OkG4I/Sqj1ezcfuH8
noT7TTyb6JXD2FX2NjTyyjUY/mFSdIJuOjmNZnLMRbfu35FrZbkXfSUwm+Ubkwxhoqj1qDYgf8VY
tJNH2nZV++WzUk0rC/mLsVDNjsBQX6a2zNin2T9HyG5pdJ7PVEWRdcbiN64YzQPZmFsGPzh7rCvk
ZsKopxTRuTm1yzyOBxZbnCdnfoBcQRuNscbwIG6YMGVBH0Wyrig7fFL3smzPDa8ICTgYi5vcT4yf
Vw8NzYT9kdwk6nPlwUGES6c9r+cCRCnO01ylzAXPq27342YZq3unNzBmlC8KsaQDWn/tb3gM39nB
2dE0j9I4eZoInS3CU+le2DaaJth70d2QjqdP+h+WkPW1Ba27K31cZU1P5UmFg7n4kuuYZvXbd82k
8d8qtAOWn3c8hYQvp8pHtdwH5hKIFDeFoMjBk6S3MtEmQ6giiXaQl1fCgV1Cg41lvKYbrnKP/OsE
J8mgNVkUYihtganJzT/ueWBydqHEE7Hd/WdslQXRwqeEzf3sDyxJYBdJNuFhpjLW+NnbvtAw+4lV
K8UgkpLWLQDB84fpHV1VDjnnBtV9cTk/PrM7B7ZrrZsbHjdNyA4zP0K7HeWSTC0G/3uVO4dkoCDQ
imdjo1c7/CYQ6uqz0bzljOd+oqU/2zwrbOa74iRyUXifLommFgZNbG7nxeDjxEY7caf1kY1SFiNE
KKjyiys0tmTzqKMUTh47QWv4PBAj0+t+f82cFZcf+UFfNzXMhj2RykKOCr/mjAMeTwK+KV5CuJl0
O6CIXYhG9/abfwZZjp1kirji37LtY9klRtb1tyKymkOChxdzcjLe/wD5q+ry/ACcCsSo6NS8NUq9
43cK08WQPgB1tc+EP4gm1qtPVOcjzbZpGRt5Qhx9F0a6QWlsxIcX+gLkuuIftOp0mx5Ce2gCdj3W
Tn9vXOuXG+r9Bl1DnSq6lIj+z1fpOacLaMNYnNceFkuxyiTiODqMZN+kHRD4cd4noQ2y5dKqrwJe
Il0biflg4NqaamFCAnuPIuiD0GQIaEzIsGw/g355D+VsYkKv//oKUvL7buYegs4I/Pz8an0nxqOx
6N6NQpfeNF5TtN0IdE+5sVKxk1RzUIpi3BejQIGXo7Wros5YRqPa3u9rYZgcuVUt7cv8a74eJdY4
1J50xeckys7USH7NrtW82DDUr5IudVppQzvEm3SdM+pEBFWm1KZKA9BIZ6Xl/JkP5T6qGdoxkDES
Kh4IHBcHKjtrcE7Tv55umIywULyTekrzxnKDHnJlFNV4UMvdZp30/u27uM7rlzYE+ZmRxO/rxllO
i7SSpym12AZqb9ANzgqDowQOLakOZI6WFYmOT1A8nJLFoBguEvPnZsR1u+lI7wCA5P5swRzSex9e
pGlYDY3NjeB1nAmG7bdIYQfzECGSndry3usqm6dwLy11iI7dYNH0W0kwg65bA+WtB3LqvcCgRc4D
8ILRBARGZeOcCot1WRcTNaf9zWYdGSjyx24ONRZ+dChapzYA5UdEAd/rNwVXb1fnNWrtMGtKDCIG
MbzRcyDYSD6isX5/2V42CF3lFl0P9ZrhhcJnbe9DBuErqIuosQVC7XWCcwIWtJ0AV4vtLNBoVZM8
ztDm/OvfkFxhh+iK9c480KSUV6OvzNYecQr0448SM7PJrEJrfOo/IN0XoLiTCbwazmCXenUhaaym
kioM6ax8HrzqhwpJnv6MQ7NcclPhOZQaVBWobdSGI87jDaieOrbufI9NPbwTFfAXuF/lwLho2oZX
+97+/TQKOJ3p+jqKTFx6xf4hdmgLh8ElWVCKKAot5+9wu88vQYxipTdLvhPR/yIPim4iHGzlwpkg
S94EubKwx5nM4fxYHOApdbXeavmyU70zqpW7hWMdKT3qyVMWe0JSxdO4HqmLoxp+cdhqKn2ft1vK
NIVFZAqCmnaAeJqnVe90dTB3PF/Vh/0G+C1lo6wvICoAF1myoMmg/mNTOwkb3KVLK+OaiP7d9bg7
gMwVRW54ctbZ4/rN8oqNGhEaqgroF8zWg/yi+WbrJZzCGgFy4OLZSXYFxgLu0ZjspYcuEgqLgeSi
0xkV5bZkuoAAaVBrGNBgL47jna/57STO0KBUI5WJFYUFxziKK0mjT9Iup4LPl6ueI/5cgCCOHpMS
7sYh0DOmKKGYaLSwJek84bycnVdvgVIjVwqZflV0GyqOxIPLPEgCK6sccS6FYEwSY/CZHW+pUFh8
pOVnqkzWPFxS1EYd7LiZGU9JecHcKDJhIPYQwyPUBqyYZ29I13y3k348uxJaAWjvjpwg1zhJ+C19
iCYaAR4WB/AqHgCzjdNkzxBQr/SijC/dSBD5rqgOi4FvGOHBYOhjBi3wqeuoK13ZqveM1HfsOyIN
KOqG+KohW2hnJ2yb7ImGZasp1/8MKhsgVJRjnOeKBOWcomk5jRJOZh2E5OFSqEnztz08C5Tsm/Rt
P3yVD286avSzxHz6haIEk4Azn9xRPcqXRy+4HPoJpR9ULATv/eOyvCi8M16x2T8MJldh9p8LxFpZ
/mKj1Dau5HCgX0zbjDIIwZOYuoYhQ/4GiFhNaFo3EgVG4SjAmaB40j98+9DaY3a68OF87dfaSawJ
qcCJi0oe6JxGJ07PuuO6mUY1gFtl6nYfuTsLPLlRhBT7UuY21Jor7tCSFxf4p2IFpiEs9CjvD0H1
2KPhohGG1d96JFxSJCENRaWlaoItdhaHGeYsz2n/NZ6vXH1Xu/jh6lrt5Ach/1DTwwlx8/ecXSU/
k/FKKhalGep8+mDQdgqUdVhH4DM1p8jTSFC5FF/UcgvfvkuslgHzDQL5jizxUmlB4iDavfyOklSl
Q2WWDlWycBggEK/Y/fbC/VYoFtYCEp+9qNIzmOx1hAYUFgPI/2yXbm6Rwj40F85JXYfJfEtrk1wF
lz8S3cEAfVN2zKY6/I1oYu+R5/XLrxgY/1mzdhT0O73QZJgKquxYNiP79cDOey/PM/NqdVSWvKDW
IX2xfjypc6Y1WOftY/aODIH43gcOGmE42LKWTYLjHaWGashs0AfwJUtw4/b4IMSVUwEDtRxYDoWJ
Cse3BOidcev6bqzthwpq54mIJp4+i83lkzn2nkslk8KAkXinbJOXNpNquI83/RPS6EElosbSbXnH
H5ky7E9cnQoXbKn1xJolGm4fA7+IJUq8vOcOm0Zafm778fBFvSjoPZ/Nd7yZPvVocuA4yQoUMEgP
Qsof1LN2t9ieG5Hi8yELsdo00R5cZ02lsPeXwKnQaZ2bQ+852HneHP9kv+DNl7qC7Y+63cOB4htL
yZjLX5x7lGxCLTmAM+TgaHlquczKrQIsWrS/275FJ5l5tmMogBaoTj0+6480WfBhfDgE4x9LfOn+
C+D55BanueGYRjJ1VmWcMOIt602ZuNeN0SY6I2nJTFJiICQojFdGHzPkjJ5+TaSfbcOZ6/JThsLv
jXDVMpafAF5YmEWnbL50y3Co+AvLVEQEV6I5Jj2tWK98SOuDkg+7IbMV2MiHdcJZR6Fyzie04Xjv
+tIb3Xf8T8KhSaMNFERG2oueH7zXlzsZ6cfUGC7t/AHEkDfRMRdjvSqo6ry+nrvx2rAXhEt8KCTu
FLawKsmZo9fllEzUxN02DjV3xlDds/vH6DShmB53i/319ICyjvNX4vAs9z5zW0uFMl7mwE/9n2iI
oC2hqqR3TsUS/3YHh9JQIVgF3hTemYT4xnPxIEXonv1CD67lxjRVFoWb/I6BXr374nrQTyzIcVcg
R9V/QVKqzE4Gqj9m6pJuwSJXqBAyqAQiU4spwTxphsZ+jWZ1pBthbSda62rfeeYelb+vhuNGz4lJ
EdMJDhDEBOwM4NlmoGfozYO8MSYtvxwwhcayh6wbOB9ANAn5q/Y6SBO9XPHWMArzv+6wP1+MlElB
ENdzm5TIoyqkTBdZ68RHe1zIqxfI00Ip2vKFdF4GnZI3ihI+AvOd7Atn/xqw7xrMT6PIqO0C1D33
ZqVPQmFAzYsnDLkgFJ/HhMZLOIswou1MWhpXbDP5xd+5DTkGnC9I/86m92HiBLuVIGe/4L483jyT
82ryKcI+4hn2922O7mGLEgNvYxbU1+kxuirWmrAxv6jjasuUj9h/sYf+o3cGXgPl2ZeKNqR3CdOW
EH7NPXejcjobo0I6K3ARSyQ5Kx3v1XHvauPCrCqmishGXA6BNWhmFGELZts+18oQ5cDSqrw2GBbJ
bY7yaDmmCJjiLBcXxh7tLHzTSB+Z3jf7Orcl9KM6QMzx/z+eGl7dd4hfb6sBNEyYbb3GYoLd3YJ2
xX0eZ5p0lJC4JkCD6M1t51gSdab2KVwTqjrlo6JGLoIu3WueIUanLIjPl6QUlci0aeG0Hyqa84sE
qhMdqwxeV+TF5T7XI63omDUhHydyNd3Oc4CrzPPBrkP/rtqDspAk7NScnw+y0DaQ03pcgVgWETOZ
9+ZNvA/FieD8IqLNBefWTmqlBqTdWxJ35mmGGDMZSfTUoI5bVBhNy0uAOBkQqJWlzC5tbLmAD3Yq
wBmiz9xmGiTu9UC2evGRT8XRJOufwmI4KM9qMCZyNT9Ho3tn9CObwvocoqAmamPbOXjtK4ow002y
XXhnBrbBT0egYeJ2zhrksH4BfMIXRabunPYtBgga3uW/FCp/e8vKjxlNSdtYwtUnYocuEQwVQrC2
6+sg+MyLrRjPDMBpdUlJng9rkj/uTEiypZSTQ5wfUUUVsw5Gd9KV465MoIupYQI9dQQ08ym0IfdT
UffHCpfmmNRQFu5KTwSX3/AAszk5N+1l2OcSjPcPwS5t/gXXr4x0ANlydtjl6qxMJm0BdAXZl22r
B31LmVKYMm5bgY8WNpDsnxN1NzpeiKn+YmHjK5Dzi9/ljKi3IaK34yTxJ7entSEiyrL1ugLP2zR7
z1GLfJYw1wv5pbWBy5SACLcVO/tq+5sgHBwL7si7k8JQza+JX5FVst3h4WBRInpKu5N3rK22gt3s
giUc8cX8bmJPtlmjN8NF4Ay2E1Hw5il9BFQ8Yvo33kU5PsKWEuwT28OP56QvvJIZcUPR6oSjBmqS
XPF9//5DX2JhRP1gYiyrIWQutcHV6ez+QJL1q1wxt+IP4PRP1EbwQXEoNitxE52tixflRl1fejA1
VeWbPz9FH+axhnJqDzm8duhllO3jg7Tge99CvAd1fNelJdpYkTuLYFesAL0WeWxKfuJTsKRUuXEh
uF8UUjrNlcJ7PazXlib8gwd7EKdztFLB8a+vZMva7e2KGPYXZ4zzM3PjVPXKljRUVblF22PHa0uT
L6UkXwKFVcIDDZHWIHYvMSFE75UTLCGxySBijZfTpJdK07STRqVFCHfhQazuVF5Yuv82gaCdgmip
OfISX3kiwN7NKpMUiYy12jhLxiLL6ZXWGGril6DVV9ZevyGgPuxzsWSZFTysFxqup4ynBS6NFQOG
fSRIs2YyqGvYJfe4sWJKQ/We1zLgn661GayrDMKdDec/lnV9LRaEOwRhl0b3ygxE2LpzzLFUh5d0
I3Z+AeIrgtTBD5fvYkCHRn/ix1RzsdAFo31PC8m6jtMTUvHEczfoFpChp2H1Q+cIcng5i6ra/7m6
gHWnFrwujqltANATv9eQZplqPJHPt5qTRLUprOH6dh6bs3OaKETUuUnxgUlnhSoUQbQt10G4Qe0K
tqhSwqYUVKy8U+XfLngKFeQMqVwO1mrfPu0HEkETt2PFZMc7pHVRon4oewzzeMMPd6KYUG6RByP8
Xtp+JpmqBZ3UIspAcPzP/02RXR/WWvoR/ALMWqr/eAildJUyo0s6AouuteaHLkDphTm8BZ9EzR0L
w6CuhcJ16ND4a+/BLIr+GKw1T1w4kv1sh1QJoCFFg0RgLQ65fnd/qzyoxMA/KWMhHzieWxE8mDZ+
pqaGc2YB/Z2icy/SWVbdRsqy+gP4paMChoRRguvXvntL76NLxam2YF9GgQU6Be4FkoDJKVjtMtuo
c61BceM8n3Gl+7OZM7+GNBKZvEMtTbrJu8A4KeLpORyjd4xDgN1wM1SkNM4aHtKqIVXyk3IeRzz/
UrCg3UKahYu4Lr29AHpYX5BFEXJJfmFr6d/s/bUPka3iKtjGXBcGVj+2BcM3Sp2gTcrMfiSZGPkN
aSZPXS4jhQdT21LZeOr83TvuFfTzAz1s4OHqeS8xRQntnCrkhnggkZJsWW3BiMrP8jcjrkLWQVF1
VgthtwMeBW8XWeromakZy7iBhEZb8t+E9XzK3andsPSWhGI7QKQKPKzCSc5JhEpvK6xe+dDT7Egg
Wa1wRu8UFRWsdy5h4DdDkq9Xxklljcla2YPDnh+WW1KOC0CiiD4QDTB/dp2d05t7WTNwQS0xg6Tp
Hs2MJpB7tvzO4Co4Wk4xKcXchQqu++MGREg6Dcl1si7+aLuJe+IrvClfD5vjO3RSEmC5hUK4MBe/
mnvRUD1/cXjiz4Q9osc6336hObxYbPwVyrzxFZ5exWY/9SBhbfVU6/O+Bvn4L/6ZcSCj4R/AONkO
BuGNkY5k+zghhavwRdy7i4E1eM4Yv1LTPtfZbt5uQRaUAgO//eeLbbCNIRtFOaVtfTCHp7uQOJBI
bhqEKcCWdo7Wyd6zwCIOzUMRCBKIAYKQf8D/TN0f0i7PE5lI4+VhBPNz2ThdlkMHGFrosZxEz2wX
7UbIbmNHF95gda7QvmGFOFEq+lcCIkLRszKj5nfymMOxKTAPNOB4tqfWTSW1u8P9FirEmqyKQLfA
9N/u/2T/UIfupB4NyH1ZgpmC6/lWuaLT1bI9m/osB19/OA3Y97DLYz8wO7AHYbB63CserW4JtoAW
d5HeCeZ/YlfifGb+Kh2hIZ2Ry8WYZ9Uy+blZiykI3UCqyy/ZOgjwwz/ra3xtUD/wZtSukxGG7b35
hi8iivn83cAPDZnWjLaLK03bKqYPwMspZX4rCUhoZIjunu02n3q/MrBXhXydE662mA6rVuFLGWNZ
SJkqvI2ABjyWZOeSSxWU/MSh3zAKhwngaYxMVCMnJUg6Es6zojpzjUiRSGnzmXyCe1YD95Ws3WGv
wdGjlRt2yrw/OmABZVVE3pA6fUSgaj8obWT8M/5mDwYFK5qoUgCsK1rF/AjX40InEJGhrV743tWz
b0Jb8fJCcFU8JSLgrBlIdKYOx4b8o2B8j0uZwk+Ay4F5o+6EKdCJLIDs+EbA0kSO6KGRBmLx2uUd
wgTfmr13Hc4swfiGKmfZqCie8DkkkWI5FLZjQ3hr+g6YbOFfgU/D4WgXoikI1LU5YXpNaO7dniaY
ZD5UQAbxMrQeCUuZCO32EMRzf9H4i1gFs+F1I3nbAwQ1zD9JQhx0wrF0lzUV/BxZKa/k/rCG2kLK
A2Ug+qZBbTiiFdsKtMXFJhsjPFMRJGBYGgHba22zigMQ9bWs1c53svXQQ9ZEJyhH7Ih+FL6294wx
yXeHgdQZF/snD8BWB8BbHIGorIZU9iuKp9Qabelt3GQ4QGs2QI4HIszEzQcug+ZRqjLhRNefOSJk
MWAJRGFtVXH31VENKjCUT4aRtgU6WlxMPQZA3uCfYXbFS1W9WiQz+S56xtXv5Ds2Y9sQqiH+9gSL
YybmHkL0JE2d/xX5gzpr7CDwPorc1ZK3ewloNLsdxFzpXsZesVrNeiztxHV49LXCi93DGocR69Wi
mabnia6Kw5RqPZX2cxlKIzTE34F1GCfUREO5tuPtxpc4rS/w6JZEOziOtu8iIMASLwP6sQeTnRYI
P2NW2s0wHlA20GSzkxG/mjHY2xSYAs1qbV3eOh0cyd7nCvIF+bRBfWNepUIy5pI73mMamHsw9eM3
1e/lwjm3vQy2ms2HsNSZAmBdAcvyI66+PTVUsb9w9jJjCD2N2FxAI94el6yMmRZT3uatHte/VHU6
4rhmP31Zmh1TtK+vw5moaZt3BjssN5tJxOkCMSJV1RPDWsL/1lFkPxpvPkCfk9MjRvfAgAmRl9Hc
OpzMbM1trhZbbdaJ3Di2kNxoQWbYjyzHqEoGDGw7B8bydXIbmE42N1uyatSfoJTAmVF3iycQtEnG
LiVT6kxrGVbLaDq2dxBnvzbPYI4act64avdOiNECdEV7ZmT2By3Rq3QTkX9v+F3U1J+38ThZ9w8n
9DyHu9KDKZSFpGNG8gyl38WCJY1iFLh4BADcF/yXEL0zsceErnoEQeaNKZCAY1qiXS95giwqv+jV
3W/MZCSq69MvGL6ULrllvDCHcUnWKsJuP3/9xLdOrdhTRvvLwF8ewV4gun1eflePN5Zo964UtGhy
sWsjxefQggFSUReaZg3tTNzlkQlWbV+8BYEw72+ta7+Y6f8GBjh45eyUm2vLZUQme8npwX/+JVKv
P0nwmpE6kYtcn/5Ec/oQBZBdlHUb0o4qPccIh+SQzMbo2uPy8DHXHVVLajRA/TjnckgM0Rurcp+y
Lc9Fuwt6g9GiLm8nGEirI6ZK1vApsfOyjSgA9V/b4eF46VfCX5jmK/udWGTQIxwJ7gf3ySMubR91
77mMCYoUKMUDqZ8D7M3BkyBwsSnJkmKFfX1Jo2+PGJIy3MoAKBJi0uJhljPvDTfvqETh04HLrzji
dDNr15axFaSU+BB76LaJtQnm70xAljXtDes3eiVz/jgMWENPoPIi8TkTBj+JeYao+WI8uALwAh1S
sVTmGf+mo0Q0aXeKH2rCHRdIF4P4/6hBBVb4XKsINDMzLqMydQlzMyRWU3Mm27QG1hxUfiGu8EFk
gefDIsdM64o1DxoZlAzdIDWfvhRd9/CCdsrz1OjE9x1jVnjeyWAZO3FHASRXEbfb7n6CwndXYRsY
lloUXTEm4+YxW+g+fOKK+Kl7RhEgWTW0pQ5u/UtpQsWibWgyCAl3CYQ2EdefHZ+PtzsWAgjCL6Ef
Hp/FjUURqwVxGgiFr6YHdNyqRMFT/2VNy17fwwdNydodPz/ZwuxYkzadqmrqJZze6RK0bC6iJDC+
EqovJ6sSHRBxFnMapKywPnKMgb9XPLaw0gK3HgVNNk6urblfa/I0TOHnNoJp9UW93rsh2TE590eU
nQpQTSLtcfhO/y2wED70ZbqJYstNDKX/XnpIj4QOFZf7Vz9uZMCyA/74DwUOK+OFgwLEbQ0sw25N
BkRWaa4/pfU4vJpPR3WEfD09tVzTfKXjLAsZGL8qZlMW8loF+xHymqvkXiy5NnMo0bTNC2/oLBj/
pOScyBsbouAHmnS4BIKGieTPQYtOn1HJMOBL6KrVnLDGKbxl6uavaLN/KWS45ehQ/bT215ANopF5
Qi1b5sWNImFxfBUSrBopxTLyfUEUC2XZ+NZZKG9sho6vA2Hhqeej/B6c8FhKgICmmqzW9w0l070l
KJaXxwGMCbz6QE69bowgh3i/HqHTKVWGGl/IbXMiBCZulZrjyP5sXPGC1FKk4SxS56rkYB7LgTil
RONVNHfk2Uvy0k7CvvMtNib8FrjNbaY+NBYTJ5tT3dW0JCrNVK1mV0MJRWAwTyKkqqn1VG4OvFOo
mqx+ZZWPscQziEUVBDd75IMLb4XCV35CtMlRVrWlo+EoXO4cdseBvdBNMuBZdMgooT3uyMM230yk
23K3syXz6sDt5eARfUL1ZUi8M9xzUUSg1y6N0CV9cZCs7EI6R1IhPW7WConeEC23/amRnCWdoI9j
geOl8Iz79K6cttzVI0X8kGICFf5Yj/i+ndogYuxSB8u/rWpnUc7eUSmzqVt2y8pCI7LI5ZBVXt/f
nHBIp1wcM+myK0XiPYvPALZqupdb7q65/gQeAFdlbhALVE2kziG/cyr+nAtI5s3qenoLrqGswfhM
uXkCtt7MYiA4bLTYX51VTFQ7Mf5RFUKe2j4vo2ZYGqCz0CT0VsZMA7BULKguwlFi13IKwRyqE1Jt
slWEysuSaU4TKFTyuGwYIM+zs7ljLovpj0dAYtyHcjLxmB33vlUcd/YHBI6xCT4DtYlGpHlmccC+
US3ly/tOka6n/qij4T6TJSBHqyHqIgiTCKr+NsHdA1UaqsWT8XvDLJKwC9+OlLbwcvP5ME3Y/97v
w1puzIpl4v+LsUJeHaLvDxvpMXd5PuhJKPkGvy8EZbiMGbZ9a7KvQpuStmTiq2F/aBJzj6tnT6Dv
M4/otydwfEM4hSzylmi1Us9xihruKvdK/w4UelwmvwCD6SHJ9wlCJ0ZKa2/RdxugTdP4s1eHdmh2
BLVLCDLXAXzBqy/JkjJ8BMtyaDrECpHNy1ZK8wOWXeFgU2aDXzj6gP6QtnRJan8LogPUpZ4kQGiM
7LQdHIiwEjmwnWWmnAoqSDSz18FN6+uS2z0Cfz12ijVEp56eEnKuEgh2+l2gacr9JEmJFPjhIr74
XDH0VsMWodN6CDGrkFyWH2zur/vLsT3diZ0VsLe1sSjT/4hHNepeiCeM55phm9lPQAicfVpvhsGd
cvTC797haxwavKz06wGUtvicQnZ7AKadMbU3Bu0FH4NU1slAAtjK0y7ogIBvsEpycCpZxuacqxmd
7gadmltYErmw1A+I5fixl5ibssoGJYaUHQp5g/cw1Y+Mte/cRHPonLGPFcRQ3M3sDSZKpRNuLeYl
iXRkgbSFc0T1HMcW6pwLg1xS9H9z1XFZ0VCG2dhiOEsEXoXbytnID2HVlLk4lwryPHu/S5hN35GI
Bp2hJRVUPba2h8w9Aefjn2EcjOqcAn7vhWCGvqv12ez9AuGKj4MAASmbDEY7Z/mzj3stbc2DuxcH
ivqLaU9U9u8yl3QFQ1g5rBr8YjCeJxz/oZ8wJxDPy1qLkIwxn/PTjB9TeSgQzB5msAuNtfDkmXHZ
bJ2ixmRjyYBwiaBMqsSm2ho1x+k8i26ND4aGa4Boa6YUyoougy+2aEr6bmIS1/X9ZC4g9hqg9aXq
J3TLd/k+uKHTsKtOY7o5pilJC+kZf/qxArw8J6VG+Ipn9Koelqrq0/KCXdyJdBOLC37FZiV9q0cM
CYwSMI/kmA53G/B/9dct1d5ZxGet0Wsu22DuiXKvRkfmAbAXjZ21L4XmzYX1RntVAy9emQqRkp+B
yGiQXTMU8NGCeh4vdYNxjT+7/9tJf0+OMLooCW4cYhDFBRzdM6oJv4xec3VdYz3I1utKc+sF17xM
T/fQLKzIdyYmqxfXbEFLT9J5zz/z4nkl7xP5+tDIRF18BpssSRMflQBAGLttLklR0JwsvI2eHOip
r3uBp9wGkyr65DDHz7njEEe5lbJJiu3M0U/P3tPcJZ7Ht9vnFnPd6qDY7Lz5dbR53K9BEnYXCITn
bJJS9sPLDk6lDRezZ43iqlziG1sFUAXR++ZrhLqZfY7AxIXYrTREPeHqPhLI4peISG5vZZ+VYRQQ
pnzgrEENrCmBrWrre/JzLRTGKkNXIi0W8vcpUhgy4kmJPMOYxAq5nVrC+gvWYpBesDzOM2ZJFJqL
Q9P723G3tsBXyNQ9BQmFsGxYs4W9L351VFKT49Nu24VmfsSU2ikV9Vtm7XEvcOaej21gqBd2DFho
t+XhjWbMOJ4TgV+AHdIjoVItirnufhrdR+qUEHdL1qpxX5dWOsEcBp1qOFUr7ieI0lTXRkY50t97
suEHUTVqGNeQ4faF9s2rgyhJCEcOEDBXM8DC/4rnUaaJPyBvXwmGld/5nPDHqUuxlpO9gIhGh6L9
OgXxUq4TAdxKy/wW49yOO58ThirnTPpE9KjVjSrhvHE5+OLm0ogz3/SmCZXrr/aKLr6x1vrCtded
ArUipHM77j5IkpVYaLQAZ6teGkhupum87ONW72owLo+NvEr31MF0TgN/f6L3p2o/FA2n7vLK/YjK
CzNvxqfbYQs/rVEt6AOxc3Z0loQ/OPQXm36Pvxp9AjzcyyqYB0cnqXxceTWFnp5krzBIbBBlbbgk
ku/fhuPwJL9SLPWQL8S+SCDRIvHevj6BUB5FGix+17+xi9dG4JH2MWCGd1kK5UwrkmUgk4aIE7AA
GvfQ2vjzboWLYHZufms250wKmUmuQBSJrPOUWNF7HDOhNB7W5xLjFfyA4dXFGh+zBm7iBTiCy0cW
DT2DCBogIOKJgseZ+HRrPH+IOSaTpcEk3wyNDPOyBxOCGnqquGWYgQLSzIz76+nvf0m5K3yhkdGh
Y5wLXaC3rxZZWgrwauaapwWjomZp7EFQT5AM7Owl5cLJQPHudXoNUpfU0d/rtQFsXuPwIpF/jFlK
l3Rx+HNiQuang3jjcvrVFAb69689yZ5Y10yMtcCvEGLFQ6NEumWL8bCb2/nNKrVvwWA9fqldSyeq
0v6sG4CEFc/Zs309269jkxq4thc24b7vUFHgSGX8ggRc3B7WMzL5vC2iXO7oXIQk0b8WJ64qxbFc
tD/dh3OreZRM9dQG5krExUwBZX26KCOGF9ONwQF4ssjXSWc92i17tXnScT3D6Gbt+uM0buBJzvjp
HtXvlyMTT3rukXS0Z1nEcB+WJ6fdOZ6sO2PQ9z8AzN1SLIzFEWrqPoBrMEetnIvrodo4SgbTad8w
QhRgqdNIizI3UOuttslXSr4SltO4/WC5XW/eQFHfnSdQA+U5BAnOUMJbI6dP2rn0BuZnhYKvUlNn
RgfIFTbn354m8bOSNc9c8PaJ+955sj5BxZBZDIiGxKoC+leAIisZ4jPPW7uDG/pzIFC9a/VjSw2k
qjYRIT0dTncI7KRAGlAOWQHpM3Y8n4pI86XJh8ERnISrgbLtAuwBMGv+nBs0z07NTCHHZtlUF9kv
HiQ7LZt4SWxnBmiVaiC3/uGpxEEkkVmrag4c5QL5V9PwoUo6kuXYUbkyFeA4mK6ks8+ea3CgOjTb
aABAsBURYMiMXJAZUZa8h7OAzyoSXPx/szfbB2AanI+VLud0wbKy7ya+Wfm0VDN3BqXAYzcSCZwr
5L3GPIKhYoS3HjQjK8C/m/H9q9l8i09tcYIgag4n/vUbisjXo/Sfc82p0pgSNw4o6ee0cRlo7kKL
Pmq5vTFR3m8O9IM21JrY6qSbpdTp5aJAAq5ZZY5KH/S6kQkcW6EUdYmE0OjMfarYh7FQgUNtqUNX
rNxc3r46k691IXrA+rMUkECXtRjlYu8U7xiWx2oVimtszzXGEle//488BveD/l8TKcIDHuZnhEEc
wU4BswD2bRJiMRWJIU6pv5k5WYsZH9sPmPEANIjDedA5/Ex4QP9/GDlQwe6aUids2CMPUEhuZAzR
rLmEN8NZ8NdjeyudazQY0TW0ZuIuAmvv50C1baP4j5wnbc6Tg9TYtTg7WeJe1RJlZ+xwvhDOiy2o
ioMNxgoVSA4tHeezX0VCqBw2JwIm+BaNGSR4xONehZvUW9NMh82xcrvbpM/kjMwSyWWvfCx4VyZG
0Y/OvcbWN7pgRZGm5FSzYkmv1fZ0WcSUTLctVNKqwv+1ECV8ymGJ4rJ744vEt/OsoD2o1XHdhyle
OpRfG3Up3ckGne3d7jClS3SpyGbjuCIpy2ndxt6/qATbQE6UyE8XdIfBWdVOuJhBvB6dtrzvx/Pa
lnzoeZ5w4Dd7jTTX/jSldoa5LP3Vs+u7OnsaEroJiN4vIjTwGOdiaipgE0AttZpGy+GTNqaCZVYK
ZAB4xH37O8mGpoA4cMwzBiRKuwyZJAxME7m3uv6uK2n6rmstBnXdMZR4F4haxtg4rMby4ERHyfdp
54VLoanu5Se/T+puWXKLctmM7BsOQJDFtOxT8v+vvziwoOhwqdjLYUka5YMLUmlsDV8Vd7sk9t64
DziEpnyjQkVAgE9Mzeep206D/pOPmD2foDVKYSf3hQRUFESbtzhzxbBbuF5qY3FsovAd8GMmbQoO
ew7loJv5cV4Z1EL9RDYLwcKllOwuveLB+yyxHdRYUDaRt3BGC2L5cG1gWRKhsDlzavOi9JuovKdg
TEXdZw6lcsqbRgJ3jTLzobYppMP+mRMUlcEri6B6taHipOXjulMtu2RV3jxLPb3SAECH/ww8y+KF
qhGrntkEIyINo1Q1a3gw+LTl93YqTf6Ow8Y0tbpoAsSH7l2LNPkLHtVdUMJuH+qNpkidRrOrD68G
gN1AG9jNHlMPkLJLnZoo35bb0oyItfml2ABPbPnNSatDRyvy78qWyECEWNfVugY6xgRFNYYPCl+9
QWu0BtVPoHu12fuZFbDYqu9/rAXBDFduVHedX4Mf5MU+JXZTBSKlSkNsW7IN5DsJ83sJht9yhpmD
qcWZ3PYHcOzEwrHf3eV7s5Y/j++jIWdWy0bI7JLIcXamcMaXrBbHP1VCPZ+87eIY84WUph9ffoOr
pkCw0dQPj72GZ1d7yAsfgli1E8iScND4UxgY5Mg9iy2dMe7a9ksGP8trWrYavl77m5aFc0aUFOzK
6rXTETbI3TqCzqntFEOEJOmV+F6OJgaSxib4O5s1GUKtd9TNtFSsnPgXzrlxgtPUYlq7sLJs2zgl
341UgpVoxMXmleXpLI7I5xCtqz8ddxbN4qzNqOC+wCx8r3jckLvAicsNMZfXL7uYMXP8gJFvHZ++
4KWOQbQpmMayLefhwkmjM75fthVf6GmYBLNvS7wZYgcYHw0BLxV7mwqLG5PVZpgFWMq2Y2g/+y2Q
bCcEjwGAoZ9w7njIY3fAsmNl00c9p01JdxMOgzV0YHDpGaOFp3eppYvXxZW1wje2XAas0FiAzAaH
draylb0EVRq6Af3fPvimmaJJ/O3SyfP3a9wCYCP3nnymDJDfLhf4W/WpeQ0fL0R5RXW0aJzKWy5D
xO1QgR5rbp1Cqcm+pFq5Yd8aUg0U5vqHGLhgyb7iYsWjSVvZjyLftxpEIssrH4e7vzID6LqJ7jIe
Lg4PoDg55v/E0ABmmzH3vxqHPhrwU6dSWnIXSPnjZxgo9EHAPeTozucREJ/TagfyetUbZwECoDUM
GKJFIKYqf8uLJw3MbYLSThpMpQs9w75RCc0J87h6lY5FTSVw1KeEF5RZ8oo8WuxFgvQQ+gbaT7cT
yCVm7yFcl2g5bNPt/VfM0cQhbMPCmmWLmI6XX8moLhDS2a+2mY5HMk0bll+tXXa7YrB13UWSTOpG
O+PsRq0ne8rAjmTPYmyEYwWQvjai17ZwGZMJrWy0CrRtj8yg5CnX/1cQmVoXEuuZ7RNNrmsnLtsz
BVQKC/y8yi+lFVxMvVcqTzwnrR0R89wpi1hrxkzMgwOxKNMV3XTnqsmVmH8fAavqCKPfApgEvmVW
/SBlxxrf8Mt3946J8dcd381iEeJkvgS8/VQ/CzLUuehwlVmaLkg3AlEa9nG5AKoi7asN6luWjii2
wQ/Gg9EKZJYeSfQi7P/9Egck8JslQb5pYUnAy028vkczNfZz7Up75w69GqSkWYgc3orqOON3PJfW
HTA8yBLnUIdVbfU6V/Z+WZARNqyaijisc94WSRop+U6rgJ/YLQ74Z4PSp+pBh0rGCRPyeApVvZfT
4Lk+AO6lDhXoYjoPOi6s/LzO4NJZ2ssu0nwX1MUrir4OvcpHCjxsCI5KmRmUf0NEECruAwefH+Ow
NxcqLkSa60l6ETzcIgBvhCcCH3n3/lck1guiOHX9f0tVv2FxENSpxAqMPQEf+ZHGImFjRDcwaeTZ
zbWeNVULkQSzNOlGcK16WV7HdEVaRdILM7jr/Ph8ey3Lh15SIS/1QmYgBnbzql145Y27i6HdcCMK
dPyQVuD3aCuz5dHBnXxO6zv7W//J7m2XtzCmchyPIEhbvNHowZsKwU82ioolKcYASgwNHI5ojwlh
lAffsqkkNZGa+2pDHMmWMUKxPbuP9g8r4QrdprNR6o46qfGw+BKaniQqtV8oj2YSTOeTbg2s9SIw
DrGwhncOV9VwY0udVOYWWVYspb8viXDyM2fUJhx6eKUrLwHy+BwSeovzwpx/h+rIV7TafSaQDYiJ
vLvoLCGYHXXbfff+zz+X9SSfWAcyITrxyo0pBUXs45+lNGNlVEY9lefDG9wa/mWgO/MCmZN05Agl
Cpe4gI5hkYe3NVgK2/zq9GEfe/T36YFcSGJOD22AtxQCAiffNsPI81iZ3VaWpWyEVM8mx0pCRydo
2OIM85Dv4gk8zMiG3zSFJ23T+u5D86dxE4HV0ouj+gkP8wnnthnvPRzrPIqIualo8gGdXqxuO75q
coMrk3zMYyUvoILuuaptaxf6gJe8LvQoxRX2Rd8/HC1vunDpdT2FBigWJkmup3dvU6c3oq6HCZ2l
mnxqpCOPxEmNkdOjzH4fFhyXtYQ4oqKdt7XIjDGmzfgE+lagDtutWTwm+s9cxQB1ZIqYpteBHj48
5FLLN7er2hmdX6la+DepSqvpmlwQIK6GmlTDs1vfjHfW9Jg8hWGTFatU1DhZIOYY0YLJ1hRqsdTE
o+mSZNKYMfemwZBZECPBgyCBhohQEaoA3sZkKZ+fiZ3aN6TaXmZKahiRIPv4yOE4wquabhuH87vq
CFuNZjwHO2KPtAw9I84+tXv7wqGyg1VjoBgubNtPMuQRZJB13EGBIUMqq4wyu7KGjoa02aKRAM65
jtB/3K4Ueorp6uUegtq9vb5VkrsgPpS98M/d3EJJagT3dzezVPieaGdq/1HAkuE9W7HQLM6ofSQx
KVehnMjq0k9fqJGrrabho6LfIW/rNWeI08wqPyrPWrwk8MbsAqPaSfpsO5TLbDh4n0Lk30V6eqPt
50VKGH203bmqVkDZZfC1trr3myNivh4O3ngiziru9+MU16Pex4NYe2LYBoQ9YVR1XQMfBAuLPwKN
5vnqQbpef4yUJ1xYI5Qt7lnoWyOr9HhGQ6mHNAIYm3nYjbdMLEAtXXooKmWsy3tKUesH3FQiRPQC
HmP5EFcAQsGJhWh+41caU3aNGOw6gpmnaRW0PrEHlC8jyVv2Ae7ekW1Ncnc7F6Cf0CqqJBRL9Jdh
GWumDPioFEX9RLGK9hsMULYwbfEuwIMWYSis6v+cCNLvEz36JvOzHZQ+ZwQpKBg2u+JZz270uYmn
CV603GZs9pFl3W5bZYr+VsmIkC8biJsicNYhgJQjLY80NDmj6BZ4sChrWKPRDOHZdI4iT33ORnYy
vFCOBjnUpFXXz42+e5HlL3NA0SCAp/Mg9G+uIOhz4WnCZGF7SXPSTDxo5ZPKgA/jNO/of4jUwFRd
NxjOOv/njC6P9eBnohNWUFZHz1hgMYisqMDfvhSasBs2+bZ63bPAUY/IMIaW1hhYSittQltEjnwo
qOVfn1RTp6eT5COmicTxghwoyPuZLQioGJe/HfV7RX8JN2z0vs/p0PrrwOsavVlKpACqFFfOnyp7
NLOnfh94olVfJTA4aaqxIWe+JCNynCZUZJ32PUyQJGWFR9BCG48l0AtMbUiYQ524s0dvpYITXqCn
780VIqwfNmWFWx7Y+aU9qYL27Vu4cHlpfSiS0FxdS+cmjycTfz3TUR+i/jxLRhbSp+qQpRZ+xSmp
M8bVBHGaX0+mELs/2NhLVr80WuD7MAmaPLc8YuMFeGw8whZr4FCYyGEf/QzL95fygKB2fPN2TxtD
klJ8c56e8XQoxXEVZrsVOjQRqYXAFE7pkmuxe2SL2Q5Gr+Kdw7mf689D4E9dfltyPt2FLTLT7iMa
Gfm9iX6ZKKKVA76diAQm/QfyKsulOkgchtAEi34v4vlftcs5LQSQqdw1IP4Kyjo+YC7RUJxTcR91
eoYE/rlLwFQmpCvCgupcBa46QpaAxQFp5ZuNEiMq7P0YRhkjnXdnbKwiiPP0/41h5fMmdnGdjbya
xecKkOAKTPkXGCo2Y1ZyxDbE+rrPXhz0TrSbQuyYkZ9pQmF7maY45Noj8tuhXaVXccsJxs+uJGzD
1G82RlM0yhWAkUvSmwOQUCZ5Rnx+pU+/eQr8lA2L9DoEJxOpXV8MXwTxoAcstWEsgR6HhkHHacDA
n9qwEuHWmMu7wqv9ozCYblUweQXGwaJPMNK5BQDrWDLgWUzalE2X/bvha5uY4Aajzy3QZPhqux18
CnyM0zlCqlla8GB22sf3tjA03GrWxEU7Rv4E2O//ueORVrRYbpCjbhjwrC5XmpVPuGt0CE9h10lE
qEqCa1Y5G1etqUryQ79BFlKcRxGxZtybZLfYIKxCmv7fkx2fh9DsJ1V2ONpoAzmeLuU6ltlX6j7+
ngRY7cI89RDdlu6GMJxOoXPJTb00+QOZYmA1Upf7jTf2sibuqfWMhYcx4K1PF9xTSnvNqOcC6yX8
3GJVjy1RCE/sV8Vl86SM9jnYm9lsiCbalpxb0RuPDrTrZBJF7R7t20+GxE16jFhvDwljpBLwupuB
JxwVIn+10kxN8OoYgNWNDwBHVzA4OKw89SbTooQ7KwxnDLPnLSyad+f5UEof4IRy6fPY6zb76sYg
EsJx5eUqqg748+yKcjWqLsdeKhP085g3DMEn7KfyP0q0sF/3niZ835wBNtiPH7vl6BRiNnLNRpXc
nOMILV2wvOGOqBSBSfRZqAOh4wUDy1ZkI159RWjQ7FL4+6eAmgRi/IebqVSVi0Ari54c035aCEoX
eq67bqJ4hzmfRb09+7pQybJS8BLyfoPLC5+a6EJCHjD11tZEwqH3sN40bPOOpKNx15QpSOMp4mX4
U14KEcbvG8xMuL+XT4kda9Hast2sIagvmPKe+NWQzih8wSlDNkaaFqntHwX2dCSvmB6Shy6HzgLd
cg/iJ+ls54dtIA7oJd99RTfTzVKAw/pPUw1k4EQIaT0QzYNWIAzeAQmtTyFTZ0CknM9Rc9qF7r7Z
2wAXmK9rXcyNK5nixFQ7+vf3XjONqH6nsdHFWXiJvLxrnRqrgSLRQ2TYJhHaMxBMRcZ+jqzF5mWH
HSGPa/WHYI0IcUtgOjr0C5M6bwcbqt8I5oVdVwpcGYt6PU0MiV037zGfxDqAY8H8C4UsuxoDgUGW
dknbYXSI6NlpemzQ+pVniaj2G1GpiVNWPHynqJlylH6EOI7K7iq0rmFbWRzhaBxyjLLtDn7ofbqW
iiQQ7KSA+1RHkanOp5XZP/IbvTb6OOtC/lmVO6hE/wqxdJ9KFyDr5RH72p79la7ismaen4oBmOIq
VUt+e1iUkRvELfNwCWgY91MCYZp0g1sHmG9QsS2CzwsfYjbm5RAduIVwfokYJ/2Enu6UgGfpEazi
rQHAxnKrpXEOjKVSXYVt9FlYI6YLTxAUo8U4B6X23h0jWeQU6VA/k9VheyuTlUuL90T8MEJy6UvM
kvRf24+bTf4J3Qnkjc0Owaqc+ozWs+fetBQPZsEYHJ9nHNtAx99UcNGhYNVao+W4/9TzFHsCNgwO
sC4s/e2s+79BqZb9BAohmwtf5dcl/iPtMrAzoGQSYsLFLas6LDwtVBunsvmf1JrTJ/fJxwx0N2KZ
EOjyMFW9Zumif5C6GBFU3uejHhdw+M4GP9iEhhYlCRppwER24VCwS8Fwi4cuEV0DaHBNUINgupgY
U18DGt1CU63WuqGmwVdRCY1DQLRuLQEld/Fec053ExhZdokOScUYWLUuLINtiDq54WsFqRe1lsDo
idFTZTkEr2twnv1m4hTThvEZvvT7putHWWPzRvoDRvWpPXfEnd6OgyzMWMTb6j8TI3Q2yR6GMWgl
RCSKCEAf+KfMrS/x+lMeBntDx7Bi8NPcZS65BgL8qLSyc3M5mYjPtx4O1IP4k2UQihnupS7Qw7j7
VEgx59dlfpVh+sUxo3nZfS6mAip+QJ3KOMpuHLLEt5b4Ehcyf+bs7lKAkM68KU4wcJn8jTaA9CfM
oWT+OPBZwbdwVWMlTCpu15kBFOdQgVqB2b4hS6hsIXGKdiHVRhpYR0A50vAn4PbyiCfcHXRG0Z+n
6MD1Q95qSKPMAszvkLv6MGMHwRq6jFLtTkedt/xbQKv2HBsVpIfNIEthhJLVbnoG0qyhcksMuN5/
JPkzy4TXFYeWBmIhvxnYcKubJBsOpelvSCn6GglOCE7iK4Eq2VSZvM0Ut83GB3AljawSWRDysf6o
5zDGPbHu8cCuUEJqwIWrhGBlt5kn7+ZLjNv99lydmbdpgVtghsE9NPMmEjS4zhiGgSJ+ouCze8Uc
IwzM5xpb9Iu7CEkHEDnPwVVVR2JVGnealyg164eRtdnN2G5BMxM6BlzG36k61ueos4CB7uWf/LKG
06h6A7Heh1rz27Pni632boRFjx98utDU04q5pXbUaKWWbsFVA6Fd11E3WNPdiNVDxNc/u4aQu1Kl
gQTCM4HkBKBgGxXBu33u/pXd9JQQpt6snej5CaykMikAwQ4aOQ4d/nUHnq692CkAp4c6HiA75QLP
MAkCX4TIdSuMUKQkD5fSxNFBUlfqsIlScpBBK6aK6/ius/MlkoOkiW71xBQ2FayEy40XW7x5VVrF
SXJxb8g+9MH7A6jmGRC6DEa9Xhd0/EY/3atFgo65G0g/rqCzMv5ET4CmV7z0/nT3sfkACeQ/5iK/
RPrH1LDNjDohkGkQKfmD+we536TXmY3iD9NCR82HavFjSQ31I+1NYqJ/FeajgJIQGIr+MIP9ye59
8IAzKTtetaxulQKVQz3Z+GnBujOhPjjWnptidzbODjiExb2MEzgf2B5jAe+qdJs+XYZdRm5q+K4P
lry8L1hH7eMNhUu9TH/zkd7rx9Re5FsciMrxMZV9I0OzRvnKfEe6yx6SUeDqBFDjY36I3wCwE73u
JKeBGSdbUqK4VaKsHY5C95ENr+tfHNeLe+S6Kll8OTuw4LWA3T8GTFYVZcU+7rpwREXKpq6GBqY8
AcKeWIXZKbI63GSPVxMtcwaAaKl/9oBHN9JEUX+zvLfoHXH7tQJTh0+B61Bf8O9Ob0kzuwDOYBtH
UcyraUfO5p/PUXtp7L3bk4AkFs5jHM35SfKTA9khipHvFhxq/aLLe/NA/k3dKRtu1PE/kltuzaPo
hYqPUs9MbPxDazLKI0ZwBW/hnxbv4DW/z6esU/8ZlYFDtHnnSHzC4+Rn7dXIl738xVgFc8erz3hj
aB9c1jucftVkYknam0wpLpc545x90pdx8bzt/TNfcT3Mk0OKmg2mFZ0GULKG6ZlQ8Cbvma6ZlIC8
G0PMb9a5Bm4QYP1/Q4vuPhHO+U3vlcm2rtpGT3Zql0QWniksJry0TH2ytWYqpzMkulq7GYGayraP
TWhpLSgi2oeuqfva40+uf8IqYixzqfXpzWnFCVNNO+44pIlne1X6N4Rn8Rv3ZX3pRicorYa56FaI
FGfMIAx9TevUkLsP71o+H8aiweYwrwmOAbgByJ/jz/tWOwuQaNy74SWCxTpckbA4neKOxWNuBXBA
jRPS2L8IX7eQ6kCpTJ21syoxzffO9VVk1v6HGLr4XppMnqDHyuO4tt2i/ud8IItGzBftsuRNuXz5
HCXspZJxOwG/p5VRMTcxkQXzaA9MB3Lq+u6ATXpK/jkHEsPgrBCgxjW7KPp2QnQ6UHpFU26jJwe/
8Q2/Nia8CiiR7qmP4M8gJrgUjVoYrvOyGMg14HEwTia4xTxiRGc1LBtyixHREXrcn+C6zxl8QeQt
CzMXoeYHwV33YRXFwU/2Mq2S9QN2Keggn9Gx6Uz1+aCByuGjCFB6GdQrgKnD3FQKaGizXaOViG3C
vPi1IUdszMtKtY2B92I5Iej/3ZzUJwIZKPlphbXb+UuMMqwPMujsfDQ+xVHcVPJrmdbEyO7UMDnY
dypD1zYZtvuPD6EVW/SMpoU3oqxueb3mlmtFmcRbDLT1sHrA8bnA6G/f71soJWp9P6+XSmWl/XeS
AqP6i+j4+IIERPyt9G+nAYtio/2A2Bv0Y3+z/uyxQiYJ5B3WNIJNESansyzgp7WbchR34Bc/xCWj
OKr1l7ECYuTkbhVmT592VEUDmeLpC4EQ1nvGyvzQWbrc7F/32QU2t5GqoyEeVIsAsQi6prO19IAB
YJv3YR9qv1En5bHms9n+q2B7vI4OGfWGuJAsOSOUPkfdyn61HrZncdH77fBhLN62UhjIBrtDlapF
U2RciProsPEJATDbPILCepwcWo0ckfgNxbymo9trX/i0pzI3wsHNnHjAJi1g/7xeheoLmSeOZxCO
9EjFLwfLNWMrctfKxII0sPzCwLpaqwBMTtOpnqTtcP7yLiDB1UFJvgyiYaNQM81QvuHP7xaPf1ik
JQ8bPsZr3wkNCKoFpjyPqzIXf538holmJUKEuGq0z8taB6mmtpCaYpG5xGj2QrjkHIVRQwo3PEwA
lgNrThOwJiHq7CmSJPItIjvZDfQLgHlSggEpFpUpI05AxPm20Eckm4Wm/KG0teYkZKTRDuQc9EAf
xIb3GekSSaUMfrSI+e3kKIDeZsVB9oGu1SoN7O3r6ALhX1uRLoVn0E3Kx0fs8oXQY5NUOK7Adt+I
0gY2Gg75Ct75zRT01TDfPpyWNcI/O2ffvZi2ilVE35LuNoch0A8iz/5uW9nn0+DLoCIG6fgT6qE6
iVkCFn+BZebPvi6EvfMlKnhQjgwscgy+dyZ0OIY1hwS6q5JZ+TF2PbIU3UdZXBkO0kKkC0uhY9aa
l2z1Mj2MN8iHkW8hCiQoakMIIkPbkyAuYey0kBUEy/N+kRWwRKAwDzp+tZjozyfpf4jRffqp7iTp
K2FceImLpO4T4RSeTSCMFpVIzorm+ZBOZnELX1yQlnboLT5QZoo9Se3e8KsZuXt4JyKJujTaMxHP
TxopCasIFikJAE+4L6DhG2V5N2kIa6kv28b69g2TsD8wvsZhzayBfrkrsEbTF781KBVrZ9mBlTdG
jqDOx8ggrOX7opOChxqPA5+bwDCj/uRzCv7Dk45zZzMg4GNHjMS3AoXSppQbeq0OeCz0rha5V6+s
EFQAJ/+SLWkZEs/7VEU4+DvSRFwGI70p1OHLbwwOcqcyCOqy8H/UI4onEpYWwTkrWMDk6XA8sYlt
HwiP38CGTLTP6MXU+ZtMIF9/saJEar/UWF22/D+TmsI5WIZB1jwIUPTzqBHdABLWmE7mR9UDsglp
PXEJoGnrOV4YU7ACYy5haoXeoddI836Up+XDvLenzFsETV3vNZUcfGNNmKD6ApBQASz+YXo4Sr+a
qTRMLOTGEZEUeUbAP2cbOEOYdEVx5ENkMsCBO5MjRl4Iz1CfvNXNKGVu762y5Rvlw1OirpGKarey
dnZhWZQKVAkulB7vhdJuBDgusg7QhaQFasy1XtRJUFT9bsXv4Fwl0g5idmaAlgs8Pul9aUUx1FPo
k+hUel2dTE9DCDWJd5rUqVpdjHe63Tt/6YnJ37i9DwIG1I0WHXOkaARWST+oNc6zahMpgMvg4Sv2
8JmjUfEX4N82dWz4WsDjXvTJPkVC3qR4OpHEoWap8REWtMzLPGdO+ela15+rgkIjstRWjdJbIoH1
QolIsZmKnoJxjrw8h4NseswFrQYuImHyoWvDDKy/duzMtvyhmbjiP2OZH9x7s0LthMY+MkgN7D2o
0+xlmI4D3bA5Wip52TFay9vmVm3EWpeJr0sQfk1t+zsQ8zDnYIMcZ0ydQY1twaWf2gSmznbo1GxI
oMko5eGlJkyYEHcHlYY0WNIUl77/qiv1uHYZxhvsFLmqQl/Tclx2+jkHylrD4lSQmr44hj4ClQad
MjvoMJSXB3RhFWJGBZwR2fQqysNtUoSaMTVKSrxoGa6YtIgcm5mV97k4dr7HoALhMbwnijWRRWVt
DYzvOSdexla3vV3bSZJGgTrs2PHY3xoon9DgJvpmnmTRGTwLSTGNrX+GJBnP1Csqby8fO8wlkNcs
jOBU0smgJsya7sZy/lkARsZjyi2OOrOmOzJtqI+Nwu2LHvw89qL9XdCYTcBdxwWaQiiGw8CrQB6X
df60BdvcXZifsUhHHJ7ByyzNlf1CE1VzwmNxZ8W84FiAAVyCQ5Chzmtdue/3wfJ0RQZVwQFR+IOb
QTISmz12Hwb+AfyzAYzgivN2mr5uPus2Z8lFXYV8DSokjghpIYb7Ly2igdV+Lk/7uKK5NrYEmaZP
tB7V0pXEoFrvFasThy18/G1kIA+//6TOTnTarMAoXq/bLq6PNImytdMcFDFi/USNWr4LSYZr5b37
ur8rz/EBQYEbE862o9iA8KNRkNElo/eZ/uhOOBg+uNO82IaO+DTBypl5wTDTiK3KKyNiazMhZSov
ZEAzSyGvP8afacfQy5kQcqmVOyadzSXYYcamlSzSp8J27gOXmNZzYXRoL+b6Qgc5ATbQ564p+/sh
p/qhE3Y6NRbRofZc5iEytfi5yyQhvHeSJslJPvPjntknLdgvT5mBTUAa06e1uNUR3/0NwdK5XMSf
+gS2WpadVMi1EHNWdqxb0CVEXePhGnRqw26rksaZX/op2i//oXpYlP0Xqj3R/R5YCkaiC1AY5cFO
kFgZGQbSNrUTW/u695Mky6zgU04Ep3MFwgYRL/pXyvYV9Mi3VGAnxNbPfPV4pSfKEbyhSEyhDsgW
Yk0zQa0GlkJwWreoy/G721cAKRf5BUG7vcVP1dZbjha4/6pbipmLKB/kCxrZ+K68y8Aal4T/aD+S
r+lJhgqVldLBD1lCjzc6WTIAKvz+kLF4gDF+ajx5zEVi6jgRp2dzMjsv6FFy747j7MdEvwSYgI2S
8Cj/CxCSrJImZ6EmZG3BOkLDZRR83AVLvj9UrxlKRoC8amOnDpqCfQu3G+IXm0TOf6BFOJTD53ms
b58Y1HWUKneI5TxRaIIpSR9bMAurgKSSuZ/iqxuv/PzC79NRoZBVb9rkRA855LNMDOJxgorB92DN
wQRGaIr8EqDmUbybrJk7X0bqNGr2j+L4XELPRc7qVkLv3i6S/SBSrLcnaNuID7mYNW8sm27LU+Ux
MgRxbGFb06yQ73tS1b21rdlVSNFRhsIC0ohHbXMOf8bI52sSYPKSqSP3+DnB/svdXHsAh4A4CvBV
CUGHt++va4Hi1bnUZm/8el41Bn0RopUnFdUrpSJb/FrQxBDx9sxCDBEL+bTzf+PAaAdzqAT0GskW
jl9jCfzPT/MF0xFErKHZgRhXO6J19Gp266ogf2VjK1xRps5Ja7X/w38ll9oBKavkUJ+cmEnTxHHc
Nh+dW2cufGUdmdyYgE23xmlLqFszHGfA6rnJBBsS9DxzGdX5fygEETev3gMsGqLM2pmsoAkqISEY
H9C4Iy9Pl/qiHVdBCGxeQKL0Q9iHb/Up7oZlmn/orJYaijb05BEXSKx+55fyyYiKmHFyYzvOvIkL
ZSBmcLU0rgOAGwiAbvCWtFzg/JAIvO7Wc+c1FyzaNeBMmoMX9XIhYGR6Uo5XZS2UYFABQaBhkP+E
clOgr74pCF9Yxg0hrL3hu8VZxekSUuN/EFaw3PT5iSJkRusoDX/289xD33WqnCnMhCQZ6TxVbysS
RJNwT0NCOJreDnxsWeh8Z4fmiIHg+O/vWQndB33wTiE1lkY6i1TzcH1vgk/VHxUddgHeRS4kS5Db
S5DIe5sJgrx69fMU3C6Ty0SKpAgQCQ8vW9xPGK0I4rILvetEYOxoDnDchvAu2b/x0RH4FxdXvTUC
mnDRrW4K4SERtlr0z/DIX0k3hfR3/X6tGQmtizbxGuaG9KrPpZ6MoP1vMq6kRDpMwGvZzwE89B4p
DfxtXfwCLhsV4HS0fhSxxhr/Q7tV1Ve1fpZSNIqt9zcYt5Xv1Y9IeoG6iQx3UbvjO3ncbn10sPfa
FQjwhI9hEFic7VsA5wP6zEs1cL3Kpfj+jFvbDX43G5GzjFoJIxrREaYbz6CV219b+CWhGXNjsCoi
X9EbSMwe/uXoL/SdbetM+nBno6vDa/+9rwzOPXVAU1dEJ0qK/O/A8Qa4kMhdyNBfLW1eCqmW1pVk
fbZAjoTunOGb/MJSlndaY7rd141DDcxoGHSO+6WJdAOqf7RQ/4kiGSFO8jPYgO3ygrB0MnRa/At2
XUhvz0Q6CerHKG0lCJd7Qtp+abso4hbyFEusvunWxPoCUoIydhW+nq3nH1BhnVrqZEqs0DF2k7/J
IBWHTEc1UJUPCfAosshUnp8wFAYQAdwaComV3v3oD9lalGR8TRC9xwjzy0FP856rGGPjSPYI3VAH
Has956uavt85fYdY0MpvoDxBB7cz09bE5bTdwMXT0hC9FGQS7RK98BoxMzZe6ckWvrDjB2aYCPDX
WzLYHDsUwmQmTeCiJGzY54humVEIky4zcURYxL9uQRaPPBHhPBn1Nr2h3hYHTF4CD0jMD+y6ZEfj
dCA322N9Y/kEcsT2w2/4nEwPOQhA4PMcf2P2rNML6n5gIlvnR/ccigw/9OT7bwkQ7bAzG/LAFfaV
eNhREX6FLB8sydLCnA9DkBWb2CFmHJ/iiV58+O5J+ckghMIWc5pqzttGEzhJq5OMFeW/9JOV1Yez
vd0yHCiKophSeScZRxLqmvA356y4/yQx77Rf6hdkTaXCC8xV6pi5qT4B+HRT/nDgrhLv52wYGpXU
4IGszfdvDsKWA2Jdf8eBBoFqQsgkurvX0WbqnYtORe31BX29BZOWe37SK3s2Y6VUk/La/gw6VgLy
4KrKAefYYXZdh8l8w97VYtFmd2rHob6F5oPiseubBllqeRZUrJUb4F1hsd40aJv/hsGu2LfkMxVO
xKb7HRjG9J1xjjrk5ZLH9dCOPYF7VztAQj6hQrc7RJj/jayKwxQnEp9ehk/DwAIMaOdP4wUy/sbl
fMi+I24GtGLT7DU3XhUHOIuKt6k41YmTQaADW+YvgJaC8tYOVMnx5Bc0svF+fJ0K7pYy29YsjUso
Lm5K10eAIZ9g8Q3EZW+rUX2btY52rGgFMprIe5x1AgTZRLkLSmfKIJfXI2YQwWV//P3R5H4e8BOr
NuHkhAWBEagiHcgZfY5MtLarSLcqyZryN5qf4HKEfGjxTaMZXMzdBusqvPVLUwLhkrd6/iVMGiSF
KmbC5708Xf77U8aJL3mu1Q9qEflaPY+NEW5zSJtShf7p0HUVw3PI3Y62r/MdBQBT1Yve4zOwyOE2
4no4jTLaYdNB8h00PoFjQVqYRm0CtEOPfa+WBU1+KaR3OXtYI+sUPRd7pM/xBEpSB4n3Zyy9qOdf
U7xyccXqzozoi/kj4w5M9C6efrHWhtrewt0drEXcK/TewTnko/chE03ZMOHbDJMtDFYQDxI8gAT+
PjsqODFs7XZ9OJt0XRif2FjdJgRWXQR48DtJhEMaUNZR71H6w8TY0BjWcKoZbF0U9DNOSufKUe21
hAMh9EF+aDZWls2dR3YCaghkasFkCgtR/kW87o67+SnFOoKuURLG5qzK6pEf/4Zv6zJjXNCmtlHA
h07AknfCY2rCJJm6wrqVrBtyVZ+6V9y/GGZo83OEun4GZn0ypySTBJDKf5hpc8y+R7KP9+L7WEqH
6PLHUCcPtfZmDoBUxn09M4JjkfSCaS3mp8Hij3Y9z6ILYfpEr/6nPQCkb/R4DEqR/1qCF04CO3Dn
ZUFy19OY9q9tUFPJrTgrbnE0zlt6nHC4dXa46AHHqE//RIngrnjtj8gmAcBCz2qSPVrmiY28wbfX
DMi9iKWFif3aIqKzz9QJuAVDwq2lvLeXHnaV5ocD7dNOungqqxBRGWvS/vrMetLTEbtOUAnAJEni
8CJvaWpCExX0HLR0i6gpXa56Ba7y3bQSiHWDiDL0j1Xqs9cGSnbiTVbqf8HQ+fZpQT90ZpwabaVI
Gi2kjZSwGeZFUOchUcfXTjT10dXwR7bHRVYwD4Jfpd8Hr4WuSkq5s3FPsbVdJUdK5k1HUtFywasB
dzZZIPpRH7sA4ijDL+QxS8vpBZQp1DyUmWUMb9uxyuh2k0mFs4eG9/ZMiOPdb7Oq5qupYegHYKEd
HiFfm40nabUGbO+mq94NDpMoY6B/b7mZ3LxTL71kZmbiBeAmyPGv+6ISGAr07cAIe8fAa1bDyCQG
lT+po0aUHPcptc37XYJRvqdZ/PMj9ufdQfQ5m6/nyQzVhy8J81G/rGizkIdkw61pKZrA8GIygLan
nfPCQOIpuj66M33MRPTWt1ywi+AdSE2jU4DVvRrjBYwxQCq/qCehWDb0IJlJLg9ihotGft+oiToo
IlrfGUPJGGR3WaBNG+KMn7t9fj2zqcXIiSM4E+hHQjDtcvBYUdLEBDulcHbdvXlTHuOoCOOcBoZu
CZnUmzM3iWIkaexcPm0kNG/DEeK9GMfg0D/NwY18fis901Y0VVrbQn45DluYOym3ygOMQV/ufQYB
5YssngO8XW8pL4MsDhIE67jEBJvOdb87jEsKH9z6xhZOsqB2ysOPK6NO/CCusJnGpxXc1jq9thz5
I/vR4th2s/IBMhYcLuX6MYFoPJjcOWP02BYNoNU8EMuCjr5Uq/QAF8YF92TtuiqomHLv80+sk5ga
GdpOfBkCFbJrj6981iRGMDrGPLDZ/uYCYm0507sGwq96WS5vRPULXncyhuE3DuvwtfBMiLrO08lt
z/gJwMOlzjnYxa8D1dccYqrCBuOd27qBfLD9u0Xqp/+F81tNEqX0Uxybshie3le9hkqRLOVZYeDV
/jJwevQ+1/Lz2L9yH0xxBL2WzQEA/ebuQTTUI1TE0mIBxFXw9HPc86S3G3dDdwHqHtwBtJq+FTgM
aYhluZyHyJgPOp+364dxd17A1DWZYWl6fBpLvr3RxpXwTlx/2d5dV3w5HJgSCv+KJYCTo69kerQU
NkIY0s8VZzH/bAqnOv0uec8wDIwds6MGMCYAoaHr4jSHveDS2yYww44N5SYkXIKxWVG/TreKoEw+
E8Glt52Kt+9NAaz8dEeOOqXPMuHSlMrpVCVTvowpVEuci7qbkWmmlHwz3WqKooTXrbh85eCK8HHx
r3avjyPd4MuGEtTlxhYdYON43RK4SuOmu45VcXS6h4MoxE1CQe9KZ24ijmNk94Nkc1BLS2mO5jd1
HuKMQMN7QBrgSirdfsWcfSirlMsVet9eRMxFKoVXBn67xp6wZMWA/TyMXknpTAXr8udl5sliyVgQ
jZaxdFDjADMwZ/m909jmCcP2HJWbaSH5A5ZbO9n353rgdcvhbPefUNTPqIF+OjvZ7ZR6leljIYry
RV9rNhj5b4g4l3aydu7qD3SlvKnsPl2fQvozTXPLx562PL1wKYlnC8dWx1hfAaWsrjlGnK90OSP0
Myd2kQfFjhOq87coWXVwV+A2k2G0ON/im8noh2XNWH30N30xJN/s5jWaHBvVXg/SbvnwNKDrORN8
pwbGKcRoYuZp+Qe31TtVgBcNATu7wA/b6wnCSwqvDPvBNdXDiiVRomywCNeuSMKc60f3g3SlH4Bc
FN/t/WrNXe+M/p/UfgOSPiNc+pm0LW2RwC8ZS4af6syIzedAseGc5rFfe9lOePVEYUdP5YOFSXVn
VXIzk2nfM/0ukCD28Hxj5CaE6v+LWjh57Cfew7Zba/NIPFK4o5kVE7dk/wtPSWj0QElo4uEbZBzZ
8rO0o18vPkRGUFhRFY/fdi9zKjO5a5Rk0yZReJfZK7U8KKZfMCaot/AnbCqe4AH3pl+CSvdzweji
snhOjLJqapQErfmMlF88VlYAvEglSyM+dgazZ7qWasZnmmzWYiQ9Y32A+F0yheezbck/CQcBc6vq
6fjatrdlPiPWgi3/24pwuxlMBLxxFBI+HUDaOPVp8kS5zTLwZhazWbyDQdOXeTwM3kAyoGeMv6Aj
Sfs3ooojD/+i8oXt1DuKa0wMuCsdFUmW0THgzeNueEfXkpt1kBqaHL2p4s5it31cfpPDkZIU1Olr
PAEAmGwvdjzG/eDrIuIlrLxuMjD2EYtKSdIA9oAQbezYOSN0GGmYRpXGhE/1owJOpuYA9xgAyj4n
LDuFVLj99pO8mR6KowVdI+eWE3nUxWoIga7npo4Rcb64NDEW6TjU2BKUfNzak5A2y0O7ZIKrkFQp
GLZV4rqo6IXZQYlOIyqKrtUHtCPmbunc5aVz0eBrRd5QHw086j8SRGiVGl/qMhBPJE3dpQKFAlnQ
MF4pWUOey8KSBDtGHeinkrz4avtiD/RgK6HdwzdUmt1yYMWhuOzvAv7ZmS9XS4bRu1W8GZr52AFm
KxozRiPxJzL94JWYIBrne9PTSZKlP0PXpXMOpgmtph0BbTUXvbT1J9BjI0+1SgMGNvM2lQs+6/T+
CBAFTyq6unyoF8xPwCxojsRA9pxB7Wi71AaoRjWAZLh/7KDNyDO7pExo0/WEY8/7OOswzMh4wNxK
pnh4guWNhNaQB3OJlcP4GN2Lc3eiBumeDP3T+mbdpgCLQy78RkRHnZ3+hBOrTdZkbxg1Ol5WGL6J
84wPX3Bm4IMLvLEclP7LcdsDNtiBB4i0UWXbrwvXeuUmmiASOWP4D6mmyBpnl5UaybbVsUJ4uO5p
xMx7c0SsaXaEAWJRdqY5ACixSyDg8PW1mUPS/tVnPDUHTW6ijTNWz6M0Z5xpFMz6glUMDk5n+p5k
w3ZKCwLz4JCBqSIwHc2fKeTvIpGBA8UHjzdvivy2CTCni/LfLVwtDKP1LVHDQ0aOOdT584YgZijh
ZHkJoGoMrtGKdVDJdr6DxldTuZ+38q7k0L28ntsBWwR8hmFasIsGMjIrat913Cp1ZyZGULtwFsmp
QkYvkiaav0cv1pXldYhBDBaTt9gQoJoIamwKMHRMMSvtug4vDmDmhEiOuO8nTh61KvkwbX8XUjIg
1v+254p6LFMUBBdQRxMJVtIKXxpfIKTjnyCFhNKN8gWNpXIpOpkO3XcpPyGK6TcwYS1GstvMYD0j
rD2zILux8k1evTn6u6H2VlAMkh+Ih27Tk120RtXhBGP6iA2/x88cRgOZB4GpNQq/dY9v2Ai+V7ph
5lZ1fb+/A1Gyod2MX8Gj3KK6QoZ3QZlgVNyB016PhYF23AFibs9m2Sa75kjTU/375DohY58eVjXe
ej+dk4Rk/QWenDh5kzvWEYQGVmKOed/yrsF2Hv7Pfnu44kLdWDx0I3u5zsPXCFc0BLX2mk2kh61P
G8Nbo9w1TeKPlNwzijnnXzYVQ8DgkpDUkJyda976Jl39QRQVHatCVhbW4JmR4rGXOtKodCQemGto
1zmcEU+ekKRu7QwGXBVHC+3DIB7tS+WnpJiw1IbsVI9EoIDsyRsN+vCxGtMwCzrCLxZlqiDAFXF7
Y5BT6ScmjrgsE1TYeJhP9zK/vjzdHpFwot+Prp47MmOg+shhav5i/7RX7lvNRHp+fgesj5gdcBlT
mXze026/UJhxMaMB9Pdb6fHwd3VUu586BXSHAyLrzEvRLJ1tNQs/Bso/LYS5c62/K0YHVgDB0kMA
N1/59Z/c9x9Kh4whm9723TLDUndfLp0mSCzzosW9IknVViauvwZ4f3TSy2+L1WwuAjFgsrM3D4fm
EIbH96NII/urYV1VOwX5RYWNt6lhFfsIJy0lAFpSfBcBP/Wvz0DVtTdSSAOoesSAc7CH99mLXW2g
iJ7WBYa2h1A+h73AhCqF84Zga0Ri2WIYzGh+LJv5EhNBT5dyC0yrOMOd5esBDLWBCj/tni3AxLAr
AZ5uRPKJk6AKtg5H4zohwRMOE4BACHSugiuUwpb01Thmr1B/qVC6prmLLiqKd+2nDHb4SSMV8yi5
o+z453SQq0+nltdhcV156P5CQrEOry9irGEgrXxHiDggfDH7/N8OKzYYF3Mop3TmTrZaIJj8+oXr
uGPfAjy99Q2hP8al6LWaENF+nYsPBlrCtfGSTUCYSPO9hW3IHfenF+rR7uyDEWIBqwucddO2ks6u
gyBuMVqvKC9J4MmmxWWXrqq1wlIucmUCXR7XqPiO66bM5aSYDbfI3qHuurV75Z12tu/frS9YkQ+y
37wI9xKHT3dftuOf+BO7IUCVBlqtUW9hUFm9yagy1Q22v6fNZdbNqQgknkVFyQqW9k9zgLsfq/0D
hiHapHLvABnHJqdERlXrAEAnA9Nn5uW1Mb3C0odUFymMu0ydZDcuh/+MmJqN+jELL4xhg4GJt0TN
zEvK6aqXQ7HqfE7Ip7sUinYmNWJSdJced0BRvnFiKsa9G6XDoCwp114Mx3COcGxgrm38+be7SyWh
ERKWzmZiN99DsybLb7rt3DMrMzU97/1QadQsEolsQElyYqboO18kQJTKAU3nYWs/aHM5Nab/kn4D
wVMnjNybuBxuy6Z25xU4Gsqtd3SEtw9HsdnmN3FC+hnOZPm9uW9+VybeezCg4UTM8EgKB0W+jhjd
VrIpl2no4fgw2FZ0cXyGClIj2fIlhHFZUWgWTVKsgpD6enlj0FbxE4VQokO2cACZwKypua1RF8xb
l9A5TRh40oeSAlxR5iYU1vzePpmdsPJ1TVhNTgkLTnkH1CRIc4Z99goG1UT6li7+1Niepubt6qTV
Mf159v+APVGdSZXVvMZPJAqz7TNMlDo1KYLLwhPoFjwfG+T9thwDa0ZSWw6VMRYfTY6ItzcmngGE
xJFxfVlAMyqmqVvmuDm1uhui7Sso7g+nmRrgjilD20PEoblbkHxZCOlKhGJUZiLmt0QWEy2d+O95
sePF2jVhagrqUB0AxQ1971VrXKzBXaIVI6Bpo7RveUAUYugv/VMHEHo+k+U6PkeOxHel2aYJdlxh
yw3WF0a8ki8plZ2JllfNAncql53TR8xjHHPbm4JiGks9I3olI0rUJvRuRO1Pw5EGU1JIt5vhM7Ks
xD3MnQxziuK9APsJGrK0FuJaQlaBL9rzipkEqOQooSk2xvPbZWcD92M94QruXFLS2Jmn1LRBxDOC
3xMsWwntdGvs2/NdOnTFMq8AWrt5C7Lmmu+gJiANLGdYSI9HiN3Hio966QECDrzeYhbEnd0d0mmb
YcEJcF52VF4tiRuYlHGSKX42M0C3i6X0Bu/u8qaA7BxMmpyNnAy4udFowEt+NEIWH0/XGzeCN0Lz
iJC6Wlfc4cXeyHOTZiFQnC7/QdDcFnTTq3E/jUyvzwE+fHmOBIr4lFnWDF6DNXoEtNNRg2WzWcNn
4N/ZQAMmbWaXU5Nf60ChMFbYTgJ1fOB3g26K0UbL5z9s28Z7UjtNX4lhtX7t4VaVK/RebCKRm2Q5
dBOVZ05G1d9mr/9ymMekvlMwstla2bNBRDlc7DSVya75wjeefjTKZ9UTpa3i/M+g4CiqxENpyWsE
nYaqMVPMwtSgnLSi2eUyyC644BwU8O9F8BHrbvniyezfEA60/WV+wISEJSCpgqtKJuj8t8we+7Yh
jo0rebk7rhEIf867NsKdIFrbXlppkxPLoOpnxA2ZBNhKQ2G+HIZvfD9InYb7yNnfLuAhYbp+gfU0
GTyECEzlmCGDtHMdnkSvouWhGjqQPnFRpiZqyh6AqnIQbFWefjbaSQfLT9ydYZQe8P3aZLa8E2na
i77mCv+cf3Kj7PeW1jgZdej/CyzktbJpc80mrC/6jUjdsGJf/Jk8Tbo6GXgBSETsZhZJl0O//mZ8
U9W91tGH9UW0I9z+Q15kho9otoBOW09/ls03jKbNnNdtlzely/NvYGilsYOMWwIKEZDp21fWaVAd
kXmJUHGa7SrHjkuHyW+0JzgusU/dK8RRPz9x5H62gtHWzNo7RB9p0yO4446LENvXfRNcNT4mq6La
2YjhH8GGpmVY79tqrWErtoN0wyBC4vnaf3BEz7gri01VfWYRzHMpQ3DI4S+PXpEOnxPAZ/0sJyaJ
/YoPybVoSKwWhDAAw8c1BCfp5uz0rJmWWBVyKM7qoqvUXU1gXVug2A+K+YQXhaThCWN2EbOetg22
S5cIV2dEtDeTIesCbzk7m/wZSVz5iqLyLPiud2TqRdpn3DmlRW2ioMVHsmpnljRRO25CJDSlvUAA
RKl4EZXFTKvKGVLxXEcgmxbxK54QD7u9jXOIckx9lBV4Ok3ENS5FIX561DmlGlIQZ/DHfU1ZFCrX
bBT3k/wYsT4bM2JzRHdkDBC8rvvvGAgSlAH/xWtZ/YNZNMYu5VRtPloWWuOCt2R+JX2m0xbE2vWm
cQ67PfyWjc/02KMqCS5L3GV93/nslkKHmNs8arrPgdmFYbQdtXC+Ke3thL/VQQOyUfug61vSvsrW
PoHBK8b0kEgFyZkWsqUDTsTVnpgm5iKOJel4HUJyP9MFfxWn+mFZzrOE2iRaE0rJq1rQOSgWOFW4
o36LKSct3yr3VLOAuzq9DFhWPD5RTuRK5oFPoDB2iNQT/UZxk+hqAzGo7OoLKOY14/e/SqzSgngX
RdqnWaCKj9kHodDHb0RN1mKQdVS9BooQSdfQ/kFVCn+e9I12YH/qoTbTqo7bE6Ux2Sn4dq+eIbuZ
QljJz/eEoHjyyenu8XdotEmQ3YLKrCeCYpr+BZDPsCYLgWAWESX16n2VfZPaqLRZEsug2Y8l3cbP
Obsc++rQC5NAYi4rC/REElWs/zTpQf0P2KFCkLnj8+lIquynz4a5hRQNgkzyQGeucttqHcMrVZpv
QEbBox7luL/LGGDjfkmsKanzL1Qwru+QvblVYZ653j/ROPNpCECDkZSx2WylagwGV3KA+nf/yu4U
TnJPl7sG+zcEllPyHmOnJtbq0SmXCKS+lXSCTwUXY8+ynbeF1dNnXNaLdvTCj0WItMCuzMVS/KfF
OMHcq1B9R7A7sCI+MbbyRELhIewEqVjcVR1Fe9yYcjbZgZJQRbp6OHctvmSuGIGSVxwkg0Ug1awk
cibJ/DrfrxGlpQ+JD0tyuN7iDtSCCsUCXcuQVB6Op303P0+dK3iBSiGtggxfHrhAesWjLmDbDZU9
ynE/UyvnliiBrchAIZ9CPO53cMk99KgOKp2EVbq9rMvhoQyG4UxDeQu+C9uyws4lrCDZc/tINcl9
rIT1GyOicLf2zz+xUkTwgy8wXvuqqvrX+Tvzz5PimvF02gnWtXjuEfN4G+PwBsLN1MhaTmo6Ozbw
A2F4uE5UrHjOEC5KACufPf7h3UuHOyb2AvjHSeNCNqZGQK+qPHiUhIiWBfQj6Ka35pK4AvpVQfHq
gD74XyPmBKSJ05CRo91Nq7gL4XjxvzBmewrn50iMClAPTEPd1nBZBrCZSP0ui6HgszYE+y60LopZ
x3w1L5nTlnb8v8ycEwRduEQrnfg8f8wcWqHSmEIO0Duc/9DYp/n7O/jS20z2uAs1nc37VECIZ6cm
+zBf49XmStfunM0AxF59vLqaUR9HRs7W4i6rLMpywGVUTkvyF1s6FT0fz2LsF479px7u51HhKrum
2J23vOE6JQycnPbjFCrf7moN+zYKmR9c3mzZbIzXGEx37+vvd3HRvh1Bs3jJxUUmKEr6PFBYSaHe
LYxWia9+Ps9kVquftUTIhrKN64kdFATvTvmMJVidE7uPxtxosszJrQMu59cXyaNzROQXWT9oBbGs
bUt/1f/URjlyT3IFza5KoixgZvtU5aq8j9Ur94fBBGfLibqdBv6CdsKjhNNXjoMSVGyzeHqYHN6F
y9ayfifoVv8feqIatks9d6NZB/PBMDU7YD6/Wlg1gQdWaJCF2qJSxvorDs0rqq58gNWK03xbAxti
aTuQSv2pNjDSW1ktP+xavlYCql2kvr6IQTEfa7+FFLtj5uyyu6AJVsxCCcFW9dLTqr3/mvhYE3W3
auJWex6GnoZLWJFAxyiGvINjBBpITjWWCIt0vk5XwF5SJRZqZbuG5iwz5kgzJFcTx2btPSxejl9T
PvBa1p0RUPY3TcyARPWPvLbDuJcvH/cYtM5eE6D3xbuEBiyb9ACZMo80NFjGS96kblpd3GCLMPkH
AQopZV1m4DkkkhuB975xm2sXXSrPC8xzOEhLAIMWuMasQMjG6UI45YDsTSuV34UI+nd5Zt5+iOIR
8d2fIFrtJwiXBigdF6jetkjE0irqZfDtEzRpeh3JNHeite6ierljGwxQNLfhMyqzjb/hT+f4ZDl4
MIPWmBGl4K/yXI9s6XYwd+YNzWXQroqYUfP+tZSKBxQJ31TmRYqLgygdCvAG21jIcnB37Zd6d7+P
oopF/vXgeMMb/Wcj0Jp/g4p9qqg5m9wWbrLylFLr2Weyf819FzX1yIXNuVQr/U3+aDzq0e+4Znou
pZ7d/rR9C+/7QmOJIGZCALNtj+tbPONJxd4eYZX2bjg55idEovnMt+JGT9bIzDhoY/v6MnEhNcNb
1F8G9b+bXz1rWq5GUdfHo1QRvs+Kw8ZcuHBh7OEkbu5nqb+zzAOSh7eGDDNE5ypnq8BO7uW+ODii
TK7RFMEJYnOgPBnn/AxrdIlb2QYQTLeH/kiCAEiDzbj6xADXnkuZ3cOjFmVZLaiZ5wXp+qAhmSom
5o1XvCBq+Z3ZHfsw3/GOjp5VkJB/2WQPcGx+5RnWKyMvyqNo5WhR2caGin1suwzQoScq+RpAik4V
tq4YC9A+xImta622bvpGyhMUVUGGacHaeBD6cG/YhVTUhP0u2GF2B5T0Xh31dNcpi8h+sUW34WGI
MA3JWZuoSrT/1xWYRHECO5Z0uwLfnMckUV5pqNmP/H2yZTyMuJ4TrE1wxuJgDaqGUo2qZe1WQg7n
/KZr02EBlgeC6e6KGRhV5C8/HHJoMEusiVZV+u/a5n41J09BMAHJA9nZt0MIelSbLIr4iEjBZXIL
5z4G289qN4yhpm1aZ1CWJIOr3ubJjv5Z9zmpLXBTz1ugvO9J0Z9V1Wd4uUD04NfLYaoVzGOsgkGT
o1lf2TP6pt/+n4Gw3xnLefDqMaReaS08K4Jm+t8ZJ3AMJ+ity8LhS/LfoM/z3qHbeBzR2cUUjNFc
x5vDZ3XN/KlNgaYmajFpOsCVMg11Xl5HPBcqdnA14uKkXkyu63iYmCDZlZVdghjwC4BQqo33Hz0H
OORf2llGEUlVkrpqXTg9TTWbBq/Awx3D94aAVXvWjoSuvtfB2uVdkTDt0nmSVUeFwjmb8lXaxtjQ
MxVsjJUE7GdzZbu186YSm/293sJn58DtXqyJGahZjTpg7OAFR6XK8r5OcceZpQCRHKv3DH0TwnLQ
UJAzNnZiziGxVCc1H+mg8WAf0jJp9sVOOU5ICsNNEQQyjmi1Ead5TxZKHXlGwDlxh/7cQOE/6RBF
z/NxDOMbFmJr9TzDYgEOoOWYdffKq+tn1XXj21VuAuTdkhmqBB/upboXKoSPzDad0r9e9Ha0GfT4
mHa5q4t4SKEZlOyw5LlaWUhpSS9CsK0akepCevAk538wU5KQl6rdcwAlaHM7fBkEiI2TMxmr2dCQ
nzogwL8J4wOzVXXhLE4ItRpFQkCoOAONPC4LORPlKKcwMqSuAu0KxLdsyP2x5mQy/AeVNcJINtIo
pVVxg2A9kiZvUcAs46/C/MGE2VOVDbxvJID+E/Y1JuM3d9IeW1GUeO1qEQ7GMY5+/sejhEZ2J1GJ
XJWEtnPGKWGVMznQ0GtgurzaMKVZ+MwVM9mH2xzIuQl9l9Em9NJ13qp77nJwn9lDFECTac6ZHJTY
Havc6XB2s8airSxPWw17NLl9MjtVFi9nDJ5j1Kz+VeLJmNp2vgE/nQm7Q+8gpAbs/NUDuyVzC5Og
doLzEYHjkFKaVPmLILYroHbrrURHu/IchLmNWQLGmYGCTuiTOOVaUqcizKkPwTbyh1J0xNmvJTCO
fMa1JHTjOGRKSSnGmFgrqeeRzOyrZBKwqf4BPHzzhLzYQ02776cwGfVcTHk5eXkE45m+DXgacuLl
9WccwleJiGKeZRFCwANMkOMSzqyPmIRilGGcve5den9WZ6jnIwR4D/Z/kc5lnkDe/RkrMCH/yKo3
tdd81QK3xP2H8gCoyfs9Y7baWbLuvLYYhbjTFZ5NIJmsYz/VOJunZ0F1cO6fMGuR/w6rphS2hp06
4P4Lpv0cUdt36IKmXQoSQhFBo8ZomFDcNA4lfI1Smteqjn+WSprrUrQjwkmePp7ffC/eDL8d1mIh
0od/iitoGSgoPDUPcEwIdBTQrJ8Wgcbw4E/O8EBKs35c6ptIeStUVOlqCZCH8w2yoY2pUp7q4Ynx
kkSj3SEEa9aj9xnq4mV8V0ibc/21F6vQMTxo6IML1n6CbDc/o9kNq8rRAJyjmIxizc4PvxZngdgw
EBQKpZICnbnVU/waeCZORRaW3tnEIvOkgE9mdJSpkJlT3donU77PwVi9bnlMhvdKyj/COABdca6s
cQyHRFnfjXO9KK6K/XtqoyRV23yq8AwlwdJC0eVdgJDhOJ0/3tAjmCkVIHqYHhzvnsE+qmE99UlS
i2Yi95IWCga3TyEK9RmWn1urwYXUmb92jfvJdTGW1FxKrbjOesxFrLTkeB6VohLlZb2rmxhisJRL
CA6vNoKvqo3keUsJI6/5BjQGZYg8gres/8Vu2Y2kJrRF+gjcW+vnlvutNxxmtJKbo2ZW9SkLtcDs
84g611XYPEjPZf+YOLSheM/IdraYXxbPjS/l+OlxcuniL0WyBFzoFVlBUWg+GZqvmHrbYTTJnpJh
NsZFtuzR5e3z5r+GSWEGg6AubazCe8HeCaGpHZVOthiRtDItiIqGFSVNonfqTLc0BlD6MTrC2Mkp
ZVg9ZfasulVPhSebkRM0k8MovTtSaRYD8N7ON/RWzsVuuZmEpvb2pzz4r0Fw5+JGm2y1t0ubjNoG
q+Gan/pUvPqW0Sd/LGawzvrIJFjbl/6Q/7bdR/3mqMR42Llqru//pcMqBC2LIsoiDTxWYP5Z8aPp
nn7r7UUqWXP18Ab7AgUtmXpWLfhRzKmKFHCuQcquNVt5tDqkJfycGYBg6HrPYphgH+Q5D9ly7gNg
kHpL7ucQucP3G7BbrN/aATDl5EhcxQmVFvquUHR0FMoMCyWnjPpBj87D7G+ph5sD5XZ/YU24vHjB
Qxc4j3YvvrS/1Lqs5Cb/kFmR6h3qmOOftH9bCjtUDis9hEh+/0FM0QbTtKAQY1csHz/edtx+rOxq
cW6QmsKXAIvv75U2Y0H72OeLYJpqg4KZTc/xzVBokrwgsW5CGsT0uQbU7Okbv/IRm54gsk5uoG5m
sY0ve6pHJnv/siwwTY3r62/tR4mDlcZLJZUxuTIgTd/i5UBQqjxVXloYYt8+XRCHDYNzf2HRy3Hs
O6x0BupuYeS+4YPe8jIKl8k//3x1CEh9BD+D30URYN/YeakzMjIhxhYV8jOZCYdIRaYoL2bmrVL2
+N2QMHx2y/I+G2v44dnGvDcaT+ynieo84eFXRLGC+byIRHEMqMQAPo6/vIPNF5FnJgT9sTpcpf03
SwIJfhnRcanM3mpOFdTLM1S5JH4p4ZUKhMtxXoqLKg5Af0Eo/xx9+FDzvskDR6h2MqAopkhNA4R+
Q5nxxxhSOQ5ljRqSClOsX1CsfkGsHrd8CFFHAO/XPWJxqRhUtgKHjGL/FGWR3fLkpec/vQcuQ4g4
5yehayQiX1ipeMf5IwZ+KMT09Str/n4V5bt6e9QzSquU+ZY/gVY7kBF8VyjHGGPmwC2uPAor8INi
7Buo0MI1k+zbEE7AARA0rQJ4iDNMLVVrjyKqPBnDdII5/SYo1y/XucsEmglIEQaZyzHkE5kDj89p
TNINXxB+GvBiVHmNwddWBSIPwa3LnnWKy8/KL4Ac02Hyk5vH/wDmB5Ksr0RQAv2BtIq5sT4BD6wY
9CLli0oVgZvGVABdm6+qHVio+hnf+7Yt+WqWJp2Hq545C4NwYIehy3DSOFUk79mG3LsfojSwO+m3
N9pPPm/1qIrDfTIsXW3QdpRvnmOAAGp218k8VPZx/a0AwS3tyitumWgcAn3bXI8kMRuYHoJ2q9u6
N+5E37/IQ+JVGLj7MDljSRHVrWDC0fI5baJDghUydkZNU0tOyE/SETv9TYGoK0DGHUVfCNztjePv
B6e08QSj8MXFqYBr1OA5jq9pLDO0TNrGaTZj06vEo3iJsXbcLYEkPwEpH56jVYr0rOAtVUWGv9X8
rCxkaV2111BFfv2pU1jK3iVVaqXRbP1LDuBSMsSxSAzIHZLYDdEQHprDElulQTJNJoDEj4h+Kbi9
18FfEJMYMDpPFNQU4byYOHpCvZqrxyEV1qgW19aitmiztl9ecfvuokJlr2THbdDrI/9P52xLBt23
jpwe9kEn96IREDceJiYd1ad/79EzsMdyF3t/QBEK5OK5T3eg10mQjmQ1jNphpDb691bTYN3Y5eVA
gGaa2VjVg7bvi1IXr0zccvK8Ur5KIZKx73rP3n9rgTjnx08lgFouDMeBpy/PhAGfahDi9FKZy0xk
Z66Cd0fgYDWY0/JSfPqfhtc0bMh8mVVPy3MfEcYvWK11VeSFNwgToJKK7Dup6/xzg4vuMKVFK0eY
0odSIg8GQC0CqAAh7lbJ13l+sah/srPaHBdqtxuwa9j2QdiORB0SdEvE4qGcELMKFeSRsb2S+3zo
4tiaZepKGv4HicqCrpROVqQDOzVyI6+SVD7qoEwMccbzS84Rvy2m25lKTivZ5NrRtqmnqZ6QmUgp
Qyv9+HVh8j3MnlbiiF2G+O4fSJZXXKohsJlRJCfs9dWT3DrNv3psTakzzTPG9wP4yQimc4woX+jv
LgeDD8CCGIB6EXOsRvJz7orRY8yk0xHOtlOklkOLRaN2VFQh+ywTBCLZUkS78N5FwJQl0T5eODdB
mCe+VqRGs/xltssqBWPq1f/IZo4MtD/HoCDW7aMb8a4yzSzzyet8JBaKnklpIhfHPPtPycb7q/wJ
n6bKyGdGI6CUxvl8zhf/7lY9DTgQ+92ls8NE19Ne7mXBoHHRt8EnJjIoqpH7X3Am22Vi7mDwQJ54
LtK5zx6AlVujfE2rUqmHf6PDQFiJ+d3yGbakJV8Iy68xqrHcXdI15g4TqMu7yGd1fG+OiDGaTDJB
HXJS5Lh59+cIEuayZC9rF2ishLwPrON/e1ViImQrj9y3Z85ESQ5PK4EYcIqOhrvfNAmII7mqeW7Y
j+pQ5sxwWXQFSYnBwxEnaMNcH1X/xY1sT3bsRGaf04B1h8dG7rWsulBkqG7rmrvf48Z8kXV4RW1e
30qt4gPHovFF8La/GaBCqT6L7VvJx268StUuHGhcPY8n0hYXCuQRbm5wsvtW98H6xlTnO7uops5M
hhR552wgDt/H6lzph3zyAwkALaeo5BcO6fV0AMNe4KafForGVEFaItazhZCPW0YMMPAICR3g8hcg
7c8/6oMUBrMWuze9W7vFq8/ha7anN881qqTg1Ibia1PCFWcwvr/GGL6l49Q1Kw8Dr1FP2fD9zoWR
IrolhhrhPEYmnX2UIb7yTdJSRNzKGM8Gm5+QDe8x8peNyuasEAaDuIvFbdChyw+1ED1TuJPIRTKN
9XM1LMlFHXVE2AVOPgO60JzaU2QFMssgSarR8uBQuukmuFOwdp0ydiytVVGEoeN1nCDnzK2HM6mj
yry2JsqLTIbiA3wr59yoRo3OfsE5PjQob2Ih02g+FiAg09e/KzfRRq4Sd6VGf6r3xGFpeh56V2cp
0wVTM58V4mNbZh+Pq6jDnC+JCnrJBfjkEbGY3X1xESIYxwlI7olv/OjNhXQ7oKWEdEKWNs9vwUty
ErQh+iOKRfJyjxukrMBzrQaaUc6rXw6uXcxVFn0B70wgypb9kjRsv0EbHbVT21rAmOchz68X43WJ
YO9Jpyw1B2raW6103Hun8fqfh5TN8G7Ku7wWH82SaSj+3JdAXGSDTjVpuzJXyOrynaoPPtHaxoOE
ACyvWsxyeSj9TThJqL4d4Ljxa1Wf+6VxpCsgPdV7X2YltoGAow/UlTCXo38k3H5tScmfQ4eVcfvA
RHIV+kgK+ILHI7H4z/wosIKSOD3x0pzrMUAzpR8FYcMXzYcu+yYl/0KJu80bgx1nrJVX6bANK17/
DjJd0Bow7VgClrfcKCg9UpC7tAv2T+12SIJIHIYTBOquymoYHlypEanamydl102E96A0VAzO0/K3
893bYnfQjXHLuJTpWXuQzPCJ/XHX3wi6dWqOfv97QzZH1mIYIGxG+moG5JFcb7ngg8Ctd3TX7Z8S
FwWqYOjfM4ZD6r03BJGK8ThioFBmpwBpZnvfivOJ5eZ1tk19NfKKNSOGTnOLMDclRRb8f2pxRr7+
qAqM0ctZpjA86YKJAUwFeFXVpjXLYbmcq0V5nnVz/fyAr3mGDxcJhwevmi2TCcPKJ4P/yRrJ7opW
V9AjQQi1dbCAa4QOPzLruT7n/Oq+ot+rWK0iEvndm/0K5/zr8va/w+5w4NOPaOAZrQSW8aVZHOBu
M2T+AgWKBesh4AyrcHILDfPhrxSlMx8bru5i9jAMk60Ha1/lAt2y+uXaDEw2KaZ26NRB28lcQiKc
Lin4cLyM5TZ2Rs2QgB2FURiUniXxhBWpRcLD1kABEROe/5tqEDrAZf6UOoPhjEGBiZKjtLzzXRQ6
cwk7/tteTltnFjDuuoXh7pVmZAciKt6eDm9uGFix55Pcmz/0yHv5JexHNvGdwqVJugndIGI2v8UV
1lQ4Uqh8rg9fffNS2dQkdLvbIkXWS3itnu7JbbekiMpEC+MeXdg3JioAvqc0Vh9Xj3dUCvqIY+by
pSjOvNVJdKvzTvvyXkDo+YNElJzZwzuTrCcKZa5fK75TPjIYL/n3hu/ChuhvRJDKfPHP8FMmhl4l
CR1qW8bCHOg4kUiSC5yLlh6eTAr5NKdeqmlH7Z7qhg1/WO7t/YTHnGBUDg79/BEgD10z1TOzZCCM
BtJ0bHIMWe+DISlG0Whnb7zLnpHVrGWgzuwp/TZdWphFJHR0Ckj1yec4GFP9uah4cwrgXUoUv8Js
8U0rRiKKmqap8OZ8R1sy1JlFn7mTl5c8bJRTYv1hNQYRHWCToQMKzwIi0a73rq0fu5QY8igEHswO
ql28Ml1ESlrXmwUGILtQ1pCPjq0JdlTUbz1Y5c/pJmygFrFsy9QzEAZTfG9QST50pk2EZSlMc3TW
lqzJ8bYpUngFHn0TmWGrHUqzu4ni17GzezqEIGcK3u4s21NAC8cmwK6suxzh3BQ+1GnVtSyTSISw
rlFqX7iRjQA+tZIplZHf10jjTQ7fxlxpIE8Hs1PMX7I8qFcnw8YXWXK1+8WIDwFgHjbZNybAKrCg
pjzn43EA6lWxYFxGsNTJQRnIpAqd9fKmQ4OFWm5N63EewOdPwrmr4vVYVjUV9/6KwE/NKxzXJ9NL
opP6bP2eUU8ncFQ3Da7QG3AigUBsP0VEABpOzRx/sKhoA5IOJByYOhoEDxLENtmOGTytIke4OMXu
WgdiGe9EZTl8vRDnoB8oyLlBmdyHime99r90+ExEmWBn903JpsXpdxRsAfdS+IvpsV50pOdFc6aP
syl/ChZo+Rqmd5dEshvpSU715ojEgh5Aj9DfovGX8EzSgF+aMnX76FL9AyOXr/3KnLWeX3QzmS0R
WlKVPjDJO/sCDS3IOWv1+iSumx99QpVE4Q5vBTpEi6/SJOF0hlYy58lQjgchz8DMRus+b3pes6cD
RCZ5qQmwDuzH0KabybEyJeNAdauxEG4PkFzP7BSlEm0Cl1oTbG5fRjOvltZ4i8o468Tuuj71Ka9V
E8bK3f+BIFGY69Wiym8zCbo8iQ22wXUkfoIp3kGM/C7/uYL3/0O0qhu6kkTMJv8A01UVXJiAXc4x
WcOhSAh75+vSZbB8cCCg2BRzQYy/TZW7iPYVbM39mCmoL0lWWGDrEkgi4+FF8jrZ2jxhYTN+yVOm
6XZvR1M4X4PcbYXijLKC3oS8ia/Ybaa7c5w4RG/pHOTNTzPxKy4FaG1/yepZdiv5kBxB+5ZhKbar
BGfkKWOzVQQXRB8NywhvMz58pw2mr7q3r8ij4nU/xfgl1g5o3Rvun9cIwgJ7UG5SvKexEayvth+X
aW+p9HSXgoY6zH88Pzesl5VqVjkAtUodJaVPm7mFH4JgRo6CkMgzJPtSut3hfFm5lOAzw36aM+1s
ZPDLVOZmPO67c9B3jeplwS1mjRmYeipoO8JhD+hE6Vxtu4gQXrPWi2Av0lFFk58AlJ6OBUcA7ZnF
QMxQhkEYw6ZwnI01XUSz1RSix6SGUg3gGq+4ZfLF2gZ2lO6vglQ0VL4XdXu7ybhm+ts/J6vf6thb
r+zxkINTr45Tl0T4Wsk2ZGPSXC5lkgK0NzIvJPI5Eb4w3Tv41jAihUYKLwvNzOCTUaMpLCXPEsRr
9gk413mST1Z0PBomTVnMjLyZ2LEb0CFRkFvQspTL92H3eaXG5mJiyvaEjyhvelcewbEcmnnX5S0o
bXLeFFg0KyJGEqgLF5jxGXcl7GDNrxmmRYvfsyXqILW5I78rMb57JhjSjQigdXsJ+D7KIIeruabN
XAxXESkUJQRXNayq8Ww+J3jF4QmnCwEfAVLGmIAlNDQyNY3L3FT38YowtD7kdSzN5HQhzZLK/wA4
6Vrw5Af/fuTbr7fg2vBUDOflMKKHiCKdIgHUfFoEfdSaXBxHg+epJaI44XBYMdC36D4sNrR0vKCg
KE1nV+uIysUM7rE4dUMt9VuEf683ZHg005O9BWZQoERwdCJKY3bdSGf/cu0WHvLdQCCBOjyln3mb
WkdiGJdXiENhNwytqC6lzla+16k3DFvJ9539VpRucjR8sFKNM4Hkkeps1tbLTn6Zf4gX73zTuBaR
TUg+WH/3Mxpi+2ObHi1rdSJNK+Js/GVtDsErr+NEiRirtvy9mPXdnsYbZZEjRHy3gzPLyekizvrG
4UG7WHd7ojmMzFADwsBVvqAXuOf0Dqq0hn5fFmonkIdifQirCT2hRAmk5kZztlfZjiLvEVs3Rm3T
HMzeMe1UoKyCC/ZYn9xho8HBuUsLz2fjrchDkDwC+CIy5FwUJjcLgZmSVHF6F0inWIYMH9PBXGkH
eRPBYkG/DgBDl0EPLXYZhbn7m5VepUGOFJkMKQQhChNsSi1UJ1Q359UTgTgkQw1dnwSalN+nt55w
5kVimYAuDgSlob+E143eoJOTBoImugruRvM64WKBih0gTQw1eq08DqtFln6GcoVLOmKJPORLS9S9
htSzIcfdi1Yd8m0mAyV1S0bl6vTHaVZm905rae27SsSxbvWyE3LZXsjyZnNaUS+B/DvL39gMn34e
hoskZSuDHXGn2DCLF0PJr6stsAWJVb6Buub7UFaD39u6zGRRD1kzClAiEQN2/9uBgYmh2OepHpoe
GK8D57DwpNd6Gkrrm+E2AYftfRsC4fy+KiBOEvZ14T6J6PzSp0F2m9kmGwhLLJdgW1NDEDvk+MYT
NL1mwY+4AmqL2y5jj+cqrOJZ7MPRcnejNBlHA6m7X9ofwBaeQBZ0RcnOHnbuIpc9kvRLorJlGYwn
/hcvnU0ju0DAM2N6t0mfZeNQHxLBRD/6CiJCT+2cCehLZ4vjUAByGmhTODo+DVDftdpCEfaDajqy
fZEs1rPBEcCxYhbYiy5ShGjhSZF65U8BsMl8Jv9ndYfQoU3vQ/L/jt0nTt18Bl2L+K91+NoWq39d
dixqYQEsvLooIEEXI71uSOuP5rDjE2t4PKjgvuCcWpRsXHmGFEARRdzPGuw7DUg+nzfFWEjPg7ew
21FBPl76gMTjgzFoFYpmH4n3SqYvJ3Es4gJE4Kkv+o02alguMOYACtnwMNLXdcfZ2t7IHD5YIRUE
oUEHoWG+OS9GH38nXtTDz4A0y70Tr0sz/hbmuiFY7nCZpXxeFbNT3uQIm5MW1hiOGylXBUVJG1+C
9lKr5YVTDHpB8NRv31d7GHHEVzan86pFpSg6hEOgDNJV6g4gdSBr/VhpKQK1a8OHqc/N1OGa4pfS
rePZ1f0uqpu8KB9E00jbvQYsQTXpp6M4knIlXcVFMFf+CgofNvGmNww3SKqeJlyDYE7p/SoGE58e
k52hjivu1EvLwCTrI48wFvWrha7PqTDg0iVm0QOy++dFe8p70Ilze5oUrWhip3SWGrI/Hgp3Qww4
B5y4psHPJ+4QCHZAU6w3dExh5gyZrRig7IgR7lghLSaiLAm0YoeFkqHCUqM6aIv/zNt8H0oS/X5T
7BB4BAeyJ/99P/GFwKF2VtE5l16muuC16Sm3HY1C5lbokPJtBswredWzR+BfDV8BR4dc7TuQCBoK
Jd1RaAmUbzpkJ0H5rnzzypxlIUwtBtY3W1hbipZ56kVuR3PUtjDOcMZB/4XrKvJl968v6Mk9DAPD
v2o/9oRZI0e0naxckhmrg8+xyDta+/pMZy2mdZwpII9zpZV++o18md/auYlDkXNF+r6HOuMtqHIE
qCg1hb8SU0JF1sdoveOSfDt7clBBYKNAtqSq0wr2sMidf2g4y0B3EfdMvaThjEP8SwOKyppXbrXd
pUV25yLxgHTSyLrxwqvkBp6NCwahTkHwUDYLTywF0o3gdCYbzsmku2Yc+yIDK3fSvo8+Lrh/p3Xo
cZZ5Z2cK6C4+6LV7hAONsJYY16djivAxK5w3xS9ircCj3waNUYygH0vnkHqf9oRVDSWZ7eRbqwUO
3r1gc8tMmas+PWpA5OnIDvwxAQfpS4fR89UJnAtN+Zya5bwNHX8MSRrfGqBfvUx0NKDEveNgfiCJ
JPTWOldnKH12QpVJbja9xJSpgLTsjnHNqGSCsyYM3X4Vt8Cohiz2+a4z60zy9qEjbBRO9o214WKm
udnN+6UVYfTL3Fq/x4ZV0ak7lXxZXLduWvQS1wETImtC6sFzj54MdbkYTeZRQZstWbuz4jnF7cPe
BglTKAmBVKZGCPb0jG8YJHp9I1sIUDVI1cxp7V1PbW5aVqwTdCH1O6JvqzNKdPuXmzpMjwCOFwQs
E4xrvkRtUGFc2u+jU+Kpy1zZIyCrBml7QUA7MQ5OzL60LzaQzCM1wBXSkkYdvnxYOFGhJbdXYMBw
kA0cbOlPmAFU4Cpn9yZXoIT457lYIFhyQ918ZbNlbVqxCAodoyoGScu1HL6RWY3BaEwxyR68drSQ
xZt5paqpq9FXDRgXSv9TM1Nb4XHkeOEP7OnRbc+hNyhde2n3AecNwbAnbdvVXY9CtlBDYeuw0Cfo
jVe0LQfO2ZCOrSIfblHvrzYYLgSa2MnvwecMzMjdtBLqUIdyCVhgRIyO+RrbyVI4NYYt6u+CrjBR
i+BOWrKP62n9Z1OBeHeEZhf89ash82rogvqGOtnbJzXhHLRMcqoYi/g0TkokNe4Skphpa/701MgO
tPauhJav5EXVGmcq2Sv3RfuZu1IcV50UC47CZ28nK3D9CSqW1rqSJ/qsgJWurcwFbIVSTLBMzEbX
AuwPOUAa6pV2jjZZYczFqLXOzoHNUfm4zEMM3thRAPXfWaqRQHZpUvG7D2xcmhxr5QB+dNFafxE8
aW2Gje1jyAYu5shR3p1RRQ7tbX1/Qe+GSDRrwnNDdRJAc1fD94bJR05xWoVUT8BBUBERzUk/+IL3
/PVdnwKNS+bplw837oOk0IkfjESAaON+H2oRBZlKc3Q8a51kwq0IG/IPtiXaftp0R7RDJRjZBZks
yDd6TWwaZ/q4TpRDt+jJSFZaM1dpo55I0nL2M6InR13HLXsK8+ihJTRcZknlHdm1jvMbghcnz5e+
nb8Qk2bRTKuUeLu+Pyvo5QCJe1/bjTUaBfNSG1YaX4dNUZxFQSNfJNWQE2CjUbdhdtu2k2r/O+ck
5IME2LTi1aqFVWvOnO9Tk/+9KAXN4ytqyJw6i2qZ48T8tk+vreNYNq1KJWCM3JVQH/l77OHE5lOV
SYdpd5BkOKDFtzPBvL7N6+XnFZhqMiVaeVyzXw/v7DHfQKPTgX9qG/3kTFP/aZENfshAWgdQhwKM
WMMU61YDDppix2abtSNTaZRkfbalhRqFzuodjKtKZQNPwzCaAwDzz0oliyMX4Y04hY8JqtrWEBHj
cr9j742n4e+nY7sSIcV/36Oqrk6vrkAxL/a/5XxEQpKfnKZ+nerNbPIKkvJOWA4de3KE3BXypp43
8snfqQq34EUELbcJYtLzogSobeCsa/QIvSUZAR4s7scL4K1Pt0WKKwAhq5tooG2LvBBdDTOS7XuM
CRZvfSMn6ae3ZzgYVeHv98UYvYCsz4JRelJzoxakTPFTbEqY5GsT6xvSLafNs0CMXtRbW+Tqm1kp
LyxCbWhtdmauZTlKLTf3YvqMAshlr9LXMc2sgWNs6wqbIrulUz4j+oAV+/zWtPH2A822ohWjDgdP
FHF0qCEG/aA1K7hFyr6+U/Us+lDexOS3Zx51CVL0RVupWB5mCePxeoU6sZxa/KSjJFrRKLxYckYe
4UG106501MKXTt84vsi3I4Aa29obvDSeDKVkYULs4YRPF05c+H3CL5zfbjas8tBgU1n/M5ELefOB
wYQM2nEmDbAp6ihf4qADQL4Ks6zz9NRM73COQCdjZN9Co8YBHtFsJxaBBJzE+rWnSuJbGg7PfCO/
0cuAxfCtXwY8tEGDwocafcoUYozrxfIMcJaWT1IiKdfCVTp0yKT+iAZMtDX1cZInV2i5Ntbbk5e4
1vLSDH3f5dmbK7rkQUQ/G+cdzFc5gEMMMSMH+ipkhc+SkPbeyL/JgWot7sf+nfvu8TgcK1Tx4bHI
bkpuU1BzlRy0TeIP8UgXQxcSRCcshgE0pOGBiOC8nAnFiYkkzQrL4BLAM4Rku3pWgm1ijCudPLyK
ytuBeAlcPl+Gp3AL24EZ+xbn6yzovI/whGVl9fY6DBXp6+wXD9XzKexuEmnyr+JfycEQWv2/UCDd
3vdS/SVnUBVZQi/ZQ7U+bRAEi5Qsug/UNoqEiNcjAYjP8BNZwrD07pivFuwX4wDp+sSZOq+F27WU
XR4jUPqHD4CgG8WN3jowCTb6SSS+MSNpwHLWMLD05mNJADb4aTpIkiWiTjNnEz4b4xy0kCD0tbVI
Mzv/lhRwJuRh+L2dVVbl/4s4Qc9WiAseXg+6Yx8jJwFprHeEkxzqewYz0/S03UXzOQj6XSGEufVb
eDbHaCXKkZuYkJ9iTD4yLqfE6BQoUoEc6yPu5moDdkGbBxghiVBT5LYtxx26aPeDEVTc1lKID3aF
hYwAIOJH+ZNIfYOehLwo5LsZnjQg97CasPKc19AD2InZAoKFmTsJSyA4K4x43OBFBcW7/Iq4VTqP
SknRKv+uSoB59pb6VX51ICvrtPEgWUpu2TIw4Qsq9KzsLPZVkRNIuMFOvXqwjCwgVzz8izM6Sgms
rfEcDiJLOLxWKdvtitfQc9EFmfDnnPAix6TZ1wJXzKRP9ZufYCID6hbUinRH+699G0HZYiOh/Qp7
fEIw8rQPLtDCgFLDm9j9KOJSG9OUP6VBcnJx2zAI/nIBz+UVt9I+YdTh9/sXuvjImvM+dZ5I44Sp
RyU4PNl5EW2vFrDtlorArkZjbmRCHotT+s2SbiJeXooXWrohN7OD/8NrcDs07p87XmZu80f9swFz
R3Cp45yc/3GS7cSSHZNJSaEle6vi4KYtinaBzogAEkQ7Z4q7p7hlQ8zDs9dgFwjlFVkZjap7QiWd
/lefdbn5mlKq1120BoZdh4qcTb2P1ZMaJyiCgsR375UGAUj7LGYJWT+p7Yn9uJJUlXFMvczlplnM
G3HuotHy4pcQxjkQv2nZUxBjnn5htBt0VjxJZnXMr2ZaAkFqv8oato3bLzJxGq6JYXsZtMS3UTpl
Szu+dIsfxRrDGVS5zdmVY4UoJv83jI3IlpmfGUO0aBX6uvaLmSNeXmRB0KF1jwty3cN1aUQ1TR70
0DeVy1D8MnGKEE0ZUAVbHnis4eMb1TpLQMz56pa99Tqfe+IvgOjTNbtJwS75YG1aAuv3wl08+qIs
Mhs2PgTj2W9+SvDeDvaJ+NwaqwAz90TknFyb6op/jc11NW7Chv2p168/kT4B59wou2oqz2hh5+Hk
IkNhG5Vbfu8v+tObdSmXYGlQs1raCVo1LnQpySRxGnKOseCAmawCabfw/Qq+CeVlW0GSCtOnTM4Q
n6/e8rjjSIsQtl7JxXNI77zd9uel/H8QWkPHOgaWceAZdd8bdpFvGev9pPpT/SfhihRRLNkMq1g/
onzLKoswsqg+mMZrx04WQBUj/MyIblJNoi1RD+3GlwcARmKzVnIaPue0J8aKLNc3FG8HLmzNN1EF
z7UBsM90QmrVyx/axjBdAyOOW/5w84dY0pdBqMMKViPXojWbNMLvJYSGaXlssJQbp4bxmRCbV0gb
Exawz/N4s68a52/a/YWDcUxJY1fED59dG8KA7n97EGor3a5g3TOvInKX1uTphHd5oZs7a2+lkcCZ
xdlnuMoQfRzcPGQo/CUdFf5N+NH6vJhfL2QY0xbFLnoeu0WyCjt3lsqE2R2hL5UzcVoDT7NBMTZX
tliMzDgGOJ5OHcQPQ/r2Hp5tR87JWdEoi0MRv9njRKatCNIHAuF6TXl6mcjnDdC41iq4RX4OxU7/
JCPDfZfaHKe397yM0l5IlssCSklsE7+wfFFvdijIkT+45CXiGtGnfrlT1jKX9czr7hQ3MG2skKnb
7c6A76JYoFnbtY9nmKqjrJjHyQslCHDGxCGOmJd1/1x0Dpg02yF+KOqsdUuuvt6cdUn3IrUNn1A/
fWZBPobkQOmBIJqCMOPC87a1rfyh+D3mWF+FXmvs9sSKVYEjR39ke2Up0vCnSsBUPIzR4Dhn+aA5
qzyXSe8kFy3USR+LYZkAoZW3HrhxSNM0oUOtmjU1AzvrUjSwDK4YVybU0+EcX1ZTSjqq7GiVQSmM
ZDWVXSo0SGlCwUbwr5wYwnBMmgXPw9WJx3oPmbDNQ45dcakXAH8vjr53fXu7eFIjFgOGolpWXYbC
r5Aq2Yz5ewv9qpbUD87XJujP1YtlIKRG1VZ2m5gMRlyShxnSXJIHDOTesR3m7m0dwezOlz3ujmFb
tH7SbqYC+MaZDx4aIcfS/oOuAvgjJLCID18lyakeRXXAN/dCZ5of0vtBmJPfvRnxfKOtnEQZTgoU
OqE7W1cFT9rCH3Pp1Iyi66T2GA6WUmEBAaX+ojnZuROEUKkvmzl8m1zPfchdusTf94tm0u6eF2FW
bbiaXe0Kq8vQTnpjSg+IR1UvjXnrG8hj9RcwkBr0TgaAudw7oocviol+YX4+BC/CscBQnYgpXJoC
pWIaAiDbNMW2PAy0za7VWx01tadTGYr3Kq41ubFZvJZL2xxatOvSZRD05wBzqq789FBVfHxYaNUV
LdK+C48sV5DS6hniCU8ez7Kw2TTtfcpwgwZ843zArp78Q0EwQBH5Vq6luyOdUuFC1HOByj3kXFgi
odaxDc9Lf9rDuBhlaNdaLRPtXgTVOKn8BkOJ+TKb99+HLjCzDVGIegR+bTn6Pkmoo30ExUtzqbaf
ZvtRxKE0lt3RoD+y5+rbGAHk598g259+tgILH08sGyUfJEbLCoIvglB36yA22oyyi2WosT8H5pW5
nctXbloOC9ufNNQNaOgCnacA4X+f+WryJFztN3AuSELZL4mwGgdaACC9S+xtG0NpXzKrqSFv5vDE
RJvTIbeCRPacsImUsjQaq0Caou1x+P/HyFlXT1OR8pgU2Iy9nT22kCT1f7eOXI+S2FPql5VlwvPh
ZBBFTsthQ4MZOgWzhGeOTiqm2wGBKHeYV0hdbL2dLdNSbUx1I/ZDRWs2DvByszrVHCpCQKwfxmop
K/ja9RYl5s/0nKaCaB6kFs94ffHTI2bB2r4MIOEjyXyl5Od8SwSBNdZuazS97hE4iJ7aMgkFFhkH
YVoD8JP05ndcEcRQFnQ3Z66cpQ4yUseB8eFjiQmU3C0YXnQVqNrN+jQhTXWlAW7IzkSHAgtI52zH
zpiLb2PHSLQj6GTiTgU1ql3w/kggfKQh6vKm3scComr1q7ootbur31t1stifL5ZQDZI1pRnBGytv
EQZ928NrNGsX8M1vDaTFM5OOghV4GEDaeLVvCV1U6xFqPrcUYAhoL0gNGgmbX9iQv2yGGzUYFXIx
mYuXJr43JhROCMAxnBhnN1Miwh6wYUhrVLBQYUf/JhGysE7tLNfQUMufxsaSDLLMcFYVEzTT3D+i
EoYMASrK1lExLl72t51S85KVxrIrGZzXVyADTQWuOGbetVuF9OpJHGf4Qa5ph5STT6TPRZ92/tyv
hfl7f8Xl5VrnmkZFxHJE0EPb5Uw3siZjMYGwAiuIc/gsOEXLQZeooBW/tYdOZPxYmaNRHwRJUW7Z
jUEikTWOG/omimh4IJiaGRv0hj61nMZHwMCLxRUCR/f7/HaMTeyIdqG0BgLt1trzSrL9ld5OEqot
vgaVIx9P3W2UhHJ1GIlVwLjUP4Jtv2dxDlibWKYMJX6FcwTUOYPDUMBfGcAQTl94LETTTv749QiW
SP2V2MPOK+rINJPy4hCAHwS+yC7xI2jEhq7UwwSnPSnA+Y956C3FSonLCjRjUTJ8tbKFUKjqBNaK
ztRqvDosEUFKHKOkbbeOmv7LjHO694f/aPxbtLTHoASb3CA5UmYc/5jZorGeVKQJTAScjqOGjJoF
fminas5/EOJj+/WYgqtdG7CFA6dhyRH2VY6xIiD6GR4JxI9AJBRLu96umXTGXsMwNwrG708RlWr1
/xR61xWYp+A/Nv2oyXx/EYL89GpxmL1bsztgOAuGw3insdFkX1D+YVNLCeml0SdYO+nhd3N+rlj4
jPZ0vntntZHYPytUVXL1AXtv2WhLc3qBtTF6F3ccfonX46Edky98VV+iknD2DscMZGeN2KiDEtjW
ti4s5T5/JWd0arJDpBWdZVSsS/BFZSF0Y/t2APyGqIrLr6GlpXcAtBFU/EyL9vYWdfcDBCfFbFUb
q1OSLIPuL1bOZJVlLpQNrWwcRoT5RweBRLS+9qprv6QmuoCrg49kFDBXc/jqjk+byn7Yf+sC+GoK
71EKFGpQdGn956Mnfu7eGj8HyWgcJWtafIfC+lNlzgU89wBSSCgYcQM9wdv25YMgsD0N8x48/4HN
UihwPHCwT/I85sQJQ4zJeqcMlZvdh13DNnHdlQI4Eg5VRTUeLFp2Ddi4LKdXnqzpnbUprXVPjco9
LhZLp0ZrLoVWwOzLuZUM8rbK8Jug2S+bS410kWrQJCTzTAyOLQVpy5v89U8FvOVOzgGYJDIGCEgQ
BGsgOp2/dqhW2RwwkV0/xYW+Cthllz6bna6BOQlo2gbnHj8s2ncyp1MjiygpJYP1UXf9iMT78d7F
+Uh7QYmS12vDiv72JCvAZa1omTVsVFOaJo3E0OG/t8vGXLp2rUMS+d4ZQAynNDccd9X2VtnlB2WQ
sjFMd2+xmVjH7o3dVj+eGiK4fN0xpcgYsmKZppgHbnQmhHaxq4P4FALIudwqdpi0U2o9oY+qx9VK
XNO1Tti0kt2EAExgshYZ7vLtJiE14WVz7JowElIEtpPGKCo0nI0qLM1ZJ+frbYGtvvEbRGq+VNbm
KBfQh04eRmsfjbeJs13YT8J4WjF7CeF7FxQKHGI0Uf4mvzDI8bLner2gV17iJ5DcVLFLbjdQ2JN+
vM/ZBre18OX5aBshN4NM1oEC4pIS4dPcK+sBMEDfgv2LEVg7duscOLnusTE6keSvbg2mKmXG1IL6
fYjymwdboRvwYMeCmVCKCjvKUMD9A1lCut9cYYKjkcHzdaUdWbifHSUbuRBfR9IaeBUoDFJ4WK6Z
bJVrTMaWUetXSkcpe3xqeJHrtLLjwlZ6VRKFmxm8G8k8iAAgvtGhRfPcDP2aMnkI7SIXOsgUTFr1
dOo+cV4AUdaoN6G4L8/PSzaFTFqbNSduGJ6/zBJGHFJ7c+PWARueh9rCJIfhEMxTKiePNNr8FMAW
bhhfIfR0RF5hybZqvNtd+mdIus2PZZkFKOPQoxxPwYp+GL/ya+t45Ok2sYUvLHUZQKuz8UxZ5Cb3
FZdGV9JJtgO4Bu1NLwGGjmUpxTmYaUvmN6hUk9/AGMykN/m2YxwzTpgLi1gmvcqOzVlZbPDBszql
K31ify74CStF0wM/236zmrA+QL3GZBKVBOkRT+6bgDPJxe65Bt34NQnm/sZ1pprkjhnndrJa/v2F
GP3E5QL/U3A4SF19r1+XrjYeC+y4UpXWUYbCoqRWsXBve3j6i0TwoJSPajoIvsFQEsXc4Ddullfm
WcH97fXMIw0HkIs8fXOO5lVFwcImleA0wPOdjfeLLZyUAD6Kt7RM1jFj65u/Y6E2Le9DyhC8eWLJ
+m16157IxJSakv/ppluFlehlcDgXpf1TsZRMl5pda0e5rZlTw3sYUb7FZqkuuUHTLRqg2o3+YlDM
Lxi+Yzvv/yKPcdfeVQEr+dQC2ZpSSj3oqc28sQ87EO1muHyNUciGVvvwY9/GZORFAt+wAzMQ5PXL
+o9GhHEdH1mRcWYqczfbtHZxJSpRRd+hV3g4+YFaqklKl+YZNwqBCNICwQQt5J3tQRQR+foc4Qt5
BloKm0d8mcxJ9IQ/0VYKdzJdf/pvnC9WDUhFF7UWpUAcug8Xu46yG/s6T8AR2EMhDFEw0A7ub9TS
xUUnLmZAHtWiYCFCIcUITHvv4OZsOhTY3fgECfFoRS9R5lO7oM/TVgqPT4JobrLSV6IoU8X4zx2/
oXCQzJFhIIU/fPivPg928mkaNwzEIMELEl7/p2z4lWH5aawUpHw2jRTTBdS0OJBe8AkLw4L4fBGO
i6Slys9JiymWli+SN4S6avQ6GFm0MwnZ/0ZkIeEfH56JPwKtqPNArUJcZzjAsK2k14KrRYCpDgy/
sDemz2SQuufzVPyBwdsgk6O5scgFVHxsN1/bqUZ6aFVnhmxUtk5MND8tcItXCYvLfxFbtWY9M37s
flokU/e5xe/uw/77EX5zhEj9rj03GrMqMg5UdvDOYoCbZWkmrBZPsUaKHt2Bl37k9CLdscbBajLK
Loghj4Z00atUJvClnp3+2J2wYK9jaVG++AH7jgPhMaZkDHGxvM6hhLYjropK7j1EtZMmJlijIM2h
FQPXEbLBCK/iUkVmloQd/iDjBZPS/nDhgS0p8zUGnwMrrvcI/rU/SB8pjWb83EFnAKlhqSjWQ8Oi
oeBUTOpfxB9THci5i2CSYhXncw+R9z916XfXDeWQBJniq1wdYfxjVXvwJ16FaBZXHV1akAc5Dr4U
kxv+G3oGqLVpzLiODVZn8626ftObhldunz3pbq2Cw8jlyzAWKDWMeKF6RjtwmH49XQ1PQ0EEtZhK
LyGKCQuPsMlMyzxsSzlko/4QpCMK6eA3f5se1Uu2nXoO5jkAVS4N1WiAcF/5Fq695Yowfc+xd4Qy
VF5gVnhJYNTjPVLYTN6eo+iAkkHMTuxI1HcexUzfsAWUK+FkKTIxJb5THXeNQY1rPawvrItl/d0V
TMA+O7forndNIXdwRhI32906NkNM2Ys0dZw4iKmLZUweV96l643QEwNiQxSxq3C4FLDcWfXjS/3Z
Lc87SSUwv/nMJahB6Ux1K0gkGAR0UXP/l1fIKIICfRICh5kawyGUXAHsWnNZWqPM7x3m8IamGX6m
RCaTogs8adAEOkECyABtQiH0DGY6vvO0wI7SZGJfhh8cCnMEi02fWa3zvam9J1ocTT520mbrgT+b
5vdSmp/e64KTfnsYv9Fyy3stKhlogIO9m7u326SD6/yzwQJ1yEroaTTKfiMpNdpmGuMA3o898AHE
oeQImedRlQmZYidztL4EfZJE503gUe+wfPrJLMLGSyU5lQI6qA/wnwelUD61w068nHDAy5U+BvJb
8Fj439eCl8iAaYJjNYqqxh5Tk9ljvc4A+sBcr1dTtYbCPc5z3u7miyxpn4Xk8gCe7FAfv/Cj/UAb
NbzwAnRmTwC+7zBy+7OLF+v048nO3pTBPF1w3QK2+WjkOU0U6A9p/5jceSGBPqPJg/xd9DivHxDe
PzH7zBMl9KFmHDBgYUxJWc5gn2hGeqEoBo+5cm0Wc+q2xcABsevlrPUOSiNptEUkw8MU2PIzw8F9
hQCoNwqqOj/9BYT8o/NbgsUBOTjuugNV6YL1sdUTu9mATMlyfhtfIw0MMSbvZ54L682wZ7uhz+07
o2pGQve3Qt2Uel83cKcMiw9TxnQUeKVFha3Y5n5DBSq2Lb6NYPVRngxosgNGoiW5UJ3yMxvxG4sN
cBJ6+7LU26CdPJijW0TOPGtGZAbcpA0W6GdsTKMxvHBVJRokSN/r3jhL1nTbiK/jQFp5AAm9lhhg
6f2BT0BlG4/D3cq+zBpJaEMXix/xLUKhYb5/v/QsLW4NJMRguaNaWEKyCvkRnGPsVeJPUuS+2yUX
nUGJOSOOokM8Vn61jKpzRjnQCS1hnbU2ctfrIxzc1NflFABdX66mnr/3aukfkcZonGWO4FRAn8zm
Hf+zQ/17ZGKGXBzlXWO/7SLAgi1aiOwZXFm9Ayams/kcmiS5XFvW7qar8awDUO182/EHc7btT5AI
GKM9knO60AfL73gUaZ6ioE2Ja1FLHK/95+9Sf1v3FN4o3Gmeoyd7+ZHqrJxp7EA3zMLm2nARb5R3
FPfhJLBGm7jylSJPBG5wDjuW7S6WTR/j6MYIrieQD7RjXKtNPsnz0anejC0HPNCjQQkgpOxTjhe3
221d+sL6QGL3r9roZmQkTFzpUSNGVFh5Z/HZleNOoHia/eIkRp9gJw+QBWQXuYiCPxsWtLuvYDva
g2kkHjFaNjLJbUtWCv0YGM15ptnxk9h6r1YBTxFEMaS41ISyf+8A9MGi6hQD4mefD6YddihRclLi
1+4JOFI30H7dxl2i6FMoyhMXOAlclsUOpbuSH2D2FLXZKVK6g+AhPCegCdd9XTWaHg0+o7c0375J
fooQc6JSBThWnAi7FG1BIJLzDTNN23mapMMeZbKqWM7AUBE+aCbozMojkIz6iz4+XlyIbCrRLiN7
YeaAIWR+fP0EMPoUiYZyNM7Uc61G0v33jGwzuEGDI04j0nvlJSeBT/6qz9HZfLj3kLCbWFEY1rTT
8iLcOx+CCpbh7nPteC8GQzdDM/a5561e3ZFt/KUN4tNTUGwDEDJVo1VoCy5k0eaH1axoAgvx3I7A
IT4rdIgcHTu00yLPFd+3cE7e1Gbwo1pdMFBNh7ay2ZNEp5cIPncBUmaRLws3kZ9jdgk0dSXHgT7/
ATKiTdwuN9toA8zr3xvAbf6e/Wm0C8bFuuVIBiFExzpVV9f3j6bsGFemHCnelnOxUuBeUnpg/+Gy
vqMitmJKtfXHzKvOMCdMjedByE5C8zKWRLT6priRdUMTAvefzBCEUN63v86p463H6/PLisiKPrW3
74ECMYDtMKbrQDpDRp1MIJSO1rp0DWKQWKcqRAYusJMzDshA+2SMwT/gWg7acymm7pRuck/fYu6x
xzs3zdfU9cbsyPuGrSmfl73ejd0jNlKJeF9g5Bqz3fQccC5KcXzUPMbbmFKDhqiugYid95VzOEkK
G5VKRqLDGVSy/vieKrYENwnAwfDqlQfgzUKvKx/eDQQ2zOIipoUnc/eKYOzIg9zKlngqBbQxUGGg
8bnN7ZQd/WyZc5K936U/JWoI6FqpYuEbHGDB1wp+ZnUWwGlSa4amCNxgGKIjpVQ7dulI0kkkpN1J
KY26w3/aaCxvZU5AChleThAA6CgaIc9qyLb8Yk1KiMnwwVT3jW4YR8QMHCD+Pjwny21WOAqIGK8+
OUKuFvjaJvp5RBHVYJAMleWx32ZXXNhX4O0mjq63a2O/NkBLk3/Pn/cuhYUAVqKd+kxEkpHWdIJP
8TVkujlEeT8IhEA3You48PShYfi1Gp+rglwnLCvN2I63A93/LPSIadgqY8K81x8H8AhPvUltzP1R
GVH7wZ9TvqTxW9fPTeW4j9PpSmc9OtWZ5SsWFgSL/wuUP8je5IOvwTfkaSEq5O0CoM1o3sTpq5/D
ufrg2yRJedK0GU9UTfZ6w0o2pRDlBQeaRDQJRn+LWgKw+hIR4fk4RaHHR0oR4vxK1h9VIlfgQXFI
6UTV/DyZqR+aTxlEkFj9FvnCvQbHRcqtfa5FVvVYMSiSpNYleEG2so5+EBJwsfKEWWdOPf+ViThW
5Qx7ygMTqUAx/+vch9xgkzjdSgC87uVQFKYLS04PM1TqUUoPtWWxLZvytyimaqmCJjd0X2N/1y0S
ny39xpCsQ0bCOd26RHSg/iVCfYuX2W3ADPy0PdhWcmBOwR55HzTW3YP4jh0uup24bXlrqf+w3N0w
aizvGaJZeaPQPHNhS56wJu+fA7G791R40BrvnUgbs6yfQdIc0okKCyTunnCJ9vJFD6EIgSe+5fSV
9cLfIOPrbHz8qm4JUaExTQZyXNZb8f3KOycZX3YkBTa8CkxsRcY7SCwuNKDznXKTndRT5Xlx1/Sw
xChh0HfKLwkjW/x1Ab0hkw2DSlALStjvu1R3CO9zWLEaZDmnT2R4xFgkT9RGwf9kYc2DnUgxEDm8
Vkilo3cSMCf2TAdIDf0WdZRMoQznfJst7QnFZIBaSkuB3+iOYx/fg+g65ZfzSB/mVgMLFcOUVVQY
72TfjCBadoglLA8DR2d6rCE61c5IWd22hSGNQvKq4Yb8l+viUCkxn3HVXDMEkl1FBKrgY57gfpZ7
T0QRaly0A4UecboZzkF4y2B2zDmC2DYbn+9z/UKDtEVtqzQEmc/hjooQFYYNt8+WVdT0XJg0CHNg
ZzxtO02K/yM4hGheQoP5Mu0ggm2Uz7k+dvQ2XIwEnkUsByFGkDmwz0qpUfJYHPyP+W4W99/8KZvj
798EQhruKjeAJt0pO1/KC1SDdc9bSsKrdwGsL0Y3OSf9+sBm3ZIDBhi2+SaXwSJybOzobG4g/GFW
Twh6VAz0mBWxXF6UCV9lrhgUvd/e0AVYh33jET/S6D3ig9cKEVpFnEZOfDNoelT7wIT2ajTGkeeD
APVx3TrHmxuJAoOWE/YK1MdHichA4UJUTxvdt3KYatf2y16R0ORZO2A6URxRvy4ykU6UvBLZ2nrC
o0N0ZOKKn8mCLnn1HyxiVA4i8PSOSm6S1UED4h/0s221EhWy2v3bJkKsO3XIuEzzJgQ1WE3lKtED
Ja+eyb6GUbthhxlchK7hAHlVO4felexXA2slmWUxVlFq85QlRtGyCDeKZ2a0SQbeUDcqyTDQvt7A
gM0GGjPAJP2q3XoHwSviDgPUlFNAJuEKIU9BTXL2wOemiINAXiuh4R2q10pu8FiTII2NBFpclt4h
P8MUaIhBcGMFGGRkOI4oGFujBYbYvAf+YfuATw8/aifGJfqwjZKYi7tbV45W95ftSk6PQQ1j6GsQ
diZyaZ/hm91yP8eA8y8DL3403ReiVal/hW1EzXNXe1XC5kgDIdXERH7WV/PZ5LLHVztmUnZcNWPZ
L2WC5L1x9dlOwkCTzwuvMLKT1NQrqH09TzHsZgGf5XUJhzqv3NklAjVSR3tRBoKeFxNN219qGyRf
8DxEqc4eRYtxkwxZzSQFuXh8pftqjXWwgPyR+YGnEpeioP8r5EmafPFQiXP4oq4VVbnbOpJb0vJf
KVV7dAsTCNw+zpxoGWeo0ifmVJc6Np3ihLirfXtmHyHmkBhkEbPoXVInZDQcuqvGtSGwYjNLcoO+
ORVnTIsy28TjxWiWWvbQiz5DIYt4bzXLwHhNStBQs1grarSqc1FQs05mWNsQf8opF5W2qHnrDI3f
/sIolIgoOwCCHNcZNWIaC2lzxXw2Ch3uP8uFKrxwtZ4yRHaTVthQFzpeT0WcSG7y4DBrYtGdOZ3n
Kw0rtLX0SqtCVTeBiYqLWXEEDTByQJokKAcuxl5ve6tA80SGf/VREsfMLtF0I8eBHm8IpgPvbGVv
jgpehHGQ9lW9Tc0ec4YvXW/+r+UPWZMnjdUSgdVoXxFXRYQT22L+13iq5JXxV0h3OuIzW+P2RKwf
GDcMU/M/6e3ovTpprQpfc/ak3KKTdU2fUCOryDgwc6hme2YGmsTS9J1hhnSaLHXXp7sNDcPb4jrO
qS+Nuc2j8xN4ZBD+0gngRCbdc02iaKTfzYWnLOBTZwPF3YLf66yRFFUOwRHRFlVb9JrPSJTe0kUz
EbxWjb67lbFCRjd2S06dfmbH0kDdGGE1Wdhuk3pXoWvpUfczC9Q1L9SGUhoOpfC6VnEYg7tVJ7pA
M6WTTkVFDSg71SFC1kkVQKVT5QyleQwMojF2PgB3Ngibx3D/jRpbuMvRKUb7cYfhu0kgKy+WEH0D
Cav9oHvK8ritDhzYe4NqAmxK/xjyhYiD3z3Vhu6wo6qH+omHc0ucoUpxSLN4mmBEBk1+aSrEl9Bg
TNESZnXrWakRcg2XHVushYO4mrUivN1K/tB0mnBr6fGWF6+zkxqa07bNuG2oTQNJ6e2nDu2DRZNf
JjO2jMTIyN9I//iiyXRckc1KZywJqpCYkHDJqZcZEwYxeDalH8alcj24NKVxHEmRj1QO8jyMbMm8
MZQDbSa7VrOKoSDBKXqts3lt17QMsQo0gddCFZgA6y/yXc0naF3PCJzHHbgzBgWEFwYxdfH7841p
FiB7JB5MEICmbejIOHvYlG31+yJ4idNlgkCpVSQKvEPECZ2OHzNQgvdP0dFxocdKTMJ+XVI0go2N
TxwJrXcavqm9THUOZjYExYlrOdY+dWTWTewlgB++tBypo9hilMC1s03zAuCg2tq8r5oI9XgJHfGP
y9Viytud2gxI2vdoRNIpNegeeXqcTP+QXwwxllT7tBI3r8nAx7wGmFdNGoW1G76rTUUVoNr6zT6R
sYyHDDyXFpXHkNpe8i7rtcnATPma+jpZW1Y3Ay8S4kC/+8kMKZb0MmxFZma0WQNtn8KjpCq6J1mj
jLOeoNC8wJVut9NAmkvfOA0jE2BaVNzp7SDDgeD6hEVS+V04kyHpXwznzEjoh4DOa6gC2poBmTqU
2dtgMw5xPYzKb5/rwtdZ9ttvN088RNIg8hQHAcM3RPfXYY6lecLj8jjxmk7Tabfa9h/OC4butjwY
qmBKPz5SvMa/avAS81IERj0hEre+Le595HJhgrMjCgKQxw+NNU9rvSt1LhQxddJRM38kSbg4muPB
kwQu6R8UMb1EFOuo4vfYkrvWrllGRZ1tf1yg1JJYkptH9Xopw1t2VpqwCUGjCEO/c+8YMqESgnh/
5lpsYvm9Qq2p8d1MwqPGAdF81eFMwYPQWW9fh61It0hCa1ADEhJu0ktH7v7depxC98K3rhqcKSgy
XorZBGRdVu/g2EeQml19V+9DUOiYnmFW3/p7Q1xYwCdzeS36eKK9bFIgR8/8F4WT455DdSjQSlSw
J2AuItqmTrvdyH1lP9b3LJ83q1Gww6PCQK7Gu67aUdg3smQ1IxoIK7d0zVIC+j0ZwfeshmNZ9IS6
xI1YpeXjkyx8yG/3QTVxQ3mzeW6Uy1CDc3AZTsQWO7L33jkYLvFLoY8BXJEBu50QrhWNBTIyGG8G
OkHe551q+HLhzf+bywts8aW1sA4eViA06KtT3buqmS6XXaFSncBlD0xGgh5zwvsatDHUG3FfufMJ
P14Y+Nv638ePYyBVYuKG5OR5L/HOs57M+wMtwG4h2nY9Bj0khHdYKiT7pN0rdgrrhTyawkJrfcDw
jf/5Ib3FRMzHMtGjnwC+RNy10FTom5TW2UDAUPPfF/4o05rmbvyRKXclDij3ZTxDr2o0ldeioDvt
kQvXr5qmP6ABO9aF7kEGA12w1TXjjY2A18CLd6nVRZDAZUm6gxS6aiKLrMqr/iw93iiqpzZe1pBy
xFyvFTHxuARCZlnjmUx7tF2obikw/SrYEoBGsciHMMCdV9MqMo2c+pSk1UbLi2ewgIMXgIHhkc6g
AyFu+RTsAALi/QyhMaLirodOK2oSr3KIWoEtvWOKYrt0hg9NUyARhpums23iJ9nsslmCR/zSSbZZ
Q26R0h0fRrUhPP85TNNw4eSNLfQSHra0uMbMigXL92Jri2BQgau5OtWiTUXjTq3zxwdPM2Hy4f2Y
H8IDZz3sZbCOu3Ai8vO9/VMrAJVRxEVNZ3F7GVv0wvXtj0IPUtABZalK/QtKYLvg0q40+TPEWIfn
JM5lwA1JVdaXLKCE+nCaEkRNCrGBGliQBzl6ANSgRgwNW4OhIgHtKB2mI5RI4O6GjGXQ468BISv4
AVbCUHpHn+v+8WksdNLtXidaKJA98B/YBdOx1rRp7c8BlpzPnstSSZOqEYefFnAO5LRpdv4zoBIj
OfnDUHGcNu4Ic34Dld31Dr9rhSJVH7rN36juii7Q5FSB9vJlPMNAF+8jDXZFLxI6KKvsl178qfAf
u77eKXqomfos10nkbc7nNCfyYVYOsNwHgvc5D98oXLHUx1MQ9y0S6Ir5vVtg2pqlhoQgKhyqrojj
1RLd+Rt/KC07IFle0T7BIfjxcCog+mF6cEiQS96OFauOJFTm7e+Z28rUPbofrM+LMe65W7IE/Y1R
Zq5RhevL8Wi70+RRiJeyLPRMSrhOUmcmClRv3gRNp29v4k8G7L+MwnLr1v1GYo+WLqdL84RObEtF
Wy29QFfGcXqukojsEdzhi9b9E21P/k49hHAbPt4kFJK/KDkLbIg8X8/l6kZUqzwLg3MDH2CfS7YE
4i6qrN+DjK+sudNeHzacstLKrhVKgh9OcjV8IDRlxdKRTQXvOHdMiTbUifU1Nq3Fajo0eoOg97Gk
LgXx3QAyeiXZAr2F7J8MSTJXwbf9KYxhCRe+/vAjyp1OAcaUtZhctUj4wGhcrl97q2IHOUr54EOb
yhWcm4h5TDnAQ7NgxdhNnrfHWhu2myNjo/Aj8e0C1VVQWHe5wbNweB2J+oMuGoOcgrsdBu1EuDn/
pJzCPR/x13gcZU+XFAxpoSWVIsxsHKqZhpyD/I1+wwa3g/QW88QqqQCpyOkaszLAu5vtp6acgmbe
QcJrLXDhmnAdWPaJ2V98BPcamKekwYU5HMvNedtu8jr9d8EKa0jWC55OZsBcjrWaQ3yLiZ6lGa6j
mBGO/Q8okxSW21Hkk5jPN7RiTd1KUty/DLAHsqyNVN7+mq1m5QaAQapBXbxUTYIwbwZZR8w8CPCX
y0Bb26M0pzZ7fwhn2j/H4Jif30I5fe0ekbbA1V8kCBd6jKZ7BOJzFaTxPqQI6TZE00BoVRarAAs+
FywQLvGdRWRRmA2PW05+IzFCQf3DreOleKmOK1oQFNG5IoqpfhIk6tJdwnjMb6QaI+yRGnJkeVrP
PT5/wA2mWE6zxk4sc2RVgrkzQCzrsm0zMmeeq8TO8XraON8zlgF5MpCJzYI91cmdGNpdAkmX139v
XaIlCv/Fdy1ehx9lSXNZAj4EKuhGmQSxFQwdXi5skVYnbg6xzULTZM5pw8odOtu6JGbc1JGJL6Xf
DoUaLfEdEJAcWd0frLYPpMYDsAgSbegK2u/VbXdLTtaalv9vtMVbxnHJTcI48zzssjdqSPkF/i4l
Y0fivHMCUUrefHqiFVgppYIIXwGksBjAGkpU+RBNFrrNgXL9B0CJtwJjoMpaXjE96Or4XH5EVqiF
Q6N6fjVjeP6JrgGJOS+EVIQ6QOJxyrEPAT+9rRpgQI2w62nE+HP7yQaIPp5hwXn8EtV8QerjfTK1
FzU0j2WbdGcBR3elc6cvmW1h+9EkBF4PsQQIY1cFpAaCDUMB4e8XLpCwzNjJp8MBz4ROPUTTr40y
DQ+vLcjwyYILYxmHNnjcyIXDZtENxTXZl2ae68Erwdgn1bgoql6s/DW5MSHEhmz8eW0vK8XEm5HZ
Eoif/0HzIaMJqZdRuPP5Qg0v7J23FezRwKH+Jh+fdpjdALJjQQ3KjR80F2PPgUUHWtOZICUN07so
Chk81G4IKyr5k8Xhpf9uoffc+tR1oNCS9inGHsrz62LpDHXMMyG7B2clSKiFl3xPfJ5vLXjo7U38
1wcQ2bv2CxHg0sn/l3ShYLU6t+lYjwmIOSFe3gzjlSiMxYBN6ZV9//TJqb/R20Yt8gvBKhKcQefi
a94UojLoBIqlO8exfTrXVo7VF6KlJbtgPiZmKVU/rcvMEL6wQlcv5bkfzVhk8/ISSc4SvzLOM4y2
kdstFzswBeRkcIc8wVP3lwtq9gE3ps+dKF/ubeka5rjrXHr7s0v5ofjOqUM8zaxGi2gXx4tPE3FB
dn9+DOQvab44KcC/V1gBHByy0FAWNkrj6tKh0v38L2ia8YX7RNzt227YYqO0XqnhZ5iXIpYMhorX
tvfnpKhsnwBEBH6/wObBaMsadoKaTs6HTBw7Z6htN1M0J+eb1PkoUGXEMjlNkhULZ61Blquq8k1U
WufCXEihFTe50FdA1W/uQOM5HuT1YGC/SRbnmpxYPdGJwhqclRMW7q2Gs+8Yhx5W+ETlmV6fbNY5
sV5eOidH3JrCH4u+aByXl1H9kb0q+l66tJQ8lVorTK6ySYAqMtbwDA7639T9TGCG77IF1id3qT88
X5D8FoWASkV1/YAv2rl29p/U4URzitw4znsPSW7UoBpgPEHBgoaSKdT9ZFK59Nu7e8qyF1SH4jD5
oKICp/Kcdcwmmvw6ahwgKJItKfEYirDCUHh7JxvC+bqdZ2zHPmW+pz8yc0f3VQDcn67LPXB1d+2M
5vVBnQL4B660b3jTDB3L4wFFTId+PEmlZ/i5VAKYVUCkxEhMpx5wJgO9gRWWmB+E/LxnXccGd6YG
HfoCLIZ/fUaDslYAFr0aK29UJ5YeGFg9uNpEInzaO1VKu2OXpz4t9b3qLLA5g0dW+wpsIZhY3aw5
WlZKc0ltJ36PXMIKNnynt0nIGFfwLOJNfwBRzWjGh+fQnxYn9zsY4Y9Jy68iz8hddfhEtQYZSs01
DSbVR7fAMc4EUzOtiGEUpcHTuo5qel5Mhr0tjGYYiC2ocMqmy8O1+C4MFnpGp2fVGISB50SSiNgq
z+YDYBF0waQLHnGEdXlU0CYNyfCD7w+/jQkk0ivV1iOdg4dMk1zIJLM+fUo/NmJwtBjaqaA8bRTO
Irk4Roq7404r++N2ZnvJziJhGOygromj4SM/8dyWbur+oA1fnO1pkqhJ+FrhaseZbVTQpvYXtMrn
PtxEGZ8N+AlNdENQOwQEePcU8vRxxLoXkCquxm7WGWT64f3FTB3PxPxfrl2MUSEsGz45CJQuwW/q
o9SSfUGDBX9AM3IyIV2bGnLoOR4L3ldX87WkpJd/lhbkMy3G++OcWO013xxMgEh2PjJ5ottGM6CN
hiLlruZMXnGusLG207xW/vp1+wPKVujpvtyZ87NZWawvepXiUzJPpmEDVdZxW0JUo1yTXtZXlrz8
2wkniJ5lGYOTKlEog0taS6Ec5ooF9iYkYLSCIesGBQEX3jQ9d07z+8gyJJGX0cw88GJ4p35oUVXK
4HVTTbkjyojH2eSn/1EeZLDH+dGCpt68Ax6QMJCGmrqIXAqc5BGGyONWIQ8bRQY4uxATD2UEpdoY
qPYGeZ2RTR9U+j9v10Y+RkxzSjVb/GeXRsrRhleelLS0qXU/y9GNBBHgJM74NSqquCbv8WE/+Z+R
XiRVQqeRdNqr1ysE940CIbLx4SJtD/vL5tyuR+gnT49HzAEcEA4CJzzQU0IqSAxBfIa/2Ctg1s6e
D5u2Bj1wnj/A4Oze+NX+itrvb55g80SKjNM8DQ4hMoprlHnQFg9ERIMjMSxiZmoAtpLXK6zwC1gc
9xbMlbftLHQJk97w4ahVKUZcwR9A2wjq2xwxELVHwfjxeZDJGJ8rHJ9QcqwNYZKulcBTsbE5DKmI
jgTNqYOYUaDhqmZs9ivwaXFjkT2/v38wbcGug4B/LInzCEUU1H7X4NwIDeebB29/kOBOl95ak6Id
0nXe414vLM/ZPaCLMCFsjZcsWIvIj3jIbgPpJyoOel3x9oSgxUXIXNw+C3kUbT7aJmKYbDtN/aeU
TRqxrl8NAfSTdNoSu0BOBgagelGgVvNqzyq3CFKDnsb1EYW6gHaVCGfLqXLNB7E+W6LXSmNtuG2c
CT/Dm1QnwB8ciKhr3p5soXJk4UcN2bcGNfFiFTEzOIxMz/LhOXAurdCZqWcbKCcflNny4ZnhE/uN
yqucpkEh/LFZ7uk6VxxZVOwiE7fs8zyyGyLGC2chdia34Luo58p1bl9vBnpPlbkroQr/ZETBGP9Y
+MRNFyUBKRgUPJoH21VkiV1Zmov+LTdXmjvQTXNly2dejBUbYYhgP9a51OoAiuRsxux4nOdPRkWn
Rhu3ascenQxYnijSz3qEk8GAjbVsAW5juClag2yN8Agm5kJMJZ/X7tg2+hCeb0zAzGvMKUSFQ5HI
DoRB6FNqYG8l6JU2YGLVuxB9AzEZ7zi5zxqYvl1mqat0ZmQD5fs1241PnbU8u0QhAntJZz1A063f
XvRIuzumgopEwMtpDnquEEtH8s50YjG0/B/gwCpUVyBIDJNGXsevK5NprZE5sMVLBJv9N1HDoM8y
iB2h0MhiN0A8RN5PDHc1INi5u6YST7LVwIqTD7DoFQZw1RDwM7kGRjM+tTBRb56TrxCTb+BdByV2
sPuktvkaWAYjIGV+radVnlMG056p7bPAaEYWI0Z2VnwVB5Xfe9hI2tTk48kpUCyJONaPBtNyOojF
Rx5ySn5V6CpifRQbyyjDx4u7Lnzm8byvBJI9A0OHNwlxRCZNUOonQArsE5Z5J4tKAdGnNhXMIRZ+
Mm+1YqScoaDIr8sSGC1J4ZuAU5S2r1U+gqLAcxuCL+VNWqQp61DQ8C0CbWskz72oITfQcs1yf3y4
SboFeQ6pWD4c3yK1ZN8GZK1egEjy7nR76C4kkbfMMQILMGQ3lYXBBJQwas3Z54zvtceVdB4Z9gs4
k4Q4k3LcOguDWlXWi1/kakV1qYp3cTz+ZXNPJRQomNjtWeU13CPTwj8TL64pPPMyoKRJwLD+Bvfj
SHXun0RsbtJXSRRF3njZiQSvzQ/QcyCoYHUo8cCOBN2wFE7NamF9WOuGca/iCYB9H8EYQ0exjSVz
6guNy7T6gYM41tBAdiLGEQX34D77HwKHMYg8dgJAFCeW5VV0ObKR28NP6FVsA+VGqsXqGxYM+v3e
1ssyfhBVMQIbZ/iZdNX+SNec1dFiDLwIVWJ8MQ/cjfVveLfJAviJ1NAz5RU+CbNTug2tQ0/Hfxw7
/cGTg0oJhxSr0f7ZnzWKutGkhL4XL+NYgtRpBnnTilUk+cfX99jpCboR7WpBv/tf0n5+bZ0bgLA1
sMeG8Unc3vri+RYEvID7b+Aei0UEkW1ZZq8XCBYZNu6YUItcMQ7nGS8921gIfVFnHp4ELrbUCux2
m4//fYVvGA5P4Fmzq4oDbRcmoU71ujgP6XmmobKcQM9VyBqarbjLaByCWjzkNPxVqK36TLXNuQ1M
Jv7l+voW6EgNHR7znYAnbWOqm9cNBfTzgSoB2KT9cI0MEH9ra85gKLIu63fl5xXEhG9KnGjIEUwe
gwe9Lyogfk6ixa4liQtP7wlS6svTuTH8cl6GyQKcesFPsZRs4xk1Hgf3xz1CZLoCy9oNMXJYfSNN
OBvDOMl6NeeeEmaT4RORekgIuwAMkzLyT7qv9B1ofnb7f7HpZ9A41mMnsKMqne9tXTXwN4Hu29Il
735bQ0sF1Omb0XTa1hL1rMUDkbcIgyrFqc9av94Gz911elKEf1OUay+w0kmXMXG/fpM8PYWLJ1ZT
KmsgLg9hXuLKg3b7rGsifeaFjzwOdauHiJwP8odaqzqvz7dpCO84cx70ISS5XOg11INCm00ctG9d
/f7rrGpmTZ0EMF9c/JPI81AtNI6/grCtHRAbspiU9Z0eImas4RiF2TakgmQIKTKA0SuWOHbpeQ74
BwSlQW2fwDIF32PIdTzPPM1WYiPFR6as1zffPRRFM0IJlXOPIsvaQgm5wZGQCA8zZOuyZQENl6mx
xN1HoqpCwAVYzSTOIRg37rvXcPtC7Q7qlX76Vw3E63nMf5TZFXyl5/wOVWTp9+IYAm/SIiTGFHqC
Sjx5HpOmOL39KvJTFzD9lwOiXwFj8r7ukzsrzjzZlQlyeG1+j0epM4/fcRXMSXpa4PddYtgu1B6w
G9I1MmmUgdk8yMxf5vRmeJupneVyBUgtUBULvrRHqhAOS7zJRlTcdNa26ylrTZcItVsDuVf65TFI
QjjoinBcpdI1cIeLNjy9oNt0ivROEDkUipLXxL0FKHAlJq3OVW7IUAeQEUp9WoennnvJka0F62Xn
WCmmRpcf813FshWLeJtjwG/tiKajpFw88WnWr6qqkymkkt+hu4tpwmiE7bfSxZC+oTypb5uKtKh5
PEtFk+QQ5aBomkA37+mUs4ezYtcIZ2/XFpGEMGgaF5pynBp/FwW10pdIeJqV058Kh7V6je8CpCzj
2g7MW2wBMMOTO/QL2zSKNg6Ju2fZeTxcPmcKU8jCyehz4qiQ6CbDFIZfaqgziOVpfpwmmPGhsukZ
7Jkmt4rPBI17yPsPKQ7x4LFcV3yB9HwhqCXHAVajgyR1BeMNFpZKR77v0qr3byxIE2ZPOKtXIvn+
/d1JE11qXe8tiB5SVufzi/s8qz6OtPuj65i6xteAC/ZR+G8xpm2jEATi3BYTkIEytisFgBVpnh4o
s/JMluo2NVKmUXwGg0zIYr7M6A9gBaQW9tAIAAoRuReA26vGhhFjGbFR1Ly99L3BFvP1wvK050lo
LMAdzAqKfSFrqW4uJ+bcrTjQioHZR/Gpjw90/1bHQZAkWfP3Q5W6k8U1qPbUzTuAP6pbCDGSJWlb
YeZjW/9TnTvGS4zd6sFUCiYui0/PvzKK7s4E+ZZqZ1jw7c7lweoKaQ3F9o/lkJtPB19phdOna+SE
8hmE2p8cikZ436TmeOH658wxFjSZVKVOzdFFLYTJ9Qx7kj1vHSdX1zljkoVwiwRghgz4k2UaOhdr
uTPgIB7hJe3WFwEaqAgaexr/OXKh15lWLrluE4Oz4BKLZhq7nEEXy25QUOSji8e0WLcEZcOu7aeG
bUGwq0QkNNx3QGFca317ynacVr52Hx4PYQbDiTyL9PHmcfkR8zCLsTluw1zrCtxAbpv00grqXtz7
EIkviCQAS3RtkNsLwcs5jLOjMaE1oB1ORD60w0/ncY0WCI4i9wQ3oIsmfDjfo0AFBs/UaQ0DOWnT
uSU7RA4Euq75Nxu/m6k6nzs2I5s0qSRNAmkBJI73fjslEBtPAwnNfBl/hg/tZ5iuNQAo41V6yDbp
XViDCb17H2WykwT+yU+J0mhcrzxaCNOVblrjF1Zk0rm6QkoMCzw8XM1Dpld+eXOPQ5Fc4IonMB+L
eS20GVxyU1r58TxW/9zF/0bcwF9OSzqyRvzoA89kAuGwbcC3T2E7tjsLudhJ9wUlnkwARJW1JIr+
oCEIIwdC+SIXRlqmXT8u5wpdWdXtX4ef1C0bRndgc0Rwh8k7+kpKz2mecjU1XOZdvQONIOCgEBNk
f+7KRCY6swryXjsLNfBcyI5sSVe0k674EybF78DcfXR069/F76iaRdxDuM4O+TjDDxbi3V5wqdTI
ngwye2F6Im0WixnoAOAuGBKD860Uh0Vg2VtnUoTp6dXuR/D9k9uXGMq0Zwwn09XIeTJylaKERkqe
G1/XQcyNV0XYV0zH0dL8tlf2oPKt+fT2FJSIvotXHcyH+KKeM3P0fiYwKOPE2/qBdFczgDyeIXIE
dkCNRRYv1ClZcpEoyRZFeRP5m+OKjwfgDFEv2UzfssNTHos/k9eKBhs0HJbQtFJMvacAIA+FxMTC
fvce9rM9nHIzOKr4lhoZ5RJVQog3ikudilV1paM54H5yLj3RxH5LG40duJyKuBXtWRDH0twYIbWc
GBacAB1LEFMADOXxOsu8e3JiG35er60cZWSd/hYBqABXS2KFisqRIDAj4+drse21XeE3M9xZw73g
USghbUfaHwqWK1TNcW3BG786WXMl2NClfTOWoFB9N7eutyGOB+pqbaLS6m61VXUnE/QQ5RNyFw1t
nOMST/IXmHs6OkNd52a6I7EuWsvOG2z3iDU5JZKPIrHtiswRUiC3OEiNNZgOIsSlTa2UgfcV/SOV
ztXi4ONLH8Dz88TVsG/LpTqlct9njuzlHQZeYMLJSbfZKnkuK/Gr3ovlvMo+2frzFomVKw0LltM7
6GqGsTGzLxKKvLx6RjI0RcVF/gR/tHVburncuVig29g8lHqy7dcjvEO/UcEkoXvuHsX5MvwkDdmq
1huhOvRQqakQnYb4BM+HKe1opBPy8Iq1bSTMa3IhpXpRdy5s9IyuYDGaPAVVFEQl5oifM3FEDfOd
4zB4zdiyTsr9u3B5YZUPTSW07mUoPX2M5/xoVVjcgseBVUJeQPrL4Px/oUx13qOEs1UC7mggfNim
hM5Sjn/CA97RfW6W06r93DEd/7bQIYfIgrccgXGnLtHA0PxKuDi02Q5ScRtmPsOwyN3f+ob6Q8dH
Foe0iihX5SB/E+lUZeiK8f8E0H4wFuk5BQ8EeVkesTdKMoDveHJyvUiLzrfC8XT2e3CoG0dgAVIi
zUuy3vJEJkYjo9Z/a1nvXxatm2hZVTHS/SDrmYsH+qpbdZImEyvkQ/aYXQg0U5jkaF4gnsiyUlXN
PFQMlU2ZFhd323C5UtJl7r5IeC320xwlHEwEomoNPWdVZFFz/1359Xy3vekiA+Hzkatiiie2TOLZ
L1Q2Zxjj7vbpUtIA/oT1oc56m8u7+PLqMym/qJ9zP8BUY4L1bsFe3yADh4yEqeIlm5x+S3Str1Il
PssUmC1Qu4nlXfLoKqm6XGAY5ahZg1AuUT000//kGRLWePBwpJUKv2XqKPYdiFyHvuebXJYuZ9E0
iB5v1f2NKaJSrSLov7yTm4eptA1GuLJMJyHScEs37b8kI1X2n51Q3YNdA0+JLxMhh4gHytIBlgJB
KCsIwHS4syukEHOE8h2DbYaa+0QICiMhaqLKU3mYqf0NcV6VYlumyKKRjA/rfwRbdN7x5LExLqIB
oQrd4zrGYQ3WtZNLCOiesHYcAmCwKhrFS+iKhh8xK42BbAyWkjmZrbwaZvW83HzSDwqFTt7mOvRa
33MrB1+ZI6LmOhrNf+CykAklzytXNa9CJROlsWFo+DbEwV+UnACLSNH9aN6ujBHIsYXVzdwW7aBX
U1l4CrE0cbo5s+gEttqkeXdbv9Nb9RrjLAFIBKOzSebA/Zh6Xt4oSTyFGf5r4Cayy3y+dovIxzpi
/VLIb2bKoALbwhIAByg6lrcZ2mNebFA/8aDQ4HOafeDg8Sk6K65QxgndiQ2CqUqZhGUIFoXIxFlZ
btrDlgYnvwONHAj0V4SpiFOkak6Izu0ZRF8GfihlmOvs6xgN/eUQpGeamxEsbBOGrXdHtuQP26Sr
DrqBRk+C0zRDowGMvaWg0cSXJuPUlPBda9uVMwGSGKR76m9LYtI73mEJs5lKbujtDG4t5B+ymYgB
f8IvAmiPO1ftDzmjP7f0nQJsg1DAFj1Br2rkSZjbW+FCfnBGvlWOy3Q1IrcS9b8PidRmAukRQKp5
F39UlYzQ8fTJJfl5vjQtHvcIrTab8NB4TSR91uoPYEeJ0ZIS35SyznL1QvKQTotb7en8CuSIfVHe
cBLCUP8+xG1pUrosyIeB1PLJSGMDZ+RTyIDfmKHHA1THpSLjmWPp2majBDdK/rP38cFJMudvadYh
+nG3vlcw/gh4bNyN+uSB6wdbzjy0uIGuKJHqxm701dR3+YVx+wgqBzPIXkDSryLJfMM71kCbUiNq
5oX3ONGrFwZX2KK016aUKyiywJxD6pujrYd2QtP/Sc7aSs8WR8psIrEzirYh3IOH1gOD2UYCZP1x
4KI7c2T6o5M3ZZ75ZmXG8u2dG7qke9nMTIiGiLfAH2Aww2MPczvEBztrzuORWkzDWsEbS1HtFUV9
OqnHNlS+NSKIKEFSEcgt9tUoMjQ26pXObSfuAa1unXURAoXUzL+xsvihYxpwdX9YJR4Fak7LV7r9
7ibg0hWs4lvRV+YUHQSom+DYqo+NvHXUUtDk2ln24a0WLEUQf886lSgZ3U3zjek0szHW5cGHi/Ij
fN/CNXbV/LMsMZ5Eaq2vBkIiuoFky40H0iSBpIwMgD9y6NTftvAqWRsYcKMuX15/Jhhx7wYzz7Sh
QtVkqt8Dq69ny/Sci9sm8jPxYkRvJMAbT90rbC6gEGmzmrkvl20L9VwFnYM06V0lDG1PzZBEpZLB
TEJz9xjc+Ulz1n9s1qE+d0I0WanrESoC3HgI6aZvN3+FAt6SrB9oP9lIoKV/c82Ku4DapBGaOOcc
qYlFu+vb1x/3juAd25yrn3zLpckeiwU4mV7PIote23OUHMB0eHuQVJr5lp5awxwI24YIE1njke4l
mfiBi61eJcN4DX0KG+/dnN7TTq7fOXAZfl8v8VBUoKRdSL0qdSuDKcSzjP5tk/2YPwVcLTpd63na
xfKNkKOJHT35siIqwGVVbOU0uyXGPIV1ZkSJbODqSE3v7XXLRJIZP6YtI82waUcwqBzEaDE0NmTv
ESTO4z3YwFgO09hGsI1yvKV5UQwPaujEnMRAmWcej1tjDTENKhWQvI+wbZxfWq2QRxhzuNg2Bzlm
nE9N8J5fKnIhEemDV5KINUxqnuvDRDf5plM8mo0St6fdWHGeyzhs8CcECPzRwXlyRpFYsQL2ZKhQ
TnpqdZCoGr5EQCqk6WppsbQHolrTmWxpaSS4T0oKgOzjwD5NI2bhly0auGXnX+qjpfrY5L2gYYfX
4LpaV2KfB/JbpwgrdpX6Oguz/rOx2an5M50tGhBa6pjIXVPEi4lZcCDls8nf4+9zlynVq0Wb6gyi
vSeJQ5Lz6vkCPx3S4wfq11VN8wAnUtBrqc1gjdIwpgSW4dHlTDICixIAfXWyQwfCjPvItpV01shT
gJdOTIwqUqZOZajO76FcqQRzorT3S4+ZsXa/ToxUr0dVuakN6SQZHMin7exDUqAADbgZkNl8l77d
WZ0/Yh0G0TMviJvwqSAvZPeTcbuTV4eIBNowVVZHWJpWbzOJ1SwKiBZM1hEy1k0Jcy2yirEB2+HJ
gjTqwr68eoGwiqHcJCk5gPSW3qQm0rtzUrUZXXWlh5J+MJPA5SNXQkJUX9bncUrT6jlxSK/iAKLc
+JSFBqAPflBXGhWZ3xg/hK7m5KQOmAN91D03MfdZftZ5ZdSZMCp5I7emnPNhCNW9ZsHFJCCvXlUi
Fz0Sq2bMtWJRc813jdv/dd4RbsuXFik7GbncjK9sVHntdJ0Cu2hR9W8QWKDiIP6VrjuBXv1FAMYh
+C4JT5x25qlRxcyEq0liveO7ef/0F58Lw8avhueiNL1o4SNHYnVsYv2TkNYcIyoYQGWDT5jLwCPs
+PDPM0xlrVUyP4fZru907IVtTboDyHXKcetrFgmtwdZVoFC/jkvWyGvd0uc8DNzGmDt4yDnJFpgo
eIq0patpyVqeeVsUURjFYdmtgOjTp0so+psoQLcRPZxnhwJXR3LSHpYXy7OjSxTZHJ6yPp+FbdBn
I10Y5287eF1QFsxAxp/lEcXepTTLwRNzYeQEK70RlcbNN6Hus/nn0SrNxdbMw5PeYNr+yR8ia6KC
F0JaYa8Cod1RurZmR6sBwAKnoyOIxUeQlaaLhS/IDLQ1eyfMvc20Qpyx/aKHpnMOGM8UJABlKX2Y
/VcTK4v2u+jFQvCL5NhpRMZLyerOJCGBsWOlvytShvKmuwsT1Hqhu/no/d5ijzt6PrnDDutUfEze
5SmtN42PVRLZ/gADZs/qmES/GR3w+pUSbBVOevMTCXqCzzq176qpDnPF40hiur9pCYxJncLUmam3
COCWUG9jupIzhKC9uPDNQC7vZKEh6k5jyixYrSNHHgCjwy0F/aBN94BZvtHVgSU7gl2WBcFqyr4e
WUtF3J1MYFxxBzTGCH+oSaNmkw6KQj9M3pg1XcIjv4xZkzNM5/NRA37AXP4tZ5atW6yHhgBdeMGC
cKe/lIGg5UoN/V8ZCIfIe3DCD3S6v1qTviowvoUvK926rv3upnmL3SIgI6VJaDGPGSF4O+Nzc6iz
Xa3yQjf5Fy1HDRiB6h+nKCkVrKY3z6tTTvGtGuVSUszz4jUnrKvXXGgQEu5HpwWVIoFRtf3LfF51
2jZPp+w99qjJqMWUSqlNjuG0ciJvbs5Fn0JE6H3Oh+JnQ2hlHES7W04yh73ake+Ra0Ix6hawdk3X
lACPPiCS+mD9fwEN8A5Vzq5eYzj51abUEkEYgqJQ1EUtMEpFBjfvy6sQH0qloLqZvmjZhUkD2O59
bdEVXtv3TDfbMlPF9LvQzmkPL+mEMAO+V54gHnsnbc426Yz5x0XFE8pA52QUoiu6u9SC/j+RIAL4
JqKNeVWCWCGfPUooPMnRsD2Ax8DRKQ3WbNSp/GSxyXfzGx838ju4Aocbdtc/aDC3FPrAcg6Gbm8D
WrtxaX2C3jn4O5ccQe4doQKLg9HrhqA5AQBB9kKsehGW1TKnOxeVbL0FH0UQUoK+Kl8t9LXQT715
dAS56Kw/q6WQ1/AwHi7rtKWOV9D8taZ7lPhSIJZgLqP+o3LTL4dMhCByZLD0jlxvmH+vuVJWmKnP
fPaQ5QG4Q1N+AYKsYN8HLNYpkNmz7Ff5kHqUIju1pTQtcb0XCPiDw7yh2zk3yb1RZ96uhJAqEXgT
m9KhCEdPyOlAV8pK8bi0GQs5ve9hsZ0aXn56OlsU7WFKX15fJco2KOOAZQJiPCefuqUGwmLy1c5Y
UE/Ov+g3xlpnBQePJIMVdSQONmfAMWLHjQXftykVvUBnahDq2eBKurYPhIVJ8gWOytIscT0qwJwG
6/TTDtWMBikBNWyPT1PMXMp8p/PrW8OFul5qVbGQDTwV0lM7HOEI8eXbq9GLLhAfH8D8AKWz/z1Y
+RxzTz1aXx61tp12ZW+DaEZ5JSWrKvtT96zxL68QnQcHzJqu+l1vawlAr7U9ynKwiuJ3vjG0AToF
Lz9PlRatPC9QWyNrdi5LpBn9UodJ52JlMCY/AAJLgB0x4nGNW0DmgCykXtm/QeHgXrw2bg9V56H7
uRMLBj6YxtGx49+VsJH4mIcLsHK5FjI82qf3tvEN/NLteYabbSBHYaIQGJGzoma8PaDIcVndDkAr
6r6C6MOdNy3CTkWgBmQjVKGBKxnhjXMxoO7skqltO0En6brJP383k/Kri9I16OfRcD5ka0TrQqKE
oXN4CXaGY+QmUgTW7bKxEBFcVJJlQKuD4i3gh80mmSnC1wGc9HEaRxour1D7PiCoAkZNxL9XXrwg
aGOaiOZb4fgmR5vETWU02/YFFnhP6LrU9Hsv7j/onosoVo5VvuBHdar2+S0pZqp6DYYHGcpCHtq6
Q3t70eO4JC1VwjAN/kzd0b+58T8x9FcuL7Zt3IQVK+IOGDDm5obfu9RmvUrhnokZAbFduwL9QVSE
NGqAxIR+2cHJAnr6cMwM25vm49n6L9OshOYKc5OHVULbu+3zVv58RiOE+YrOpeCNXds1zf35+7bI
lokXct1uAEHWKQVAtgz8K1XVJrKykv0C8TCF8zJ+7zvqZaT2goXP/i7rg4SPVd0nWxk4ZZHc/IOV
+V0cCPArUfBZBUgaLRzUkjNdqy9HdxTs6gOmS7ozsQxfW+f3D1vOpS4IdASstpR7j/TcNp8Lw6xt
xcC843Z1LCiReHFUCg6HOmy1bLPCJxKbI2YE7gdgXAbtW8RHuOLJR+GyVEuRipnzhqcj9UWemwgA
sCm2qYfZROUGoSk3i0u4v+4O0TGfguOIj+XNvW+4j4xJJZywm5A0RK950yFe9ezmft4itfeBAK/s
UxDtp1+qqkjR2OhQQG8PmYYL1bXSW/m4Q7V9X5WPP8vuPzB2B6G9nvPd9nrhHBTe34EMhoU2EjZz
FhTPW0YqTfdDo9uiViId1pbpsub2x8WS82IFDJ8llMetAoshaGSCQO2LroBfBGdI8StqsTEarGe0
QIQ9CbWgH5AXO64R46B/auWix2tokK8F3Ky9D31/3mq7QijXE8Io88tZOWkdVQTpjQkNgZv0hHHA
/VwK13NQ4gQjhxe61jf6hugtLPHcC6aVek0T78Ki/GvRHs6V7qVjd0B+hvDSb5CNzkIqxqhi5EyG
nWfHnw0GGEq+8qxM+PxEdVS6aQ6nYKeyzkrbPF212Tft6z6fN0UIpyEL9OmwKdhQu/RQYZjlHFep
O65Nr3xTcD1h9XN1XQdW4XVxC2riTAoRY9QPop2uNoWHMRy0f1XLqfjykWat5OVi8YD4NbXsyf5Y
1p9AKbZ6taSmmdjMl5fr+RayVk+PRr78zXN3hP5L0vgQItUrjEVgMhxoS9sDwINKIiQsvP5ZbZuH
6DFXoXtJzMrs29+/te1GFwCVzcIxVMb13uNeIFy0WOTtAyUxkDa/kXRoQ94O0PCAT+FOvt68FVVM
89qrllFLU4mjw5ohs90MG9xJVVO5lTX+WXKshRA8cykO93eCrnIuyUXS3A3daXDIm0uVymok4Ova
ShEXK+u9rO6AnagJRSMoUZF83DCFmOaJBNzNKHycHEP6kJcFzp0UOYWWwIWzo2TDJTOUpA5STrzi
wJKGWs8xZIKn9jTm2qSHAvRIbGKcuLtQksRJwBB3irklFeIpz/RVkkCGa4AsbANQJ1kWID0Tn4eu
m6iaht1qSd4Nx0ULSg7ASPwA//OAYTqtW8yGYLKcB287YvnudcBSFkabjRlM1w+wLpiDgp+tFL73
5/QUT7xQlmWru0CA7jLShPgTitnZ4e4ofqDeypNnmfhAwv+1BHnVoBia/DhWfxEYo+IKP8S72Qkb
m892z9CkVmtdFN8YHl4VjNnySWjfysBCAzaVQRvupHEiiWN214psA5OiAQ4xWe6m+yR4eJVXBb5t
Zr/ICc96vQgBoX7Jo16uhXOctQAKY1KrCf30ZVnEKkqWu5wMB8uPKZ3GZtpUwvAV4zcrV3ITwVA1
K9jVjIOLTpTX2QRwDQk0Wq3y1Z2KRrg5wm3cG2tu6dlEZEFdvdZ9vgFz3NFZKMvpfAvINcRKh+d4
mrey0YkXbcWFNJxSqk/iMTQpQLkXPHIVGLFpnmilxGqtsDLZ80tYyq9v6eGXkkGj5PSYY0flS60w
bMpAwKOR+wDYglOuGJQ/pHHEtsHIvFaKXUUXnRpYtEqBONGoShEdUHT8rmJZ1AWqUj7rGMSgox4o
rUrgIxMFKqUvKB9VIRYdNdRVpFsQW9v8ID8mw9RP+eS0I5j6QwR6/wi/EgOOtFG4tv68PeDoy1ME
vJ8+ccinGhpF95Rvbq1ApyIKBiYhDr+j4jLQs1E2NJgKEVlJz+qPXYMClNaTG/elk+nQlsLPdJSh
siF9CJ2D/1TlDudIucraQFPXpZvGGEllskdX3FFIFpVWzfmeak6x83NBkc5dZvRvxiyKrDsqRdDi
l54eh7AXwyp9De2IUIhBMm2AigvMjl2cblOEjFUfAyd8Qt5pETjzuYZShrFT8kqElj4X6+D09TNo
QsyJFiUPmuA0oZ5GSzuMeGv8gM3c/l3isthMqOsW/x2v4xwAb2+j58Os3AlltdTqJoGOvjhB/MHj
1Uw3tRQB9j6aDxeL6ktGYS9bOFPrLtjOvPd+mdM/3iGJW+wV55j+dYqWl9Oeal1Ovvq76Zw/eWnj
/ugzjLBGQez3+GWmey6pTCzklD9W4V1wQxMDjoOcwvSaBRHcFCSycz0BOSLAWrY6BeRrMRUAX0I1
ZqLMcb6AxKhhYO/XGDPGS8MxU+ekV9F9gsI7H0xLnr3+oHZ4eaWVHbX5hcCNxHPp55jd/4sTG5qr
hIxt2DJtI8AWQaJvA+6yfei1Kgl12Qf+x7qwxQrXmiGwJVVNQBvWhv7ND5PVqtliOqyXKtMO04+P
pYG8vbZR3NOEQhP7rK3cNACBCO/ZU90n53m/dRXPKoq90VsS1GCuxhEx3wgy8TXJ4E03QrLY7KM+
S68qEpjG7EbvY98sLgDG6YI+eNPvHk0pOwsoYsFoGuQ35EILb/cfNm9GIW5Hg/+3QSovEdADxAig
vqnPoah/dBQkspqJ2iBN3iPDfDjoTmLop/OoVerp536a0aZezD2VnptKxeA0A2ufiKH4ufveDsxp
EqlLq5RJFqsvME0sXr5K1QMe2ON9hoIudSdjklN5dQ1toJ4saV6mMWXMMoujArC/ihPXNuyVmMtY
ApTfUnV/3dSrHYGL6pT/E24VJy7bck2t1VymR/nJW6NIgjMLNOskVqx49SvEnZnu/A00XpsNgOeK
QaLnxWQV3KIraKDB4AqHP8Epn6mxgZvHZz7vwaqM6hf2JqmunDLXZnqCiSWyIJU8+ZNSBQ84rJ29
FloRsYUlvtF+aRsXr1xdPDjVApJZo/UqadQmgUY2C0+WUcR5syL97TEi2kRmOihBzgRN9zeSuFKi
l+EuhEBDDLzQKQN1mfxwwv6RnluSO3nhCo0bjxNGWj9iZJGBMg/U+GXFueHPouxrozzQDAez8KnW
p5gNEFr+Ka1HSd7LLnoDpmwFTP7mj0VToNXCHPfg1+WsfHoH3xnXaTTMn2n4XG12W2f3aGZu1bA4
oz2y4oOcvMwjia4+iHksti6K1JGU5TqrYzH5cru6vo+C12+qD9Rn4ZRWoQ/TiY7VRfDfnZvlCXJY
aAZBWwTYa04FhkDB0BCqCIyULBrop30B9rEJWS5sCt0UVTnHJQP/ac/9XcdO5H1WnmN59snB7dK4
wR0zf8Ywu16lYRfn09HwsTYUQeBd9xCnY9gxyYgEq6CG3OeLbU3io/c7Nf9qE0MEpOryUBeVErrJ
ygMjAx8ntpooGlkn17KS3WRto+hy0OJd+JCWl5zSoO/wV38+/7TMN9k8AMx8ksJpifNWF5WRaJCq
qDgxWXQ6o2sg0E4dWZDCUhaoU9zbIE3OaEfB/b5ug61CHyZ9I/9YXVUWqXwXboBJm0hJl989YYhQ
3QMMKeNwXLcAtcXZ1QfrGv9XzjSF0+V57RtuZgw9N7HJfTyGDrXI67n1IoChDtRhN8SNbuftvJe8
WwEtQif2UxPQaMDr3TCB55LCOk4Lq1FYH/SyuiiTRwObMUfkd1/3AmlBo3WzogHFHMmphU0123hT
t+62HepqxXzemOL1kRp6z6JdCy0D0EvC9BSJfbzHidVDiFw5gaEEtO6oHkcBH7/f47W26W6mfnc5
WWR9u2/JrCUbgjvoLadOL3AAQ5lMdhhcR+ab/Qlvq0ZhkVFVi7+h/npeQCd45r0ZXxfRw3hP0Dkt
OcGql03vRFkIDtbCnLo2+FcVye1PYViCHGCRV9t7L+QWCs36GYAwKRW7xCaRiYpzCFFYSHUm5kJj
+B9Kdqm1Ch3ZRmXqXbAtD4eABd4q32Q8KCfRXPC9u9m28GDrmuhPwPXf6Of/U4s+58e+ZmCTJUj2
L6JUAAhIU4OsTqdAchI+mPcNn/l6lJBT+zNzmHN0JHfaQZAs26ysPrWpQjHfdPNralh+HzKxdLFi
iUUABUTUBVUyj4bp6ENIJoxWqIsJF9Bsf4tZJPtLJ8O4z5DhPjVfoPM0XEqog0GppHEerO5ggBZb
cA4Up/CF5UceSbJ8ncorgIsYFf3sv+pxr6tokkrl5yrNYJKVe41pM2SfJmFyBXdl2fbkjubqF3lX
meNGxkj8NYejvKNFD47otOh3lL7zKbOL+rPqLhQTZumkwo5B1LEtcjZPGoqq0wyfEvGD+DvK7ede
Wzy+PKT6q3lADWBndjDGuuGTBPSZSAVTxEFEFRLPaL9SGnrPPrrYytHQNujknUYYBmTr/nHYNa9X
Cr5j9RUpT2XKkT17CDVGaWlpHMLGFlzt/PWRpkt/M7XDcnsvSpBYxSziR6lXK2Fbm9DB0Y9tOYXn
OFLxvh9aXZhsjwVyHmbrGjD2govSM0balY8loHesqzXvLlcRQX+QVn7ADoQCvBKUNyvwb0rruldn
Z7ByQZ2w9E4dQtVVHat0Dn2WK1MLHbmLDHMAOvvJxYdhmh7Ire4FWrDX51YU/bCBqCOKOP7t+8tR
s1oOtKIUEOAJKtBSjx9sHYj8qdobqIsni8AHvjUicAyS2Ks3P0EiPKiQsJbnUnXSLViPoqlgyq5d
JAks2sgkX89DWoVfr+cAqbmZnb/aBNufPU4mj2Io/wle/DAbfyPhTKk+Glr5O2f/znhmlGmE2feG
Nt2yg+yTSuLle1phNKrbl/RwcBEQFp9WdpgAGB3TwSZFSVxhfZbt3HU/UvzhauN6FBc1lN4xUpkc
zNDEifUvcoOwsd7k5L2kRod2qTDU7rDauV9FK37eYCatIN2j8fDNLGcVd8011YmNd6fkacVRmuOL
9xWnqFhBYd9cpC6E7FNclDHkmYVY9wrZ8gLkwDcUN4XIGITRN3CmjxNZBk1VLZdSvSp3Aymc9fe8
2w59d9O6ml9jpz6Nxmj/rGyvqrbAxOzuBWMePIUZv0fFOxVWtFwLLGzTT6F5WD7PKqK+A+5S/TaJ
yBh/KVce1b8dZ+7wTj3lyHw3u5rpLK/cKEOVKfUrTOccymDAv3mYz3h+0vPld1Ye6kqp1Loqnxk6
uo2+iwiuo4InCwvAWVeZGioK1Zkr/PT+B8Q8fyXsGIlQPB+x8S816EvszzGipW4icX/0OvCAEk9X
3CoDOWQfWhpdJu5vRiIsPgVcetnvPa8jO8Fjv52TG0OMcYwv/pFanu+XUBOAOELi7BwyQlu04vEa
+DPURQkCoOPNoUta7xjnaMTsqghv+gZuoZw+VOlJZE+UkdE93dpEuqPiPch70iMgpk1R1kwnzIVa
iVk/92NimfSp4ZC9P+L/t3ShvESpeuDOW7ALrsrtoV6md9uTbyHhqHauLAy3yLtvWRgr96tWaRNu
1+45MD230uZv/7ddqmLFgYtt+HycNKcMsKT/XFdMH8RdyOUIlryLv712ECIMgd2oeiJkWRjLr3+s
tN9g6zZsQCFI5L+2VNM2dIvu9VFMFP1Z3ywgkyhgHm25JGJuPjvcWmzyhZfj/XMZDuinpqY+dNyx
TnaYF1NpV7JTChFIeJQ8wKbj3uO0EOiEeIkK2r2Ug1TB82bu3gVrFnbtOV/mcEQakIcMMGiwpMTP
EeYboC8f+dEduP9oBeqAaiyuhhugM1GpyhekICiLgjjlEfEcAk5pjHUQkFGFHPtIeOUlgsVEyIZM
GosjbjTGRONGkSQd6k846GNITKIJlLELNDgPMn3FkiXGAEcPzcxvQNlaXNOhoxG6nCz6iIqIWA7C
HHQV7osuVC7Z4lV86zC3e1b+UIxB5uTjl2Ih3TcooQB5eHFHzm0jGpCYJUBUJr8KVVmtsenZ3LTa
ovi2FAovHQmllfyyUWxsh/j4FuYkklNDrtkGeTfP4SO96jbm9dCKcOHP9fEzrawbbpD7S+CAE7cO
yYg5+ZuaqYT1sjZpJhDKMNTgfE/Gkt3QfIEpYqHqj/Jcgn4Wl4WYmPLn6qOdiPjvHzYCL5hMGafB
519E3cgRfYqu9ViC03E9hC6fkA76HN772Xg+x60cu+s8S8kKYtAgUkBQp3716CIMDbAeNtLxnFIe
SU5sthTjNmqkqggzoPIIyItNLCCVlgJNN4nVp4D3X/PFoKq7OmbtFPha0USKvAvyM5nrfht8+kx6
OESvnVLLWiXcA1U/qqk5CJjmTE6iWlalRW3+CY9qXryZk4Lh4WycC9QqN/o2w6R/ptoGpQL+Jr2c
fH+ZyzshUl9RZyx8PRoZvFqo2XnYBdVtiymGP4GhP5KMuvu9wGT+6qKf8ZXILsxy/H7YLYUnurjR
AWhqnmXtJ4Oj44rVOdOGjMb+KZpgQJXX9rwS42kPokFUVgDXLtNcO17RYITfGvi0SxbbBUAdyMCY
jXyviKXNm1MV4dVZSlJTdKhFrbeXRA1clx392qix9v2xDmWJFNF6nkzAy1tRrLXSOf2jTbwkWHIX
hAYhzCHRMgUO2e3bDoHsrv8+p4Ck+2JJ2e8wylbVk14WTVbigTnuBYNMWz7lM4AHxVZTt+VwqknF
vjoJBKRSB6ZF7SzcHeKcAwruYdHJ9vJqGrzB4eNfyECPTWqPJM/U0EGwjAr56n1jRLI5OCl8ofuw
Z1j1qCQiO6RODgnS+pPskgRoauiWhIBy7WQt42OVm22Vk2WTGSTf0vIlttBcJN6xC5f1fh17hgfu
zSANHEAmY7A0gpiz4mZ5XMpmvogmCkBxhmkB8EP60nCoXk6YFEIx1anLbCTioaE9CMhytALRwMMf
FBsMkZktJrX8QV5gfxQI14BJn0qXvbFJBDot6V5xAUimMOJ6mLRD236VzL+7S6D2/eqyon+Oc8U4
AwurHWwr9dq7XTa/NUyQAwAqGTFCu0WO/MV/W02umgCD1iFXbDWI84WxjSAjJOd3fXHCgJDY8Nc7
X1XAiMxicmFxeGsFK0cdrgzBFLUGa4KYz0Bfkdxhpw/waBSyn2vjA5N6NbfOFOEWsx5Pfx9LlyfL
Ds/2jvgazqsMoUsI71TJivvimSfCpQI3+NXryNeD/1ThCRryF9TqoG1DtMYzzJAa+Z/VlDuHxCHg
JU5YTA0D1ReTLFud/7O0/LyJ9yet0EVdm7vB+HBimIJIaZHAD9sOy19Y2FbMEkKkF5URnZ1Mt19P
Ua5L5k7ftspHjMnkCYraWjC/b30yKquj163/P2Dl70X2p0WqkdDuYATIS49qyeFSwCcKnmZy4k8p
FMDxQ3CGQQYkD586lI4ed0VYi/GnzbnJFZM81i5E/w2z4eU2ZhumkQd082ZDkUH76UxKdUx5+OB0
RJBd5beqZhU6410E8I5AEjIKbWXxZgatHYmYldS++diilaVYpjuTTtWvmKY03vQjpuJFM1OZZxQI
duntTd50PieFbR+FKG1WNO5+4lsZ9gTbR/KXwWSLoX1bYHRG1V0f5Gic0a9d31DQe6gPO/coaDpr
2JBDkMqM/IfZrISEtMfw0a7wLjjp/zV2RJdEeygIKyS/U6iEm5pb2DCzlbnjssvcVGTEDm7H4Ov9
b+NO9hXvWp0UdbsM9Fe274nkYKwjmqPfcJ60sfg5fgZZeMOaQ8ZF3EtnsNUNZ0vEiVpQf2i166X+
KORE5vBrTaCQ3HbRr/kTsETMooISCvywmjJWypNtg0ZXmVPDZbnoF7I4Y0nKRRwFMYFIBnTvykWT
uGIf1eUowgy+abysXiF5bxw8QQva5pCTRUSvMDG4at2rRYUjt96lLPWN9rzESmi5QXXBv8UYYVzk
9RM4u9135RmnIE4g+OhogrQwNHnDb4+c48WWzO894a68RblUZNKgJZ1xMweovtBPLml3iWoP4zCT
KjpbDvbguEzwSmbBxH8bZfd346r3uqsUYrhhkGMKcu1lp0s5MhPFD5mRCgXQgCGjj87lh7tuH0nr
+bb/FQMkrmikQT3/K/ETXWFlTWv3kJWGFxIS8SLTtNjnhEjVNTPw6UXyRuBzNo7k7ploUJtkEvbN
U7nh2ZAXG1BpT6Y6BlRZvcZz0NF1kjOZvqf/PLuAlhIpoI5nhAv2iZhaJVQDahH8pHlK5VtSU3tL
kP/kP2GpJ/U1OSB1L6jYAzn2DsnlJRKynVmWYR8zy3ikSrXyHQH5ido/cDXapJ3BItl4wgJteaCR
LNYr3BfFnWXEk1mlf82SaGfcWdFKT0XOEkOGL91P5S81PcvYOrI2WYMSGwUPkGUWOdnRALS7QNxj
hUGPD1fQRuef8LA5kqM8dY/vNtp6K0nYQuVXiac5R8R2Zp/0y88eJHCNoWPq8lbUuIK+89G0nllC
gUFpEDdYF+vhr2dO6+GSOH/s6g/1nkB7K4Doza1pVsyHux7BB17qXnXTwEf3n6igPOjGMY8Rissm
0VpLPMEh5x7T9dM+6EMMZfiH437RXaJIjobbKEe0JDVTIHfIHRNKDJL+IyNoYw59CQO8V/08ViHt
aT73bmIxtdTUDGK1qULI/LNCvr3MzNCjHQKAheMf/ddgcRYNz6YwjmqPKEFRZKHQg/qwbSzGN9AP
6KbdZ1a6Btvm7XIVKvm0ZMzahlTjHpvtOvBpddVlfQnC18E0C13x3VdnofTI9KLECMagzCwd13w1
24ZxqIsr4H8ZOEbLuVr+WLsq5qbi75yrRps0GYf3O2ove2Jole+tcoGx7cNqNj5ckFlcv7BNBHYQ
9a8GKLEUvPyuMb8BA22KBfxC0682OlN0Fv/JbGLV/O/2BPqsZjMvwRPP9Becu1zKO0PfZYf3gD5S
SHzaHH9e5xd+Z3n3Skjk2ppWfDZI362s5nYPCjaaVbcX/Yeq1Wo1GSRK4Ryv02C/ya/xBMK5zw1P
14BhzywsGlKOslf18gSojQxjNS3ipgwE1MpIT138XvzIHeoKavlrrhgRTH6ELd4UVQuCE38qy7Rz
UKrhJvEcnriK49E8m75l5jBlmtW7KZgsl0oQu4wSfs+su9irZFvm4oykasa4J7yE8XFSVP7QGzA9
Z89KKJRnNW0n2f4StKZSrQLpGk0rd45c2gx5MKldxD5fZdL1s9kXCrMpOnzjGxjyKqegLXYvlfPg
/iRBE0ePCGT05GHe6+8czEpjRhRhqMnU7dKndjfReE5Waw4RtMyQcbbwXk9ph0MD+h6JksShR6lk
sQg0NFbJgswruOwlX1QJmUAnQjFH9io/1h6il2qXH3IeXBSEQpszBUF04+UW1tsqnleL+5OS+cME
lnPZvG3S1s+B4esHyJTEBOR2pdBcw3CukpTL9PtmJ+wD8Cc0Yuq0jPriTci2TLysSSzw091Mcp/+
LYmTfZAxZNmUW6d4GehJz0aLC0jgA61Hm5HYkZNFo+tflg9cv1LCULmFD/pcX8JBBx8SkkLIUONJ
YZuiqEtiw5waX7+ODUGRR+zLWc0X6zaaYwCFUW92WoWBGAq0J9t1JzNqk0p6G0qquOH7uPRQfs9B
QtZl4a8KyMi2yDQrsKWagemeUSRWSTj8D7LAuZPS6gDLTGMB4LtGypOqc68QNLN+h+Q65zGRkzdq
/MK7xSs1I096pdjposL5biOLVoPz68Yn+vAyafC0m3M02JngghYDh8xnQvxJTmHxW3T9f1S+IDzc
sEEjsvKepqjr3+hl+bBIfn2NlOXxDlUb4CeLdA+TItM7jd1WpTLGAv9peiuCSut3u48DdOGGirbV
klc+RrAxYBT2GiPB2FgwzdS6kLrqoE+l9YsukiB09tK/QGK9hiLQ8ptWF7yK2LpTQqaA1FoWcf+w
FX0bAGT7tyGMrmZrJvoURiaaLLFnogCeOX5qu2IwP0L7ATmQCEGJvCmFsraOzSvvrhYzDNJ+oaZg
TQHTmMD7Km4b4cE84SCSACGdC3buUHoUGbc/TCGRAcDcgibelDq99z4Hs3dwgR7jUmrS/TSmDBH4
5ijkt9f1UNBzaBUqNCJVf9rhY4zWgYbv+CK2OvM2ye4xsDn58N4wloSHUFU4tsFlbPw1LZ3NJ+DY
xZKkUfj9YeZgVkU9C+LR1LVF/W3nNRdol0b0hlzl/lpe9PXY0YIg0LETwl6tr03X2cY3GSe0JbS6
eVHE49XgpbgYQl+xbFgntEM8+tcFFm/cNZ0iyIgQf8bfpH+XpyCp4RELD/bSwQiJRcyj8ynxP/K7
jKUNYREZiW2zL8GTa0qVz53a7Xxh6BDY8HWq+gMp+/wyfJrRkWeTEbdhAsNkf41fduKIjWd5wej9
MuTzfrmYoK2Mn1ou3X4E7KFFW5LjEoTR46pt+ZyC/7BjZLgYLP4JxIAE+CsmXsPX36qJjdz5xW8E
qYNjzftDOfntHj0mJCmXWr5S5fj89Vx+PhaIyJlBEwaaG5vVouaZadl/OiKiQEJY5+UurD++SxO1
r4waiRdVeAA91MUIa8++7j9ENIoi5KV45L11CBE2J1kto2N82PEe6RhcfL8sR5gsFLF1BJbey6wC
io8hLVWDzEdtoeKjd5OlrBBJCkENyf7PTrzHaiRbnNYxu5ePtzf5FPbKAzfM83qVRcFjD9iE1Lxq
5iVdRa1Jn2qfCnO7RJfaDFP0obBxSOlVtyePBIUZxER7/fGa7mi9OmUgzj52ED3xSqdj4Ig3znDE
Q2XZa13nj+PYlAZc0ONzOISjcFGwC6PMWaYHRuXpRIcvzyk2SXgr5kwLWl82GT/sExAEu0T61ezV
yVa/9A5WdVITc8eKhI28wQLihNRttG19zI+Hfe1eXrvhrYw8UBGaoX9BbzDd42i+IgQMLkodevnh
p0fYQ0ZZHQFlbOl+1DpyqtZeN7AT8fbgzZwCzlPFHoLL2XI74ID8MCEMiXl21LJHd27Es5uMYsI3
5HwL3D4WrdiCxuzO8q7cm0iHTP4JIy/1OnbRLeukMHafobYp6Anzybp6dli9ka1yR1XIs0LnZzMD
A3HIzm448NKtmsLqHZngzr0fkt0fzmxLbHGxlRkM7yLlaYmHpcQQrZ9FGzpLvQPTFa9mPCmbdOWR
50ggLSlOEUyrD9l8EZSorz3Expz0/wzGQhG2R9bpjbuEMmKsTcISaMBG+DRKtV+sj7jBPr1JrPNK
DHP5Gvnrw4uAdAM72e9h797XLC+dFHY23F2XzYkoUJnsU4Ai47u8vU6dG+1qy2HHB8iIAWgcd2to
PN5VSA3HoKNey2ctdTftLw9OKvJXX/g6EYjn0etPtbTu84hFfXbtaWB2I55WsCvjdxK16HtdnJdy
cP9nvj0245sJf5lVWSiWcOXCQCJVDRSVxF3QA5Laad40qVVocVx0SzC4R5XbjJyc3wV8PppqWtb+
nxUlaWZNkE/YSN79csgHSKmBd23KAB0FTApLQ8rJbY3/qA+NhmEkHgMelvRCTib/ryTRDSunTrDs
t8gwAz0jSvOX5oMGlRqojN/b+Jm6WLfqkKbSK85CW+TRi9tEQvz0oDMC/+qkT9eAoxqf28E08TBL
bfgjXGzb3r8C8DvmS896RA45B3V0lqN17ZN8ljz2gqzpvjKn5rtQZ0RmPkLY9MjBKTtG/d+x8ae7
81AcDOCkUCOr3EXwTTP/EHB+jHdQhDLoFxY752++dq9npTVmEFAZ8zLnpdRR/MXbRyGx7fvLtZ3n
c+6GiWzQZy9uRmVzR7+EsI9M2wueobmJJv53z5iA/xI6fLsg/sRX5JHz6ErDzucossezdQLb2zY2
x9KVhY9bJd40t6hEUQSKqeBwDX/vod8mFbi/6bLgur8TVq79FkfW2d8vynBk6Y03wEKafdFrC3eA
4lk5qfeJ5hedNhY5yDpeJxwN7opiYWi19qMaFh0Ewz5J7/97fNaeIrC69TObG6x6fChrkie/P65T
czcIATdiaGR5FfypUHfKUi7RG0kpLvPXQmpAIiJJB1D1/iu6uhPqbURhRltv7Ihj3XTQXKuJECS6
Tv8amgP4PtONQFjAeJ0Affj20/ZhNa6lziwjr50FoJF5Udf8SMGm06gfvomINBwQeL4OQPnqxeZ6
AOp97jRZgBi0XRQCN+nTC2Spzv3uoUQZBCzJEej7EctCdpvVh2Y74hjda3COWY5QpcP3BGTWbAAA
P2a/7FQFbA7YI7h1nrYoUN5ZU6/BfSqOBnqIDmWaBJeFlexgb5SJKNl7vcifmhBm60pbJjA4dskV
57zTjiMvJPZe0fS2j4egQgS8+SXSDm8eysMO6ZZJtjiL4eU25K0anbwZ2WTnxWEplBp6ekAJv1BS
iyunbbgmX+i+3Hw514oA9zSU4sEy3tUzXY/HsitUHoDLAWUXgBBfURms0rtEf5IIzWpFht5jLDw2
K6L/NZij9zMpBJdUOYnaH6o6oGj2mMkcT2l9Phgv8VOigB/D/sNPI3MM8gjJ/9lTmytZspyIwtgO
zehn7qiPFzbftgDIVj+GKky8osvWJgx0tV9KDNJ0p+cTbI/6bFwiMFVoJydGhSxCRxRzOmZ9lfuJ
5VyFaEA4IRnsRwM0e6RFbvspjdcYIF/Z9pRXoiPDMCfnrq5pci1Hx2P8AC4nN86LRHDiwOqDayr3
e8blsc5BGsqW+oL0f9qdwb8/xBFQJtIOg3cR1Y1vuLeS6DEcI0U6LP6sImU+M+UCiP4VqeGxcPmh
y+M2dr08zk7s09HBxr8x9q9pr7OVY7OofxZSFhlg8Bk0Hhc2jazavUpTDZGnR+NVFc9yC7nqJZsj
sDdEIk40f9/F2LyP8JWBJDNf9/XrPrtvz1CVXXYTg8upGKZpZf5fpIqnf09bAm14qgMhPT0owTuw
bNxM1SQGYjHX3yGXdVEzgQxLDPmAvcuBB39x+KQMwlLyuIs/QndWl3XbQlI2194/hRTfk2O8pJVH
/RqgppirGxftu0wO21wir+GBQZB9oBE4r+EbtM1UkT1H5L3KhQfM6HniHyORQzZsYvSJTqc7KcCR
t126fVbc88dEWNvMnafl0fzOYNp7ccmgFvxoBOH+C1FVBrwtyB0qXqaG6TVsScONv8xz5vKui5zq
0Z9GW4xyCIkcrFQZVs3DRyPZUtaZ9nER4Hoftjcw6cFVfazSZLT/YZYykhwWGAe06M3FVt45I60h
9DHqVYDcE209HOwS/xJwc857ScCN96zLoTB9Lkvai/BZxoly0bjhsYtkGtB+kd7GExHMQAZ+XCKQ
qtui5l7bwkVtIcDjGR/id0kVVm0bHrp38nT8iYSIhGcNY3NjAw3Ko9+tnEfYfS4FmAxKsX3TuVpc
UV0okTBbHrK891WlIIMlcntv8B7PeAiTzSlxpd44wqRCz7OBKlbpE2INhmJoLYaZ3FJB5Z3kcMy3
lCOCXZxuX/rU0XJPpAbvvKUW7cEfNPb90GLq8ZUUwaIJ/V1WyvVOxATX1CTsCGDFHgLGTXisvO/7
+rcEKWw96CYfmdE83a1G2DM5EvzYHB7RA91yNSyecPIiM14BlYQKOeVOIDyDbCL9UG7cIlkY9HXS
+bJOkZUcjaFzZOss5EcHaXKcrzqrmZ1Y/seWV+fyOdRgG3E84w7mCHrkCkAQj96RGS/EAFbLNOHz
h4/XvRx3jAwcV2jXHs+PN+BcJzw8NkqyrMArdrlxM2uieUb44Vlt9VOWpOx6xItwZnd5R9Ivo1ll
Uc8d3tb73CPAW3adr98t9etA6fTGcKWJMSUXr+k3ZqRwpXYXopTFQeoM9IwKfHFAkcozNVRlyGqj
A8sFTKA7dPZkxrkEDLwDhSWvaj8QlW3Ev0hOmFu0v/VzxxdRwUAzsQ7LaulVx7+hs4wEZKsL4tP9
2raiJwvWJWQ6ITB04vAGaYjbslOOR/C3zXrNGgNl9ESnrXJGDDRfgWeGQZf542QWPmqZs30OtgZi
oESeiL3I2F0ShvkCG3Wgz85QsQIyYtc0aUdTVxueXbNDa9JWm8D1fhYGU6G++73rmaCwQ98chQqb
8eSZnFWaElC5PMxLxXoWKl313eKowVCzCudyJtT5L0TetOJWqPSoRvKuojZPtM6XajxeHGm8JSgF
9lc7pcAvS6l9EOrFvtj4OzNVi14CNabvj+XF/MwFQAdrBoTrYgyJfmu6e9j/HKyHiBJ1rjnXrsh+
an2rdw1rgb3kKgnAhoR45ADMWzQrm0ZeaNlw1yr6ZIqNmpehh8jdjuHhhvEKY8lUtKP4pBgc4BfV
CrEuNeAKuLrDyGZEIm1NYOPygy4V6MwzbJIuppGQY48qzx1o9UuVnJII1iLddmnNiZxz0ZMno9v4
HHPIgq8gQ94MpdvgMIeyyOH69rpJGPtNDMJ+5lXga6gShH55TmJfxy9QPpWx6Hzb/4E7bjj6m8N2
D3skorxA/Dfs61hklLrIyPeUQJylHTfD2Era9etyzqWcWO+V2uM0wNMJJbfzjG7VJkzMOKLH+NLL
C2JTUmoXDAtKLad+EbDfhcIHr5hSm+D2ZTPjYEPOBQGBsTmCGYDE25jDB+aMons1gpnJ0jpY/NaH
RYSeVTQpDh46kIbgE2Ngh07Vi97ZG2Nj3f8IIYZ339NuS3AEoHpN1cwSeSAM63g9diCii6XmGhKr
y0q0+rm2Lv986Nml1uRkwLNzKUWTnourgKTbEGXHnGsz7ibprBtC8eljBW0mfC3hwaIuFVbY/IcD
qf2ro7Qgm+Tp6ctkTYgch8pItDrNx6iQXb8H1n5Wzj3nAzbqZVc26894d6PiYsUSCBMixFdTz3mt
6s1POyMaiVj0Z1r8vp3SlmXRopCj5Sk4OGNg/okwHjKJY8PtPyMbYuWt/gSQc2tq00mzbkIjhOmc
yNeoJUT4BNXRbZewczW5zffi1SaPyJgqFUQHTlXe2zUnBahDrf/Sg6hMeyQAe8znOOe/03QUblzD
pvIoLrgEpeqlcQY78Q7tXG3bNQIb5dgh7UV23pkBFoAe6z5WFzkx/t5IBj3GQgi6QKB4G5urkJ7Y
srpu7oaql+H6Bd32ik0b69SFmlbIf0vcOvU5HHBeVK45T5bzrXDgmbOMvPa7LLxlQWUtXTGaDu8C
oqiWAYmLYTaK8PV4upa/G40pE4Qm77da6LQj3e3u5zfuTj3gLcHcut48Q1zZ2XzZxaQNTrvjlkFH
Mq49Ah2sFnbPjjkn3VOU9MCuCqCCs0sEplpkvvbxyzB0CSGJIR5QobtQzjZKJC5VijTSo0QjtS57
Rq2UPmP8jRl/S02VPA5qhqEjrEjwKskijQcVbkgp7f6mbWgj8qDtZ36uqxXLHqEmsDvzZfa8zJxt
0qUhP0e4KniPHs0z/RtdPuH+TOIwnSti0RZF1faeg3JnmN1QFrMZyI092V/OxTUzU+MJMRPj70mD
jhBNKXaIOvRvSUoBlS5l8nIqAJyjvBZm1iuRffCAnQ9Dw+n/bnidrIUEiFyXY6gITpqPJLnKIdUk
3UezbZ1ilTnt5mzNSwfmKgqqIumT7R4+Nhnxebtex6SDSUmxeWedOD1NzFTe+h8eiDI5iwejPsu6
kmFktMjP3k+4PQCzfHBzpb/XnmEXz5ja7I9HRfqgmtBN3bwdXt6Pd+oVhZEpmC8Jp2rza3xpFyZ5
8UUMJjkIhT4xzymRH9hCMc81YTIXVPMfa1d3XN5BweQGwdahhlPXQstbhAErCPhp6S/JVDyjPVYF
J1FxW41Nhu8nzgLb20BlUmfBp08WIqA9J1PAuaRYPiMkSaIGtl3024VkTXBdSunkuqwfDOcH8LaC
A6zHgL4WO5TOrT4GaqKak1dxTlyJy3K07gBrFgVxde3xLCnJGEeq9+zNo4Sm7jQozcu7xF6aydF6
Z6MR5Qi24DwtBEW8FiXoTOk4wJASnqMzUVXP/h483+vS1Yi/cNnnoTL34eACklS/zKofqD58wv9P
KSdvpM++HNfK64D1ej6r1v/4clSNJgDDcM3CuMMj0Bwl3UeuHXhQIfHEqt8IKZs0Rxtlmf040Q2F
+ZBw4t0RSqnmXQcxeuLybOmucBEN75qjSB2mwAtbqGPLZykVECozJ15NLQhkDudvk5uIqSemOag7
t3/OHOYppcF7nm3z4zVorPO5iOFFF40KJc9Z1tPj+ucC9vlbRa/u7UrdSaIfhW9iATXKPofj+btR
bGbTbHAt8UDlVTscfJZRBMGnXfjX3zKQIJYdQnw9wyVGmeVykAy9qI2mYgXQ/qnIuDE3tKwRV+C6
IeCXU639bcXRa6p+7vmz1mdFielwrI+J7aaOGj0Cf8BiEoB9qIzQ1uKe9BymhATwWRMg4b1a/gIs
J+IIeogjC1DHcygbz8vP+GhU7UUw4TflOk5QXCoQA6zNrJqSRoDbw27WbLx93Pho+Hnw1Szgded3
Lb9ANZfhSh5F56acqMyJRLY71kiI601YAboOwYqjTm3xdzxPMbnX/xPJ571fXiRdUrVVNf65erCg
vhtbYotjj4tfWIip/FLq9Ctw4V7K9tTDTlBQjyIxhYW+sDS/RLKUxuOJAQpJeFrHkz0vS3l8ij5B
kM1dUpqho4kGJyfX0RAkBAIUk+eDwi/QpAUL7oi8WVp1kONSCGXfzCBkWf5qq92e0SNrH3nOL1rg
AJtW30P5pKgF3VztalAW0kUWVKtNtjdqPqXX1Jmhdq5yIfyhluM8Bn9KHT/eHuNcS8u1ijzmlwcq
l+hbWyB9jn2AuT782+33E4+58ML5O1fDsQs1K+TVF2VyMOIRXyhok/a1YJBbcD0//dRYBVR2ZxVI
HLOFDbllqp3zNYtPT6v0mw1VsMtWa0oRRcSsQ1q5yKBpYZS1qQbWhc1nEWG2E183DYMrdPBF23Qo
uNfYMrz7t/ccD0VImx5cQW+4NWpzbxMLOpnmwYEc6KLZoVAxMyjNXunGIsJDxfYaZx3DiVhTsQDA
b8Lu1vzQl0RDGf0ytpmHCWKl4fpM+Q3FbzxDJCKfRbcM9HF39pkIF+oCQzV/7LnL9dnu/d/AhD6h
NUYPrNRljI8b57P8QqQZI8PmFdcgmWqFshgQfkAv4OqT3Hfjyh20YKk+yJg2gU0p5XVFBN06KeBZ
j+/7pIXi4Swa36ElQt5l5HODxLMcgvt2fag7MTcxEokq/r6nj9l6hF7fSo63rvpZma/sdJMSFOTy
JQRBZ5/cP7Dh14sgsB3gpwmt9CWn1lSS1AY0w8puRjQrzJYZkX0Ey6uk+gAXKE/2jwutRKyyCaNg
IR+3QyePJYBMhpQOsWkp/A+Tz3ZjdzWS3pQawVZYT3uFmxDH1AilNEdjTawjcK2/OyOaDiMgT3rO
mJ6gj/sb6nosGui8nXmgpjO09ifyIerzygZpXhH42cQBv1pVwjUmNrJMwbZHwurXVcm6scIco1wz
iGyLpPlhKJ4MGcSdgNC96Ly0gJHQOKBi4yLXw9KN2U0BqkZt8lUbOk2S0nYpDoqGbyRiD3h2yxTK
TFzADn3nvL8kfqFiECMkuAfOW34Bu2M8xkiJ4+GNGx1yUgbjxnXTQojabbUHXAm4ZAc9PTi6/TmL
9V3SxtQoYR4opvQHaRY+cwIpj/x4THIQAtxIVzQ0rvkJQBTvBG3o4ze/viy+hv9bVxKL1qyJNjbN
LpHNp5N5VSd1fMH9KA2jn/c8tQbUNTsbEBgmDxh2U7i9y1g3ZrPkcApZnDyPXX+vUEZ2RtuIlWuh
yt6OMU4KoHCxhja63ANLPHlemNwxxkqiGdsqq0Fmtvl/n5iIrv3yHanH6v13zqEHYXDcGzha+gvi
e4foKEi3DchciEmYF9qVYskUasPBQlifpbZWOAwwLhKweG5Ap1S34isHEsbj5ay/yzICcgX6TQVZ
QJuYfIgwFFx0CXOhUeMUd55pGmi26Z5+o89iANWkhwXPBsJUbKJP+5lD5qV9Mlv1GqvDnGeUa4dv
ti/m9et42upL/87ukNovIxz9CUjam/OwGUW9/GduncqN0dDKGBm+t6d9FgTzhOngZhHnZ7SJSNkQ
w6Qm1XMJSOLiqIPEyGNG32OnsN9Zu8Ne3199ewnAnrG3w3QAFYBng4lDQN3Djt4+V3TVdzPe1p8F
IyRUEXSvE523MohBcZi2kjY7oqtAmJiOcxEjfIM4KkBy4wiKP0te0YaQhce49BaNPwRRL4jel+Ek
vqBQPhF/PTWvGG4mGz2gm+i1Ae7quyp85T3WSCG67YdCVjsdKoO2GF2zdMmcHr9ujxg4cSeK1/iJ
MR0+6UM/IEhJacGXMD+b/FfUHFY35cV78/7c0b9/rDk/qpRfmmLwo2G0Ya3xrv6bJdDIYIwbmMbS
bBMC/ZC2p2P7z3iUKB2guQUwIdPZY3ohaLPnN3R7UE5iL0SxGO9fuEjY0vw2z7272To5I4xpa12O
9dCgRo1/rno27v4dfWFt5JAXxHlmPOczs9095vy3eRckHTMqQijn7HoKeas0qFcYD2YT6mnJ1nG5
5EQ4CEMAoSIj8Zg/lVM0Xv2OJyrchPTNtJzi8XbKXwiGaIOSE3/kvI2dDFqKXpV3I/rvNmQzjYxN
k9eQZUfXh3soaPiqd78lpaXA1VCB/nuPi2F0jT7008yrDgHuzX3NVpjZ7FDY/oATb1ZSm6jYEJAV
/dga7z1UUOypPxDOoSgake9AHOR7hrxLQs71tDbjaelsfF4i3g1Ouwx1tWTAs5Qw/ap2u4054OFv
2oauUIHWtzfms9XrRJOF428AvCyVuN0Xoq5o0oZWsTS6yWsh+h6YTvKnxB/7XyzBX//I6dmYpoZf
Ke3hUfqf3pdEAdC+tNcgBCpKbVz+2VFdzakno1B4FV16uN8zo+a4v0IOs3/UJlh+LP8Ai+rtF/Q/
rNWbTGDdscenAV0Dm8zerSwxIcg5EUw0fAqcHafUj0v6dWPzvaFZ0TAZWGyOuhxmum4XKbABYk/K
sOWFJQkjkpHH8ryXJZDu8zIHkXQWuBDUvru8WKYTbSYSFeHQ+rg5jZ6PnUJu6g1x23HqWB0vKMj1
0bRCmrK5vCS9Wz+lOZmb1wUiZJiQvDYUDtgIStrMnKJxPt7YsmAwAEWAjj0z2mrVg0Pa0qeSA504
IXo3IaEHBm18BuW6ivuAHtyQIpfMpE/a/doSVaBgcykVTXb6GzhUoYR5h3VUWTqbYyt8o0ufZsBi
eWNmdMaHnzHtelrQO6NPvzyXefIyiq7Wh9IHq51IvVETrv7nGSqmYmYVcz7OUVeraQfqoLGtehO/
N7pD7NLo24tOs8N4JGCM0KGmpuCsklZdWpYZX0jVmWkyFy3mFaen08abxPCripl4IORKdn2Q0b5i
crwy8vmvJq1EcI6emurS0Ac23rLc0VBQ3LPQF/iqV9RXKWIk6NM3sNyTarRQBCjSLEa/6vzbY+NW
a/Pu1Blj5THrzMNhVyyaEVIXPRe36a+5gn7OnkfrIWHHXc3jxmkAxwscVLZcD2jmQVEWkrMW2UoT
VFvYqYRbP7Kp98fUhpkXcrhavpuYOAj7P3ST66yDUD21qUz5Rb1kxiaGC9nWhD7t3nEBfayUeV4Z
GG1wbsDpmPCN4+UCe+C0NEreTnw36WZjrvxp/xaGGYTuw3lwHTeHLKcdgcA+mSML7E0va4l/DtIO
OVX2s1rsFwvZh01OTJoeHdPQUbvbIc0GggvEPhuofGlEv1BEkSfNcPITK5JMeAN59DEuZTUeUTQZ
C+cIKVruRVQnmnVpSjMu5w2rTlwe5wF/OMS6/BdKTXAQpF4GzjthSwkpKrmArSs/KfSEQKJ00JYo
1pmRFlJFidB4COHl7lj75iHBQPlo1wytu5BpLlRq/eDeLmULkHSjW6++ISYixj+PWjSBnzFj26Dr
5whDJnKlck1o8QCYm/4ITiytiSW45Yj+cug+LAsRguC4KFbIYq4EZXckRHVYNR00g5Iws9ai5ewC
6/eSVcu37Ag1aJY/CoXFZfI18rEMsjuTCnwexZE9cgcTwiyIQ3tVYOOySyM/iy3ntqn7ePkiTCfE
siVSuxxe0Z+yzDhsRO2sURrwvvh4PKmNSavX0iSIyjdwZqdhh1AZmROHlbWh/rtGk+UpPBrZFR9i
wO1cnyEcREa+ifQvNENCtQW2dN4OCepzUvraaL+7Zl3322wKtQpy6dBG/kw88EHADzY40DtVihVw
uNQTKKYQoICr3swjvs1c8bL/Jfgb1BGXhI1eYBH5tmDVlYK0V7f20tq6PQIN2eTgKSGa3TOgOvIt
P6i+Gc+9IZBxU9ecEA0qLVf45/EZsoyYDic+d21sb47Hw8lLOfkjqASYS6Y+QPGkzpvBlSyHzPIb
J8I9DSP50DMzCX8/obZi9zh/rs12tFP+fKKsEY6l41s2lM814iH3/JdXt1u9974L4DOwM6/yO0xb
y5qXxs9vGUEYnR/pkoXTpHG//i0yaaYzJnzhTQx9jT4BSEFStINFHszUgK2QhM/qpK6rdLKrpyBw
Cjn9kMJxHQCpfmNHl4k8lDr85g2fdLL+/vlI6R9DG4oi5ABcnFeRWBtHbWl9J5QAUcHe6MPubIIh
btuKTFqfeerMWgkq/cOgBONBO9EA69BankjwXnn/D+TAedY2l2JjTUJBF/rE9+zCIrxvOPPCmtNU
ZEfmM0DAjXrSvwRuxY8KdWffxcEtagxnB2gkbOMGNC7drhxz8xrsQCKBt47DsUBEoSEhJIxTgcoi
SjCso20QYGCVlB2cN5lWXzirfXVtAa2iJAPtBBFj2taUnJXpDQra/jSIMLehNLjBdLb4qVUOwSN9
IvkBT8lr39jfDBQjaNNgBrsEZYngkq2461DrkEK+aVwUXEikU9qV10Io3kM+bAhyFfZN6l5V5E2z
eSIu6T9nYe7CHH9TyUrYyr1W20Yu2j9Iir+xpnz3Yt5/0r3Duld0gpGYDN1jr43SYQWx6JhxpApQ
xFByokIAUMC0FS5xiZcOs49AUGF8MJqBPd/6lFHUT0BZHi3Z/dI+qDTeSvMB2pcKKLmYRUlsJHKd
WduhEtO/CjgsvwuxFMwQCCXEA5Jt3lQ4KKK0vf79OTQZQfbEjDaia83OPOEnXwNnHJHPpOKBgUnu
C+wdK1/eNzY4I8a9uqwoS/frFV3592aL1Uhgiiq6kj9F/Hqr7KsUgr+FYWcZhIDUzT1qKWDzjcmi
UWwRrPhUoxixZDj4g70CxmS3njzu7/JqxunmRb/IXnco2NYe62z+vMJSDPtvp42KtdA9VvmIZVjY
03iw1Sll3D5RHef8Xgw/XJnyTWhKerJJPRQgEWkAasTBqNTMJ5ukZXY23Wjr2vRl9l3LHEguU2FD
jR/JI6aGwDz9BF7C6Pitm9gnX3atlC1e2b/unbN7Q0hWu7VNXPyYE8WYsyDCbd+d/uuupS9b7cZ0
HH1ezTbhUFofMejsHBvxL0uPAKqsxM7F+/8RUWJ6gPwGpAWSQMmHQGwDNP+xtUXO2c7Ep0HYO4wA
QoFDGQ4p7Zx6mWdLwMDsXjtN3IBhQbjpFIwIZGu2AcDYP9lLrTVGisVPQN1uKPS+fa8B26cO7hKf
XRRZEYTqfV6mDRhfgs36O/yZcBwyPP0mpfMv68ar8hKpuK0C7XSFvt36Ve8XTDMYGdZTxBuAs9tQ
2x5c7lC7JhWhXCzxv0TO6sDLL6+Ex0CxUsNczzujew3aJUEErVHMqjxtceVMNIdDZdrpjkPMAA0i
I1kt1EYFZvkr+kYT+O+ZCH2qRYtirMDAXNtguguXdB+INF7jsKE74JQ9kugUX4GbW9mXESu6uYi1
NArzDv9ltClgedTnosI7c4cDHl9EwgPescnZf3C7tj3pAm+AW34X9vjT2WcdlJixV5qitrwKAWcn
OR1tBe4XcjU+zMuMEMwWftF5qpH15V0nqTPyMdntcmv8c9QutbOX1Ix3plduCU48fnp8NkMFZ5nx
Ogx+3V8eeeoSZtGpnRzaQCQdL17LH8DKAGUzvLrQ4TKI+tBpIZjeiyFcjzdw2pRgAbI/CO+6UkHP
MZu7RZyFLHtEWBP8vKirqu8vrx/35M9FN88NJgm0LhHLSquxWRpm4/79f4xMWxTi3Ksfs2TWhmTc
8/boNWebxbaaaDyv5NLda21D4zvKxdB22oIA2kK81NB+H9aOGuZwAwj0n3sg/16NzReyzq88YCVb
SGuiamz21Oyn7L8XQYZGyDNPNxDu8HjIv71xuc2uY4cmxXJCIQOBxStsNbnglXnhibu9ffMRirxo
0h8xMBTOyrR+zcgGwu5xMh+9zxn+jAUjHrnjz32J3ibHsgmbXXA26VL42rNLiCMPszGV9wBgnkjK
/bXxcCEDAA6Vc6iOPtDv0Y9BvJ+FeRrBSkjIMEr9u0bXnL7cDO4+979un9rauNp2gfsUE9McMuyJ
vXY5DIh9ZGtti/yVloRIoIbNxsrUlpZO3742/K8EYC7SbHXZaDXVJNP+LpAQxySTNMAEu7kgpLfd
1Q6zgvVSqTHSZEBRCscsiWh0gNYyPNWujR8ykfypbDTmARvLnqBIFEGrSe/H8mSgPtl+5wNM271V
lxmdmmgNsBNSXoU3Mw6OsFoY097feYiYWKr6zGGDP2V4PxR5oV/ABk3n4EakGV0zKQjoKBfvni5v
XiqYY3cjYAC653rTWmfgTQ5dzu6DQUR2H0ChA/bCllEp5qawYxEWeAA6mHDwBKAqz0n4RCl8BkhX
ajlP5mM6GIyYk+kvjorl/PHQrmzgzlVoT+X53aJqSyb6+1VC5PbpoOR72tm/AOwU6kEjbP3VBfQN
PvijZshvJFbKoEKgK2B+G3OVHzmBe8o51PLrpPtd0CwSX3YFOWtT04tXWusG1gaoHOoYUTR6nUJj
pmAu6sdd/Z0euOJfzJO+BYoX101rLPCkPsWFfa5L9SGIXwHJ6SmyPQaUtJRXQG6kqcEEomnYOYwe
xWRMIfich0xxoGFq/hoJFMDDrv7KR9pxrZGmGM/ZnKDkn36uKD3veXpGjF2xsoVp0HWJL194MjfJ
TrfxwbiAJm1c4mG9Nrv18V8h9kQtFV/pfZCJE1NgrehF+lTqer3y4Gu+qvV+46EmGAr1MuuGUhPg
RsXOFKjVJ6GCo426CS0PjRJH3ty+sDU8zt5VG7vE9J+2D3WXq1PdQMYb1VeOqNEPbrEzg0jAqigV
6zYHyRmINBeTH1t6asl0nkwGBVPMQimTh9qKHxGC0ep5JRqa0FyrgzSG3ZUL+UlSAIet093ty7q+
Wlk0F8BY6f5vRYJFEN637qRGgntr60XqLnPBQyT46CGUD01f+AlQokSLPsvFdQE9KE/ZYhfCKSH9
L3zoBkW512Xh7XOjlE1SNK3wYdo62PFZ+/Rn5Zg+4HjYycWGoo0wnu45s70ytkIaSNMgFPqvb8cw
BeV4J52C1hsgPB2GgqvvX+dj0ZnfVH1FrfC/hYtTDp7JSuaD8b4R3o5+Vplk8ZNzZDgCsnJA8bR1
prvyJfIhSpfcg+EOvJNu9ClsvqjhPDSqKW+AIAlS8lX5TvDxC0s6DZ3p1UwNR6pt2WNWW3zrf5iY
2N6ATalSsl6tgRdIkTD5nUTlGyMYz3b0HozbK4g5VusuQX7LNzomcyRwk8vYy3GGj8ni4qdj/+bF
SbGBmTw7u19zBmOhc8i/FNTK2HUsAhNzvWtYf+okXKR6Ww/duWksfY6RPzfezeaPd6tUMcAi3tmB
uiwXjXOHEDBVnGoUrg0ZnSSgF8SfwE2qVkgq+YGpg9aoP3RxQehXNm8vCR3XJlA885RoIu8SgZ2k
kccXbqWYMgNEMy3/ZqDbM1mKqbOKH5UnkBYod7B4jQ2+PyL0wXFPy22Mqg/z0u79pnABfe3o367M
vZWhuAGMGvVYJOslCagynsmTOP4UD8NlcfK1mLxVhoSwxRoJ3v7vTVhclXNPKddR2KwYHms8lukr
TuE/u8CmkXwtkeF2gF8bQus+7zdUWU+79iCjaVlUye0ju1slFaU4gtmdGPO1aYK97jm/h2UOkyiJ
9EBFglLX3624U7fF6RzjbOxfJnILiYtOeElxs3kr9Mtfz3NaxWhOpIoTqX1An8IzaHuB7o5OZE97
ud0CBS0z0V7EB2AHnIRnmX9uT8yeSCwMMzH0jlDMpzTrh6nT0ShNyMc/lEruH1Vt7zHFRVigg8dF
4u7K11zO63av8oxPfjJY8KeaCiNfKsa3UHzj6YhoTCmnk6ecALWom2t0faUtD2p8xPm1jomjeg1g
5/acHaMqsQz7GA7SzxnX4zWLRiIj/vHZSnpRGWfDNZevKiMHihzLNLw9LmCadBqOkOe7x+a7a4oh
Zdg8NUxkKvEnwpNMzVOy5nPHpg3BP3j4Cq9XH8nR6OcnLbfbvVoW93cTIQK0n8LodbWkJQTzagRN
bLM5grGnvHakfmiDyzesUtTU/MCxjLteQ+4sVrAD2N9xLv9OWH0/bYHTYBGSpjHyPkADLcALtzk6
SBvSrykyACNfWXQx6KQMVOAcZjNAWlamyvesO1UPbWHbjM3Q6WxdrQpw2SLRYWvnSvQglwQdWhNC
PND6cA84y4CtOrncihYL+WDPGk6xNIsv7OvmWwgvkQar6F/n/Wqc6eA0mltX3ErYcRFjz3FToLsd
P3VoNuIURPuRMAVo/p3r2TdyCPII95/Gbnagz2EyYzqn+gJaIfTp1kNM4ohmimgmro7Q91ewcjjc
TlTa0aC5NDpUMIfSjQSlj03c7QZcQISvnqy1/kSy9ysWWpakxN86YvfMExNptyTrhyynlfOgc9+e
D7MDVlsdOkFuB2ixjWfsqKI+A5lk2Pics2g/QtQLYbIWkur/FNfC0ad2/QrGnUQmuzr7rn9gBp9z
FfjiSbn8iKzELYZQN9VGaxEhxlSnSGqR+vn7sUcAbIFZWNLClKhvOequGTl7XEn0h9JH1teT0QOD
frq2K8/8n9WZt48wFsEDdEp6BWJ/8dKZcEQBl7dt9wDce6zVYIwEXFBMKxdQmVXbuA/HzvCVOZ/9
EFrsiE045dOm2BDz8xyYZ4/WLQFKt1WEj92AWlye4xOYLtQm5AAkvxkFIMEKz+ElUct7tzFwVHhP
SWcabX9x9eg6pWspG7pJtIxl53YjxhA8r/06tw+gwd4v1OvpDD21za7haYDYuxIgNiXxL/R+hCEa
zOsquIOypRFxtmvdZdcCTlbl0c4If4TSSdlIoy2oFmjI+f2QhxfCzAgvzzooen7ptGMxdZRCr9nj
uiIwNIJx9rvyseiuNHi5DqCaQxjefSpXx1BIrgnGXHyKOnnDnvVPYcPmQETpGrX64u8X3j29aNjZ
Yb8b2hrvQlMra893jXOKdiSJWWrNqbKC+/WcqN7XEFewYQJ6NRqAAmZtVicP07eckKRGSHkP3y2X
10nv1oonHsH2T9/BULkZkLrdnRGFullByEwSY+TO3GUqM1b4ft8OduQ6QcQHM9k0h9A+/L03sYo9
1xUSk64pdNpPEZ3DwiEXtowRV3FN67Cza2iLzO4WXD2QDa6u9kabXuTKz0OeDIuWM2HFtq0QeEnR
kyqQ6bF1bKSuODXp9s6Qe1kC2upVAcAHE4FEoXVeib1OfqAKYfoDQ6wvQPihFc/ZMlOGx/2f+NHB
go+e2vYHJYPRCqT19PK6UqMW61+zx2dr63VmJ3yQTXcu3kLhCtGyAMSZJzJojM9+pPLxf374Fy49
S050fzLdaTrjBeyygYft5V0mhkhNtNZCSzVTZ83wXtkbkxcQ0vg+8F09r0KTsH/J/TakjBVy39HF
8B8HZgmXGCK0FUPi5aildSaDe5hhbWp2vbnu8FiufE2/WWO/f6jAuIAEhALKO6CpnD5h0YT8M8m1
Ivo0bg98Wa51aMSV+iXouvxKXjQMlpAVj1DaRPCdhA2fh8yCyTxiBFsdr0cvZ8souicbucKCOvqw
oqKHEygvuzWbzxZK5lRYQDLaJXvAo9b1BeN4cI84twh2fFlTcj/ZHhOBCAMPG+iuycYDMLXRYVWK
nDKAETD7oSJ+Z3IFFKFLu6SHk5uSrR1QbswyyXJj44wjEbElvBsXIbxMrDzdemTPpE4d1PFuPLbi
mRARmNsAC8+YCJpzk6i+U4P2p58ve5tYBHxcc+c1QI3wuI9GdOrPwNPXa5U73Mxervpp/KUdBPny
un9CbWIlXqhnL0LDgF9yRP7IqgDhIGPtz0l6Fg3NT5lX74niSt56wIMxIrjpxthKCCvi34dHWz6L
foFM5p2EptIWm22BiteSDg69pB1ckIo/BItD2KaNjDxxhy5Waa3gVb4+TLL0yIrGXy7lavhk3KeJ
JmhY1yL19WlCWK98M8f9hAT5dpzoDrkn5ADU/09hQNlfzoQ6FLllZxkU4loAw7HmYT3ENLWqrrxq
d4fDCJZpeWlm9tRUZvE6req7EtC1DfI+hK24tRLgJxa0RCTQDk6Gb2zSOdomUXaEVOyFefKB3txx
Vte3q2PaRwcFg6a8opVQ8eGm5VlUxD27LJnXRTk44Paa65cfRDDLJ5cwiqKZpihhjSal+idcLQJf
iqbbdKlx77SyL32KzGG0uKaFmdNdnKsHBvWbpeM5oBLFYCMLaxUdANg4/muFqHUxABgU3/2z//K2
BzED1tjmIIBiiBAarF3oj1ynNx2VuDITrNbtOmzwJC+Q6fC7OzDiYRiCegw1gYHDM3PxkgwRHEOv
OnKEmtqNIZEzPr9wspnNqwRn+PvGK3ZrIEe4GfVHcjCKWotPwvoosKDBuJyGHLJdW2IOwgIe1u4j
kFeRxrtj410ZRIXPCdcIzaRILoOX7DT1aHVrPgdbDHOps9t+NEiiBCrrhzuY7sghuJvkuwAweiyP
yytTZfnT0q0BuWr2TRmCpp840BgeGz+miumJFI8IHp/p1k7Ost7+y709ADDjioVl6fxKUQAsFQ0A
Qt3SJkXrcbyshvm1UNKDaT9QIWulChLfWHs4Q0Sjpayhc9H362gJCHuhGbVEjlsvQIjaLjz4Z2XN
Td7BlpGXYqMTZB6ga1nCOfxzaauS5dg2MeknO9bvJ99EwDfbkRP+leD78o4OugkFVOri6r0yWlqE
r4rk1xo1BCq8DwzQ5bspJBQPrD2geLTWWUvbZ7lCBFEnNIc4DXnAQFfmeVrOkI454zzkXFw1Tt5l
7M4LLpDHi2L2R2aZqAbhVntxuJU47D0lT9pzpwRVSUnacmi8bYHud++4wcVZks+GCKWhMJQwJmcI
wGxh9zb90Tm6+TQTE8S9ZA0xvkKLkqqKown3sZzu6rxZMwNjnlcTYj1/b0RTpWHw3Rq6HgY5sVKk
pqX/GsFjHnAVSUmCpAFEzCOZj/X0hIqcZgYspnrP1hx361b6F3zrW61wWqilf75iAhEuiTXcJ9/R
fzcO6lnT+TIQ7LzIhu6JkmParvJsdTWBO2BqK6jkIxgJ4ocXe+aqpthp/XDUrzdiJLh8tu9FTMNb
aV+ms5+VbktBv3P5xkoR11NYfcic3EGfizaDBCQ2GgLItp66eOtGeSz64dJGxHR4S6EZdmmDs+Ew
E9te5z4bXDSiXfFvVg9psJztp9mjAtnqHxQ/mnARwnQfDurcAv2tHnnhlLob1o0mHNL7Ya/UoOAO
7k1G6kd+Y4juIm0SJ/YYG2vq6Mh+ybGh4zID102CqHFapv80ouwe3kGvwpw/M7pYf1wGs2e6vdjo
C0ZicwjohnTkkCP4cbpXo4erjJmkDf0CLH1jSoqOORCx5+GfxdHuuHZ4UVQ7SLJne8kW4ZRgw2lr
V2pE3ChWjY0nxQJ8ock2kcDCMA+GwhmPfSJsbG0AsL7ymG42zZ050QgYfKsr0z5+4FLkWlZK4e70
inEW4ydOjhM8EBKIMVOH5Gr5kL2BNRc0SlLx0t2uky3F8bZBAh08if3wPSFixBK9pDjtWEiXl2UJ
fchP9QteKGQsruXaWHxV3pY8ZntXnTnR1L+TyuI8S52ToKSJuC4l/NtOgWxQ3mRXIlxq0xrPumll
nQQN/UsMxQxR3uf/6bhRwchjdcZgA5btx70gWaNitjP8Jb6BbRYiC0vWhFxio2J3tyK2IO9OU17a
ROML77fGOKRwAzrwWCSsMAd25n4St3t8JLEbZqWJw88JAh1biL7tRAsYehoodKpV00F7oUECFdN4
FumEj+tKhzsgAib+0ff5eCzAiMfqJ7AF0cMg7td/Dac+Vh9ic/LLDaOKCJYfTyr/I8IVbChWV48c
hrF7YM2BCDP8HZEHBUWfX3CVkIMoTNHoT87KavQYycoZE0JIL07QLpl8IbHlSagINssDGwThAFJu
/SYeeWt71nB6MJxZgdDcPuKjeoWMPSGy8/R+yN+eYBc2JUMJv3zP6dFj5jAaGHk4bHVEmqY1ssYh
PxYiaPUnZYVEeffk3OcJo6IRGDHwXZjvq1s3jTGt8JdSbEnGWvnmq0e0UT1Y6k4S9BfS6XD/AaCb
UDKAZhQyRYl6bnbJktiduBTnmRlvFB8YJ3ZMB/tzWON+WbpSpivhz3t7zn7ouLjqt1bXri3XRoT9
bMBaAppaBbBxVqAc98cAr+7iReq+kYiKwjY7J7DxZY0WpOMfmAYFR72NybPUE0v4TmCfcYS66Be2
ov7GzM24jAIcCCT04oMgW9mVicC2GzWjtzFsYrXHWRFVN4i/rPsmo24hUJPhyvt0ktk5ZEHlXQPO
eWQrRn5NMrrYo0qu1pcEJFvvEgQzF4e47NwlEpQgVH8W4NB6Tc0IITIZtS0OlH8BNugp9WDjgUHs
OSnkBd3m6+yzgnqILjdWep38wGEUvZDzrCYNp/IOHGiUSSRC53oUT6eLxpbX7mQmwb3lxuF6Dp/a
BFEpnIczXYsEBLWksMZtSp2w5T5jgSJ2FXA7gqQuCa/3ko5/958p+yfkGtkXY/2VyMPvxFlzpKYj
K3USI+LoHmRU+/p+E+FwALGyCc1NC1H46gOu4LZ7UvPA0KiKpysnhrKksuZy18aX0184Xlzb2rnl
dUvrSZLYBmcN41gpTg1iatwPHulmm/zFCB0pMs8W8uJmJ7w93KxLICpB1BQ5ECrCbnfFdAQbeMdK
nnCJBjyKrJoCNC+dV7eSTJhDpKO8elG0q9hgiEdLnJJQdJ7EMSu0RcIbbpqwIOKuSyZH4Mno0pAy
lBMMnqlbNImQ6nOW5UwdpdCV3Jert+rpGnjbvFXmuZk3N1tzxX5DV/VR0UQCERwk4HVZpN7D6RtK
3mxIylPHUZQTnm8vLO7ht71lLYXneKzHvMsJaAfWMJDZZIdfl0d1AnRIC/+g9+F4DKKiPcUEayME
lPUI3msXUx8eRSY69+kKG594vr/3VTP6HLvfgk7hwnQX9ImPm/EXY5+os66zBZMcieYuLGOLOofq
0ec+pbwA6pHriIJoFyXFdOg2HzIge6mncYk/Yex/sT4uz+A9lXNnrcplNH3iovxJTuSsA9rxmVxy
pog1QHnhCpxFFtw8gNNPArOB7KPUBFzS47GkBmZWoIIQR8DyBPDtsqU0y5g3WXKYZtLFnm54PuME
pNeMVCs1VCPeTzslHy+9rAOsSbG2fkwBH+0Qs1/biTW+idGk24Fh3nxBDkJ1N2mtsHeXtcDByOwe
l7lyoorm6lauTl1xdSOHwbMlxxFe/4lgLQhCMNO5syR7AtXMsi8lI+KmGyXj5QnsjVZ/w+nH9nLR
ivVw0TWg6OQaXfB0aXp1C0/bAgxJ4+ZOvqP3Ft5k10kYBNHZaOaNbYNzgH505Om3g0P1aAxpmrzw
z8ubveJs8mhk+3KZs6dmTOcax/UsOv00pizJyJkosfozAh5xcPXxN4qcrRLbPFX9Us0VHFPRNuV2
nTPZx9Q6mt+3crBvKwtV89THfu5PkfqdGUum4HxmXCQxG9/wyt/9Z9QP+8Fd3Au8J7XBkFCTatnZ
u1RFhLMnv7QPTmnokRxMvv43ucGn8zocVSxWp7SB/ScccGAnm1HBCHRRAS8/KseTh9iACx/Umf7/
DUQ5bVrLFBfknmXm6adRKI9WiY73F0/PckyPWKkQarGjwXgbsRJXwRquC3Vxs1N1pJFs+i7k6JDd
suXeA71xUMpw66PVAZWPr2V/j/3XE0GI2rl/TRSCEstRSe6A/hbay/xWmAdsJ5QpI0qalQUicqAE
rxxB1RVf+6xxvVRj9kZpL1Z0L+EKy8m0FezaxhK3M6bioi86Y8uCVhB7GeNxuKFe9YObeChnHeC5
pXmMePx5cfc6NPDHrMSh01WK2DzUPz/cK1IQHfaWBwctO2kcubQVfziA4WewvprDhUJ/LB6F/5hd
bgE8uaV3InXbBwDlNhThs7vbLDV/TTN5x8Rnu3qtC59QXL0qWHB8U/a5XISwZQ/6uhyqM28grkzx
m7VejCYzp3BHf+4+I5d571Twt8yrZ36oMsyrlIDNvRArTctLgsEXOCY5NSPcMKaZ62I6HxmjNHtI
snEKwwgwnQjSzc+VCMP92xWHDBI4EPBvNJGNSBdVJxewFLv+APB4Mpx4p4TJKBc++YIilvX1KBGP
rmRoZymIDkmEa7/Sp9H7/InmlKNmKzpyhftUyVpcOlw+OpT6dWoulZHDlXdi2cHdpYvP0igJbJAz
YUWVUnxhdnv4JqOGmJo5W9N4luHkf7AIiep9lGUsGDWzPjXwhB/R/eCX63QUTLUjfqLyCLST9+Wx
ym3bgumMoe+ud94cdyPLzCgrZXbN3XbVkOzn5xc4e06nYG/XnJjYC6vaEhNr6SA6yj1Ic9lnO2+D
KFLW8T1mpIAVojvvXMlaFl9zvaRLWlSTzCwLb96GsS/KAB8h1rSctLWe+Uy7SG0ROKL0qHlKdoN/
cVRUdI9UZTcZbZDha75rwHTePAV9GITBDlYzZ/kRzA4GAni9FFI75jk4igPuNQH33Qn3btW7FVYw
gUMcNxofyMq+vOPm1wMopj/tdW9G7CS034ZiIGY5sOhI2e+TUd0+zeQp0v7faxTEJ6WPdHOkqUMz
VeGl7qY2UAglrr3uREyRpkmDC8B6oW/y5N//AyPey4NglAGYF6RwO/smhnl3eKglKIPTP6gquxqG
siTc8Nw6H99VDqjYanFKlaScPRKrlPICcpEXEXcD09FA6zm1i7KBqPs+hCvkG7XUW8Q+KEq4FdUb
wOU6WGk8FLC1vtbsQzXXTfnNoVa+p8ArP798P5f44hKtsLa/6hxG+xJzi9CcC7AaIRqiFbyF5CAK
5iEBtx0GUDBq2JXXT3WDzqmpAmpaf/uV8ZBuVPPRewmM5/5qG1fJIFMkgSgO7eEwAVRPy0Ayz/r1
LhVZ7P6yv4m2tARZV/Qorwqs9NGbX9AFQic9usbtwZ6ZrV1THIOuHcRUrtnYNZnoZ6d3fX7B0KAo
gkgs2pwxEIgbMSh/6yiTk4DEx4aXo4ncJNCjzozD3nrvBzT78H6p/HgjpAoPV2dYyeqK4qodmHaT
meLhP8wvpYCGc3xLia0vbDoqlnGGbr7Mw1DQN+2uptW+bTjetzDm8/8fYcppOPFFPlBDJA56oxov
f4R14XE73FKvqHT2MQ621kHjZpl5ZJ6+KDDIgbHmc14P8bixuRtDsPqPpT9keXP7SF7zoJzKN2zN
v1UtTcAamUWpYGvEcyqi6SE8SKFxv0XUx5OB77DKVl+AUBXjNvM3BzeUOH+uxVp7ABcGj8jitEws
vtVuQMncsfjq3CEK6jaPNKFmkz9j7ODxtQ5757vJlTbPfoguDV8Tsgh12BtwzBFTBiw8KtNiOBp5
kYGY4emYi0PR/wkARpFsYMKZQKyCnoC+vlxgrfLJciQsnOGIUwaoLHSrcAgQrD0HreVugosxKMWY
AnEdryfjpQb5U5AWDNiqOp7BAlgu7CPmL1c9mEU1s2MrwN4FiZoljL586dQMBnsRdd7/hG5ZGQj2
6YHHm+LkbXGE6XDQpcbCE7AHPzNSUGoG5zZzoDaIZsXHICQWVN69oyxCDiVaUNkqlywqRplzLSDU
lwcBo62EyAazvzf8+Pt3B8gsplB/U1QPbzGYccUjdIrzU8DsrAY0b0LPQkRlgM4UkbpooqcYfLn3
OwQtCPYF30PsVUrJSz21rhFtcW115HIcD8uYMnHgOYHbPdTab6dzQMsTplheMF1mHtMSwFBHRiBx
CF2RLda/lkgUTOtPFJgDAxxHPcTsY0lRIDXtxZF49PsYVRIEnIGjJnd2OzCMVeHPbaO32wXkf3t+
KDmYoKzKoeoorEraEw8HT77x8yNy2uFLQsQ5YOXgD0LYIjO8oJWYTjAYkrHbbUf3ipXeLgftvPTw
Ixi41O5EGhEyNcMsb+8cahdRgD8zl9zGVHSJCp+VO0Ho1w2W5yD7O01btEMAKCEjiD9jBYRzia94
q/xzPVQ7BMf8vkH4/QEEXCXDQ2Z0m2DK+S0M4Kkl3L+9ehXO7mhsCDcoRMqQTKYQqEzvyS5DhGk1
yTopUiYeLLC4SBv8QjLEN5PLypbn5ktH38ZQJ1rEXQ9iqZ2a0GBevk17M40BUGQF3+f3qp5St99d
Ly1qNKSepJIMHIETDXLfh7dHr+bJoZcIsRWUKnzL1/IkGtLisbUjPv40r7nDIQdpe2ls6v9QF4O1
TrOKF+OcZkFJDWLM1WvmHSpzV/sK+l6laTrvwWa+Kg86GLsH6Puxfox7dK8JManDtJCY1EVBtx6a
ofGM6EzkAYJmmSBgQq94xMifqE3IxyHEaf/iG0Ot6wafps22ihSu7QKdIDaTF28G/rzY0yKap0Nl
4eYV9f1kAFcEPHs58Tkf0+VIpiLBUQwz7y4Z4kGuyKiAXpQQb9JaKGJL2e4PJPobywIQ9DrIYMxW
fiHaWoYaI+Fbm5p76oHrUZPC8xBpKlQC350856VP27N9MCbZ8Z1XFY3UrCnbVq4ADvmIoga1i1lb
0QqqZdcFxaZKxdf2/hxiLGmdIk8qEgRbA5jpMpwMl0HPaECHEIf8FHiqFjLG78z1K0mA/6aYfn0S
Q80SSgiudSPEJL5tnO6VVrX1tlnA/uUDWnQGVpbYVg6pDh67g7FYuL8HW8sLFxPHSp4eeGnyzdOF
fJuQx4YsXEAchGum+d5+hdwQCurITHZw8j37aRX1cnoe4VNr155GX/nuYBUzepd4KXUa32H4SXif
EWAO5ipSOsw+r7EEKZOZdjOqU3B6x0TcxpOG8pAVrEKX9FPHIYSOqecoQJX/JZrEC/J4rV139vWh
TRpwk56ElbB9ZSBd5YGxZdoS2pe0ag9TcKM82tXJwmu/2PkY8ZoVnQBRMgMYbd+ZkKiWUhNGqrgZ
yZlQfJdOBUwGufURsZehRttrArk6qEyN4GlhTmrz2JNcDUf/kMFKvH5VPBusw93ykcQ23IzoSg4+
hPwr/uFPzezF2yZqnOMPKLaixOzAwjlpk4S4pScjfEHxTgVB0sqQLCYgAzsEHFS9vhrpOEJINVVj
6jq1aNd3tgbPlmgQBIoSAS8NPgS/agMHY9IS89rocD0ggbyfORIDRhIvf3yuzv1Is+f/vnBawWfb
Hvd8XXyIj4+ZfAKeu+GvFkJVy5iSInqw5Bu1kg6VsnsLPnBz/WB/toInSOob8PBchlBrJhNCETUT
sZ9dSyngmG26GMuS7zyrnxK5Boj20pXQ6OIRthon8OgfsltoIN/wuw9E9yne5rX3jJpviU77FpVa
Mo1hu4refSbbDihKh0sObhWu4ZcCN0kK2eC77pSK0pH6EjJ7b/M9+6AK729luV3OvishPS9cZzzk
mlpXNFSJIIcqT8IpdSUI4+awdtWtGzpFw35cgu//KsS7szRTFZoF6y56mbBKecmmhPpvGw8rOZ1d
IJQZVl+paYerZgPNSRhMSf5IWS7CaGBDhjQUWDak0Bjx1pD7Lz/4CS8O4bfZtR1UzTgBdxOJqswG
fTtgbdnzcZYY8X85ih+c0Wf2h5RQoJrFWo5wkvuNq2au9zdnMvQxzLh5TO47uVAmfZxUBMF7hDGa
/59entC+e03pz149AoF6kzy3bmpoO5EDsv8TDVZjqdAijGKcLN1CVlBEhoGLpbWuI7IFsRJEJd5d
ivZHegQlyhNppFaNxsK/b+RGAUk7Q4dIpU1UneG+vXi38btRa7WS41snMf0CPBA2ZagSltmlmOUo
lZEevGC7cr1DqFHUUfdBO3Tc84eWyOBItbFIe2ZD4rlVD9PGZvhL9rn4kD3X62mGOTReDxklIMwo
FJ22BHXMHDj+177M9PGU+gzjqsTWmIGac04NLc5cGsroiHZHsHAJmxGngMhS4j+urLaQlgot0TqA
8V7ia75XqRVxj72OFMZQ2oazLcQG2w2OeUnCavRc0tq+D7gD39xgF0RrwiPn/CVyhXYj2wFGVDST
Ovv6AUvVRHUBZIOVPkolUTGrmZQ02oktgA0jiwLt5RQI/jHENNtRoOOaNWKtQKeCGeIFd1h/6Frp
clql1UBtzfivRBPB6kxMIcmT3u5G7OTyoFVea0+qz/EUTDZeOW7aZ41VtWJToJGsVEgOSYS6bRKc
glajmo1oSst/k6mDYj/4v/NroHn8EGhVXuDmcIKfROW43sgJQZDNjPEjI5a780yxTR2cHOMRocfR
JVNIRieYYlZvzGMy36XasHfpcaU5qIS0eiieAWdDW0x0bPRzH5pmbMM/Yv4vJSUpOXVVj1aSvDhG
Nux2FUyc5j8eM3i4r6pjuFihThwo2v+XH2J/2sbxBQntACxHVTRxe0K0tlJVt7d4BTbKkJz68m9t
YFPPhI6EFan1lwQv0YUlBiRKUYmGCRhK6xeIjtfUKa9G4Gt/yQyTE8387fVWopA9csSETc/t2zZK
CLF3m1Wglt1+OoGk9JhScdPQh5kumNQ8j9NfuAUGo7bd7wTt2GOyUKrLnvPpMn3RkqNHGBmFkOFy
Uw6TtZUhjVdoqHMO3vNQtQjJWVgGz+eIyvC58GRHeqnBXV3hfLt7lDgiWhDj3d8FZlwMTJMAKtQW
OKX1yVVBzqnf/QrxTEbyhGMKMmko5pYlaoCZHcOTAf2Sc3ZnVH71ZE+ujErNfLu3cNe28LWN5QZM
LKuRq/Q0KDcbUK4dOnP1hM6nB8TEBegXQB2VShMiwjyIBVH7qlt1IfZX4eIu3KzMCC7+TY6kbSt6
20SI2O38sm1srGHfOaDrYqEwcrFauxLiNXDN5055cxOyk8Tlud6lhHe1KjljqXVJm2Z9/2b5hujl
lcNybd/8DkW331zsdLfP0z6fBSJREXYwiP4hwAaGQ9ERMWRUZUoKzwwbl9tbChL+gdQ9AuaOk2xQ
qoVhHOeb77oWle1yG2lamuf9b8Zriu+jez5AG+ESz/r1gL13965aSSMPR3CRWF6Jt8XuG6l3G3fx
Pxvt08CAk2iMpCpvfMjNCgk/E6TezoGdNTfsKng+rhRDKSmFvJPhHft4FLxDATRM91OUGCPa6ogD
hz9cOeQW7rqrcdtpIHnoWfbHDmHIHmqy/AUJYeh0c8nT/lMFarMBpzhJ4Py797qdEEHQeX7Bnp28
sEWf0ezVQEBFGcY9WqTVtT1lVK7mZcVak54MGcGhch5TcnwZlNUIMOrXoZqwfOttCuTTRG3gezS3
h9/L3uZ62+Epll3Jtzm0IQihL/XGFgsTQYVR2SokdWsdYuoa8sQICOBJxMMgt/9iEZ37/C39evEZ
Kmqz4UBpWP2YoK9HGmrxsijFrjPquoNbpkXkCWwiGqjugNKA5fFEf/mtqYCmhBja7xTIN0nmkhHe
8PyF6SiiWkldyRHw0Z/q+5xyCdr7HdGLhhzqDaAc13w6gXzwbK4433+OBwQ+z4hYYJLpe0/obzBe
+YLa72//8AtUhT17TFcMMfTmKKGxP4Y2RmuxJkbbP62HpA9i809ziWbtk00OivntC8I6MHLZwUX1
0Xelxe9TOXS1OkCrhRmwacPE9ldre6QDtsGwBAB3f+Pmvc4qv53LiGzWZ8265ZJ68wztjThHcVyJ
Go2UBfqnq7QYaihfqUfIDOR4P/FymFgay6MliKtOhOidiRW2RZmwGdB6MqFdZUqoTs4SqrIp9zUi
me3bt9qoCuMNJ2WbMALb8GwCg8xYfhi/LVE/m0wo4FvcHQTqmhpb6T7r8vUsa/GXQFUumn2WJ3P6
0T0Hc4P6AhUoTHGjZkaUCuJ0Q9wds3m5qHwjUGaPnrevlSXcz8hXE+GxpdSD/+S/lGShddo0cHNn
330q2x4EVEcQmUjt/IN7eD832d/u7diLOt62nD3QxSDZPdb6q++pFSOOCOL4nfGwcMPZEa4A5hVN
09y00Al27d1jaRy7hqL7IMt14vsn09YTnJEBQ03sPeMMY8JOTzvOhzqw7yofLRQvUNvogutKGxBV
riCKcVX+BMKjEBOMQEQeeJTsJwK9mD92SxSzjHYLyRUWgnmizrzKbecdSFR6oVDeX386zkFu4vc+
f5nZT0xjv1tW9BEVy2IRFBES0tDjeWhxTgwf6NRSULH34bST0Vxf9vaPLk0e7O6edaPVtY3y4sWL
a2WwOW2rz8reB2TyVrQc+qsmVs15MulFrCY8f8IzqoKK4Py8wMPLsgKJi1jexHWdYX7TcE3yODDe
EDZgxdU0zb/XzO34Yf7p1UUaFiCwvpbrb5NWy2+Q6bbuqTyqmhY+mp2G7/5NcKBMlRE87GmZ+2ez
ABSOJVPjqaIROs98NP+Gezj/w5Zo851iTC+n/rE5PwhmtnYc931Zoc2ql949SsyGSxHh8BImmXQ1
tJyN7yEOEAZGu+iqXeYRb+/1fMltKYfyplsPPLkEQkV1UAXT+Jo5+zLs0fRHJQ1OFJ3VpKJaPCG0
4t37IjtWIMJJOy0QIi71luBvhtmr6i2ZI2BewpW7pYiDu7V4kehWwrx92UjhVkcjburdSyBBy2re
P81ufMOV9mqxYKctIMrWaOHuI/h4GFLY8+giTnUU7QDmmgEWgNKdOJloVWrNAn1u1O7IuARhFsnG
VAFDgVxkgpCN8+6coAuMeXlh01eRFS5hQusT1JKilq3HQQuYe30GXesTebYweDfKHSMs0lZ0NDH0
OO7feQKNWjH0fJP5GmcRJqRO1pJ1ixo2/G6l00n5R7ilewnpulll4vphz8h/7ZhHzkhFH1OURnkt
EYSSNhEzW076PoBFnCXhY4AU3e2U7zPd2fJ6szTwKhrgDLRGJ7EQApoY7tyAOFRnp8dpR5MH5VK0
ZNjZVmbj8+X0SE+p12hj8KN84dMMeGZ4BCrYyvgzTFZEO/0078P37N7C/nAe9vIuX4CEVoWOJ7Ib
TvtG+t1dXiEAn8HimOc3RZ+44b4jViC6ScGQ90MsYOxcsta2VoHo4vttkr5ouR6dqoofolfqYvO3
4HTONGEQiAI/cOJp9KvRDnTqqsBBt+DLV+zWRy42uMpvw57HT41PHmCOiiL/Js9Ib474d32K7IsG
xlV/xKMozsZwRh2hEtESDywveyDWM6fCT1S30DKyBnGFM8GAlxWEsOR4LJfc8wRqnLTmoIGWl8Gx
3qXHeeVvDHGLLzfSyrYBqbZoVsU0Yf3POZ9WQfo2S8FYSyMh90UIi4Wywkc/1SRNm3Mal7FQJiDQ
PygSut8SEYpW8SyOWXo2TWkEhccLan/A9Y9uiHE1cMvjzGWOH5yoN+zhDDuWrhJ4La5isDt9FQj9
aT8ARjtUXxSrv45zvOy1a7FjzUfieAcfGyQt4l5D/lWEIsrW642YlvHpp1yHV/iTC4mc+ICoPeH5
kqldZFZHnDSdMTHRFFdJG0eu3ZXL5y9mYMhtp8L8g/fo6d8Q1qiBRVHozT0NrrLf8151hzcHacBr
KuRsVGk1uK8FB/KY6Bif4UDqM/XgzxN8lAMQmTnKdLYf6ddAbnX73Nhwrjl5OWdCQoiMWeYJsu2B
mT1Fqgwse6kpkC6zNODlYKrmO3WNVvbYWPzAuw2XHGZHSde2eqHqoIFE5DmZUXgKQfdyojVNlfBp
h+pVYEJly+QkuEgU5amO0y7crm7GnAmTddC1Ok/kySI+6XGhnEFO8WAtt7oxIPP+wmPSRi01VyxE
UgeKgh2P3VmPTYOadYagNpKOfzWjNbbnFux2oxNiz4/RlOs+UkAe9i2sbNsyx9rwL1RJm9MCnP/c
+18+xHzPQzMVRyaPFytISmGZB9ex5wQ/o+pVgASoZNCYKxYYVpbxruWjX4ZW/vqFVDkQGPPvw17R
CiWn+7bI+hw81vzW1U+3NQ1rgVV8P1gmefyUojXnHxLT2kilvwJv1zvCDTa6j/+6sP+7Rv3DwtGu
GJD25gf6VNCzZ00jNC8HxNhe7U69ta+4V/qDZkqMK1aTsOcqM9G/EFcDb5BBQbPOByWhWoXHzHOw
TRXVa3hkEr8Qf2OCBA14Hmn32prPY86VRd4IZBg6xm0qzODzE93mGFXBqnBRhpCc7/lBkLENgthl
nU39lWQDwVgtBSbZm4w8pGI54SGQmVj2uOkP9UwVl7tQ0YUatfX3JXrqFw49OH4Jj32MH4q1jo1S
VDkiEhJirTVrlQRdQUYdZHDCEN9SAtPJMQiVXUv4U5nlTA6qLDDXU9l5nG/0iDztcW+XWaDJaE3v
jMePtSg2cmXJoef2ezZRQHr9F1HDX+IEq2NrEwgiiNblCISxxRpaseYxjQN4yLzO0NoMvvSPHHLQ
tdnbatsOy5zDTKg5/s2XbMqzYXJF/BXJO6fuW7MLaG2p8TazXCgnZJ27RE3/7tvKg2cKMo7if/AP
azhDoAB85WqbawxYgWL0XRvGW9pJskGSXR4dyFYf7k2YWyp7ik5NN6VI3UVXSfIGwHsSu8f5vhaj
LgJ3rFn2JzXc3Ll9OvvMJW74N+nvjTK5BhRv7yTQ/FqTbGArc3JHnYxA2IrYe4nkiHtmjhCMaLvS
WSy3qFOa6iFPj5QvR7nkKS4yBObBZ4h7G6+NfP6bTbo2HhOQzfOwz3Es3BOmmQoIJFqOni3f9RwB
at1TNW3lgnlxnxWpqVU78kGnyPi5kD7Rojua/2FwQZ83wetihNr7qxvYlUH0Ax7XaqsSEndBmRUo
BSkKIyhjXV1lUgBfZW0gYjeG7ntTqG0OhDXkjHF5MZ7gr7AtZF33f1fVmsTbh+/yIeS5sXewLPKA
MJBuA4eKnOQe8Olv/nK2Cpn3/WHs66Wu1uHTJevbWs2Ofi8zgazOpRGhhtUBYpsSNWRpeOBk+Z0Q
HCZTiyz2ywy5bSQCzZraN3TdVN5ROfAuEPZGkRtPf8FfslMmtafsTEfUh3bXbJ9zkj8u4soE4vb5
8ybtigtW6fkELqHiEzndF98+6Yx4mTMorTy2Sf+K2lOFaqN7DFSP4AokfSdRuKlYiP0YDAgen/4G
gj4FfOhO7fvMqKv0fLn7Hzkm1fFIl2vGjvAGLtgWYcz80L/HO8k6S0RbOS0n/pkuGsuhYSYPYhMm
VRPf98oVm+CGwOCTyLtO/LEpcudRypqVK3NjGFhAq6GDP79VqLiv+WwOpodsP3JFT65b61+Od0vt
bzJczVQQoHbje816KhFkDU1NGWhVkFav2EtGvWe/Wa0CNlMflZJKgF4Qb7O8lhz5D+foWIEm4QJ7
PG475tqz3uHt3SZwo1HWtGACdM+iA3iu6jY389yFbMxz+ZH0k61jAlMg36f5bkH2v7lDIBHNdMG2
ZQDEVGkm3NcC4UcIWOT7nZKMIePvGbPjBWqxyfxu/HJSQmcdYmHqcifbI/ohhxSNxMNQF6rjt82I
ksXICm1nHm3FiFY/8NDobZOU4Iep9VaQxgpcQUgD4RydgiUsgNLii3EWQWRZjrAKH5hi0zrZU4tM
2HDoGQ7SQTrbF+F66A6+7iG3PZyqBKXWfyiQkausttzJYXX/WA0+fM0/Kr23oOhGlF9LRxYwvfHd
JrdlKBo6491bEDP6OCgLQZ0IEU44/4qwjFh7o+LuRKExt0pKOoc21S2Wl/86+4RWMPkYWDNjfQO+
kCxusLC+sAkOEDh/i/g17ZOcAK3yaAtbUxW1waQcVLtBWa7oIDjVWW5AAq7dE2rXaslEmMr9vTWA
N1LRSCiULjObnV7RIy0MngIuOMAx8SHzt0ckGaH7fVprAPOEk3FYt6Wd/fIJEyFuKCR5OpMNQ35Z
33VO4f3u0mLu38rUBwiiWz1O7R+huiKqMNE45/92gb+mcYtJmjuNWkXDpdo35RrnfDmt5QtDmu1i
KySOB7Kq1ch+PGfDeUxoJb1dilOGLsiSPv8SwLyu86qEYRjBWvruNAE86Ub7aa6/4ZasfKbLtwIn
30pRx6p+XJD5bkOFKN1Kbi08Xlj6qAQICnNeqFxwN/eruJUoHkv8SGnrO9pLsddtn/tPMfQ5VS69
HSv/VqBInP7bXwW8AHXSOoQeLYgvlHEcmvtMjlV0gvcWH6LbiJg7CQve9p05fQYCX/e2iXFevdnR
MvaE14wQ7NQuOP3urHCF8x3Vpvfnnguvpjf8Rsp0jMC94E4TOpIAT2KElw9N+wb+ULMDmdF2q5ky
QEPHip4ikj306/GGHT6WJEG2CqMd+bCGZSyZEr0lMWQwzSWHFedOfToKEwRFBZPkFzZvJ1rsL0CY
yi6BgQk74To+Wy9tiXNSd4hhnnioX+L74gApH2kr0b1JVx5VNCaUICMns/y8LWVqki9vTq6usaeF
+NYeDwYrzPVA2SWCEti+6gpNNSaYyiZ3zVj1u6JR01c0tWfEJwUg+A08w7+RtdBpsSJV/nso03Lr
NZ56/C79zVEnk6M0PWbVu4hv4Ww/bZ+XraapZh45xbHFPj40d5SvKqwN1jYdXwWRbfWLJPgHwihS
dtKArUpzveQE3YYiVqtTML5Ho7xcH2jyGIr8d4wkviULlu5WlOQLiqwJrVbC8szLnADlTfCNB/E0
qpeRh1QwEptDHOGHtLEq/GyLw9X9BnFqGu6R0UX3wPuyURCQoqdp9UP9nmhq+u/D2KLYDmVRjpzj
1INKVIandDYxKhl/27+D2mZnGEBtoVDwWZVl5dEON4vX/59L5wfXm2AnxlwF2JqTU/CNwA/4Xwor
L8dQVY9xktMJZoQdZcdx44ufRcVWSWqwYVz0y0aw4Gpe4jPolO7+PXXgOk0LovUPMNAEVk3H1t8t
8o6OzpxOX2PbGXLxr87azJlRIQvSTY/Qaf6nGakqYnXwJQnUK+NHSMTipMscZV/7n36M3iLR8l24
/qsyVIjLjYQ8oL5pP7uh3/BmpBHV/2hPJ/Ni1m1WzfyUAyw9gYh0/3UNcBgZ5lW7NHkXEMjvOCzG
7eKU4ZbfFaC7G8jqBN3q2rezvcjnUPIiqFBNd99S63DFUEXWx1MhO5gu73qjSLEqebQDsqgY2YSg
Rau0B+ShBh8AJaExpXLmzbwHyd51nMX+6y8xNzdlEzGJEwut9zUAWejkG5xGDhaa0/eh7ssOYcZ8
8Du+UnWBNYsd1O9LtE7/7fjmNtga63o1s+rVQBoDrp3kWy1d3d5AWvMikLTYBYjPNcuKLoVN1fsK
K3iLwGztuOj3YLVNjmWVvQAE42bZwPzqKZFkJbNwtzeZ/S2uM3dz+fnyxwIU8ewiES+czJdK/+zG
gwwFHj3fqj4XN0Txop6D95ftBI2tGj1/9r2qQ5huDTQ4mVk0CuISmf3WmZwHwqEzXJr3xsQyHsXn
umuukhTc8jnQeJ1uRWMSg0Wkv4jpsvv/c30ZfHB1LZQW8Ahen2VAc04Ha75pOhGSTLNbCD0t7kAW
B8D8p+BKeUHXAvdSmOnQdfDg1Vf3RP3uj1nAI4oafgWR9HETIpJofssiQxjhrImRFwcqfhopJc4P
Y0NH0g0E4/rR2P2h35tbpJxiEMXP7xUtQqZLRswE2pjT8rs41W98cKtpyF7Z1lukQ6Qqm9FuWMcd
i6GK3olaBoT6aeVUObBCsNuAp8MSXdOP3AWAyFpSUH2N90fi/eRJHQb5umBLl4x+t1UH+p2oh1JN
DUWDi43QOOtgnPXkVQf3ymXSMKWxbWSkq4tlvrgcWxfkn3XBaxEmPbySzLet7w9RF9tctvKNjtcl
brwKbpZc0MyFKNd2An4N/EWaoy7ocugPcCv2NtaKT+BV+w8AxXnSbRe+yJT7z/ViMoQUKMSpsbe1
oxX3knofibD3BLozMqkIRqGit+f1fMjDVTwxPnnFE0+gdveOB+tAEKyK3ZTYQZATDCJyFB2CV9tD
dG2orttpeaYHOCEZEWZCF0gXd72nFbWmiYvnmuyDEudkI2IVnLilFVe1VU9tNRsy7uSJyYnw8vnN
BCV7RCDnZWLbhMpky6/70Y9pQW1OTl6GG65aGrBCPlt61ugW9RqC1RjF+liF9+Z2siCpoaMkhuON
vU1brC1bLk3ghXvyAytkywvCb8GpskyWRrlejJe0OLqGFvITxviES8F+m3tWltCQkDkpbxJDCHh/
k7yfxGgG+wLcEsBOj4ccl5bmC2nVQH1gY7vxYq4xXV/6fE7lrP5HNoj5pcFB5pMTT7+LOeL8oVsG
rYJH1ANj91gzUKfT/tTYoStcj9cvX987sAerVaSs3gBi7XuFW9yFdbg0gEae2g16IZHoxqiGcwqc
s6znubh9KWny4HLf4WgXqNmrteSRF/+jk0xbSPWuIPSMAPOWh0+CjD02PND/SQaI+NL4SL/cKG+z
YkUSNVW8zwu0D3TJnmLjl1dRCnd7AtSVay5J3UaOhJtVJcDjqAxBDx8xp59HyDBxYN6GDqWBFCxl
UtYILWSJG/OAjn3IG3alY09yxhyh3K9uLq8Y+U+rBUDTYgmZdRsNHWjvR5yZW8uLAZNJIcsnfrbu
qIUNQk9EgNcwOPKn1NseyaALCmnAyZe2OZfuCqvTY7CFkBtMlPA3rVsILbu5V7Txd3YuBE15UaJs
BHL3bCdRum5/QRUw07D5UBMjgsit6tHb5e0Ex+Ig6rgt1BqIZTXZXeMXHPtSHX5v+7Xg6XwLATb5
ALLOVE861bVRtukJV3fZanWSqTyA8NIznR4tHJl2i3fiXcudWBdI5Tf3YBe7/RMIY7wMWNrweUbK
67uH5UMLyoFxdRIXdz6KtwO/rFSOSl+7IgaGqcRQ7HDrz2XpjShtgsGLMkhMqZ2Z0aJq+K6iIN0s
9VyQgjvw4RReSV/+jwqdNCRgTMP9ScKRoTOG6HID1Cz7iSC6pgyhzsa7wmMCcgkK7GjE+5Lpl4xt
WJJ++i/+NnBeLsF0Vk1Fw95TII8iz1hqMmDSbFQYewjdbmU/OjTfXrCTVCTHNHmmqYnj9wrZC+ed
ezWrIsbr4yKpxJmcez/CRR2L3l+yq2JHj71ggCwzuCJ2FSmaBhfWNvHEFh5smUx7p+Tkf6AKYAFe
ApOG9I/0SFgNjA7YyiF4dGrxOcjkgVoGfj08tW0IqDWGfY1IgTN2NmstGmC/TJ7se5ly33PZKS3u
QY5pxFzlqPt7TikMJAsgKPmHX82XwBfpbn7dRSLKMddOgU1c5rmGVg4mRIMX/t7xEjZGJ2wJMPdR
RtRafQM8BR/VgSfgLwi6I3xrr47ZBCW7StvcgJvNf5YP7u9voSUx6wKF+wM5DIxpTSHYKf9mIHxp
GPfrvXrmtLJVL1OetpLVhc1ty4h54EsT0T0ePEMkS1jtTcSBPMMp6815jyqRdyhwL09TnxXWWL13
QJKNDSXEtvQs+130Trup6Qyp99G0RKh6Oqa02H/3iodCBfGEr2xDrDLR5in3riQjQpUoBZzaaEG1
BRVhecyp0dSQEP5jIpmemPbSRdew4NBrivk/TtNzul3lHrcBcQk4JYIzEjiCILM9e6t7mISvtC0u
fFYhKfu+i/qMrHZSNtkapbrZZvkSG9Mm3UnNNI5OT4ICQhfEzfH2jntjKha20vk+ioc3r9I0kEKR
eK9B5kx7tkE57eyeek8J6mkjMBk6cD+gtRw54hVHMC3bbDMX/H9qZQdvEYhwg2sHyycrH0px1D8Z
rK9aZyfQm34J0+LJs5GSGbo8q0eau3+YJkITTTEy9DWmIOCie8xc9MZzc6/xj4VdLdl5XAJIoPO8
fWa8BHo2bVLqXCJP9Zik1oncsmgKSj+bl9XFLZtr8dP3DL2VFT5VWXASfEmrYndWRhtEhmju1aYC
fsBpFqXsLuzku9mxL07Uu39Xxdk31rZ1I6zLOLhpZ/CmusOaVW63UfRjrl45Y/cOuXYJd6t79ER7
XqRMJUhwxEvUAmVwHQPNhaD7F/HEEsg2PvkhzLKheXdOkVCaNHBbGx0VyTUfPvZval+yqy05Bbes
GeKVvsCNDJLaZ2ZzcYYBcU3xapUXevEoN0uk29YWjt7jdThrqtzhbQQBJBEe4N+3ryTjLf0cI41t
NRHD4i0h9Dv/hhygnwC/rN2el1KuT7NVNz9qiADk79OCH+JPjPQ6oI5xOCS9Xr7SxBPCgfFfEUzh
F1XMbiYPZmRgMgOhr5yVHqJK8F4Z318dT0OXzjKa6lLw/Hj6yH/yq3l+T1NnlmeOiGlXQ3ZA6p3u
Cm4uNecYh44lzt+L/Kke37c8dMw3QlJPHihQ5hw3bty5VWbcAa94dxEnmFidePxO24oeX8L1I+Ba
fHOXscs97KrFOLHzw0JF37C+CIomNQ80ByLsjzpN6OSOSwyVjD9FV4WTm+0e48l+IpGtlfob5Qlc
Sqo8EWWs4rS2Pph8UQmxyD1fP/L4+3EbXw72Ww2CLisv80M/5CdlQgDjbBrbMAR2odMtjF7O1dSO
wOHuqrRLju3KtiOAcGWH2zvjW2d/0F6qBvnQDca4ARvHu8BwtO5tTkofxkBJ0VXnCacLmsTd8DTA
CT7XHLMF3AL4iN6SPw5OTnXsw4HwH3LDYGGMDTJGby1N8PqkkbAjJ8DTl8E27htdMSnRHVJtiWWR
tPIyHXcrmtu+H2C1LngSZy6Krngu7b79lee0Z5OQkjvgHsh8W6i7EjF5Pu8+GWw7QjXm2YyYtT2C
O3QSsl7gcacShIpFqDDiVpyqxW+IIQJNRPC6X3NUW/Hguc37XBV62vTUBdley51yeMDQluiyfU+E
AAW/NCrmWqnvOHqcITGF043SEwdFITe9QgLOiwr8mlm3VCHIGY4gqUMxv8JSrA6V32SKfCpH4CGG
HGeSvrVW7IvNsOjY1dlF8oS1aUzh/naEqvc0s5bnUgkOgNsZnhHPgmTCgMuI5YH+jQCUVHAIuqQ/
Jt4uxqZvyr1N6LxE0+SGMf+6ytQMIyubUNvk7N+91D+l3/lRwYE5YnP5EhOxmMCXlORCR6s93cEW
AXIh5F0XEHKP475zIVaxpxez7HMWilLEBuzswA+oyoy5zPY6lUc3PH+hVbA5rQF00EsDeIJfPbSv
JhsnUMejem67cRfMRWTKOh5TjuPbQDHg3OoUfF8GXpBck7WoZRZXUDb0uxFvEBS7XOfVwzBmaBJF
jj2xez6/QgLtO2yCsnOGqOLQPHDcLcuYwbvhdsNr+5AwYmRuXSpHCYgxkCeBxSogreFSFR3r6Z3a
tBCEcl4+wEUmgMDwyuim4yf2iWjT62wT52xLZ7mCNxJ51AhYWkyz25eigaBn6xe+fOmKRwhELMpG
8tZtDQUPybOFFG2nJAK/yO22mz3on0Ghb4VrX0QVtFMa+3iYw7SK5aQXU8GWd0Jr95Rx8oClC7EJ
7JjKK46oo/U9gesvZ6vkexydQ8GP/OTXKQG00hMqmu4NPR5NJrEGMcwAab9y41iX0HObdE2tYLU5
7o7P60Yd3vovm7uVtI02xEJGsPyfzqjSZqYKH2y3XqfNeH+sIqQ2mfJ9nxh800oc25GmiUB8QE8b
rNVrhzc8kgw2gSOC7pdJknLroFvYW/GH9R7OMakJv017VoLDX43jpXeNsN4fRAJ1ZuirNSMCh31I
0D/uPVRQBxfBeDcKeW5fQNOKd3BPF0+5ZaGBlG+E1SqI3oyEO8Lhtjwsj4Jr9X2xzTTh1vgNX5S4
7dQ8ncnLztGhNeUAVppuvd9YzBvGtWs7AgiFeFtH+Ph7DhB17tPGZ84Sby53RlA5HReCsiTGZBjs
sDQ5XAJrr75ODmMz2KLsL5paKqMTLRhVifqbX/iz8op5VkOXzfLcC34PZTSO3ln/CXj9bh9DCfCd
rS/ddXX12wx24cR8f2BUnulcSUemvDhEuDve8T1BYkXSHE1QdexkOFgW+++yPvk1W2nQ3IwEYU0A
ZyuMMICCfnSkGsI+WaoP15Ni9kj66mutAPjNkQUTcdbCjbjX7uRXwg5MY1UtMMYrNMTX3IZ5NTaL
yyJ4yhQI132bgnm1SEcmeOfwHyG2BMTjt6UJcT9iX/88xyNKwHdwe13PyLHwfOkNgFDSIpGKsUD8
kPC74LOYLs1F5ZestWZMA2tpaopohOVTHsIFrQcrKMhOgtr+qrFABEU+Z+5WjJ5Xrj+CC3vzgWdb
woNvF2JDywctqBj9eZwsrn+wSwq/+g/wY5AAKTiWCEZOp6IFtpvoaRMv9e7ANYAuKxxssc9b/Mgv
f65d8ZPHGqHbiMwmb5NORyqFBSTfpClbTZseFGPlfl3Xi/LjwrgIqBBiC9DmfAi91kl34Pd9VqfR
ouzONoIGLEAm42ohLIlDbUiPG93Yic+OX8+d0WbG2q/tkUVU2v77waHLFY9H/x+pzIpnTEM6T7Sb
Gh0q2T1Ndm+sgay2qBks6MUu9xJvdRYVTa7STsC9WbXU8kAAYGqaCKC24NRllSa3q8F4pzWQK3a+
l74S+5xqBiACYGfTuSQm7btsqIwE9tnOLgNtUSO8SriIDB+7N8SFQkLRb5FcpViTf14BDi0CyEpb
cJPk47nmMySUz0SOKgSKEwd4wXOWqXuHteeRPgSLL5OpubB7fSFVvUweX5BFGIRLo7cbaCVDFgK/
SGhvIsHXRf1GzyvB68FLLT+zneEF+kA7pjzoaph4CH1HSYemDuAE9e1Rv282yXbaO5Wf/eXWO+1E
7NMhsEc0XxZoXwNDmeMLRTFW/3C2ndArwfNFZE2uD1EZOgdSEh0/Ma31fq2edjf8QOfVNUWCnL1C
cortwJokz2UOzdFnu6Ana7mw/GWsek1BEFjsnEDiRaDUBLKGCg//DDTFd4JdsFqWWvZ5sgw6pU4R
dTw+5flCqwzO2wzf3yvCjN1u2+nxySJw9w9V+nL9+P06g/MblbBRqV3uGLezpCJkqpLrAObBCuam
If5j2JK05rjGXgcggvu68d0qQyDggEDN8dHMDASgA4qpM+7wVb3sLEo8npTtSFkm2IURBAxR88Hv
rqNujW+wG5G6YSOfzC/o/kujO9UZLP8zgCeOVOyfzqLwAhoKX99s8f5Vjopp+eVXUHyvBOfkBCM+
2xeRQpSEsttPj4TGXbV2xCNLPMKDKljImmqluXd/NPAu8fIxB/xXl/bCYzxPtg+LD6gkhuvt2bmF
kQPQQm1fm9aYLY+ot3v7vc0pv2Bp+JK3Hy0IDakQ8ME0rQCpIBjVCCDBIIco9p3RfExfTDUQ1Nmn
dRt/zy9UeN+rU/X356lN6rMsWBHYEs3Fqshvw2c7M/qLsLKme0R5SheBWLRmc/V8+Z0Ke5P9TLEP
KAztFWPq5AxYC2qT9CVn5KkoQNZyN2PfcP2lfqfea6lKf7pAJKtTeIKYncnchk2+rFcNpjKD00Ou
YjA+gcRNcMUxGxsMRN9xPMaDNRjwPmOVkDHfhuXwTqPSec8lIYtEnWjwU7evpHsDjQ94Ad2ZXpXY
D6aheZToiAOhRZp5BgjPNGY/LOjKgT4TaYKm77B6A/6jg3vbIC5WC368wKDnNgf+YkBb40c0ti1F
eaN2bzkyBr5mM+9J2Hfyc4dhtm+KANm1wfibP6QfBkxf0Cg7ah7Qbii7Wo42yFMS1ktjtbAFWczM
Z5FH1wNRBwNmbiqwwxsu1I60A7oglEKpdfPilTdn0C+kc+giYh87cWHRlMfFHipZdWQItFS3VgCS
Ecuj3UWMMhCNaQJ/t/OHkvPNzRSBrSqE5qwwCGICwM2ky/OORMMjIjNKUd+rbKlJqKU5AF5ZtVHy
smStynUGVCn/9LvsdhrjmcL2ctfNQEOLS5SAze84U85RtZS0XVmnLcWp0V6pBPyoDbjwNPS3wfpj
tYuK0cvlJYeZ08v0LTwLAdEhIpRyp+tD7m/7A+IZthoS3NJtli91iHUcdYmBuzbGyPJail5VObAa
DsHo9vNI6zYTHngO+OF0xLZCarD251jZAau/+oA/wBUb2L8LNItQYkWzllhhuIIbnnz25J3g9gPt
W7iK1EZIKHy6+kiwcs1yhobn6dRAnnmXXFIW0OZAyd3Yp3zwVYpc/Gk9NPdrWPU9eIlIrEH8Z4i2
58IWGHOdlCZtIBG4odxBybID/wSIIRQWbxSrY9BWUJSmRrGbOZwHgmubyaHB9Bs1VOorz8+QVGG1
jgW+318PBA/Ij5oyX9CRgkisx47ZId0i70R+5EAte6EI5G8dz+XqUvGBJ5Mh5xGud0jxriRidgKb
bqqP5h4O338aKiDALSflyI2eDbsCd5ogy6uyIZZ3Cs3ubg0RtDMwF6sN7F+XiyfPBZrFsTe5WKYp
dTlh+KziaNSFK/ciquZ3U2hMNFFwVH4jtMV+deYPiBoRqlT90CX2eA7gV1PDjPYJA5rEvp2jcOo4
b2qaQZr9bGglMVTfS7ck2pXDvq3nWTAopt9hxjpZlC7CZV29E/fxm9DJH0mqArpCKlMhRvKiKMe4
nhoILYDFacZMfNss1Ydn3Mtj1bjRrsiA6XDpnmOMz4oGR0KLmPkMaU0KSazZjFzv1ZhTvQuoNAUe
wmqytsB0YULxQP7hHFj60g2UPPrTmsw+1o4DKnBZHIJi1AsmUy4PwCDeyTPMULQkCrIWZzCTtcXJ
ONUOAm7Xkgycd1mYgpTTTw7sM6BO5+au3AjgtuXWFNnKOnlbPGKmvvoDkaWKY67EGQDlz8kscSI9
5ma8tAHENLyUdsoilbtt1Cz2GgpVzmbv7Cja82XUOQNX5Qrvy4qXTYxArbaPWN74opQ2JRBDxDtz
wV9Z1pWd/tNEPFBtOz3KD093DuuNRBuOPgLucBsxFl6w91OrvhvB08jvRaWeyCuDm+KE929EYlZ5
MkjjsMBOlkv64KaZ4DvTqiQwUKDkiZpfowhtlsQfZwk07o0dL0MK3lKLWhNxOvQUY30OaRIkjWNY
lL2HgmitjHkJEAxmEfyUcORLdzPoCwYxYs159Cye44LKOHq7gCoXiggu777FQrff92GhH0bXixAd
JEfS3506XjJIQ1Qn8hYP9rGXlSJe1pg0jJNwsKUX4YKNto/Xs9coGMymY4TjWj2+w4lbgngesAfh
dkGLAa4HrAX0OVTaR5ns3XWEOaL61CLCS7BWYOuZsxhRzpigxL8Q50PaeqgOaDxPxXqauFTdcgV8
IiEjK+4bkb/4M0kAOC9QNYpd4yNuTaJ/SSVlF3+yXbxk+Qb2ITcsYzQzelgV+gfQf93zLpkjiz0n
nzGTA3v6QIwfLaFUPsgWLBWxGirxDj6cNb+d838SZTc0kYXQZQ+LZoah9Kio4k/U9OdCNlnmN0mA
kOjP1+EtXNY6GY5R8cl28aK2NztZuufa/NdI6yxtzLoSnaYzj0UyG5L9lQSlSGMgpj4iB0UhiZ8x
elpz2VwkzQ3LUqm9nhay6hRi183kuvZ6L1H91xBMN5K6ntaSkxXInPk8A02Rg7/zbxDHqH80fiID
Za5m8lWkz4z7mmyhIwKjAW/sxWhG0kudxFAu5+OzZz2NGLimxgTPBMJHiGapCjKso5zE2OaZEXWz
r+hjWkgVYCMJvhaheiBEMKxg/7ni+7Wbmf3+lsq6fabSNgyxUhb707nX0G21rkr3B2aOI7rpmi4S
s6ibdYmXRAxgAT2sogMDr3bt6Hpgs28Xd7H/imS0LC9ED9ZRcEDNNVpQYgWTuzQYgTsjRC0nQHR/
dROBSf7RIrO3lBqwj1fa5dOdoOPCUwvuNzWQREz9nRuA/+C3xmryACV2QgTfj/jePx1bIYCft0fL
MApi9YjwPzTBnHiJiK1iLZFrJsC13LQUIUitNuVnXbaA3CBfjhCXXZENuRoo8j3rZt2GL9wo3oj5
TyHtoWtLeY8V76y1RfLIZihJ8e2yQdhoG7oxoFujt0MPptSy/mNOpuiy1QXX/dG/8rVM9isA6Ppx
qgkyzVmmMk2X7IqJdKgnY/cS6aq/EqtKoXAWXsPsOL2m22VajDLAlS7tUmie/4PwnzrujlKHiPYe
ZiAQwALnh0qGNQMuAhAy72aZuNgJW5HdWZiY2IRBiSxjs837QieuKWE6tLdobYxmhDBQ/RoFZInE
6wpfbv3sBj/TQVtZ4gFojI5PJDeIXe1f+1+I1r/RBAGH4fz/CCILNvYgX6FNENng4nNoh5zec0O8
3DJ9AHpPW2A4ldc2l/GrHxblPdP3nMP4Nna5jTNHeoNpRtO9+U2vg0qGEOCCocAuoKbx/3Q0Aq30
f62R1qYYRBU4P7cBV8DD00P43ia8wgOhIGhX3c4w9ZlZng2kSaHHZ0QEis8upt1vg/HP+18AO+1V
/2qqeNyV6R9J9mH+4OGjvXzE9f+4DWQoo9dhxrlfwpcbRGC/p7OQaRP3ISQuKMZYVvSTPeQv0XRI
F4ak2+dgLUu6/bQE14v9Op4Vcr6qQu0KV02Crvc8gw6F11Au7Faw/jfZr8xRTSXagz3rYRApyRYG
FivBBrDOzHdq6C3J6IFid4iNZcM9nTkGSYCoPTNprG2GJnClOc9O071+dpIGLmnbuKrbFiU9YIpV
Qt8/cx1fA871OsKjwuSPM2a804MLjG6UwlYWvDG1vGExKgMCTXy5IfbWaCc2ixWhybd0wVA01YSA
Hd4SJDDxSEX+zB7Rdu3Vot9R5+bEdFfx+rm9yotFejLpxywz3wOblKrols4Lp/eMxBEfwWG31uLP
EJFAZeDu8dSLjLoIZEe9+SJjrSRGkw9B0PD5uh6qy4SwhOoa3AnxWqe6BgxLXHIJiixhKRhGI5fw
B1xoM2hK2Ed2uhZaCdFi6tUGGyJ0b4yZ3VVscUKeiNlhQa24e93uwQVcZ+2Sw5UwKYRLuiOqgl9m
V0hJe9WGtKFz9ee1sDZrWQkq7AQJJji2T+6NOroY3w4PXLRjNFBQpbAlbCPlHD2+CTyLSPCRGt2+
Ub9dnFzeRgDCZW4vADWzzh+LF+rM55ubX9O4Y4WuGIx/piQ/Fs9EtYn5D5xi/rnqfPjUc9EPDrkV
D5ZxBCwPYaZDchtGn53ShDe4As51O4vFGNbcD2VGhGvnE2b7If5A/K0C06sP8sgyO05YXIoYi+9/
8a8Jdx1y1GGjApWDaS3SBqwZ0Fb8z1Tug0MwR61b1P/y2sVvraeu79SQgzVRqxMUeAsDRy5fdVyg
zJ5KDSe06z05TPx/hH9lhQe9RYROBiDGJV7hHM7YfqavJ5I6Yd3XZTHIuxysLrk8yI/M9kMIQbSa
89K86onEUUp+hpVM8uYTyeRAqHrEk5orW4r9vp+pBCoq7+d+QBiHfJSQXgPTQSxUOpeoRVQUfCiz
fufbxI3g8bHjOMDF6o1TC7TF6QXWU0cWrwv9vEuKWmm7QsD0KDY7aRCE5u3wxoUfVTn9LO1mvzJi
Jsar1Pm7QeTBPYbzPiWBpHT17kPFStW8c4tKBn8qGZKE+p/yUVR6c9/smZVtqRqhcUMM7ZuZsffL
njqSAbMkKR435zn58Igroxo4yspIktT00I4Yui+7tBTdDhAodtd/Ntew0A9IpXw/oKUxjAg54Y/3
nG6gZF4zyKA4VbZZbIFudCt6QMQIzZV0s95Wifo+JuyznZGviYzFxU+41nzEeVftZC18gfF5Lvae
8eIJTyFUutqZn5tR8lr6r8npalLZrEdwahk2hwgTexVFlKmkG9SKSrhUIvog9kP3ZlfajIpTNVXI
RzXmVol7Eo0YCmL+kOWzvtWpk4KGMvpac7K84RzV0uUYPB1qDn2b+TAm/YMLjNLGSBRQ6nMxtPVU
e6jksMCiuX40f/8KYJLfA3nMrYijYqYjjPM1YFdnQMWjyzZ+ePxHddfViIj+9lwKAtsF+pA5cJOy
rooip3ILoR7Ek1dLP7WJHKfH5+QpUwHy9GgBLNx7xZDCCyp0CVHauAD0uDl8UukMvJD9DLbIfG7o
EYV+uW2PmWC1ifk6GfEbPkqnOBIOQd5TeNCIs+w0VYtdiYs+BnQ05Rdi65m5Hd2OzeMgSHKg1EtZ
ea9OG63svOXcgYFZt9RD1SjabA6jS1LGrgrue9hLOBdvneaI2sktitJyJW8U+ugoFeX6W9nYT/v4
Y4ozjWbSKjvErHWhNQ2Rilhn/SHRJlVH5ChSiARMtT52Sw50JEoTKycsyweIENMZsnGhiGI+kp+P
z1JOEd4H422dwKzoZrQoGX5rRLFlspbBRCIWlpOXXYPBS6X0IhmyR0H50uXE1Amxyt4IWCjGYRAS
m/jy+VGRohGvJXCZVyibho8Pr8YCWJ28zVtx4weAMHKwibTiRd6fXdYWoCV4OgDbhWpG0ag0DY45
GT4yci2SeGlc5MCHLIVLBSIREGOpsJVFjjVgroJs+O1uQn9cYIqqcD6gnxbUVhgK39ZSLh94SIXs
j1x/3/j4u9TF14OjJrUvd52x1+xkaAQNIhbVEVJUGKtSfxuAIhpVxhdcf88y2U7nZ/D0WZ3pGeRU
eKhUKAg0qjQU5tfi2lM3vyFuuXztG6W1u+071PpjtYAOaSZTlchtz8zbB/ZexOCEm6hIqmBvS1VU
w6BrutPqaKACtkTHGQy7uNC5KvmaoqrxXhT+FXY3a4hCicO9pP+BWPGZX0fcxldwr4q6ov1+Htij
wuo0yx1B1nnzOXD/kqOrpsRMQusyq7i4N0G1QpgVlVgcSSGdiBLuL6NNvMlo7IxtjuKGWII8GryV
vIMAtySgcJe5c4Gg+wxxN3NL8aaySCpwY268BwPV5ljWmLvTDVARKaozF3CllI/fDWYvgNy6extt
5TpGVaE31VnpN4YUxidpAtCrq+GmH/ItbULk8T/xcYQ8f8IsZWZbe6udweOvPyYZjW+Rmf/iCivu
Pqw1w8f5HkOUSkyAAnO6eRGiq1A0TBAYfkdxGyBkcd4IadGuj8+fVI70ohaoxHCaB50aNm0C9lCa
VTk2uQiVQRv5eqIn3c5qY5KcVh0Og/kb863oy0/uC5IAAIApUxp9nW4NPGIqtBNOYXpNkNGPeGAg
z/EllxWHIdQBhQuzI7tqwIBfQ4lXALa0HaBDGGOfax0xBAzLzQWDYAb/80S9H2AjZiomJ0C7r9be
Y5HruH3xZnXankEUgzjljhY14DH8saChXHneP2OPK2giXTT/5IPBVUvJUT7jTA97jVxBmgaBR/mE
OJbQmteWfToa19WtawEsskp+bywkgnNFCq27mFI6knyNcJPOYEmbwBhNOHwJkAV17po2Mudmc4kg
DlkFM3Lxo7n0U9C1dqBFV6qOXk2jD0vgKiPdNVoO83OftRR/rv56IzOj+FpR43A35AlWLOb/sHTj
pdw9CkjtqYCYE4JFObowl3XH9b7zueJnoiPy38E+40sPbfgRsk/B/p71G9AVZNJb2IhX9FvhUvYq
Z/QsC8ImwMglFNjRH/ptqbs8iNiOo3OhCfEsG+rtR4IvzMTJl6GJyWK1fCY13oQdEAdwlmu70VuI
ZUbcKbLxGri17Oi8bcyuLX/NhHlNCwfWE0lnduEc1pxoz0T4uphytfb9VZTepVssurRV1ixiWGZ6
JOkqpah0AKtlOqcgyOAWYj07RgT6mHa1Eidq1Rf+fNgybsmo+wElqcr04NM7oSLe4EeGHHrpYo8P
9eh3X9/dEw4ODjo4Km9HqFrscMzsd5iRCdx1ThLgasy4csK11FWRNEBwDSlBa6T02o4SMPwwRoL2
WTimLxQNZI7JWxpwCakVQI12EdT4fINXMG7jIOqeH8+d3b7jRFE2Pp4cQS/csZVB8WKn7++zp/zt
MlnCncycPAecLF3/O3mNX0kcR4/Awp86thJzl2cjCamVvNkIvyQGws+0iRgyOMBeR2dN+QOjtLZY
G9Wd7WqM5u0QW0QoF6WC58F+2YUkgeCA+GAlEpJxNciw55nn/Rwa1V/7rBg9ZMdit1w9n8zFjiMC
mQkEp1CJuExXNYKojWwPqJ7KnNhZgwNXthyE8brZnEkeyMTHnp2aZLKD3RXbiNFvN3iQcxSrEYuD
riPpeF1KnivOfPjRTCc3CdXWmI8on7Ur/ogoXDp4DakdalZfT9XFoGdeIlfe7W7sNTAA0ETMI2C5
6OQXPPFgRmbS3+ZEPIJdgPnGkADvUo3nWCZ14ws0MqZMbSfCGhL7DBtNnV88ayK9Bv81MyShHn9f
FHjlNYa6BnqKuOPyIV4DX6KhVef6yVMTqK4lrqH1dPGOe24DE+ouAeTcxvbYJrHYI1uy7LYXhVLL
PYYQAw9IUH2W3bzUQVqV00Cz6AmF2gh6NlgNZQKFffMlkTyBaFGsZSKZIOtXJMw8VRWWAkBnLcOR
jyw6etBN/OHv7lSxbrfcM06LOZ1ShOPRQEAUMjwin86HggnkuDleID7Cs5AMfUuUa9uafG5rvQfZ
TpOFs59pA6wF98HlQOAyJR7Myz90OhLfyFdUu9T2aIb8BNSXdZPlomP2qbM35LHFj3rdi+cNvz5p
9tg4VZAyVnsvxvzECgNTC76VhSzfNsLHM359q++/OprOQMzkr1W70IaDGnq9zpLxzN9V/Vog7V3P
5zaFM2b/IqXCyRPCMu0tMgvZuKfkKm3U4LwK4EaBJ+X8pRVbBqCRNx0crHYsADYVwa/4ba7KlKhn
TKjxAg5oFD74KZobRKSBKFL8WlixyfjQFrs3xgXei0FV6pJiHIgzHai79oCNy4hAmNC+lm1OnEEb
uYKKyKL03zl+55BHvMfRYxLZqOvXuUe4724U+rydxzA/pWPnVy07vyeLqa1A7SMytC0hnoTNuuVZ
vmjmwrbk1rJm75r0w6XKc0Y6jb5hWfSS5JaFA9O2cWKNMwRvefxlr5R6pCmaz48e1sHva0mmBNby
LZERkYIUB1lX5fG4BGnBXN5ITqROl7uChX1BYp5eab0snhGgJUj+NrZJfog2dzpTElwonMPOJX0M
Kc442MA6UI4RgUguxKg844RvMkJganUYL9yIySurf6SPpL+7dLqnsiDTBitqDYI3lgxxufw+sBv3
PmTE7COTIThhlaabYCl7mLnduwPf1VlamLqo65JcJ0owHcygmA5kwfXGEsM1/19EcIJQK6YrQmq3
iQMDlMTRJQBnUD78auvq3FL5iAv+d1Iva3f2s8/UPVx346KNb3J1HS/FWap6DSK5/Vimu4oT7l+F
VHqfvYJGXIzcuuyFm8JAkhcHHcR2lXqXaHmaDbFQKiYtse/Cxt6gYNa+2SL+CyCeikLrSLxiLx2R
jpY4k1b4lH5TE0L4R7yG8vhuBXvckZETnisVYELLctFNoDT+JgI53YaaBBtxLVhG2nu7NYF5Citt
weUjlr2Blgf0TCWg3W+CK+eDxW+02lxTrGvNIW2p4ludnzFVkMEx1MmihZSMDK+noVkD3bzQQJiq
iDDJ6m3Oyr6Bs0fIAP+/QTm22yYm/Pu6stCeVtXtnocBNyf8NvbLdsFS2kZyV9I5hFoNO7nSQqH+
HR7eJt1JPHsitqkb0lUnwmksxDFs5cxF2YyCX2enlgrbDCmQEuVhaVWN9iGhCEwXtWhNqSB/upsj
Xq9BpCrB/qRU2YT33b67awUSSZACeo+NXUDcw6ivTEg4CX+nlshNqJc2hnmyfxlfVe4crijym8aL
czv7dCtukObAPErM3PVtox/yshFZx/OEenqA9LM2nPVWhJHhNb2k49nkdeNjJ3RX6gJk9aOoZHw3
Gy8l4tu/POBt+hLZvpFvInZREa2JLNO+P5yxOXd8ySItlRO1bMeombsb9sgtIMIRuxvXzJSTQGOA
XYcdydRz80LSs0UxcLVPuBB9ijVyXCftW3BvZLyrcoe5MDUSe2Kf6nM9PTywjLfgECvEcIv5wYyA
a1eqsUYgpUjy9oV5InS8eRf5m1UjJHvSCvhG5n6iInUv3K8wJ/6axxP6/p14u6Yj4cYAdshdf4st
f/xPtDNMytBBJOihNATdOwz8H3ukbzNk5ziiX2l6+v3EHOpOPDIVKHXrdgwFhE7VwUapE8CFBpkI
+0zm49V+MtLoijXuNRxmAiyfWmMQo/Uib4kxS543fQFiPgtKXq7jmF6KhK8/CiPPAOKzzuAO2q0x
ouBuOI+CV4QIkI/Q2ZrOX/KqoxAJnhOEPEg4KojLlgye/Pm+Ou/C6QzW/5zRuYsFOJFXKU31WxHJ
6wDoWFbbGGGRtpBhKcnMh9AbMhjewnD7xkaYtt9ntYTGYt4Z8xjsUUfJctTLcJOikM/nHBBYI6jY
cMHh1MKG6SvV/bnIzJjpFH5dZ/Oem3Qxwyr+r/KbzL/VLyPIH/RW548PwEG+94vThF+WUvkQeBqF
blZC9nJ9kcJsN2fTDcsTfDwNSyqRwwNR89NtcR4BiaWJnDvYOlJEkpC3aYXVISwwl3bpMbxaCA63
rgpgrPjsNIAVlvxk0zueYLKrZP+RjfVRc+sPHjqqa4LKEQY+tmJb9yuV2MHypAqrsCOwbPczHKaX
kKwZPs7bV7XBg+4KFtTNAGH2P1fmTG4ixK3KVherUfzAk11/nuZ1P5nsqK3LFmZUZbj51L+dt5Wc
3cqmk+DeVoWMIOZeKgXJLFr78swnu79FEPJiNM79yrPf3s9UTVam16kV/pJ3SqUMbf0SWDccZA2b
zviS3EErRG5So3rOFoyx08sOzeFPn/eLhA3LyC4OfBk/iHtjQkiHn9sOTquQcARdoGgi8Pc7iXRp
f7DFcwYIRnt3BlamN6VAsOMgZzzAm0hcOCGUB4830hHiuH1oJFkbIP5y3zoe6cK1wrVigENtX72V
kHHxTo9KeiGlEbuzdunEPb7k2bTsFuTz1tgkpqoo+TRqZtiIRrf7rJcvgf+ZUgK9857mOi59jDcj
RweQYgOCaUEBMM0e3QaVqvcuh8tqAtoBvFGyRZoeEE/z8dAtx//Cqfsv2qvMP7sOq3dkySgIJK4+
maE9vnERtsgn0ujXkup/qQ1MS78r0O84ZBDjSVtREcLN7uWCms7pFujum0PFA41+K5usCIQ3CCDo
rbYRJRwuwLnPHakqnC96jV1Yh6l067SFGpIw/a8ppsZbi/YEB9z1qcQCFax4mxswOMm3K3tTsuhm
YPsbWC6B+Bq4iDYc6xiGWuvWAhT28ajJPhqoF7/wqDULqxGE+kgECQp2U47+RgUwKXuCdc850oVf
Lf7/viG8ueQ4AwFQVAmftZHNtgaYzKhc6ZTe4yeKyaqXgLN0+pA+NIFDHFZjeH2+BfIlnji8dfGF
dsDUMUnlVTTskeNi1UHqPhrsBLaALhKdSVg6CklNh+rwVEdLGDQb8av0zxTMn3oEvZix7PpWlzS/
p0S2CG7FFHtPu7gGT7UrqDoapT4vjNJI1uD03icXQ8TdXcoRXF8Q6UCbWgxaNCXXSuO2JotP28T6
/VXp2+MdtTQESVdv0gqiE0DCgPcevoHKS7QxTBeFgx3M8YVZYq3cvVVEudWMFqApQl8N+6b6Gt2O
YmBqqR5B+gmFQLmik6rvTN4Ga2+6kdZ99T9jGvTr4ppxlZJChQpDjKcfodFctqOikcYmZaHExb8F
HC2hMekilH82DDQp3vvHxqhEpJ4qnZAMvcdAXaYQHOrk8X8wfNlb+DDGPoySO6/i7+/Ti9SUW5c3
YzmA/XdTO96KYV6FlspjSXg1VhAeDP3bFOxdZ+vTadfmgHi16p9+nqob+5ah9Ixdyx5d6hIL1jZR
aO13Ww8AnoG6781FC/HcvODwya5k5sdohrMcRPjJnBtZAUKm3pKmkvk+zIgDe6qsvqhNILYxwKS/
d+2eSDA1DFU2sguiJ9usfBjC3ZwrwU3LjDY574Xy2+H9dIh4b478KZnf1N3DVqBURHrlQSwhQ/go
2uoUfY4scZvwIv+bssFBBJhHbEdS8OpdVwt5hI/EWxCPd5T0g6BvxbrLmdhyrc/0/O4IlVI0CbfI
A4tN7KYpH4CGltTepyagUGuDT9l6t4FIzuVIW9knLNjHXDoqoO8RROkzDpBLVoQENoCKQHgJ0H0n
oG9cHSnBN8giJw+TWk970wZOF3Ckh9ur6DPsray06HAiAuIpl1W5wZvA04uH01iCa2J2PO2od4gp
oBlzJHjXBobkMPuBlI7P4VfECJUrF8jrD2KnaehAhyznZvJSgOdAUrETIDXCIMb+7WK7VfbPBEtY
0pQwZV5W76otOK1KMWN9D4Rg3wEYeNuvKMD/5pajsI0A3mlHrUthDo8VMK6frAdHc4+jLBkQnhqf
oHS1uMnDP2LUOAsdjCaFe0qb2AR7RYkP+ouw+up7iiGdaw0BnOvw6Gtim06FS8NWp7pYvErA8oni
DFyFbeZxL6IWEwmZADU6A7mCW7QZwIRgjl9AL12bJXpEhg0CfLvb75/5C4xsKCzMlyBY7E4MpmTB
UMDYR1wNB6Bi76gqf0a9ArrwLyaKVhjqEh1ePSqgS6jjU/DS+i2BLKBH733LGLWKRmT4Rs+KcJmK
w0sYFthX9wnZ5Go/JIkDo2zE7LlN8NDb1FvCee0bFwdNz8X8FvPqo5Z4vxNowLd0j5aLDx3UxCkM
tOiKf7IsHCoNWJBEHdWtl8yYsmHAUAtgIEio9zHvyOSg3601ybC7Rayw3tJynelHnIUgz+wFxuCK
8pBNsHBZ7kN9IcVJIvLimi/gRND469fGVDUNsUNWTgjnNYrP+jerjMEexe8vhSEcoG7dup7GR6zn
xbq2+7J2+x5ehl1d/xnzOIDtc1FZndx3vBHOiaGFyc2tJAtP5CC1vI8Q4yD0vvoEJ37+qTtCUYoo
o1gSbxR1gJoRdzHxW+qMrjDJScXmQdKSR9S9Gx7sPkkI4cvtEAcJJRaE/Te1D+lMVx1j6DBltc+5
urg2FzJuD28Qv9oSWd9eB+VeLz2ixfBwq2NcOFvc3m9qi1ZTnrsfXlsgySBi8WhZvVtfMavocZ8B
M/EeA6zx6mtECkLlZd1zR5bw83eMzQBr0uK95Yk+4qFFxn+nOb2tJCs93Q3/wh68itPsIWkLCa3Z
hTORz6EEeCflutUD4k99cwI5KIdnGQj+7c+02JcxNHmp0DXoPnx47S2bdLp8kR7fur9p4SXqdAMD
RiUq0lJLnVxQYMvzFJcLqtezjYspezU34yyniJg23iOjxjUEsZIYUNVuazsio8uA731e4fZ3OAG3
BQnbeAKT7+W7+UKv68Htq/IadxoiCgNmLEbZo5MzmRT+xAlZwOA5+BNNfXS4l2aDv5re1VwerHM8
+rLkbcKXwxN6h2Nig67IblLIpFP0K248L0OrjTLIyMiqZHSJHd2FUa9XNW1oKzTTN+nqG1lsnUKz
kz37uwguT8FgYd8c8n6Fdh7aFzyp4+hhF5yskSL3lKdKdpTi/DWtj74lNUDtVlRZrmXM7EvO8IrU
ptXYMMX3ohZKdiwXbboM9PYiASCMDMsLnIGhnv0qa+eT4fMdlah9WCj8VS8N4YlLh2ZhLxIqHYwo
YqFanJWoLsiy598xGzURMzt5OHULfKOB4bQwLsn6ed+1ccJ1Ay1FzeFVt85FJ2wVDG5fIWvX0iR6
YV5qatmH7z5F1sjrVwrvfS2ZNj+aZWp4l2pUCG7vO/LVox0NDazsFypbdT2vFwhrCiKyr0mcwVim
eeUBclvQhOfzLTttkLRnl1doi5joEteVHtCjOJIeQUeQAgcZUIixqOIEnHVi4v4CtWIbX8hCItFp
3IxGlyxvQe/FvT67XOhWWKMMwhnA9ibzSJrBIx97fAVE3GknPPxSE9HqiEW5XJOjNOc2Eum8u/GO
zWDZarhjEW8UVMRxoxWTm+aGs2pwhWbCFrtv6Qsq3CsUR4GAr9CO6J3XMNfmWtnMZqgAHbqFvYY1
uoheoprBH0sY/tZn+YL+ZxNqIRu3nqZgky67mgrH9awcofX1fqQnHw08uHIr78k+9Vrk6XfYjCOx
C2HxsCKKyufXlZBOVNZjuFct7QILm13WrEr1s6is4Go9sKk9sixnF2vBfOdohutw9FAu4mkmxtWD
1/ElF+u1oA7I16WaeSal9Hnymx3irPtgQTiFUpKW6bXFvqIoTEsmjtOlktVrCbQtTYTyPpAmjkdw
6PPK7yIM1z6ta55AXEKal3hAyBNUknXe+a8qsNcIqvT3ZmRjrJqr3u1GpZMCvtTMMbzpng/sh7w4
uApO6Nb6qca5OJpB36tbV+E4iZBIfxrR4NZAmKIcaTmXGlxrvWkrl/93Uq4C7T4rZLJOxoGbffAW
vRQwnMxGh5mGgcxptbHbsH5cZR14JM04dN6hyxXLOt6auw0PhdiXmIkaGN6K5TYYI+hYLHdK+IR6
bRuHiEsBZJVBfJ/AAoJkcCfA0SWHKIHccRGPFoDt/q969jlq0JZJa+JrXhwrZAj5xio0Ut09B4QL
w1mKB+IT9DWDHjt5eiYeBtXSCXbqfthCAC5jddt3B2Ey0zEG108rWDdoWOO43FkbzHeBQIq/tl1D
lCZ8W0xfvC+9fUUmK2z5kWWkcjastpQIBIi+61EIDxiBC6KXTOxfKBa3Kwyjyp9HQ60qbT3Swwbs
2+5YxHkmTe+Ceg9Yx0wytOUQfLtKguxtVapRW6HrkSk69mkSDwcrTelAeQ+LsNoBDaEmUgRYAovl
nKEmhjaMDp3Q8I0aHI8EZnjg9CabYqi/A6KlWv1RMhPMxmb1Dx0w5P8HmipHK1om9adG/DXbM+Np
oxhGTiOKN1IMylc/t+mCS1yz4VZnQFDz7tnH1KCO26wRrCrjiifgEzT/VLZkU7oIw3slVdczdbcl
ACYVMN8yRNO6lWODcDPMT80wl8Qn+WmQ88OJEAVxXbPhQkDhnDO4ejJdSy1DYet+RNJepz46qJNt
TOrsGSsFH/mpSaFcW+mFKED9atRXgbfw+7ArPiZQHwzm6iU0+Lc8+mp8LAzJE4AEtoThmYDXkXXl
SSN2s1ggjBp9Jny+zd5zZST53lA20bpMm7aAhuppy7/IV0JFFxcX7l4EtgNhEP5Jcz5ApxP2am1D
wQCl4KhqWSHgm882t4RaZSLl1XVe4ISVYybYRyGVZ5hOu+ZI2knP+zX/zcUlPlsWGdiTPRJMFuSC
z+KPNLFQN4DoGiqduIQvq93fjso5MFLl2WsmNaSRuHxWWIrZS5sZUvv8fnDqu4Lr5whX6bkBe/0C
EFZiQ3ne1J2SdMsIUQbMIzWvIokTCYwVV5/Paqir/F8OVM+g0bxFd1RiC1aRDuanar6RRS2xqN3D
mN5wu/4fvUbNcNgW4227nYqjMDfLDeyeNUz7S65/c0PJ9d72sHGjxvmYGGGsBQhxRRci0aJQ3dus
zJm4oTibsfNvmXlEMf5A2vr2z5hCQPjz6v/EGoVNuzUsk/CGtsdYYv6fxbKN96ubolEXAc/5NzK5
suSQRJhfFCR4K8bduvAAyu1sVOBnlZCrt0IRlFbE1B4lFQ5DdxTKikwh97WOfAHOILpTrGmp/fv/
MqlRjeEUVSVwDGuczkJg9+YsbdQq5U3JU+U4X9Ee3FJdh8Hjd9Oe+La/b1w2xP/2EPRt3ridlVUR
ctNDQKcGrwCCo9TxWjvhcu+usuGe8ihP9Ty+ANN0gLsXvsHsGzNlXWv6N5k/5Dh08vzDED5m1iNt
rV1nb8AatmIf4cbbVDLUNlwGw5Fmz6+m0bhTO26MhoV+UWXQvKF0LmeI8a/LHly/e/v4bGFdZKcr
aHsXl2bVF+MBH+uZGJb0toZA6cYt5raAixtbg+LfmMO8GFvXzofHnS3bhw6wHioMGR5QvtGNzVOO
ct6T/Y4yV9i1t5ldEttZTTVZyh+Jf1y1WMV0wGoN90yWwVAf2M4NyLqsV/+hZkAj4geIPimOGX2j
7muuJDR8LqmTPoqTsWMw1xfkhMPK+ewxmoK23tcztuuJ39a7coCNKDJKzhO7zEgoQc0tFl+Se1b0
giD51TsttMzWIY4l5lzyAdGTN7Ee3AX7RHPeIr5jKkWImlLCslbKxQYy/V0pPu6/sIxp6uKQ0Zmf
nkgVToWKOOUx8fEbI+KcGdJ9ou1I6PZIwW0k4mQBnLOyKaDVFl8W90wgaAQz3sV2PjJXkP2aLMzx
Zws2AoLWzLRQs8uqr9uHYHWmjJFN0RQjenQJjn4l0/zpQZSl912cLLs+O7WrtjAqwbt7eSGsuRX2
WD+aQUG92ZhwYjk9VencAHRHHXqPMLb+3evpITWwyA/dGBpCd41W1MX/aKI4f9f5haMDGU6WFyN9
XDLAGB6P7aLpulmBan6t3Ct5xlwGWAvDfgZkINlIqJN8paullhJNVZMvp1x7oIZNRPyJGIF6cdp/
R02Q23C5eN9iqqDHBDw93E+VY9ihhht5U/c3w5GJKNMrA6iBg+6zd877x4AbaLh/narP7wo7TxtP
oBpm7HvdddArds2ZvffUxgv5FDWTRKytTSoxoSw9fPinHVteZIof+lWF42IcaInm+EZV9BJsv3yd
1MrFCUiWLvlyoVrOhwWDjvQ5C9Qqs16b2wscDj3Iv2l3eaunvMknYvhPtElvH9zu6EbogMYZYXKn
Ypewevl462mX/Z6Ww0Q8xvLRfuRUou0AcQF7f+fbu3uUZy/6oK7MzMhbQbrTwAZZQUwCnRYKIhtV
4DIe4DiDk1wz7EZXmT6tirGEH55EZkIfNoMxtq5khpWOZbVh4vIRfEFTPJ2pLe3Fg67Bt96Ed/JX
hmuvLoWUV1vx1eyd+XkY/RMoG29yX5Apbjj4EpHj54l4ILCFodUoFUW9Sx4RpLfgt8ZY+Inem5iL
6Zi/kiVMoL2Pnyj+gn0g+XgGCxPs8SYyg5giA7WvccU65MxGco5Qshqso1hkRCrEbCApTuXAU5LN
wO1cw5UzUViqcp5/MV8wIs+By2gvEoZ68eLORpytI8FG03wpml67rlqE30SnFElrKq/srzqVYErl
yZbucTAhBYPD03wy4umx1ME26ng2+Hq2x80nn00BvCIG2ajiHkzPT4u7IvINifMxyGo2st9/cXaI
QnldFj855woBs6RolN0xyoz0FmYefx5tLouqwiHCTVEOVJk4jxiuCzLukBQw2/UIVT8gvCg7554G
Jtog60IS/GfKOqS8nKtWmmD2zrY1cf7qw7pz5njgVhOctYMcFmbT8CJUxblb3cHBh6XtJLUbI37p
pNvEpj6yDV/Jg24t8GwcoJmZ4MB7/ailRfMV5ln+awJD6oVxatMPXuI+abkMSstAUnymNEOaEsAJ
s5cAjcLa5M/NyWfwJXh8OKGbYHu5jLNp3P77aH/a0+eOdMYdUiI1+VIW1F1PZGhIHhAv09a/WUHQ
aSOgiPGI19AOqLyqhV6VB1wXk6ar9hlWNJ+NY6zngcAoWO7thi4p4k3HVq1pV5jWOjomLclXmRb7
7xOTBCX+djIBbBgXbvRBVdnV0rfVXjzbWLWgvSqNEalrSGUt7Hl6QtOTHAIoezZgPIXPLWKUrLha
yQyYc57EoZBY/Ryz4KyIKhPaeO08pFIG7Zb84ILMnaXDyjJ6Pje68KScGuE3BdkzsSGHtAeVUHnL
tBcT4Tpt2GtzoTBK9BVQt5q6X5+bf8EIEYa52jIoeHKup/Bb6t6V5CWELGsI7sH4O16P5pVEuMY/
qj/AcJG7TMWk0iNxzNRJLfjLN0G4FEH8q3dh4aKAcSaFYRtCH1janm6vyZ//dMtwam8fmN94kWrS
/N3MstE93nHwz8QxXoLr7IBL0C+YlNlDVufJsKY1dHe/lQLNAmSsSliQ0q5OnE1JGzLdo9OUQkHl
sI3R5Rpv0/B5hA4p5ApQumhxbZsMcKuw+ifNAD15FaITGI7Dps5DN2xivtZS8lh3u0L689t6U5Mo
X5rplDC12FAmIlLq06kI3WW3KXwj0vLWgk0NqvDr/Ny6gqfpSiOVpOWmAUpCxYMKvusQJ3fC/qSh
cU2swvRjHngseKBYagt/fIt/tgWkuWIXncCu0VuwZ85DMrotef0b2tZ56IvYgmpXgZbZaCk94XCN
gKlSQtz9IKA0uczkqqbemlj9JRolYbMxhMvB+OgUOfrlaXqj6zyx3dt97ToiWRGhL9JKeo6y0MqV
5HPeOQNacelsfAUwEJVx3sJKXT72BgLVP7/T4WznXnPQ8WWu5s1pGah4+Bri464+ynWZ8GxKT9Jn
laPGa1ku/QW2A9iIbv6kvRPd1vjoSrPQuw2Yf7akQzdtvHWof3GoEeG0H0SriOISlrXv8BFg89TS
Iv1f2KzxpNq/iUy1d0ggSfeaEb0c2CDxpxyinBTJcasql+WtdYLB2CfPZ28GS2b4lKb7TeaJKP2X
zn9JRfhzzCx33lj+QtNMIS6KtdA4yUGmIXI0xexajOqFt5dtOmsLty+NsU2IkyWAVDBF5gZykAC3
jeqkkq7ldbI343jCzEx4nuduBYwA1cpEeUldtQC6pDz0/uKZg2qbxFT10ndR4on5U4p/k90jSMPw
gyE6Q4Bfb51xDhjdVm8k2AEBkNH+mJHsh8MMjfZUy2ei0p2MfFHwEukWLKXWdixKuEc4o5hoooK9
m8sgN3eYUtVewMJIQ6Z/Cud0STSAGPCrbNUGTbzJtWnfPXLGs8bGFbI6IPWs4ul+hYSye3Wc7HyK
Cg4VVKu5o+fHRRZHWGwwsgUgssaDeadfk9DhJvVsBLfP1ibyTYODdCgkk3vq91FpH+CAMtEi++bV
mePViwl5Iukoh4XzxE1t5gTEdGHrV0qj+n5p+dpGyMSsZh9MWD+Ir94QUBJV38d7+7fHnzV/AQrw
jqXP7Xple0IHCnqclPcG0DuHG9lm8Yf9KiqxVkl0s1z9/CHCdh38JlMj2nBkp2CV7wWfkN+9Hqxx
yPSaVldLZpMkvUqHM6kSf5lyEQwHtu3HRu8mc4vYE486LSP8jxxdXHa/mVwP5LKURPv7Ft67KI9T
CyyKoK4myBJEpZFcfJWvKxDnSIxrCckYyZQG7kQjw2iAk8ySlVALRP93aLHrHuL1vaxkohZR7eMV
avFNHFm3lAa8hp5kywHP1+X4jk+mFHFz9fBd9XdQQIID3+eMRQ3FMW7T5C3e1zWt9eKDFEI2oMKN
VTiZY5ZJVcWwmqnO9wQOnUBcPu++zgqzfR4XShrxiDKgG2ZXcGLkX6G1bEy2PzIIRhsV2c/zcLt8
//ZiVB6TlAE5v2Mq85X8hrNCI1076aEdK35Agp+s4fLn+Bk0vDNV4L1h82AXQQT3u66yFd4hbGxk
UA19k7wFI3TnB+zsWSyKSZre9Mn6nVOKvh7qwYmvNnA2Q7pLchoDMCRIPLl7Yg8U4S6zIxMwzcif
xvmc/FBGnafPoI1SIDwgQONawD1Dzw+FpAFLRw3o7/I5YmO0RgL4iLNBbgCaE709ZPvzQiNypxq1
I8w0NuAbc5c6CbaoEVPF0LYmQt8d1W8CwgSH4CDjQwXfXxdkr2OiinypJBnHfeB4inaswOxdyv9T
GcBgBFa5DjkEmJCPagCTHTGYxiZd6PgSLNRUCI00X2E4SEHGhYlUV7o81VMfd0JcHCNVKNc7aq5w
6d54iK4AaEeTp0ZXeoE4Pn9wSeBmISdmXqaFKL91HT0pJjNwmJDd6z3SRR5aDQvERFFlnQMYUCqy
SQE7CnLnWBjMlxoX9DCneEs9S/pxFaHnUwrsDAUYliHuw1tfD3ycVb6+GBYkkxB6BiQWpGsEmWyD
mvt7umrPUB8qCeM/Kp7Dt+7zhpVaC2ZSIdhKxhXBLGtEnV+/Fj2sx/0UqDs5xVKHrgZCqiNENl1m
VdF1yujSBNFcXLseXmSlYiGwxeLp0ZSI1frMKbrBKYr0bPpECIjS4ZVdFlP2jB8738rCXqUzro1U
9eE8v18uDeuoA/LRdyO3AspF9vmg/qh9NdIIBzGgMTVVX8ZwFdRXbofl1bUpcuicLGgBuxIsD6BI
cv+luDnvbj6J7kb/LxCGc7ll/8GwE/LiM9HT8CYp02eodl7I9hQpo0zbZCjp1A/EZ4lrdSjaOp9Z
R5QNz9KtPgSGZXDrChzH//Ef2oloX/qmH9/qOqFfY6q6yaqLU+vSWVrJzsr6alaelsEdP9QgMRfx
bjB9JiIhoq5U9aLveb6zso+Bib6TjOCBxP7YrfG5FMHHx1qV5OFZIxHV6uakm8LF2X73Gkp6sCEf
Z6V/1tsaW0iubowjjqi2M4I9ZKx1VcN5ZzmB6zm9Stlzdn0ttQi/zu9it/4kj4ljGfsnPEP0IY69
JQ+kjX6tQqcjpJc4MpaJvA9nrE+GaGCuqClvP+qn9mjZf6eZ7lcBJi1/8KZuJqdqnOH5k9BExb1q
CZ39rOmZTD8MF8I/Ktv5t2mp3vt7ixB7QD3nYDMumRzeluLCEeede9E1xHtG3VhCHYoH2LCBqCQg
haFyLn4+hRm1j73IG+i2gFiIqG2wZqA6YThtLVSZJ327aV0qRr1FCX2KsVPfmfGFFJrFFZc9tgZ/
BGdF9UGKzNrQkHnP7sTj0JiR9VqH5pPUT2kZNlE8NHCtJxgH5rxEBg90bPPfsy4i3fdd1DirwZ76
X8j70sixVaUzewgtWke7o758hegLPc//PZnV3oR3kmPM3Q2jsjcARY8y+sQuGKuZgkXkFYq3qFCY
zwnDTtPdXuVGMnQbnRWT6137wRGbfBZv0xIIyaXC1DH1wicK5q5SpXGzN0uvC4cjMbT3L6Y593Wu
esQuQtu7kID1Oh0UdHxPLt2ru0vWspDbVMxw24ZowLYQaLl5cuJ4FDbvYrm2GNSOmRLB+Zsdk1zR
OQONg4zudkPCp4RehwNpdVoKE3H6fo+EY/TIyDPAJ/yiVk+6J1AHfIBiSviygMKGwinNpB0Ll7XK
JtnlEaqSWR84UAcJo6pKeUlXIjgdBqJSbk08kMtmiT3WacujlyFDHea1fTsS8KsD6G3t7HYivi9y
U5SoaJp3ZODLpb0CGUYhpn3XIUf+5yz8Df4OIb+eOep6gEi+WQeQcdUKY7vHv36Y8IvGVkzCDaXo
yVyvCvqdFvjpFl+q0YDtSXQPChhOXJzOcMrUIH/H0bs6A7ui0d8Y9ljDLxLKk8TVaelXWNC0HR4G
5cAJdOEvGUjZKnBJL4Elo/ukyOSVJWQGfrTJpoO1C91iYK1YceObETjwlhqiBlnymzISTpe7Bx3C
lNZhIgk27UX1myl7SgRGZoLZA492dyhj8/d1AXLFZoI7jcRSY7f/c+eBt9dreDn8MXF3rJ3dAtYc
WVFXOBG+JVoVgqyFYSljVcNQpJdutY2lIu6S9u2/7emj6u+HpdLv4y3b5kJd+Ru3RbQGpR9QXA2p
x1wKP3sIJ2ZSbO3J0SarFf9TldkehGHsiK3QVxqGeUXARLS/OoBjcrKaDDBHKuo6yRecsaZBgE/F
3+fITS5iruXB+dwJxnR0rts2FLyo5riveorN5EUWG0vHBL8/RuaDz43gI41E9l6SJ/OP3/n2UOCR
D02tOjJtP/4L1u0stqCYQs29v8etd2m5ajtxhrqqklypJzAE54t3es/tBZWE6Xq6X8flRMkqFSXv
yXgq7DERj4wHCKhKLE+jVoh8tUfcbH8XW7cWgAQmqSuBQz8wuf5gvDKlhSCcQrhj8aOjfebQQGMR
03QUwYFokPDwYEUb7c8Ai+toTzgXc97CGZn2oIaRArCnh5dImf5/Tl8R8QeVfuCHGJmCqlfnzUCh
OfCwZ/sKq0OrqrEBvALcy/KYd2ghKsdXVY6HNJbfLYPiTFWvdsmMYlsvwBkCo/CuEbawJ9WmUmbx
InHOPnOpI0yZQz3Fu4F/3jGBAogq+26xSGxj/4DoBqjifAO7zC+UwjAuOAH0q5MWRKS1teYWXobo
mdgyso8NrQnAzmDZ28jDuI1It+We6WGbs+TLZwzyxdPDhet2wTX8ZBxU3ZlS1b+Xk6fdtF0mMtby
NKKYjFmh/kx8gDGdfY7J/MTFfZdzTtqvnhqJedtU0ma58REqT0oKRZZs2i/+FGFsQqA8WPQ/CEH6
3hmYmSWfZZYIm91Z7jhvlX54rBWdgnrsHgi+WTY2kDNRIcSY1kO42s0AffY8pvTi4tlBKInJfCsE
f57+JqUHNvacbYEa7PGuRggMdUZ4i7WVFXFqg93QC9toU0+1KKi3PiFUN0wMu4ojbWse6vPp5k/A
5Gs3Q1tnoOnj0FF9ODoZbBi3dM9LuxBzZC9ZogHcRcTg2ghAzxXdbSeIMnxLe0qsgYTpF9OzAgVq
vhhcqQm8V6kE4/Ck8fjgJKxC7ereVScT/U2X1h1Axp0kbiPiYnxkJvVceJA0VoVoMfY3ps8QBSaR
Q7g+P4QPtARhiFPk5vejc68Xvr97ymxSTE4DveHD7mNop67fwSxjHd0qSupevRzqaeC9WqOtbhMM
iKlTV+cNq/9oA2TYCZzwwdmlVzEtX+hEMt/AfTzVNdzDczWRrfLsJ0UwU5yMg2UXWaGHiHrgL8ML
j1SEkM6j0PeNY1RvM44/Xk/ybwng9PuwOW403mhSTOTLVcd5U7mvs+zqHhpmBaJGrDf42pnkkxHL
s38dV8a0OUXQ/rWedSIT2HsIbsr9a0Q83BztNGPoaO/28WaB9KgBrOhZGVEEMA0astE0pYyFV9U1
zFiVwSdOeSk2TqZ9Px4xxkbSfq7Y/de+IeSSQCNatRxXGHYZ6H4j2oB1ip+2w9J1JwlOmJ0hxelv
NpURp8brK7OuPjKJU/CAGEQwGVwC6Poxt0crzJGyGnta9Rp0dost5OdE8e3rO86fN50A+/IXBT8g
V7psWs3BgVIGOjx+T+LKAhuzr5r5/pG0wGCQ65m2TW4tLRY2Zv0yEJDZYOrRKd+4/i890BvIhoDl
hbsah03UxGzIsspxxV/nuGdPnv+KCZj7FkW7HgBxax1Rf63BFoVgv8kUYvPq8kBY33gM7lQysbKI
OHZgxHFfwiO7nCMxZ2lUeD8RtuM0Rw+0SSkjGQqlgBGnsbAVZ8lh7X3kSkT03N1wMBUcs665BArn
N/wgIME0VmIwfkOiVwdKJPF3GgJrm7MjA8aYnXGDJ98NvTyLn+ZYa9LrMMC6nbbx+rv6TPGiWBoG
qrmkrCcu5s8dSg/VKMgme170vQq/ND5idRI/NQ9+Q8DLt5oBdhF1CwyX/iC4k226DSRvKJdiQW0g
PRQSSt4SHcP/MXnzY4jhVjbjZh3T5N9XAks9cKq0u+Xg0Nay+HuClxFnYQWz1yAPeu8ypgdANQke
8Ot8wK8huCuA94yvqkho63GXcg73OGfXVOyu93BF0m2YrTeaIPWB5pmcJjcZPICdU+PHi2MDDqBM
khX/sxTA5+9+49Z1DYzKFZ9NzZzFVb+5X3YhkAj0Nbp9CG3dGS91oEPx5zpwKLvHVf8MFq7H41KR
luLYZeM2DlI+s3DaUS74khKsAWJ8SXC5tVkFc3mHGyPcLXvEaY5yYmwkjFTtsTVshxc+GAvNUJmQ
Mx381vm+65gUVMMK+X2AIhEzH8SAU2ZQ6JRD+vatOW5oQPvenq6Qg+6XgIz+gGibGQOhRVZRKUHU
x2bzTltsRM1Vtgge03qSLDkTV8wC+3g8zUxMVqNPfdZ9bPu0lDlqheM035+x88aN+iSCGhufqeNX
DfNy9CJce1IFTk0gEAmGrimjvSVHplMbCPp9c5pzf3amk6tpzlnhk0kGQtck6bR3cKizkCPESQ2R
aJgGbr/usB4zgSfoKFSmrqEA25jcNWVrK8+fF7dQXxBLD2XAsQYH2YmDLm+qkpFHO0axXAaHh6yi
YcksMrPmKvGrl/2ICz8GEimEFrUeeM+tnVXUJsQ0BT4yAkX/UYgIj9Pef8ET9158DmnRey+55LP0
2Qc1PluwjNLEbxq+1P1/w3XJCSuema5Ca5UOlh8J3Hrl9LZ5AdBL6hprXf7PK0eH0AtBMnQXJ+sn
CS8qo0+GuMi83sHRZgEGcz/VTarkICHKNlJD3rd5Ani6hEeYI/3qiny/bp3vgUUacekXjS41qy4y
YQTB+cjDAu5+TlcCTM3uVFknBalN6wFHDOi16SWzxGSjsGMFgmsE4ZkcLf6tNvVAKa8CmsuPm/xc
Urc7CySWiP7QYfKQiDOPDHWx+yxWvsiaFNdN9C9yAyVV1AYAq859/ibMfebenshNW2eT8kZlSBih
EqDDKiE6k1iXVl1HF3vVn/AQX+9ONPlkwpHmUVYujzxculp8muGPji2Id0ufwPBKcoehFn59Bh71
HYuNYZVerYdbkY0ivo/2bPLj065Y0bKGYFLl9nEtrtWQxdyAcXBKHOCi77RLegGcbWKIqpQubXxJ
uvNFMBgJ+jEY9dF/WV+hGj81ai0BSuWCevleMcGL5toJsGM/I1SfcJERSVXIAHPaIdZ05bCV8A41
7ieJLPZ1597MfT26bX2gxeBno0VdihgR4rXo/jZKmgNbyBp5KUXm90A6PGFzTAqRJZPVvDVpbWYA
SJgR6ki15/jz0qBNjdieL2/SSKTSnCARmyaNPeQYqE5K4lh+tFpT/9m+VlZ55wLEhhyAfzsv4Ni/
PPNHytg8qSG5K5On33chTH1SmTSvwICFxiZc9CjF+sFZDNIv+qGCcLRsWv0Y/9NvOks0cnGlh8Q+
q9xs8386D0GmVsY4wuMpGUDDq1sv7n/gt+IVcZHj1ae7e/Vohksb9BRrfkavkGUaePGWDTC35f2S
M1WEoQUHMUqFJwrUUZbPTK7+yZWEjqVKijbGtchDF4UccIUvjEnF2w77jLEqVR7+C3R/HV/kTiFu
0H8mh1Pni5dNW1tN072RBKw/E7z6Ei/O6jGNi+edKpJqR5AhhJXwqnrZaWrO/TGFYe1QZrCgM4vJ
YucYN01VTeVL3fdx9SS+fJ5vjR6vzXLO7Ras4ifgMOl9d3xx0kJid4Ym98xKI9T+p3jvnT5NpMVJ
6Qgv718mGy9xC5AGGAYpVdCME3l0ADQmoAlph15pv2hWQCEWYhgAERC5jIKTtou3wRyyYFFr6Ewz
byEPJXCfrkCpqqa72CeXDbKLzuchyPCPiaoYWRaeTM7yV9PQfWHauYQ4g5D6rj9l1I9STYDXnFiP
3Tq0IWgjC0OYDdIgGZv7CgWChnzRP3wJ72x65HUjUZ821ipCoNUvorFc+hNsMROCL3bsWhwzNvj+
NcPnFPw7z7Ccm5Z7CdQjZCaZDuwV4lYVAXGrTNVlwoQv3CQFfTfL9nVtwGcZL7QSz+d2tng/ivyo
CaOEHVrejWsTaWM4H3ou7q+ybiCU109djuzhXs3z/QQJTpo+P4/qiiI2V7XtmV06yplw/hkPgGNk
ox04LTGTAAR/uyO5UlfLs0VrtHx60v5t1+rY0Yrc7fQZw1Y8W/7WYnInvNMxuXJ0s05Ty0MHnrNE
b/WC6qGWf5N3jD16ej/9CFygApf8v2WXuB16f19cnGLgf/rQ3NO+mU44RQug8b0ZapCGnMmGs78/
o5nyxWb5Ci7+zHSYB7NM5rQPProjxxNVCteTmwwJPjD96hxqt6ugKZWH60Iv7BnHb3k8RO3Nx6Jm
eN9n6nLicC6gAek19nHrZXhAz8AGKAiP5/IIYVWEd0gFq0FeLH5+gIKqSO5MBKi8vjJUF4FuKCoo
BgEb9cyA64JT74Y6qT9EwkXbOE1YGwyVy+5/os7DkCnisBqGthq3CYX1qL1Obqbpm8brN+P3B/F2
9xqdQkWwfzo6oeIf1QqoB3jlLpZGYBWf4VU2sW7TlmoHmv4n0v0W8Sy/fuP6IaOAoR1q3AGwJIx2
r5WyTYYU9FeEj0kaNontqUUOEXH5THDVs3OYRmkN78v36Qtb72z8PSR9UvJSN6YVTfiOzPg+uQO3
wHJxD3nb7nNQIcJq3siXh/3oHdJdvQO8fhwe+Oc8L7nDbq9F9fHsOv20LmsVzswVLuRc4JDyzCX3
YFXf/3qglizE3k8mnn+Dziz3Mj9bkspOvyWKT/IrsiAsmJZxfCsrl37Qb0qFUBsmiQ/mmWwy7rSx
K47w3MjtSH/ycvibRQpnbfEZR5eq7h9dWhuOpOjxVttoVZ4YuEO4HTyPK51RhXlW7BQ730XuWQvC
wKhyeSjjlRYxAm/D3Jk29/6wXySYZuoq5iuRxtCYtJKhAUAlP6WsTPpUH4/XUe995Cg6iWUADTJU
cdl+yW2mNMf/h94tO65p2bGhCsSdXKyjJhW8/K+UnlUiDbUC7rnwfVTNCOulCpd8r1mGhtZAzSsg
1eG/pe8WfjLuz9L5XLuKy/7kTLDQtUd4QSJUSlsIu9kqjlvyynYEOqr6+SIgETXUw25T+8ZLFFKG
fFGLrRU7vwLKytrFTyISunKuv/Juvd60Nd9CBZdvN/hhrSamjAjW6OF5cMdbo7w2Zstx3+wFcstm
2UdD0QwvSsklLqO45BWd2lV4zlbuVlfzejiGtYj03hgw5Ipd0syvtTtDd0VzaZlF5I6VCWsdPFbw
5Mv6Mh3WtoW+tggGUaJoLPj5H1RVRXQfPPfNfsRhffdkctlogUg3t9uRuhCw6t4npvf/tOGDC0J3
rq6ryELLyjRUERRMcfiwCbjZIAbIJW2qdqLh1ugQQNq1t1ErLJRrth+pPksc+YtDKTiPKgSxCGBs
BP+4W7MciRCif/a6IAH5F6ibubJA2ydb0R/Zvc3DIzyojytkuR45K3I2oa+pNnqjxf3nTVmdpm3F
Xg2AQ5P/GwWCwUw3YKbZ4Idl95kavEEUlEAGmvcwo5QCg1X7mm56Fr4gy6S+SSmfEp/wwMwWdwYQ
22v1k8e+pKEreWPtbK4o+wTW+hKvddabK9Io0aURGt2293buCOsKyo/33QS/qbun1BNmwcvMtn9m
42gxyM9kfnd58OMJH8/psZHseoHtCce4FgU3vUpa+WVGtD5/CZ0vFNWZbw5C55CFSA3Y1Ycv7FQ6
yReYghRrjGaCv/oj/qC8nrkgsF3i6KMdbj8Carr/uBeBKmai8dTlCL3BwGwsE5CSkvfdPCfPbqDo
eBSYX0lZvLmZGD6bZdUviFly4ltnXYit9RbLds3wMZKehAz0Iim4VSI4I3H++Jc8KKpi2IMYxqn9
pvxVxxR8fS+Ayz0/26ZjLxtNuutDRQghV7HQyajiaUFvHTcqR4pqKQV4nbCsJkZfC737VimmADiD
yxtMrFaX9hE0iPgioT9IFxkpKUL/WAcqd60w35PenFj/6X8R557LjYWsagTzoUgm2cb3WiPgHsyZ
V9wblANr3q2uA/4enieNxT2cKFmRIfvgVMJj8UtDKpx+UvLWD0olm/JRKYYfAdWdbSF73YQgPNvr
Je3gGEqhaviwHU0L2VMIosDBFp9tDyb2prlrhQgwdPCU8wyb4lU8dgVD9EqjiFEM7ftAP1w3qt+j
XO0bOGJHGMxB/krQyrVB1caPqSH0eJQG4bFuQm2yTB+iEYV/5RsPPjmxY2OCDbHrTEl8+ifJ5RLI
l02KVI9Dx+hVad6qtAHO8mz+3oYyclp2BVsYqJq9p+fIr80LKAzqu5zX7htvaBsuk2ae/aD/gz+V
R95HuIDWQsGLA62IFTIhxLPuVN7YCms673H0d+CqgyQsAWgvbLFWn8wUTEsD5p9l3HTyh7rHifBi
YGdlgEdBmSm8gX8CnpbZThCsMI9wIS5F2bk6W4lvjg3D2l8Nu+dY5NdSXtnxm1+Hph0Szje7vEzV
ct6u4AYi6rIvvzMu9xkfUaFz8b2UOSnnWmY41NabcmG4scwGzHpMkX5q2Zc0JLu9Gz51DuLbqzef
S0TbddPauzVLMoJnYtDVJbzB1bDpS1aBJNx/IgMU5fBNUcVIpd+0MBYgTw8s3NvM41wU4jhQ78J+
m4yBPwjm1p4lEzX2grT7mRUG3eTP6PBKnJZwt+ENS5nxFGzgNlgMo/KhrL0rjv81j0VPs1qjjjYC
+142TQJHII/w/KRfcFxmOJgixeE7fsyy+U2fVygS1W6YoRhcwNftCkDUdfWF5mdElaHLWNfnb+Qy
nzt/nm1inO5IEwK7ZODAEc00ML9vJopAiSmhWeqdTJ3HtM+kE+6a2qJlzaOpUNgMJOQVGUE1QCn5
STKrpGfWlDcRv6n7J5/okKUlUbn0/Jz8YeSE/5MyMHxhhvWYn9JRniMzkmCgKw8FEwTQfJFNkR3K
DjVyS/jl0eeIc8yMbSy1fSma3RZ+rdrjVOcfSCFXswtn14e0ipM8RPVyhmsDlvR1fOdGhyJf5Ogc
sa9WMjbJ8KW1/CZXmFGbwZhyt6dSSC6ompHqmrB7pMnZxqhju0I/X1Cg24tnE7NRXhuHh8FQfs5e
9Qk1/p3KdOxCcspL0Od58k516ZuIAoPqcEY3pKZkpgEhg8vfimSRjQXg7b54nJdIdToyhgiDTZat
6GjhpwDuQ998talVt2NK4GVLJ8P9N6MsuXOki3lzdhPWyzmB1NGAr0jHVs94kjmfpWgQUwEtOblb
g1l5fTFZ055NlMLPQG/ByMJ0bxJrTp7+WZ9osC27gEMhxH2IfYm/DUc/h9AknLJhyX3ViyxQrZtZ
wP39/zwyF3A1IBSg3otKipKODZH/wxRW5mJS9LJsQRTI5Zrc4+/zDdQ5RML2nTGn/9N2TV0NKLq0
yAUhGtcw9wkTr0heMEX/qAtwpAn9ojQcWNKUNNpWW5Zs/TlcORI36ClNaPelp9MQZw3uqrSMbVO+
98tkkW8+DTaiWUuXSnDd4iPR0rxkQaMjM91v924F39MOzTdrOH9JGBVo2yYK69Zli1wrw4c7Tw8H
h7Iq2imFZLfIUUZOkuMwQv4xs8cZUD6JrAEOjqwXwrOXPgkKYBRTKVDkCqEtmtb3/2VgUHY7VRL8
w/m6wmV+8A4/X6G0eevXBphLEjA0QbRaFv2MVwuIh+m1f5nIwNAatw8oYUqmDLE0EqbvV1E34nu2
OD4SgvNRLTLPpFOWEdwQYQSuuA4lIPWMTI+Rm3zPP+A3x3F7+payqWjb03uAxKmzYmZOOdLRf37N
glMElszIlxnGwyV4IAemqRZepGkP70qSAHV/yWsf+9jyVMt1jo/cDGn724bRks6JqVAcc79pUWax
+quz2L+q9cPQIJjCkI/fOtjnNwSgItEu+20xFhdnCZvoZGPMq2n909fxJHwHEnvOZ4iMXsI0bv4P
MzBr6CZlukrfo8ExVILh4K58mf2JPOcXG63cIRj+YJv8y7dP/3gNMbRtemakNUXdQ4vq6pyesLFA
aTyXnfbtFPwQnAztSJ1UYp7jQK4qgxF/ULH3jA+a/QpirIlrhUYfvs4GAMcAyjzZr8mL4T7QLMOz
ufuFUbZtwWdn1DgzibNIVdaFPWOue9YcTzGAJAyZiNkeJGi/FX6bksgvBjuW3iI4mW7n4Ftz7KaJ
b7aaf0KG8lGY1BduBHSreFROpMRlfzPMNoT2LkTK6Yt3oxwBq+o0JauvOwFVNltT70kTGWuwu3Jy
PM/9/2sBX7Lu9Q4A9l/v9ZhEYauV0syGGxBSM5S7h5YCoMAEVfxJX8H6k0i+TPjfwU027oCJiJm1
uL96zRkLpgfni1GrhkgEa89czQTtDaJNeg7CECiPINWz26jZAJ/KnULxI/vY4XtoZv5OIG37jf2N
6asl6r03haNufOpm7jIBw/uQr7UuMNyexVsklsPSO5ja8WkB9OaPArGVEpQMFxQ5YqUd2uYBpp7x
stlBWBYuWkexueje18wRvZ/8RhCjCElJ5MMCEom+4QwghW4oJ15kypFKipooYzoAB2yjI5xpkcZo
jE4zEtaK8Q0ZksZUQyrnWz/sPHbHP7i8pK6K4OCCKAB+ywMw/AtsYO7/KV3QWb1UiBl9Ycb31QgV
nEQ3a7SbVbQYeSyecPWQ6kfknHszi+f1WR34JeuZf8nCiesysUziIxlYjuST0SvzaBeDFjOX0emu
WMUKZo1b84Y5v5UNNw4kjtV5igfcqrvp5kGHwQfBRyL4FAaVweKWe2uy0VPlve+dbG1bZppfG/TX
uxXr6eCVc3NfUcarIJ6G4cMNJvSgaC+p7oJdgbggb3YWUVXfjAlbrSOlcdm+Jy8AXKj/neR1sojc
k6TFCEQ6ElMmogQzkGhHmROds52DZ9nMn+I0LkJ+OXzbCu02Q9LzmzG+26Fp2Dczy1P5G9d5JNQB
96Wr8/hV/dzkcAvAjXy5HWLmN3C39L5U5vZQcMclO7ViCka3zbs/LqKzmYlj6RO3YiVaaujavyJ+
lg6uFu+O/+Or48sydRHNT/6oENi28xrF0rYaHyrEBfLSq+4Bh6Yt8t5mttWIAYo+ybecvofKbroL
CDB20zfF2dEkAEQCJe06rynX7jPmTGu7qmm+NqtovHuEBXrFSMSupBbOBRsQMaAlft1iKQt3ebyi
0keUau3bv7JDp+pJDkTEhWiIBWmWHhEI1GpMAh0QPwIcEVbZ9fI9Fao6ol6FqP6f0WlHxZs6WXT6
EPtv5kYbCeeMzcyxtn01HvhMa55P7UD3UGi5r6sEAKkDZKb1PFFj4XViA9Y953f5bqV396BL1MzW
9p7FT+PEVnIwkDDSmp6aVJTJ04LCmvRyORr3zZ119R1wizCdUmrra2ORuVcqnLUfGEqow2g5Rk8q
4W+9uXQWM61wOfQeUqVquWrHlihUpKdukyMybclcm0GMcsT2vN9B7EgiWdD31oDDfT6/llW6BLax
UGcbHImXKch8YNf0/V59YtdlV+7S16Ealo19cIVm9gNSQrj3cBO7zDPpOIp9gK7ZmPvOeIu+IVR1
M96UvYQb75gTT8Xm+3oGYwb7ryCoXzyKObGgq489Q6WuvwzSeN6K8RucumDk+LzGuHoronMC+OfU
xIBFPglW4/2aIdqpopZY5D985qEEtwDW9HrYyWgJqn867UlXIhCe+a7s2OcomZCNP4g8a5KjnKkU
83ugGG8NDKNwbjTHR4PS0vYAvVMVxWzjQ9DdsIpKDxbcJG2FmqiZdJt8wZVnvUD31TnJDRfLej4f
hldOuuu0ArnbV7ZBn9hpVzk2yVizzjCZDyAoX/Qqpv4HzUBkLcErwZdw5e+3a6z/12niGlOHX63q
X57WPcs2mhstV9RiOPOx49Gt/e/fjYX9ZkIM3CKv4tB2Bd1PDdjogMX5xwaiTZzVq0qYjPTwyIBr
DbhrBc4uK0atlEpyIs8gpAgYpt4F0mEe/5waDLPD5La0ZKkJTcRWkcCsfAVZeXqWtNiX1Xamd23l
p6yG/cwTzs+V7CZ42dA+PUHwaqNHeQiQT/VEvSNglYYyrFvjpG9CuK+0xw6g1LTIc5Df2NB0UosI
JZeDIm+jzLsZK0/g5I/C5/IPTcsWqfkPNoX/ImNMcj+QCPRYErv8uwAc35/ZGn1ZSdAqFi1KQRPN
2cbrsbRN2z6YMhB1uZUxbm9IIbERTqx6t2T6hvelb35LdZgoTnrbfyegrAqh2Tonp+iRStrDh7a9
h+X51wFPlbCzuHZCJqA2Rj6kZqajZ8eUvTK/UCuRnx+lxMgBotam1oiq7zk2NDhaNPy3kVDRXkbQ
eOswrlWtNYNklrWXiDu02ZdxzFElA0liQQiJXcl5RvM8+1bFsuDT+u+QaNt+ILeh24Y5lpVkcAXZ
pJooXBjpjZsQdCh84iykiE3QMJ1M7h7SOGsBXXQEBRf1j5bG3G+Aa0ux9cvNVIQlLfPqs6vjMCTy
jfeNxE2RjHVsMgicUZstHj2NT+ZG+tH05CGM4CBYzQGHXHALRX0NAwzzFafVcRxdXs2f91Vs8kKW
viveWfPjfjqU0oH2YV54VP3yW6Sy+ZI1h4w2H4K24l7fuUzVAjVrxnUj5eccBZMKthgRhNC2NqEx
+5hpwBifHqmzC67HcnPA6JHQXA4E6ut7u+gkB4FuMd8Hrn1Pjktz+VH+EOkSUxvcPSVDtU9uhH2n
HJsUjJxDGEUriGLmiqwLcTP9V91o3vFjjtQ2LzGNjOOOQpAsBozXW7VLZo5jhsBCldnyYtSaoI9u
4dybEE1ABGQ8JJVhIrWLIHvDC8uOOS/BEb49/0RCNQd7mTWPmqiSqt7HwvPZKg7uwGt0q8Cihpzq
CoikewEtZCP+ro6robgrplmz4h47u6ngra13dPo0KceIE6z62ia1QwuGnlJgVvPvamQ5MCzi7ac3
tSngyhv27iAvJLBkKo8hsLeLGZM+9LbAhYzN2oxnBybWb5kftOsFjOb5xzomUhSS2DQarC1uID7i
hqbkbhP8TEV/aScTSa0QkQfNSYbJidvKK6eVXfFbLkpcrwwxpb/WV2hqn8d2AvdEKxUjjzds9z1P
a6ELDt/nBmm5Uibz7y6uVWpO2RVXOCVznOk4TOfK9C6XL+dRA44ELCSW6JCq/HTnUqwZ4RV1FxTs
Uo8i3PJQJA+72bcFcfsqRUmgJFjojubQrN8xG1S4K4wUYX53/4WPhSTzbzDzHSloxl5r0XdAzyA/
vWXL3QRT26173ep5umHeIJ35BEusxcTw97fNLHDRgwudrnmGCT5qg6HIEDDTQceeCglx85PqeASh
rVzxpUo+ny80F4dF8su0S6epVHgaR2ANAUq+H30qAhlSNp5rp8AVJYtoyY7kWZ9DJ5r7052CNjN6
Ox2QFbji9IBWcz47fg4Y6YSPQiV9AUHxZhJ0vWwxAC6XHDIIJI15yRkRM2e2jLsaI9ZQEc/ZZZyw
MUbEG1Mw2+Cap9CwQOYajR0ehC3SRrB2ZpEOO020J1QR3Tu4k20WhVZkkS/buTeO323kvXGMKRJB
MiuIRIh57Q7LQr0XGTZuRnV9c9hTG/EGKYm5CG5fl+3HKZM4b1t3sTCehiHcIaFCgd67jvqLG6Zw
LQYKgldpJiaZpwjPSsBEztNCyBwWbtEDpO/KX8xO8tM4aaMD7m9IWzGpDd6BDBbh/eYbFRgNH3vb
kHpNMROE0KqigQ8v1AbEI4qxMgpNSCbldD+wpAH4uis2FNC4DLYs8IkQDoch9VeOFacxdmHb4uTk
bh/zgmYemqYibteTVG7dwI3BzsWS1Zl7osDuA1L0vsaNMMUXXXeVgPtyRV/L3/9dlbYXDzv1RykA
mls/mdkVrQh9wczT+sqNCrxaxDNuLr/HlLlgS2D8FePalOX75qZOV5v8nGvXKvDip1IwD8URX+gM
5hL0Ahaq7wxx2RvN7oy/XoisSVtqCPDnOwuBUeCJybNq3o/vpu+DZDggZXqkJ44Zx0QlGc4ubR/x
8/UhM8abe24x5c7W2qYzSQQFzTyORjMC8Sm0nVhRi62nndFVE6IPKNGkmPD5g4NmJm/Oy2FQ28vQ
ji7HaHf9/9kT6k7oreZlnLndVofBL+egR7HYFdEDAC4DNoefsSnvvsVe/GPEA3AUjm/oVw9COfts
O7BHhLTQbDGLJjUb9Sh8p/EYqgWxGN0WxsPFVpgWq7HPxRrqcv9fqrwKO4XBTSRszDJxvnyg5XWr
Pfo0Nod7PZuhRPMfEOysWo2zwqyup+biLPKiubI/M8PFRkyYevQ7xZHab/lUcXzSJcXhMHPb9P4W
3y8SXTwspYJikh/w3is4Z0T1nXo15hDW84/LR3hboIADaqKkKLp/j55qen/OQl6kWHMKRYsPhYOJ
FtF5pcs5y2EwDM/HNbFUzDkazSUjK/mZLKgX/Y5V7UCx9TmfGqI14o920UHszfXkq3qtJwucxOuU
xV5M8H+SCGflnzzlP1Xg9AdBAWRZ0M5jCBckoLuxXCn0xOkLvsOsGHY6QBYWoEfP0XdTSiRACD93
lPQ7t8vpK/aAXIYok0GiKIRy9wzKDTYUY82RtDchwNwg1NiSoaRWftFR2qvY6fFW6Dx1X7YoBIzy
Zo8eCUOf7WVPr/mvOuq8lxS6fmKrB+0FS6lx3rYqsYI+p5oSbWuCm0qwnlG3EpwtAxIxsY1kpHU5
sl4A8lJcUk0OVAT8CWPHB93+kDt8EikoLQdK0KVVFi8SFn8ZLxVxtjhGbXO2SmNoy8S8qS06x+Ig
L8/tiL3rDvfAlME1WchjhQRZysJabPUDve8+B7cpNGJb/r7Cf3yL/By/wxeAi2WPVwYXt8Izpmwx
CiB1H+qeBlMAqx053aUTM1+Y6bMWR7ZzHlrD4aDheyxW8mFelrA4oUAC8fK9PX8mcCfHV4NQsu4t
pgIYV4C8FddOtDtNtu4eFacMPaXeMubAjOsnS+GyjW7fkb6TSjkJ+798Badd3vyxe+bQcn11OoSM
MJYRSIMdhcHYTQ/oApqGoONeOKWNdYbOPFXE8ln1L/2/TunnI4srh7QJitvFDUBQHfaYUvsGBb7Z
PYUCTwNgWgJC8j5LesWRsftBRAe+OE0QuYfFzYDhYKp1I5wbd2EvZWq0ze1qrE3qS8OpuVrsZ42B
iE7CUUC3zQOY5zFD52thIwPZBn3y1t1he0YiNxgwB1Zx6lPLBhCVZeHOqO5Oq/cPtL2LxFLa0IgB
YNFNGQYQo/Rm/T58xzW/fjnEyspPo3Lzt7FJaQVDZEnN4GEcqGAgIMGsuStYh06ZWyKhCSG/34jp
sLHJWpLVP1A43EVK8YtsL1U5nqJZ0d8pgr5mITalSF0QTRrIB4dN4YPqBrH8wMnQWK3GJ29DFd+n
wS8W0vXhl3pJQn2yzUObxcbRAvB07aM1MHVBAVL6BQy8rNxnS4Kj2JQ5avjOYjsAvUhg2pCOZ0iz
7rSBXXcJOyC64iTXesmMiyEB4rdvQKXPjGMSVRvNwoEII+9DCEZPtUqxZtq+k1GtjiB7+7KzzVnv
kCyXPmuWzsqhOB6jCuc7PtkZuMBhUPHRaeWmxEU5LTkm6SkhCSFSTD/h5TXT8sm0x6Uu02mtZXMk
+uBfcH+Pg8wNEeMLSptkVRS3Ar1Ql8b9pbhYT0DPzXAdrrMMd/EudkVEIXi8JX1bJjiGUD0N/3jP
scriEgiu7phWs72ZhZc02rENBtB+YskM+ZR79ElYWNGapO8qE3BfmvNetGORlfn7gikBaksRU6TI
i91XzQbmA2xoGE0lNCzbtR4qZwMnvTh3SlW2bWpnUA17//G2/xCw4u9VFloJa2D6oljFy6SKxHqI
VEofvKJ/RIaqJJ36eIfHUDaC4XbFmFiwKMGykPv68DjpdCvVSoWa2XQd83hPYNkPK1nwDbyDLmxo
hmc8TYaVfr0qTmcn2ayjjv9axxBAEnXfifsh1AMnB8Nkv2K6pi1qppZS2JDHJ2OOf2ZsQjvcX05U
Uenr4CuGspoKRxDMpU6uCj1yw75fkOj1iid6llLrYCB8WzBc/4R6ssvG0C/NGZ2YNaaGeJQ2+x4P
KhJ7CAbRrOsySY3dQlT5KYcg4I4qqLoArZlg0Y7YDlhk6NPzVk9Ks/eitsKG7Sr+vj7dWWRhxMHI
WtgUkH1NXTf7y+cOyxpL+L1i98WO+E8H1cuJPrvvAtO1774GqqRsC2hNGDHRU9mfti1VRdmcmjF3
GENG3ecE9NWSr4W2Iejoy0Le4dvUBy9RayaR0qLvLBq2gMQ7EZxGMk4mPUqQdQulIidKWoihG6z8
tg9gyorA4duKHWGYPofNDqp/xVNdz1fIBVvY/Mk7Nnhn96gjtTHnTaRDjwqniRFJxL70kjoFhPQR
402xpQq8cM3vSAVuE/BEW5of8qs1FNHgfY7NroUdEYs1l4yJobdooUugXKHrCg1k5abELIA4+BZc
SyguEcCHeVSrNeH9s9ho6SQ1qLpdaljk2SwmMHmtD6CYvNtuIi7KfNoFfviUQJ6cBAYNBtk2K+oK
YbqrU1izfYE7qeYuC/Fili9wQPMu8CAaXGuTJqMxOtVGDZSgEjCvhKgvBpgHJqK5J9hozvLVKvl+
HkW5PpQQgUxmkrVQJdmbjyDspu9slE3/+zRe1/hDdFGbDalRf0kIwRmuUZIhD6kBlfDIL90YihMP
kqKxFD1+4vrSnNTKM3ywr+sCEFSo1j3M3+AHHsOu6Lk7cJBTZS1cr3zGqLquGDsL/8kZZn9V6znY
w7lyrE7THxlhEsMF7CSOPZSmxZo5sZcgnSp3xWtW4X/YFPudzGtUv75UADYHgo4rTyzTNBhFu/w3
fIliHBfyQNoktdvkZvkaJJBCWYvHaCBkRFjfMwhLzKAmW9FVv7lv5Z7rY3fK7Hl3x5Vfk7bzk31Q
+LlliLc1TJ9jLxSo6S3lrzJ6UsKE1qWBjlW08nFUnzQtqTfMy/RT+Y5iUaLjcZONwZkRJ2/6jvU/
2xUwRxE3Y8FjWbBMPUbQKSO17S6e+hEs0zGftkX0i/u0CPQUw5GjfP6kVDBUZFJZlgBZ6WTXFeJG
fKs0yVlV3C+CchScjbNenM70voHGHinOhilggq66kG8pykdRtAEq1U/SU1ULL3HtxVkNBCa+R+A3
n29ag8mfLwmwl2al2r1zfs5bx1DoUT9HRPaPPQTXnmOCkRRmYfrX72lGR8iBE5OoIO8gQRcWLBm+
f2/p6IHe4UbQzaJ50bRH4VgLdt+spRcjQtnXGiHNvNN8ot54wZkeWVbwrDYV2NwT0lta5KiGX22I
2Rr9WpP7sdaR2e3Y3Y+mzTJv+a7DEKYJ/DV/kykst3xD1+7m/lrAUfUmX+czbI2z7puPhRaQYkYy
TBv2NuZh1Sd2ykQLXCRT/Hr/XGQrjEibVdKca8Bx4zKMEuAiHEkL5Nb5TGIuLXdPskrjyrijj/8I
OHTW1aHWrnG9jo+Zai5S3Ar1uCOxynyKhMLr6xfuGP5ZDQXh0bRuMuRZKA8ncUm/TJoGnojvOc0r
L6GbeJ4OQacYZYMDJRU0vQPQ84mgKoVPEIzc5n12IZNtLped9v1aZrbr4/QIrRDy8e/G0qWOPQyf
Er3ng8q0rDzXiNznYS88feeo/P1uImfLs3oEh+qCLdZ6pxc/rNryx+SQtnpU06CBP5JAWNqp33OX
J1PCH8ZE/gaffWzkgU1lBV1h9cYa2n8xgae8jLLa3sWKEto79kSyEmPKIGREWK3wVlvZWz5ykB3Q
ycYG2DOLDAyTcGkzWB7y0qcn6LLaVLFZLDngckvRtwz6LsuJTT//7qGM7YrAzVYNAe2sVRJf8pV/
qjy/L3DaJTd2rdytO8VyAb+EI8ySjHNfLsDQolaVZxtjB5qI25SPnerHHZ+S/8B1eIMDiKcMO9dQ
IXLNSpdZXwJGi5EkEkxcxd4ZJjN9VeKZP/LXk1y5MhKZHJoWBUwevh8xwh0R8zRpEN4GmTCYRqTP
5rXAz3aTQFgsTxKq8TwWPNZMLzkqSr+FeLlos0/YIhPzTf/XrkcNVC4OiCqoEuRdISRNACBHecuP
HOPFRyDQOdNP7EHoixv2E5MyFWBen4l0eGxJUxAfQV5ukjAPwwMAKvbmAjmv2JouODfS1kp2hIe7
Svu3WIcoLcyVFIDSY5Iw8WPlXJsfB+hSakFVkym29H7EDhZ6d+EIvK0PYB03a7bUnDeZ2CVsbRdT
lbgdXrPaT6N0Ro3HMzs7cDri61NkFiBL/yiZriNzBGZFuqFlBpafVtj5icKknYoZKzqNbNciFnD9
rdEgsdf77IqJhC4+Z76Y0i9+D8MqlTBsxodxbz46qVO9yXw5gfL68mUcQeNw/hWaATFaZVQ5F+zu
NTPjZr41qC1AQt5S7/8SU9guyEFkaIa4JleUVztwxI2/H/8TKhu1wOprlbZJ4R1DaZUpTFu4463F
17xtMASWxYQq5zaZlnqqlNLwzxzRYHUEQrLH/DjkyOSn8CnOarvW6AYMCfkSXVvglml8OysAUTMP
uSHa4bCM2lkxZgJG/pAPoOobrlxBN9nIxOd68g/ik6NMHmbUKkiSM+oqu0etuRd7IrIR5PMNOoPm
NwN5yrbd5kKYzzSqzTp/4Bv2xMwgmGSMi7PHw3zn8/QVwvNWxp0JyVh7SLtTPDJGhuw4u89D4Tle
Q4c0AG024BHKrmigORwjHtHO1Jm46n2q2SFROHdAe7vwfTaBIgv0Qfbp8VxaE+X6DUAm4Ea1LUge
taRzj2Af+TYNvnrA9ieteKdkxhsncPbUSLoOMlUoKxWrZmEOojd7OeAmdps7KdGGhZ5VXidhGrju
Z3YejRtEyRU4dz96vtQG/PKZ6yuOMEkVlWZSaVkVo4JjNHupJwNfHOmBszAbTL9Di0ZqkPFb9sGg
IV9JEWkw1zAcrtvb6mO38ABoAD9mvVDPTbCSXz7/vy2QFdoKIM9bneMLul1gdcuOUK9k+QTQnLWh
8JTBNunXXCjnHL9Lm5O2Arm58CRefBL8QTqze2HUYYkaUeEjTTwkXXZVXPngJB4vq5Ladl7dYLjN
PE189/HQYSUU0cd7KsFY4JI4yBjJYH/Om3TNG95AFhwdXq4LMV05EwhNeiDtmdU72dDLtxLu7/Xi
Q7cnUxCkkkcisU14YvmgTAHWa9a3lZKCYTMrjVQ3Jsc6fGoFtGakRuz9vJnVecCxSaoTWMWNp8dq
oUEph9xoe7Szd642qEecDPoLYhyTQBhPILJLqpSWQR8LJ4uqyjxaXXFAlF2TNzuJXfoZx38+/lcd
Fo2ugR6LvGlg9UomdOj53XykCOtfQSmr3AxxuDu6mPFprtdmQrV60Ft/aLUg1IhPcMCVApOkS7kF
q7ehdtoGVDg6+EnQoODbgG4bUfen8a/s2csSMTHlqvz0+DUQaSWOUD+iUYWOts1jlbJ+KbDsnbJ3
Q8rHp8++2Uk8eAcyHukq4YeE90MMz7w8tHYiZJ3AluQN0nxMec4rBIKYegHiEOqobGJEt4yaVu3g
Vujtbj2TQdSWDmh5dsx8OVFe5NIaUjSQNEhs7+eVXqXuhaOwOLA49mTriWqpP57rbuRatX6MhwZE
fT243cWirRmDKQEyMmzY5oVRQv+s6OUlOgVE7zOvEtYxzWHVqzlMxwGkvNr22xJw4o2r4yRsst9f
nP3ysg50/k8qBNRuL08BRPz5uYdIsntRAKjKHrCQeJPluVzhmoAT8kzc/WDBeO+p4BfdzN/vXrOD
Az6le6NrcVcTRA76E6OZZpy+NInpBg5YkRYU0zvmqvBAuGfZRb8zBP/juvHMNWKK2lwTOUmqexX5
POcqLg9pjuStYAQkGj8vJ9mF02HZVG/9YvVMXHh5k+zl49RdioiSuy+jlUSKOsUJ13OPaIWxBR80
tLPSOWVB+9vlDGO36tGDiv7W/YPPV3qgRJAOpB05D0WwzoS0rinPqbO32XnReXFeSt/0Zk4OnxuQ
SjP2LaFzVUBOdRJZ4xMnwDlgux0sMJzIsRAKgnf2o7BasBRIigiACgOPQN7qc8IcjTILtVZC6D60
1rIV6WK011rk3Ve/qAWPHu668PyE8xtR2QEBR2xAAE3RVQMd4av8LAXGC1jhtJ8CjwFiaEJuIMyY
Dg34HcAn7/ihFgWa+XcbhiE1gGi6vba9Z6AU/8JCqmoiJXIt066Ezsl8BvlgNicONHrbAbLque57
n3yI/Z4RRsBSjt+cc72NejpHghjtEU7jOqjPU3LrSOqR3mWKrbs24fyqRTt2jeiSbXpGS0+iMkU8
tDhfRgQcxyXJ4z7DxuscqN6RTL1w7ZTXfCkZXxFxQHrb51i2eWdhSIxL7NiVZDzgxhOenHRz8jks
4xiNHymy1ZIDbkrzDQmXDHukkwgTayBTQ/cRuAbpBT+RCI5vQj3xARYiZSdZwt5dIruvJmroll0A
ikid9hDptPxHFaTpIecwIc4hOUMVVdoSCd2MapBCPmtUgp6f/2HKLCq8V9UFoPUkTCJVtz1tR7Yq
aeQslUcwT8ChYdkSWGFwcQ/IYmRhZn0JKOq547PfiGpXDi4VvOtDiYxg9coMdx1sSgaEJD5Qaljk
9dsy/OMNpJAx8cEICoxu4OIYJ3xUdMd6tAfEwKiqlc+scW8Cini6AcV2eX7K31jdwYAPOz9Mv3Sd
ux9lW6bTiJAdjgXfJzHSxcoG0qorrkSAKgYo9188LVizl2afBB2qsOSqTnHNUccIr3VYVhkXfM/R
t0uFzgSbmJ/SExSn3S0n6RyJ1zOck6JpVPeiLah/UvW+2vzLMLu2QnnaHe6c4v9r1eFbZ30dkOxD
XtV7k2RfBvY2xkoYxN3j9Fzj1RHmSEkq00/s34853LFLj+Kmfn406Zchwc54pTh3vdXkH5ELdhOo
J/Wh6nJaqQAP1q2hZwJYAgUX6LiOzeSo5QPjo13a7dxbibE04qoqyQtrS20Kc60EDMk1Tsy0Mt8i
YOuHJSg+2OsmeFU5jUTq84pVkyjiEHhrO/prNEGEIilfPeFVG6uFogCCx99TYuaRdge5iwyhYjB8
BilbepJAgtkVGlw7+qUjjtjbmBQhaHjSQf+i/c8kIXaX7KqmCq9KN6GTlswaLo61AJtsDBLJ+Q1s
DEKUOvUz6+VbDytR+C3HNqNJpjdNNkJ56rk1wcNY2fh9TugWoRhKmm2Fk90p74dQ7XKdiaVhKqay
sLY9Jq+LgWeOQzyIqUco1kPG730C0j0Ut+8nzYifvRGZexLzjWAul5MiJH7X63HV9GlfH6FiFgx0
P32z4WeEMhOiFpYnY41Al+NMeQadGOF92FzLC1qBrnelrR3JgKydJXKbj5VvK7GosLLp66+vGOut
w8h1mrdCl0CBGR3aD7TF4iKytPvY7oxU3rZJoZYCv+23SnlhxTXiOVfuGajfCJehGm7Q5bDKqTwI
IyVD5THJOFO8VwGGtXsOfnWNMKfyAfCIVA29eSXC8Q03aI5GJ+zrcEU5nz7YcWRrYEjfnaWmHSv3
dryO4JWWa8VM7BMPVuot5ixyNsV+y4vGaR0oXmWVj0N+VBx07YxEdKXeAGOzkGlks3sA7gorlymi
075Cdk7bRXGttLlFLOwS3GwL3WHO4l8sp/kjawdYa0FrusQW/qqZwTmCRDB8WOigQ/9WWRqbXTty
j1YYDCgKZww55Fm/F0uePOxi/RcTaXexXtXsuedS2iUrL25e8j86yq67LNGHdKYno0kh409Zo/9e
VsAhoG4t35b21JutOpeueRO23VRID/wUpjv8HrAnjmB7EOOqa9taGpXVdC9evUIcCn1JkvD/ilki
aLgVwfeWyR1XKEKcJsK1WmxWkyFYGk/RVL2Y/U7InaK8/f7IUQFyq+OPP6Lv4UkNPCmp0DqsHYGa
i71UG8geju1pcOi8tUjqqYpxcFFBO19QpymTi3L1H2cuyUkOmZcruvktkpgqWWCED+bOdqY+czWx
qbKlzsbCu9ULh/fyRbkZG7YT6PyFQ/7upDyXwoFxsj2FSMKUqU9NNFXo2ZBZnI0h+X57sNVq2UWB
6zUBGKQ6EYObMigYqDetoAsEMf4CGJ8l/Lw+trWpbzotBEol1WICvDmJjrAaliDKk4KySTDGqhsP
RCeRXloJmOOtgH/Ti9Om7yNK4OvtiHpy8Qmhd87U4GIxSuNM6AduBfYNzXdo9et5xndFh5AkaxHB
qeP5ULWISHMSl7ekkHp5WeHlBu+hhl2oLS5mBrhk/Mo6pCGasGVw3UPqNBWKYGPm/kgn9NTuQNWK
uupsOLEFwBvPvd/qDrnhxHHdrkHqqAxtz3ZPWUjjqpXhOrfHveL0ArlD4mGRmOs+YeXUcvL+tMBk
R6moNDE5BX8ofKCo+XzLjZH9Uk/MEIQ9/KiVyjeXH8IBS+QeoN7qn2fyb/6tofi2VHdC43SHzn64
GnAccPZhpMb2OPAlUrckGuWPUPZMPfX0/0nEZCXvRtaPgCa6kg2DIuKyYE7kLUckGhLbqsY5LCsH
qb0ihDVsViMIE0lxvnU1wuh6y9txSrqTjPYNHpCz62aRmyOuTuKiiNOesUy7WgftwTtXe78m3L58
rxGp67acBk6jtaDKZ9BZc4RJisnf6AJ+64fkhy4VVe/Z7kJB8nbp7S0FC2dv5JSf2MkzIp4KLxhW
twl+zENKB2N/yurGjhX20d4Jzg5n4AL+17OyEXccCRwe3wSOX76f6kZ+ZEoqDbvDZHTlrFEJx/NP
9hk5IP78EVe0zUkVphEJyinhUQwoWsftd8Hsm0bqoO95Un5JPI63UjFJXGaqG9j4U2Te/0JWl5KY
4wv7Ob5aKfhWlsDHEge2d05hy5HaKn1JlSmhBPSpvTlwRq2CMluKpIErMScKW+VBnD3aBbPI0hJ5
5ioSYJKs/U6Fdej4b3aeOJvLMRj3TU+6O8OeMOsddcGmXjFYyvQf5B437/LKOnvZze+uEYRjDRqn
Vmo48jyLuEQJQAf2nPzqKsn/FB0JyX1hzB5klUhroAqE7iS7o2qJo6OFFxJQSEIeOj2UssODKjK4
BFhxWOKSnAhvLHITSfgh3ujaBZrqSziRmeqU9hKWdkU2S0A5EMdINJY0ehOtL0nJTOKC8djkGrkC
XMxue0XGTOeS37/7Z2tNfOrc6zXUeVZAVatNIYip1skWLYD+55Q91YgobpC32XLIwxOSIEM31Hlq
VLj/bQF2xz9cm/hbJOqLj9C65Uit0TeqTeE9/UrImzwKZeID/k5zQz9WbXwAE5cdn+yaLMERG8z2
1lc4Pkwq0f4YHKfwu8S9DMCAGG1Rw1dv5dxinvwaPSCs7MlXJ7bEakyrr+blLQGaS4ha9NcRvXS/
kj0A4EkGCQqMtG5eR1MfqqR0ue/zC0KPn9oCcOeaRiHHkl0khWOPNQXN/+aKGxvpSOloe4+p+lg8
9MGeVj6aRwDGXQng+AtFEfzzcx/FDSjLis1fE724pXtQz8TSP0/RT8U7Pr/9mhMLHLL34n/1EbXT
QEMA583YTxAT/xc0NEa7l8nmh4p9pdFtucUsoCO7c6W/EiLxQPFfTAi3qRuHHrfMkGhI5hRgZdUq
DVXg5uIEdEQN8dzJLhn9lsBXR7S0Z+GriQxlriaHWx+j/SUQjARrPmo3CHbo/vsCSMTyCzmHPtgV
dEmC0rN2eVi2Y4FovOs+XhKm3LMMEOJCB649oP408+fVI+7qwhydzXsdf6kRGhB6CypZGKKerHVK
b47mI9I6weTJ62yuV59JaYRkySrEUlkHptfSQga//ZFIMftoX27lhOcaqkq8ibWpJEQD2cWK8cX2
XC/wqTeOeHF7osSus9sbovxM1pnPmJQfxEbom9j+JMrPOhkRINLKmk9GTuHesu2bIZLo2aHXc4Fe
GL+BnonYy5zI3C286Y0PPDqBPzpfodz9XwQ2y3to0Ztq+c2T0Pjg+z3cEEFBR0In9A/fHTpOwxco
x6A2iOoWdC3c/sdPe7S+oB9soBdf5fW5HMxjZX27EhwKxobzrUJu2szu2gJujSZwXTQGkPyrhlAL
d59lqFn44GRb8Cn5UabfxNHh7M9vhwWl/1Y8fzgrtD/f4kUrsP5o/8rmQUZvQ3mIjOK5Yr8ZkOfL
TRKUUY9wR5a32YJBPTp0ANXKQV2kkqbRlm+ZMEkJbRGbrg3EhDUuQk6h2I8lIDQpy7LhRUGLsyNz
T6wvQ24Nb9yguN6wIXlkNXIxmkgTqUUpLIcl3n3hdypwWKpQZwOrN/FzmYeHEhyhc9XOpKOOit/0
YbxJh3oca+7bIfADDfCSTvNcCUM84o4g8qvxlZn5/5WNA2QB3KoXSzvkfzKXv4wIlNmLLiby3/6N
v0fOLx4sonbu63IjYmW3JwGFuQePgJemX+U2mi3Akop2fNWUHIgj88UseJBuVZo3miz5g0HKPKYB
9W0Sp4KH8cgnrnQrGT8aj4r5BM6eG4gdSPp0NmTpd/J7CETVJY82JTGp5ibhN7wvOd5bhhj8Q6Mn
SQNw6Q7Qt5OLQzEqd7rF2xf2xA906pttww0CAmCuCwLdyWGM4EAkneUGP5aw0Z8UvirTjgmK6pXI
WHaqj4ugZ9YOXOJG9CsnUoxVE7z5Y3ltPfY/GS/ItXcKILmjisrD4s9/WlGX4BNjpJYygoFbV9Nu
Ols0mxbJKcXVj/2m7BqEiC8rartN3oeGprFveBfPxDUTxdHOqTDtcY2VPbo8mS2MZnqcWxspRIVa
c+/chFXDsD1+gEM7SOdtTjsQFJAWQOlHOND2QKHzBaH5P93nwh5f/pKohnNn6aOlFZJaO1d1qfze
iyrIgfrmCZgCC9qmuufwRdZfuxXrcj5KnGJmOBs5fEzNcYhAPWHZEWh7eG5iVUN4H1DUtugAuVcr
FrTboCxx175P6vwsjL+ElNZeQo1B4Fl9fgjy2KxadelwD9ugoC+zm4T/8dz2Of+VoYUKtYclPEzR
3LGqzIipVtXkV8118NpR8iiwKa3MPmIEQl3fLT0Umpq2cl16UI0F5ndBxbkmz3jPvfIKDjOhEx/g
r29gxyMdqh6cVPgfosXAl3nlQfG9iJDTkErfqElPq+36ZcntXuRUouObRA4uqYxuMll06P31UbWp
ucSAEmUhGFX9KNud+Um4qr7NXbYuuqb4XoaBnLGqwRVU9dcGluWkk3jzB6CpYyZ8588XHei05qmz
9OBYYvLrkQfLoJoqcdhs7rqwFFwmRkPJHVyAsz2R18WWxJ1aOGqkiwUcrQ7gKQaeu1doaWirCAJM
Qhnhxy16cTYB0FxEmJiL9gLX5c7PauCDSXj2XhpYHe/+NQqEd94E73cY3Fqs+K6Gg8Siy7ntQzX6
Qvdz6DbLypk5dKMZy66W4jveUgi/XfPLjgDu249vB8HdVTkmOBQ3qCqSEcxd4s8R+uJbvrNhiqex
DOnxZWL2odm7zxBA3uYzjchWtTHdb6N5TN5Xn4XWm4NflOcAkYBGSyc8PDHzQhUD2iYBKPkpKmPJ
0LemFeflqNtCtR4mQjgaoVCFPeSzyTO1j856+tY7Fwb7wqmGQU3g/PV7si9Nck9ijbjU6XevCdVD
Z3vht7gqPEkuw9yU2dCBTQKldGJXdZ/HTRaKD8QZiwkpDcyPSSDI/GH13Z9OdbewLsRkpYHMAAqO
L9lQMjsg9uf6abtFm46E5k3wRCahLzcCGvQkHSAlWTQV4JMnHtz5/ZjTCQFtND7L/c3wLUPVTygI
3GKOpZerIC+2tjspZvrgXtayJ/3ri1QN/tqGl8ZWftZTbXNipl4icTvugWW94yn7x3k0kCuzmMUf
l2FROh6swm5az44u43pF7sEBJwQGCpLFJdQGM0j8V3WUaHbTN4zDM7e5g5M0u8+vp5ZDLFt3vVRB
gn0ye4XKB+9dDfxHNPibj9587vJuZGgE4xV+GaB1cxpvd9OZSH4n1a0aA4xM/hRgqrxVVKrLnqOV
Cy1CsjEX4ljAEVfRJqBUVLL5EhkDA704LiUwknsOQLCfsQIpPVR8Og/R64xjoW9jeIIWzjX+NNkv
WWQbg62d7o0RmH1AMVVmNTZHRRMR/JBQxqMBL4bRZx+dw35BwFHXo7lp1MCcDgRYQFwsfBGGKgPj
V1eEj6Adtp6vdwrjoGYFBfFL9fNzl/vIyamlD21l4GwLYDpQHGdShFyAYjLspjgNzJrLNei5YeV7
vwSb17apkZuycfUj2NiZTliciFveyys2C4B3JR/U8JPRoXEZQBBY909Rr+hx4idf/BrJ4cYFmukk
lq4H8aq8EQJF5uFpU/vToxQ36RsFiRYsBG6begBxn70l9O0Qwfhwre5Nu3FlO/oX60GglDWGiFi9
wRTSC+pLbxdnMYxdU91Q4kxpEVlycOk/jgi5EtSeEgMht1ETh3vfudAamxcs96fGfunw8/95zI7z
XspQTjCpPXMS+aqry79v93uezmzBjri3v4U+TfnPIhfJMRUmx4xeyUipK0HMEgPyLC/2jyJmO1Vx
lGDf7+6tqPKBCzC8lup6u9QQdBmin6YSG5I33IZng9tkp2XPfHyl7KbM+vqcOC2++oHilcS76zjw
08hQX7i5jjTFdvKF4vpo+tJTUvv50VnpQFV0YZTbsfHMeFKh2I/LoPv7IaHQXWnkjvfFpdMKVD+/
8pVZIUcFuVrw2igiMWBR7dIfkwVjwSc9vZddIPNlRlR1WyFpG10b9anwQ97DRbW90D5MMMNA2QZq
wbAPMem8+HBCM8ZyjzzNiS+WIWAE46jby3LbKMQjN/s9lnIz+5fcty4e9JH/ZdarRw6cJAwSH18S
QalPg4k73sGIajF8uxePYXEEvDJQkui8hGAms2hS+pcPUVA9sjCcQxjn9HJ7FQpUgJ3W4CpI7zVp
8402t4lK2M7F8aXI5XKqDda8oDv7wltzifXEIEVSC/S6RQI0rP0EOvo2Hjls6H9dAJcQ2rlalW7c
G6lGyTIyPjtvc0lHdtu0TjwPVBjuU7hCa8GVYHJFbNbB7NN2ITBThMcvDbkpuxPqrmJwv+l4Kc92
7Jpg9Sv4laCN/iZXZsf9Jt+VoIRuB7FHayEX3BLUEfNlxgdG5JM32H3NWLyKywqYhTd/LAdMXYOT
RiNf5B42AY28ZLMYPDZbrzVr5Wjt3AGb1xIvHPtR+kh6cT0yoXXsukwtL9EUKhXOmNK1QjginTSH
DG7anu2rM/TtY++BGloCFBcbAQzBwvNOFFOYYXsjnLA6+nB3Rx/WNq9c7skRuzO/zMljCrWRyAKP
jx2NhPxJ7Z+B0F1PdrywwQSyvcHTQto7xsjfAf85KOgxGep2IaffkFttRvD2Ro8Hy6GCwvcPjeuv
xMuy7l04gIL2HyKFU9ph44SJeqnZ6lYIG1gU50d6vVvEmwOSVbqgd8fdAETRdBWb1Wmg6QyKarf4
4xwRjkIc/yjhRdhPjIEbFcUM7ATkbIFN1HhKo352HAzapzNGB4RlzCGMa0/C4DTb02VLGNmivKP/
sjvHuVilYTAIZ5rE9bZRdieB5DF2C7sK6mSPX0tk14yMyQlFHiWcq321+06zShvODjE5fgxyf6jP
wIA+lnRPoqiQqrFI0DR2bduG5TjuMWqqWWQmxjyeKiiM5tUgwf8TdghHl1MZS26rJGntqWJpSH8x
sbAGVa26Sf5X4OLQCZoHIep//a9G/gobdu5p2OeW9bpq4eBMbfuDLt0GVScfKYf8iJ+8Skh0lA8A
v7VBAy+ooOBLojAbz67hpqi8nT3N0vG3ZkuuBrhQjEiU459k0h+wnGbau3h2CW+lYr5k8KR16JF3
xnnQbWGLE/POn3yNLkZo8OZJ2L599i8BQj0btRkfTm5p1bAGsuvV2OOWrCfvRbuPPFCsub91Nb1p
DtRUlzh8xol+PkWVukARchUicniA6+wN6PT1vbjoJtl/eTJSXjXdMe4ZUAccn+0uKTuAKefoDM3J
VBcUoqQ48rtuyaIkjnCmhfcDgPfBBYYQO0l6sMf2JGwtPkY2lbdXSZEiLPtfkmqfT23+Pmxe9t0T
GY6dgYMxl4Jxzm1Kid0tg4uTwcREvcqbID+OBrz+W8+hNxc1Cgc2JkvaQpG4xHXtFRsJiT/gAX3+
e8xaGp5iyeAyTm4Ugz6+fvq47rO/japVFYtm2xAmIFvSJFRUHcJWVEurAE1YQiK/uj+4h5cP4zrV
TUCYJsTxSAof0azD7E2vwUhuZnNd87JrNo9XZxjhrMAssL5N/wPWRrQ5lKymHqh0jCdjwp94q0wE
YYkoinlNj7OZOW4hW9yQBZslLhZCV2fLWuvjH7X4o00Q6q6e3CwrORVWbBZD2/cQC34aZaMZjevx
sS2veAb/t1+Is32Wg2zscQpcezSOVm0KpztM5JTZpHkNQzWb8NucTuoBN2ysB12KF1cc/6/G33fR
VVe8zhVfSa9T5tqGJ+sBwuOGxaLnoBkuajZYqx2BCBlwv0OZ/Jg9UC9AayOy+a4lYwKVvCUxYCO1
o7JwX94ibyrZAtesEk3vaGKe3s5BV42p+Uzo2o7u7P2z7gvgZXQqor7Yr0Yi5WP0bgMhVMS+mO4Y
+G14yVuK1Bf5hoaWGOG5NVn+pgG9BnGbdVhEu4xY4JBaK+U6bXUo/f6UfbfZa7EAOe3H+OpPmoR8
E0VWaD3wnB2b8gRwEc7kN4Y4Va9ZUkoBPlpnmFGdt3QHt4kn/MHxQGRTOD/KgSWsfjp5LQ5ibLgN
hFS1lUs7vfpYUMIPLR9r29Gm5SknvB8WuhB1br8spLzFWoOGS3zFnffe3huPuzOqDF0h6l0jyk1w
Gw7k5fTelpZXwnsEjR97RFwk0pDBVcsfQZc5WBNsKSXlX6B3uCzghiA63ddcp8ZbsvxiTn2se8hZ
UUo7bTOXGaJh8Np/vcg+sJB92SRLRV01zzOW/HqPDvIwiiit/IhxeMSwD2mhBgp1FhAJmZLmXoRf
CmyXZID/Nycgnn38pUDnnTsTwfjz6ujU8Yv/RHye6Fa9rF/Tth0kCt0WYjaOIrDC5671l1Hsc+4s
697TMhRnC/cPAUG7Sx5blOExwHUpaCfZORwXIjnOES7H05qG2SANpj6rQfLc0t3fABYB7v4r/Mo2
H5ZiDq8de0jtOTrYVqXMm0M875mwtwcn+e3LH18H670h8HAQ9EddPeP0M6e0aMIUxiZgx/o6h5FF
yDCWwHSvBYzuPEevdr3nN5Zo3ajDglrm2mDwpWV9Bphn2J2YqkkuM9STswZMy7Q53rHkZP9wetFy
mZIyGg4ZXDOk6TgRZOt6nTPOlqPXxbKuWqyoKLLzWtCF/yyBNuFZW62ALgWHCNkvoZc9QxpD1bBV
MqkV/32CJtfd4ztAqt+5L0GYlvY9Yke8cv+HU3PsIH6SFDJ3hNv/L0k40GZ+5UEexVFxtsVEsQoN
LtMjVI7nT28fKIAluElEahPpjfKEubOUBcpnfp8Orh6SnKLtcJDcXTCZkRhRx3ESmN98Nd9hu1uW
1GKIoRbPoUSsxruOdsXwAMgCuaQCw82z0d68zvkDn9fVyMgXAVSxczYY0/jGvd4R+n82JWNxG22p
wRwMHTYEG0slonhOJa4BzOFJTrZJ17wlVHP7jXO68AhUcfJEVAD/wK36uPfZ9j/z99BdXjdkPmCh
14Jv2wuV2QrVxLKLjHM3jR+hcMaPvyCGRBogevfhnKtI1fZ4vXFTkYjdHH31mYgUospXhbIfZCwZ
bliALtMHVzgxlS6kXGX3VK/rkt0oSbVMYa0aSbp2SIgDPx9kFYWiPq0d3Yr/w0u2YWzWxsmTCpRl
oIpJ/CLvUNUusczdRbneXroB64Ym1XqMpFOJCUYVxTJUVVnMs20RLNwoYtKbMOeDabJ5NRzc7Ahj
ZiARsHwOxUohpu/JjeNnCgu/kj4uMWl9DB7RfNliCdoPJtIi9MODHySbpOcu3a7QsB1hE84AVTQS
rUzhjYlN75zLtiQzwRhB7dMq7Y6SNxto+yhB+hw1oSVfGjTKebDKTN48VzR3kqeF22hmA9yiLB6h
UYtX9r/hxYijstUikgcinjF7mxRYMFpCt+OEGgQjHkteQKozFlD6S/sWw6UtC8fwOTOIZuFl4CZc
qhniAaDcTZ4nEz3xsImbbB9mst57yseUXyNIuONpXraLgLBrCZ08Uxl35keymahNVVErmKVRu06b
Vl/6ewFmc/CN2gEi1FVruVa71E1Zt7gXgBImqDu+oIcRFMBYaUu2m3hxe3sJz3qi8awQBpGe9SZZ
1wH1LdRSdMiyiWYd0GZHj4E7EbRNp3GI6xZvgf1OVT7fSygystj2c/IUCukHYEn8mdVYhmevGE8T
cEFhfJv2lLcun5n3NXUdRHwWq92earwshspbjaPzTTgX3fA3sDWUuqLfJWrYvl7CKA4QuGNeiwLp
SVHwsNWv3vjwBX0UldIf/SVguSod2mFUboxaPJU7MxW5n//YdTITDuQj2tAQ5x/wyccJAWsSPVxn
6A5NzxZt/9bCpQjsBwb80bpoCgcKc55yCPtBoVtgY+iT7MMFv4MKVnqo30FDlvpXwa1tZR29fzjI
O4VspVboBKLh+l7G60Y11Y8ggYGgI+ELnBHU1st1p32ME0bsqAt4XpV7i6cml9gWilGHYSSBiFqX
gIoV5s3lTspXWb+VRmLzP1OAcf4fK/Tlm6KAZrJLaVYgqkTp34727OwCbF1pynwTEmxH6BuRlipf
gvIfGTJgDsXMHwwCjb7cfaz9lG1R5dHzMiLyl6pEiClAuXpoxVkv3j1O4eYbPa+jvKLHuQzPvEFd
uCFwV1F3MhFmk8TIKduuR5hGJ3OKrTVZ+Z5Lv/EqmB5NG5g01z99gEC8eW8buCGpJ8tVTG1qb4dp
4i5VofbU7QoGicHwccMsRVSoHXkSw/C7l1GI8oyfuza5Fbez0QWD+FXWtb+AG1nQYPWLMOUoLHaX
m+jNZVDAM1phn5Z2a4reiUMmpy0PzyLrkpeq0dJoVbdB4DLnzC7V5VoVSq0o3Tnf5gPe/4w8Skzx
UJTAYgKIuxT85AkRQWjWdfeQT+c0z5AIAfIzP4e5uJyPtb4pL3PYL2Iq5R0Rqis0og4QDRGlf/Ua
2Jbpk7txXWQ3FgieRn5vBo7tJ0s7SEOX8jgsLwBcQyb+lXugnAwy908IlzOA9luB/FUQLnWxsKKu
CpIPNYhWZMhE0PsYDjfCJmue4UFjFbQ/RRiPDMAZFOefkocOKekELkKykF9AtDqMOJrTUUvEf73P
srvEnG6ZW36Fh/g0MnUR9lS/rVGuVOJdlMJo5Yi+TxqlAPEdTv5sfoFZwaEstJnaW31GQP6vQ4mG
D03XVCuElXdQNtYYLomsNmyofXhOWOQzs64Od0COlIIsuQm1TQGyP4ulBkoL1Y/Cwczgz3UM7QKn
pFDMUWDTV3G+iVZqoDkm/sVbF6z3nSsFirYGp89pDPOwG6L0dBOSlLNcECvvq/CqCvPpT2OJKB+t
IZrJ+ZDXAxlPGkCiV9jFoGbW3NVsOV/LRT7nAQ+0AY7f69VDllhey9A/TtqFdgd7kzBZT25CDkF+
sNIruawiEqLhlWbNMw6jBG7y3ynGQAUyiQphmB8E+vSjmFFENT62i9DUZ42CRQmGjn2Iiw7NrwZg
ALljQ3mziAVImj9KeultgF5E2cEdF3OKlZDp0TNpsnX0Xt5XS5Qe06++xZ6wl9yXC2lY215EYuKP
cHlqS3jtAAeXst+ZT9kQnmDhWB3VKxPMu1sZWfvleiygDBwcqa7rU+IIB1DAADvib3/7BguPIzEr
X0mBggYDmfLF80y9jw1XbjP8Folv7nbbeCNfFaXoP8E4MJuAqASqjQGpQhxjVqIbmcNo9q4GXprW
qqVgmaJ3f4TaiF/QIa/FUxf/36M8z5IzbyxPBRt8KZNLj8XlOR/5PCv734N6LeEf/PQpqrlGf827
VMy9s+xJ9svInOUGIX2a2ovI0UjIja/QCNYpBIG4AXYlOOqNs2+jQj7e8XjJsNrtdi7KJMxLPP3P
AckRo2Sq5A8puU2CWXXMPGsK2m3wg5R3gzDbmRSR/BHQU4Yh4eFs3XBh0LcJ38oTS6OqDowYd2Gj
2CfH985pW+9zLMQIwikIZDqOwty8CIKELw/1iPNw8cVvLTMHt8pgD9aj3bzLADMrZuzhkPTrOjpZ
zKKo/pF8qMnNbVbV/r4f5IedsQ38DQYjitkRoaZfg10r9PVapT4A5lrLwHGmAAP+ayLQt2ZhiWco
7dttgh09U7Nmf+ozD7bmaJcQOGPh6CsLhTFM0LRPtvmVwxVR1w9s1//6NREDDJow2MvI/8RhK+8Y
3dB1qyULMv/ebayL0AGbHePbcqEnYevP5d+k7H54wLFRcCHalxMdQnfsaE9pzEraxHeQYtS5CTIR
MQ0WP4C2DCJ07ycxxKE2FNSYizjsLTVR6E8jMiS8jj+eAaju90RCiGVT9j68UEHIdTVJaJJ8azLr
xJoEhAQaBfCBo+4MKsLJtLpNyDnfISmvxHQQQ3h9DSPtDMyXqymRG11U5ugFBAxGEGI7+tzIMIxp
AlRL98CGZogHw2u4CCA7EbHBP1YuYWWZVGeAPlBKhieyRd74tU9m4ATOC7oXiwQMJCrKOWHR1efn
p3GqDI3crmifttcIydeIhN2X2vCrGL3mo+Ir6bWj+1lNTKEqSSlfwJ/qmdfgaeCrUVWLTQzOwPg+
IWSKUy+5L0ZuhtDUS4B74ZRBjxeY5PyiyN1xbZudhJ7Gnljpuw7IOMT62U+cr26N4pB13HYCgQC6
ICks7DtoXS/HSYALXMGgnMXGn2JPCtAmkfBRdMQlpJMwhKbrwmhInXyh22xKOAbOcESm+5oBfaSh
itU9qGZCdk9XjB2ed6SwswwBQUKPJEr0r4MjgnXjNfkngX1BqKwlxxDOS8pooK1YCjehSkSWPu6b
6+MXzXNEgMFZmYPDuXiYYqi8J3B8lpWczEHJ81RiF/SsiXSUIQxvZH2XMDusPKqUqFAscRCDkNsX
xMkCQ0BC6g3EnwYGXVmGFJD7vLAU/E70f69v4pYh0NQ+FaR5GaMkSDwfJep6zvL1S71lycHGFY+v
feDMLC2Ql/W6K+8YHhSqy7bPFSZICOTpOjdkV9vORqTqSsLhQ9qZBiM2ZBpQLuFy6oUUdOgmDjTx
zh1KFcml3KFhTjWQkRLOLK4vp6SAsjDVtBzrkjA3ONbcdOR7BDBHKLfZXfpHlhCridlII4/9c28i
zeiwL0gj7SHg3nKqLaiG5JlhkpIn+yMa/kV8aQLd6uT/aA1SiJnhVTsjYnvx0li0W2nGAksa+adL
oauYIEDV8HvrhWp8h9IPxEgGUKnq0zX+9cL1u/+BHAzD9NKyaolPm3NEL+4cRHLYNUeMctG+pHB7
TaT0HTIILT6kPxchFvntX8r/25PTXqTfJoT9NSy3GR+3xfvXYT3qKdGkoDR53Iax1T3y2fkvlR/v
TNEg3i7WgWIkGqeCTL1jibnmE5BZLaRXar9P9nY7l1jKFnqf/IJjiDQCW6O+1g2UytdnTdAfhSCk
kFaBucRNKKev86N8C+1siNGANPMh1LPvMdJE5D2mrSQLETseBGRNYHCkiZEI9IVy638ISCirwepU
mLy5SbV88WDe+FfsfcmLrRl5dk6Sl4VYep3YNR9iNywQBp06N34FRLb1RUGnKkIreXAioE7Q+uwK
w7Kc8QEUrP5vNPYfPe3BSOmWP31g6MnHC4lLsb76Q0nG/VA6jfkU1Ahk7Kw4EyXdxn4OIudpACC4
8XK6YELybLG0C7MgtpI+0nDKKYAHiNThXUXjslqdAK5HoBi5qT4ik7z4w5CDCma7a84/UQimhspG
U5vtMS79vKrsiDudh8U/MPfLy+RRq7SDCOZ3nj4aSZeVZpXFFAFKMpidrPgUHIEgDGyYqP17HNpj
jmZtGFXAIWvA7SwT2JzuwxOxIUghQ/OffypUciZVSV2iOBdXslV+0Fw87M6o86sIB2S+aQ4xTCpO
ytReRWDLhHj1r/ZPBtSEaiW1Ui45uE2o9fyaGDZmQJf8Suk0F2NgkQT1iDdWTJM1cXLwasXN4Kao
9ra1hE+bztjM4N2uLPgmU3BP3q91/4W2WidLNls7j2wtD2hThjbiy0x49gqKuHS2XxP63+Mo6NkD
2X7AbhisWyX2L+HXHnZ8OMvgeECUZ7TNbHq+1jhpaaR7YbNcRla/c/jS3eo/QD1rPbaBvFkfS+JT
v0OqjogMCRw4HI59HJn4j82qB7XAHLH6Bef1O6higy+sktYHzinek8Gr0yJ0MZG5TScO63ZOFf2M
r5be2sa7OIZOWumHlN+1o+O9rxKo9wE3OFQRAS3EfGDuLSgECmDwdd610Ob/Clkb2bbvdd/Uw3Sa
kPmRGwrcNxbil+m9636pPfhSf2hOcXflxwnj3P+I/WUEEOKfDYHvUV9JR6F50RzyRRqGSMDU2cvJ
dwNJtG+bpsj+OUSIpRARTOTlKg3Plt37B2umv9j9ATpqnQx7RfIJ4N3cCkf9m/JFTteKFHUunTJ1
zMLctffClTW+hcYHWzo5CC+B6r5OJzSxLu5aqWgtGaOFQRZMrsw+twfkubK9gOzC6g1A7ThxcsWU
mhj/To5YQyiqPQX+c0uLXY//GR6kQvAToe1B87RR8iD9gFhwwIWeFcf3RX8pLRWGKOnnd9c4vSr5
m5xMnAsr3pxJIZqzyPp0JhEvVhZuCDSYKgSW0XJ/gKHIfVQ8dolR8Nf4PkmLEx53ABcgBjLmJPLa
GrgyV+EcuD4zc+5hQW8C1ywfostpFXKqHmbtUChiKN0kacjTOCOWjGFcJyPUIfTM+NLnEbyc5DiL
seE2+uw8zbiLiWaYvvUI+oAOwrVrMndtu0OWqwyXlnHANbUz3ZpIEbiV+1CdkmSLaRQlJwdPxu7x
/0MZp4xZpCMFI5G2j/+vbHVFzBR0AGvPNUiSDpnWQnehluqDZeFc5cOfBzaZp6ctXJgagdtLyDLG
sPJ2AEcLh+nzeqLD8jx4dwV53MpBV+96CAOK8io8AkWfLW5oUWMs0YUCJDEz6nSK9pfCxzrVN6zy
BiTVk14pZCuRrH5QEVnm3AR5IvG4xlIUAquMmGzep9SDPUfNufjqzm8PuhqJ46mDwwhoGbuPGMFN
bpYwgx7qTmNvCAAY45wAN30n4gTQq8OTnLOXzi36fZtalfs0N/TNhkiWHQp3DWB/xH7Wz9cRFgVU
SSCy6oTFq2V+uafO76Wh9ZCb8wSmLJitMtTw/Dqh5WZ7VFC6cKXLVaGBXBL/nS0zVDQCvs885Swd
zqtz27bsFTy3R+XpyT7xdcY9nhzI61TCcLzSambvoa9Cumkdrh20XivZk4JqqMC2MCKVbx5qIn2G
vvV+F1ikOvWaOUHu02UDMMX2aw9Z+Jak90sgaiwDCL/JnLCf+g5bCoxaG97XMs914UEY915RI1ke
4nZxq8VYM/p8b7CTpe04kAoVRyynTqTSRPq7vnlTqVAZISHd2xeOMTQTo6yC9/z2p7VSm5icdP7y
vkli33Ha0cwErxUNcqU3b9Ryz4lVobaVaPs1RVDedDQGkPkCFpXRA05Fs3gVxb1EWYqOq5FkOkjK
02O/PeC5jlggf1u6GGgLjClXfiia3ohX9JKm8TyKWqTf7js6Z+CqlXQCmDNoJ23DJx1DcLZZk61U
HGAOkEGhsBOEiJm9LLxiVExwPlZnPzSurHHzImu7fLS8fHl048XkwAW7i+g1dgtOh0XWGaFCV/HY
rDmxBz1OAoT+UjIaXQsbwP6fO53ndAJ/r/hT9fhkq96CNDmhdGwZY6KWpOzppxe7T0S6QSDKo3zh
KihrtG/jgP+QdPNZuKCsyQTWcEjhNF+fiMdHDtEmJG77J0ZJ10yBi3+MYjJd7fg/0LS2Y3agdPME
keU24olkWu4AbTm4mnZncvYwkQbENxnuykYWUv8M6Y4d9/tVPSJS6YP+ZiMBu9Yv5p9IUQydSUia
SkKqhzR5q2/2H9ykZuUJrcmxPyKXLiOs0N2JQ3YRDzdOnZNtdsRNHL7aHtZWbHdkTi/ROkkEys3C
IK72pKAMKY16G2hw17HghzPm3QQ/bFH+ZLJscDNuGfCnZejpFIjtbUt4mLImlCi1m9ACdZO7drkP
R3atvcdhDCPUWt/UBuLC6ToKegNBZb1VeD+BJfXplvopFoKvlf1nps9Rs/HawG01n1sSuCCpLHmf
NrPbTs2n/Uea38nLgtSfsRHcjPw5NcLhN+ZOTGr/UfBQD1TrUtGMLNBg77gNl6bbdIRtCm5LhVMa
zSpIIz1+eSbYBT+hWrYqHfnOUAHxkknYgoKNmfkzSPsz4/pS1p40GrP9XXpl+7EmYRUUn4n5hSqd
8ZpLwEYwq/pz1Cgpod8hPdbzzVwiU25mYGvLMnYcH+N3S37mC9y2KRVmAR3JxkMQ3W2laXyOsfbB
4Y1O+Be4nxAZs/Er4S0PtbMtnVnmiX5P5UC0crLgEsO3mFVDDxfZ/yHPm0XKa2MnsSDW2Prghb1G
UQ92c33DQuwkBEJQXQnITjrGCZzOh/6LNZVMkRu0Vvgeb2xImCF+J9ZBQvgJOyTPO6j0Xk/G49sQ
b9y78L9+U7yWKpM+nheHTNpXI9ZJv5BDEE7fyr528aYe+0FcXT+dTPAohBdNPF3TDiL1OE6K7ABI
XlXmHxfDz9tDifqrzhhk5hVQ0ok04IItUPmfk+aSMlWQHcxpHQDKMjNJGErcrva8y6NBeR6Vi3Cy
/vrb2Vlv+l5s0HQqyTeabZbROgrnvdEF5XFY+TXgMXfTAX/tCPJfpanksxmMPqwnQoVmWx51J1z4
qhaYIVUcX8GoFJqqcHg1POaQXPXWQugZmieHtEAeZSeZ9u06/Nay0kUmm5qb2UIN5T3Wu3J1ZzQG
1C/2O2KVAYFEIb+8tgLBzUzuNiAyFIBpSrV3q9USpCnsVQSrYv0ukoSGHvnqrOeg/LtWhPdthYoW
vlbo32O4b+aYp+kWC1iicZmArD+VzxHRmeZPRK0y5x6gsds9Q8GTacmLSwr0SkxJrXKV0psns+Fk
mtXpBA5du/CxpGJwS4kHCBUwNmOvYxZdS1sm0nQUarnTQEbp2mb5XkCyH2SvRdaCl0QstUx9KOEc
V0cT1RAKVPJR9kTLCQ0b4zXbX+dOvvxd/KbAIXQv2+zmlD16qu1U1TEks2KYaUrOKHYsrpwJx0Ir
c5+u7ruQQ596q6Wei1ZiMqXbmt3i/n8iCzmOk/Fswi11VcVMG+cGPGdOO7K/ABE2dk024CWEvEkx
RUqrpNDaBZQsPSHA3JCmZPY/XblRAnxrW+R63NNis9LY3S20au37D5s3dpE9IFnFYo8CIfhAY9UZ
wUK9r3KUVIAGDBjkUtPwJDsRUckm2tlD+jio7U7B2165rNlSlKjmF4d/Z67gCfJ4iLRRSJialaS9
wAJ78DDpl0J4OCFXMFun2eeoXKSa5tMMFszZ3z5hYWD2MGvEQ4ANT4U8KN6bixFv3BuTcZrjERsd
47h0aGQJ3X4ANfyV4xHiw8eGjWx3gtHw1Le5XQzorYeLo3cUc1dr6qHAxOOo+JsyRz7Q/8nRog6J
uk7aSCUw+Njxd2uhGXsWD0VWqekbPfosvZ0+HXkvsPQamx23UkF1dpjhxC/ZAAONeJ5nAfR2OQog
bGYpU3gzv2lCnClPiyKZWqvKsKGzG5r7Wp9GOO1E7W9TcIIpGxrBPSVf3Xj3iTrKuAMi4VrDZ0QA
GrKrJtlza60YoxPdLihs4fSFtCIVfpXhv6owzE5V3cC3Mmv+oPj4E/VP5UsBLzhm9RTn1x2zYftq
WNX+Hs6jLlCuNCuCLYL/SA17G4MvxDg3Qk1P1WzngKrh25T1ODwEjYBjdJVccHlk0pqBwiUnqNij
K4VcQj/W3Yu3PhCNEEyeKJNfbr6Dn/GBEM34GzHwaYJqjrWI2Hal41XD9pNf/ZSlvaVGjUP8cyOl
Y3tSq9sPaOfZ+IUsblyaBADoEVe7mgQKs+WUld5I6YbMtDirYQbl8h/tZZpx3XYdqaw1LTM20fzf
5XRqihjFJQjHVdTglOs6V2s16eCVpgTuUbHRiBK8t16Tr/tKQWsXmaZQTV6xYMLeNSVAhoXsW5fZ
XUbJTN9JkDu5pCoTcmyW0RBdpHXpEVz3Wg/nhvr40IZSgetF7Q9UuG1ZrAcR8HAewk6GNi9B6U1M
Jyqt+0qC8JIO18izdKtgIqoxTPWGCoiJIdcJwRuOyVPlpRnbRzNS0SxjwPDS99HaNRlffH1STTGy
M1JED3EC4eegkz8xxMVLaBZAwaHpgGT0ErKqjftLwrNZvkPhrL8GQL6Lahht7Kwt9jUbaYHduTYa
bosAeos2/eFukaSBSX/Vy04YTIArhVK7h2aysINi9cP9nEzOUTVRVf30KaWLV8XWHzDfaJvoI7Ke
s3MzJ3i10r3DOHWJzIPVjYB4hO3CzWgDkjPhJVHvUWTs//JjHCtz95HBLdMjIeGAcN9yXR/8Lwdz
giRuVe7jqi9MEZs2zw/ToAWysNqzF3Xl1yw9YEyqhEhN8B+PpKSliaUEBbtVWMoNyu0tkjVXW1Zz
X8VCDIaATVR79qv6N7MBykHMMtE+zaVNvyJXQGTHLLw6yQdt4j98NEpOCp7Y/FbeGfSVEPLWVznU
M4Yv4oq8DtEcsyHpx5FbnUKbJE3QyW0fXisZOQlbndN9OoiQvMvIZgxp+Sd+s2cCcqL9JEDrmbh5
JL42pgbl3kNfzQjwcEQ/k4W5zF5QCGbelXrlsyLSX8/xTeoXToow1G5J4BWjPOsa4QYtyOpgPjVA
VWsNk5Zrr8up8Xdk+KOw96DV3ZVuP4Rg22Ksa/Vbc6/9XZ8uWLiPVvUfjyVcKIpVTTrACP3sb7Hs
oc3SgsTdCvK40C7H0R7R/9oKCmj9JPohAPiZ+vjGMfustWXJiXrg8tNXGW65U/gNFKPpIge/6wkP
nWWDWbSrZidchAs59JGMWheJ6lTMbYdC/aqb1CwBVchOPcvz3chj+XPvcjYgOfdBOUEizk8Ja95w
/TW4OldfmmbjdBuKllP+PiSPqQZoUYnQwQjzfjomS8lv27QQF/nkKw5Gx7RVC6WLMDQeXyEDlOei
jtWo49k6qB+i3HIAli+ZjdGP9c9a2skft36G8/AORQqRyJBv4zCtAEXkwZ6Jt+m77OBSoXaPX3Hw
+quxq7MBpk9jbcrYkZN9fwtyxG9hmTUAQdzPs4jyKc1nkIPns9gV5CcmoUyL/7kQNUd8MFM3gUui
S4DRAuVKLvB8e3VUJhBmkyAZVRYkp/MuO4wvpQF8msvdgpKq128RA5TjZ9frcDFww5/3yWH5rDjf
vxbJa4Dojvj4f49s/Y02TN1tqEWJzpP1rQks9zk6A3aGEN13OqSCXlUAJeG0Qd+bx7dUaQefa/v/
1PTLKgpPPMroUNXqZjBRxx68yP+jmYJIgRu2CgVxnULkUj9vV0k+0sCQ21YUT/CWLJpviDJT/tMY
UFyutq0qfaXxy15s+5cNPLCepOkMDvmDL30m8FUbwRycNbFxq9G8d3CwC1nPRVsGn+2fpOHkPhD2
LmCRcWaY7u17W4Bb0cr428nQzsGjN14cAh8AoTNTIIPD0m6p9LAseWn5as6y0AcrTE2PY3zjI025
gnMhUd5eJZ2/h/wiR05jNiaqSsGTNDHq+sFujw/Z7Yq9B2B7a9Iiumx18ie/DOHgjLYa16y7IdTq
ppDdn4QniH5dsFTixhnL75zCRF9AC69A8EkvvXDN9jMJmljw0NKiJ08cTaPDS5sOFEkHai506Wpq
qWOjK/HdckbyJiIzEf760STzwJMNJeGucI1bD0mmKJ5SKX/PvIyGk0le81EstdxuzVUlbINNm930
+OXQ/zR3HeXQ7Snw46IbLAbBcoG8Zwrwnq6AxBflOYAaGUGYPQgcxVKTU4Y4hnK8VeLwkO6vWBfs
m81cyG0Pkj6qFVBFBOU/MJBD0G+0GyyEdiQe7R07DeHSC66WYhA84XmEb2+jTvHJhlZYfJZtrjwb
oY0DM9OPsbB9+RIayOoVdja0LvPazsQogA5E8m2eI0984Ue827jov7rWjCrxiOpkwHuiTmkvW89v
z+wkEj1HeTap1lpnyFsX/8UwjN3b65VjsMMCqH/CpQBc4wjx/JqWu+dDIU/CS5uVuFZ859iUu8VR
KsuOeyVxRHyAv1/l0Ju9zgQgH8jtm/rpsYyeyIirA5oDy5ci61Ekh7Gq3yyyaxGvIpUWT46lQ05S
KPNM7Rx0YyMnT71XVcv0V0FTuk4315ZZy6A2cAot39RxDre6sty3Z1WoVyYsbbF3kKY/1bUfljDN
/JmsEk/PwzwU8czmVePFugwSzkUQMAlBiBAApxzM+vKFK3dq2Suut3tBbqwD8ANavWsiI1uXIE7H
mZ3nuX56bi7P8fFk8btMTer32Co6ZkGoHQgi5VbxZssTeX390sqvdrYhiZbuSRQBFZr4/vGVaLnD
4+65g+wiM4JuDFweyO+gj2IRYWDx6GTf9BTXN5ZXioJmgvh8eLc2iS+LdwtK3/9yEklaw+BzUAT1
AIrTE8fpp3V6BmfRmM80P7osZeRnnpeml3jzodhQSDnvvXY/EXEto9ZuNmwauEh1B+rNR055zJxA
kEzqw+U5v0DNdJ7YeihQMdO3YZSs0+MbHkXoy31KXHoJ93I6rydYaltF8Z/k60gVivgPnSTBPURT
S0oDkRsDdq7bOfgqbj5A/n9x/WSyuUp6NaXNPyWC0fDOQR9AjtDK3gZ2bh0DeIwIlIjFYRPXiZKZ
YxjAaxTpqqNQGitDWXWi9Hw4XtieHmED8IZxw+NMYFPePA8ynWe248CLf9i1BI5Zgfq9Qav06YWM
StUQjYj/zr8QltN6oVqxrZ+22a6wo7t9QtHHHrA8ugL3Z0yZFdfvgzk9zu74h5lu4vrJIavXFGzn
kQ/P8m7hx6I19vejxzQwh0rs/cukLuUk6B8ozDtUfndrcNU4kamVUX4ZPJ6tbyYd2ksx6+9JqBY2
YDzkXN8qSzAX8VplIPE0LRVIo0+JCZN7o9LoC4xgBUw2hd0UWgqsojB/FFowm90Ry5n3CPOqefhB
TJeDkklArMoqfBSRjkcojYn0m+G10Ar4Kpsy4TPMmMgYTrr/UD3hboin8Dv85es9i4gChzuRUOcZ
zhmVUhuCJne2QAKw/rNrSjT0sxgN1x3DMRoOsXqpdn+HeXpKAOOQR51zkBiQ0kM8mvaxmFpIQGx+
mMlpL+8i5xprrSVojDBFL/VHBWXQ7xdTpw82sTbEaaAgBAydbzj/dQeyTELJWglxWdOwaJftOYdb
hM7yGm6FEzRD8xif+2aotlBawkWS3219T9TZDxAXG9ePPrk+ooVTiR1woJLcvFP+VSxcBR7rfIPc
YOO/ipW/qOJO6dn8z5krXHOdij/C+Tpce6C9YILB77zftYPa0RSCHYU2+PonJzeXdPFkf41gSO9I
JMWz3CwDeerdoK+knQBnVYQewQ8YX5DkOp5Iwfzt3X/APr1K4eLHlXm6gkKM2mDiUK1ol6zF9DyI
TRJ6TuDoPmVDPESpmGyfr+DbBu/MPs0TOZEf1mavLNTyvnaDcbLxKXz0vw18hV4h6V7QJN0dIlV/
Ha5L+EP8gHIs291FSXKEQTzsD553SsEtSYc3mCUtRNpP96RhBLocZyk6YPP/YSmxhkz0X2tBoszp
d44H5pMCIeRlIhosleYbMSp4PLgtlc4R3hWRowxfoD4IXJVNZApEpmV4retIt+A8xTY0hNJN7CCu
GNUnZqIht4L2c5YIBHPMCNFiA6pB2x5pHXdIXBdT6fDBuOUOBSDD+ak6/hohdtWOocTswhzQGLv+
umBRnzErGFA6lJansfxZkGTJGfp9NA0AQbp1srTLtawLiINuaAKEUaB/CQVOhuTO60l6xCPf6pYf
fQYvENZOEcbzH9wgdqtn3ILB+H1oaw1GBNUio5o1N9QAin4RDF3DkkDTSdMqgxcl5NbbYMRzaZqm
8fxodae2jd8pAIn4uL2kqaP3iwPvfODxWEE27vKd5dR3PXRq+14LAZughFLfzgdGjY+KEMdkPhuu
pxb07oKJI44ctZTIoVFMh/vO1LqCDkVEPMcCTFPGs0Wx43G92/6wn6QWxfklZdMPv0zG3Hqt2t33
kyUfaRtgEP/o5mzUL4JEuiqgj09/oYpzuPE1atKTOPFp9NqLFkr2AZnBzKnFbwCQmrR41vY1FKnW
3/BdseiAEavh5uFJs8LPmPmCekwLpL0Wv2vdz2TWNZysqDM0fdzOoW3C4OWigXXkPtNQefUwsCZY
AVbYOMpAB+g/2RC7pZvhEiwWIATEGU2RQcv8p6R24M50ThsfS9WaB2WbNq94B4FXmgE844syeqT9
DrKbOE0QH0bh/BajG0e3fPJooQ8S4+Nopp7NcatpcB7MsUOiOxsgWIuvMYuTtEbrGGONdfktVugl
fabRpNmA6Rzw6ZqzT28e2MErQB+JXR/2PkAfyB+tM/SCZIGMbdxtEnuYcE95BL5x+TK5pjNMPxRz
sEAn7Q7cw0B4TsHZJ/O2U43FIlItorp3tcQph1rcMi36/5KyZ/1W0X1PjHHoPiVm4UdwUGxkyOUj
rg4hkYcBDWbN7612a8iGudMI61J0ao934fEMUTXj8ji6IOKPcxMmZEmStXeR3yMy+zd7ifIS8UVu
L63bRazqySGN7dFN7L/IrsfKqHXmNW9vXG9BV5U4wiHLmaO0zzs2eArWySNAx77YHrb/erdWEt8v
N5loAZD7On4o/Wztfk4qjTZtkdS3S6q2h2qCzxiFl918HySXnEeMwTaA6yyKr1Xhg8/SMeyht5Lm
UddF9VZRm02O3pJ66tddmvQJkk4lpFxx/cQ5XWrpMirfs2DpXpqEH+gT4yegDHq/0T1/KRwKIsMq
kUrPq/pcERBshvUbJc6TnmidQ7sVuHqDCJSnhYsOVNUib2eERHJHNs7RQIhxCdUtazGu1Zg6qPQL
k0W33K64j6IxcuKkkEx13XpWEN2W0kzt7gF/wOuCX4mjrw6U2rsUrmyJmMkHk4BTj6UFBRcgd2cP
bu4wlwTWuiKoTLwpOPqhcvCX8NBhjBhZ/RnMOGKmMRmZNqT7y4cqGLrOGV81mLnszARJ8tVbKKKZ
11DqsqJ/6GyBsYz7SppLlNSZLxGll9FOLYrzLOmLd17urK767DpU4U4Uou6vdG4AhsDv4Cn2a1km
ZT9hemMHncVcrkn9CBAEZtXYfrMzijLvlOD/g8EIS8CobUVaVORlzNKTptT6U+3Qod5QFIN9UrmP
Mxgq+hf1MQ6j2SYgpApz3fOASuHet77yOclwJIxQLXsn3cwfZ4IsBniaJ6lX29RDN1diwEV/YS2c
s38/kgb8pOCqa3K/cZtwzmq9VEPfFE1AVs0hq5Lt0uYSiKS1J/ROCelPWImMijQuOJfXYZdAjwAo
WUkN3Oz0Js5GajGcSJJMPUv1+TBSviFMbP+vsOK3Gbc7ioBce+Uo31sunWywpqSg95d/pjyR6U9z
7gFly1mzPkC+SQiHvs54hS+1eY3zTTGH6NxRtu4l1mtuNW9EghwOxiA+JNOBLFGkk8BU63PhPORM
CPKQXcUAPT2EQIP4vhTiBd8nCM9JzabQwuhe6zEHz/n3cT/enckf0RUytajopSUM1A0fui4pQycn
r8VffLck803dvEvewamlNQMHNiuj2cGEL+VILsnC1qZ88zaaOLBihVoeiY0SFzdWo7tn3MQSJyMW
3rwvIQnf+fm/F5+Re/L2+KMxXOiyNpyXf2AkXfQAFsXeDKqnWPQi79FwLbYCOTE0xA6+GoyYtWIX
1NV0g19ISUBWGbUKMk/6PFw+W+ksO65blZBWO8Al13RSVu3u4HS4bfw74iT+I5kag8+rW6H+DX+z
ySV0deJLfP5iR8fIlv/f9R1ZjqolPrkWPaEgt2pftuUDHsZ2vjZodf7F49SuutJrDXlJqeMcuEAM
VNG4rSBxaAX2CALhgMKEBZcAOV/blgRLZZ9BJCPo0ib9/gkRYTJ0oexG1teVdFlTrFK8MZF+eWH0
/mGB14ugyNKFuCePW2ZB2LW0np538LVYN0TAO8x8y6RjF49drPnk2rOzgd32HkpUCrEeizzoaBLM
jTCdIKS9rsl2z+yfFHuG022sEND72Ch5KxAz3s+Q5Eib5jcU1ZiNMM9MPKmUQaL8SS/6ZT9yM20O
tovsrQz7oJZt1LOtbKnFIgxJdR45xdxKA5pxn8RrPEXjXgHxpw5RUcojzHz0Vop6ml6rbjYTngRn
9cnYXy3MWBaOWs2i0Xu1EN2WDgR+MK97Gbl22xuFKc7uYIAYZqn3pD1xVlvU2hiYXsPlBw+Xbh1t
X7vs+Awwhc+Z+pZ3nAdLurxegelZnKNPVlnLKJQLZt8Xj4RYg9xdw3JKYSZIoQl8gvQ21CefIbrR
XSSqBcl2Dc8LYivsSuq0hx9oKSUYuuzdJYTgAP+Xq6WkH068UjRzk7G+vlW1jBaPJE5G8XEN/92T
Ljw0X2x2KIFqx7BYSzwR4v6slrFHyoyWAFxr9/Lrsw56UGhMl3NOKCcVqaldHbHh0sScptjAOMbe
ZHJ7P3TvkDPg0etHejjKXfP6vFELPqNnGrMmJDVNEGXeAt6iIfEUfTGOeSRPaMX3I1t0p6Q/5H/E
JWRYOwLUo+tOyyWBSrql/rBvSezUhac9ZKarUV3hYIbmap+3CTPRF5zXm4pELilAoaWLSRWry1qH
gHs/fB/nQGbqqmxpZzynpiIExRrYW69n+0I4p0c/wLeHrxTISKpgUyoBBp/NL7Qz3vjBAewg7sxC
h6uZqQ+b0rLWFA+h7Y/SBJ05BcZsbm/94rlPYCjPAQfrVhFU/REmyfj3OMWVJRKQ4nua+6w2Dzr8
C+akjXVIkFJ8DuZtX/f9cYMwi72jydqbmamv50vNpbKJCgfTt9pPKW29/WGbd+Cy/unFcjUn2UXr
oj0pkZDFDp7HLQnJ+7XdCcXueGoDiUryYHfDN5UvqWRvvTdJASiuUCBVxt4FoacwomZ2DB4F92lc
nNhpfb4xCqpXY9ddwd8QeOFAmvUvSyMYAAgJtVUte+OpPD1O3HJZ+MA4YXV2frX7DkIvdDUw7eUL
8Qgm5RcEMs20LZDDSXDbsd6zP60zRD5azunCbdjn0fj9lGFdh145OdZiGJeae08dkqON1W52oRIT
Gkdogso2F4NSG/DzlefIV/yqMqou5rUN2N3ihx4SOlXW1IMUygHXlo+XYB7PDzR8IhOycWsLlVNL
ohqnhJWZkFth2tFmQw9V6rCJkRbizzsvH0zthYR7Or9tRJKtQIy3FUnuCB8eRaqYKaFb76YZRwQV
cKKxOWrzlSqJa9ioujmjbpeKgPp//hZkIesm78gU/YHbYgkhr0GHr15d9/L9jGinhx1p+FgZpyyM
hUCI74NokhveYX4ZaylPv4oVrrFwcRm/XptI4gd3VkWAcV84/IiXwN56SA8dZP8x5ApVxOg0a3RV
kKGEcJ6lYssEYrc1nn1cRROHX66CVHZ6HtpLLuWfw9wpitYFewplPl0MaL63ETikkyjul6rDzOg8
HDibkqJDQkM658JZtIPZf1Dj/uof+DksqD3LY3EnUwKpwuv3jNhOH9SQXi52/NizzNwi06qc8mn9
oAIj2JUyp6X81dw5WmO880FujDH2c9A9VkhpuICWfvLNcOJdv9yiRrO2az0fpNfaUtLB8jyHknGF
SUw1P7e7uR6o4slwgQNsoLoe2Rdfm6IZxJNfaALwkX45m4f2ChCtT90acuYuXPi9jlmQaBrZ+bFT
YJlAYadVNNan6qOFXSpkJ+RXMmqWgtGkML2asLTdt8ex2xEA4XMN2N3Qa1v0emnlN8M8cm6FHDCX
HDLWJNV6LX1FhObnmjjiXo2t76F/Nms/qFbO7KHCSLwPf1rYwUCYfhTCrHmM3IpkkpsUm25rsI+F
qLx540PRaIRMWeGZ8RCGUp4m36aa+0Kg49BP9n555S/kT4KbNWGjEQEtmFeRWM8IrUlhX094QTID
wNc2GbAiG/vIhkQJcj8RsOLG4jmnSwEvicVruxk3aqTtI7HGQqvb0EzNykHDtcMhR0EsX/2zornH
lFJkVl229mvU3ox6xg5TYcliD873qCrsfOGYrwbhy7qRKYneHyd37qoL3ZaZGlcSoas0+xpBBCMO
gsK5oTavHALjZ3UfB4B1bSoza5vRBxPcceS4KAzmmCy1xDbb32QYm3TVVSSOsWRBxv6P/3/GU/+T
6tIOAAvqMgEEBfwFrzcw93ZEQrti7IjODkG3NKMWOmnkTygNw3JQGHSqMBUUByPBdSaZkKodoFtq
81xMdDU5nsyjySh9FY98gOfc+qu3yeRkJUBIFsrp4lToUKe1TS5LSTzoOKdo8ze7FtKgLR1eYij9
6josgaDa7LKTtGkFqVV0GJSKqa1f/yPw1xn/hpVgzHh4zwnxwFZmxfazZIdCMUYTCXaWoaFShB07
uRgXRlcIjElC4BS7ptIrxs4eiHjDVw9Gt00iVIEbfw9uFtoAuw3qavioE9DRLxZs50wn3i9uHvGg
bcc9tDbDgur0A4B3e4GSVxFYKF30f38BXAkb2rNFsPYHsf0eeMnyACmKf8jSVbvzvkBMfA8N7hro
R36/J8jJSjEjR1SIBAupVoocEY39xpChGC8sc9vhrArFopH33WCIr13FsfNb42gnTbN9XGen5kHn
VeA3uDA4/ppHHmp05G2LQFYdqHzfbYPuEHMrTcLrP49VLmLQLlTIkZhN5mSw4e992qBO/x5bJtpa
kgI5l+NjTLL21+tbONOG/FKDzlDpNuQ/XPblC40LbVJmO/oxTD6Ztxb96WpsH+Cg97Kd0I4WSWca
c3LRziUor/m20fl8uM0bHPwzco1Vk9fmwEFjbvLNphWNvT3hHHDE+LR4N53hmqDJi+0O9wNAgnrB
lOiQLONqyjIghHH4aa9UUa7P/SXoD0jCMHOxStpGYU+jMRXC8i6zBqpAFpxVxpgCmMue4ks7ulPI
CHoCbKY3W3855tTOIhGd/N43CPX8OXjJc4XnyoDZW0sELofyrOM8VaUFqAX1BnDYxq50ayHbrmDy
aEans2pXL4Zoul5NBjiwvG1Fw5KGsdoBPshFpQWfswJrydICnUAv+wRuEjtmgd6aOJdl0h/vfE+m
DiOR07zcb05l1wBbr11XyRMEMAF3cFvfpwG7Fl67vJUXHKxf8YT30manx30Xh3VAIXHyJocSTwoD
8Nu/Ar4qotWqYK0Oy6m21BtnCRFoH+Od44c3Ly/52oRHFwe6KulV6kz1bXuLvIJI3v4q3q46i5r4
N8vSzAo//k8Km51ibXlak0OQGporIhXz03S22fdXK7m4tsHGj+OpSqITtEWjkEYSEl3zniHLFnL4
CQvg6PjIxuw4NtKvOEie3SF+hdLK9jn0l6ZlirD9byliSIZfnhL9yH0y/BIHavXN4xb/ZWZzkV4a
2hkTadOEAU9uVSMYWi4q0nU0EuBExMKPxE/V9YLhom0UZ52Qwkrh0dsRgWIky21hZ4eROjlAMUfA
LSp9hIuktdUp9IaNUZ5UhZDaijJzXK10xOjdU5d/oTMXCRTlzJgHUn/nyTdnqJlfz0MT2CmteXRe
2v5+KsbMLJMwVICaGBNTsGAUbJQijUbFH3fizSF8rhqzvo3xJ18Sbb8U+odSLzgDtL7m+V5CHjim
WVm1XDDn8YPZtH6DquIt0jaQ7tXnpzVCg5mBZLQzPS4MxcDISJZxqiDIq3oaJ3gVMb6HFk4ZIc+M
gNziAKlk1L1MaGN+7k8X1OB9TFvgHTFo+aTuKlPZuP5jfiPT5HnyprEccW3hk7EwEVPrLj8P7WWX
AlC+Wuq3ncjKJgAUVPGuVWAioFf9dwJWORlnfR5vUhTDu8XvyjmnT7cs2jyqonA380Dvg2iBqLiE
3Yzj05KY1yi7IyAkBqlkpabzAGzEK8MWr3B6pzfjdoO4dkeSotsOo3VUTqPtsOFUuNonJxkT4evE
oEx3e5AnbEgS2Fm1aAk1ql8uV6B6x9vUGHFPUDajZurpr9RwVKccF6bJ1hGLQYg8DNNKEYE4Y8y4
rOLvFhz6KLD+xC+6KEPbtmsItZDYO+OfyswWt6pSgz0YWZLUaq75LunZS8LZfOwCkqn1PANW77hj
obwpHiT4Y/l7lac5z7Vyl4ChuYm+vYeC4/Ci0wdLv8bMa+B+CTGGNHUZ+W+lBK4wCdH7JPqLTPd3
8+Qs0rKagqZ7R6lbNG4ECxUAqn7nbsO+4BxfsDw4EaEGFxO/HXQaAIJhaUUMfKuqAXDrmIHAJXhW
+FsoSqnsU7Dp4Iw1mnolARTqvvu/wAqnL5eQlfU+BXPJtGcyih0j3xXBg3/3omzvZwFmOI/zpG9x
U8BJHgbj/QsmVdUdA3MCFqCHbzdX2SLxCDMBUUz77NudBr5aN6x+Bmwahs/VVR65knTqf6gQVfDO
a1OP0BmaqrdoWZc2O0Ar8n0qvYAdfvu7hxHw/m0S95qmWuPol6RgMJ0efRyfJCXcl5mldBSeK+gb
HoJalzFd2B/IONejQqy73RD8jOBWXX4TTRkZy7butWNQERzjh5W2ODStOikwCunWbNjPywvIPpKh
ZZAkvLW6rkBgECMjlDDJDJZEaiHCK62LZlPRqsZHnJSrEl7bL8mliaeQgyq1izbaN1+aIQ1Y69Sg
IIdQWZfwb/qgDBajQtuu92QTKTE5+0N1ZtckctPSxFdG6bJFTMAE/G1C+ylTMufzXvBsyvJsY6N/
+kWjSEblzP3z9w19z8k4+sXfP3a8AskRSw6S01J0gIWKkd2mCpIwHyR3kowHtldKarK92afT+dIF
zHOzJ8VYQp49CoFJ19O5sIROoIp4t0c6MlGDNdEgZYpJhh7I7v88QA6olE6BnpokGW87k7l11/Xb
qyx0hsWwhPf3TJbkKHinHaN3m+i1XomzX5pZ6dgonuxhS2BZWILSQlW0YxqOpV6OQ79iqbMk1YCP
ZiBZsHcDafvJr34wqnTYAwGWymODnL7Paxh7bP1qMM7z6SBujOGhqslO/6QVOYTYsN/C0eRqlyn6
DYHc0P7SuDiYLhaPwrZgoo5vQ/BDJJEoWF8NGjGXIiIlV0L5VFAAPNntQyHkkCLouXC17FIRHYJ5
r4PJ2mV/XY64HUQaTiWQezuaGCH3mwTCaIghecXErYYBRPpf4fiTSlruhyWez1apU41R/SxCR4CK
qOSMnJ4fzih3po+DAi0ZwgfQYYAtrwKR0rKTFkCf7XepT/+8+dQGcBEOaEXTkjTacN0v9j0CGwD0
n3rS7BF71z63L7JIKRXE3c2HfQt8WYeMn0P1IOe/wH5a6VoZBcwktUbGpJQjOwqvUIi7W521E+9j
pKhroEslDVOF/mJ29gjuCaNrUnfz7JD7AaB0AdBoXcI+GI7zbeJD2D3fUnjzvgTJMPfHdz1cBZvZ
PVO/6HfQLPxHR7vKgXEGuKoiEBElUvsjLNVEmZmi34OCVhu+PoCh9XYkw6KzBNc5aD48mxnN3KtB
gY81QiHaavINs/wFcfBJoYwvbQTo/zD/6GcYZZKM+gU3My61VulzBuu6PTZKzmTTritkqc2aPAFQ
htfirIwHVYb0LVWfqQzrFo9BYciPG5RMGWNh/2kiDeiDiXiWc0joIaIXYpn6oH51u+k7PC0lIlXy
pjUCCkvWehDm8sMBcVmOaYWdhhPeztkQ6j7AAbYfcnL+fzGeX5hEgIInPdEaeaoWF6GDlYL1LHKE
qgdXbV39Sx7jFcb09o4dKU6kGmaJeictsHr1qlw/oZMZ6tYqAl9tglfu2Pxwu1W+ys7UqW60xQwg
zeo+ReW0Py2ixxTz9Z1b2wX9r/M7JXvobLwlyq7QjfQNWjmHaffwflLWcyYn2qdTi+OI53bV1McT
P59cA3K593l+qBVOZsI1l836qhIBS0Ongc1gmQgC6HsqeTu3IijOSPhG04JSyw/Tvi2lxybuyZ4+
M23AsNMpZRl5FqDdy1D1q2KD4mVRyUT3qf+H06p0y/YEevB6oUKVoAfhFO6/sZnDy0DJSc85Q+B/
sA+2jjP2pLi8R1wL5zUn8Im01ZV7oM7/jZafMqLViq1oHc0jJcAOxVMDWmvYDvn8S7apsZBlG8HG
hNGcGCUTh7BuYhkDy3SKtjbPKUy9aYRTEJH4d9j090PyVBmVcez30WbPXunMTjVDiGJUZLfugXK/
bkz4bCqdu2tYuh8YBa7vZKa6p1sqLhMTCFUhDAm2t5HWuVT10v+h3Esbq3MpnkRYbVmAXiC9rqJM
wlAxr5Xy/oo14Q3iSvFjcMfgJ362Gs8oKDj/v8trvWP3VpeZfm3x7w/PKmLAxSBomrcTNt/ga7OQ
lG38Uzx1EwwOxLEbjc00qF6L7/zZyvlCZUWBpbDrr54KplvRgTEz5CbH+0DlfRtn0BRa6K4AStf4
TIGGNWBHvG61NBdJzIwG1QoYBjQsu5kvfOV7/YxcZYMFGpqOa9zulFAOADYKDeP2jY2M+uSPiQer
6ryXGZsM/v9ZZUjii/XMuXSRkNZv4m5E4tcUnmePOR8hJcsev0CnarI6lGgRx2pnHOheJb9+6d8K
rU1X84hvxRjrPkV7dn9t54Kx8qyV08vTZ6LiKdKp99vvqBU8UfkPUSAHCacr5A7JqeLRXAFr6pKz
u+6XL+7raSjNoqPmaTnsLdevUhLLhiXyhgHCv1CghXnhPzoPTllwTrhyj5h5aX27W05WpWQZDH64
Yx6ttD660c3xD6YmR7pzRlhS5oSclvnL0BvwpreZq1luqn8F1E685IVEBUvgknwLzOXcW7fG/aRP
oVufV7NKrY369oajeX7CKzXG9UN0vDtRsr3upyegd9g5sxqQ+PfBosYZlnpv29DzsplxtGCeXgV9
JtvOk6dHEDpplMIwVQMfEXxJOimLKhwSRzx8agbr/Lbt0b+7PKBFMPKqrtxqXjhlY/5i149IUqTv
3sXTMsMwqBT2BXMEc3esIYdp8JC2tEvATCPAdU15IW1SeEXBMm3bFPBwHFY0SfQSf4dYGUUCjfwF
WrwnVsvgXlTcvQ6cYjWXzi4aecCN3fFNeWiU5D6gu7NPBshFZcXeIB13FqAV6js/mxVYXCso+g8n
Q4Rx2J0jH74uk+yc/VcZ9XtUgYOubMQQR3mzV2SYtiZ1SNOmMzbVNY6pSmE1H/lLhrRr1RxQJ4Sx
Lc9Pn/3hINm9QDABUa8j0PJlAR8Vt4zzexl4UY3Aqlcgxdv7jYE3F6MRyR7U/g4CKb8xF7N+YQeY
QQHgOzI2k/3psS4ysdSaIZ01dlXNmBC8SgOWHb5oqUahVdsrWfEqSzLQeErrjlLlNF8RfN9FGFKN
BxD+6/p8by4zvD6J0+iFTZ6nH2Z0zJ9np663+tAr8bYz5FrKqskydthvmO5d4VqUOByrzwmkGV3M
y4wGllr10Ieim3FDkiw+v5hmI8LN6AZVWgixZwf433pGzWWN7/tDN7F89yFYm3WOfx3b6WxptS/q
AGwqLw9qic8EgBZkmfJFIAKoSN3KG/D3QO0FHc14YiVk7lppQtXxgQk/wthwqgRG33fNjYpF8Zsr
dit4Ywj9UQPlJ1e7Y7o2a92sxDpZHose60+GVEgZuxnh6hT/XsIx5ekvnsDx2GazKf7RrzH8/JCR
WLihB0wgUnHFX14ng9CuSbJK8aKvGRyarv5QbMzR8xAKEQCrUijmUIUV1oOS9bKkS5pHGP3XnGTo
1dwLaZt4N1l5m4BrGj85Vf8ngLeznWQV8+7Q4ToF3ry7G8Dj/C+QR+KK7PjPXh3b4PxcHTjXDfSc
G9OoSnk/p84+FLu1wlyNYl9va7OqE0JP/cC5EgRCg2ieBIjzrgqwQ7bT7THYM/wOXcUfX4OmFlmZ
pqeYfwxaS4NaRXY3C9+LlyEYnVynBnIhaMb62oRlInfPtLMVy7EPQNu71227p+Q+bfWRg+TTcY/h
4cwXIftR8PtqWwecVdfpZywooM0zs+6OLtWko0ZtSQys6SH7FUhSrGL7srF7GwJi9TPp2w/GBgAZ
C0r9S1cydNLHbd4YytzPMu3AWpNzdbCELPmBfEQ2zCh1g90A9oq5PXHOmh1kQSqSu5e9a3K7+yHR
2rT/MP7C9onSnWeETy6SKYd+5MEO5+gGIs0yQkolFE0AbOuUyguQ7sLb1fjvfEBvqqTk6KICb8Aa
4sunCVJaaTTx6V2vuiXS/4TMY9KRBvs1NumDGMopnI3or18IJTwDI97bpAe0GvyLo9dtp53zrEsA
TiElSUFh6PvWUiRVjc7dLJ1Uiori4UnQIp/1xZf0as/i33fHC2A+g2t9km3RYBVMpedvv55402He
cNsc+/KrWF3njpAiwmhLDuwPKB5KD1ytfGGzfsQA4e4Zfps/AgKF0Di/hMekaasxrztI47Svye0v
Kng918fKnNntw4PmwFAdYqM3dU0NaiNFcT6q7r4UXjE7IRrGED08QHOmPPP0rnkKs9ZyadHIehA3
UV+kjJSQZotdi81/H2449ceVBqyVVjLQ4HPZDfFtlCAxsjLywJtDes+v6uKyGIu7Yo90SVoRmZkY
QXr/m36EwIyHasqVr/1qWEvwxelqUBblDjxjX076rhWogW3SJZkToq1ImnYJBYcF5A3oHMo7DjdK
FubhdeDV34FdM8pS/nWzvSDEBUS5jREJb5kZXs+pZpOvc82z7/f2xDFRF6H7R/4Z85d38ML8c5MJ
S5Iz78ACGwE8gZnlCbpfZUXTRMRIyv3OOmdk0pl9/jyKrlOBCHMu+xyN3krq/eFm2yxYJm3/RvBT
puUsqj9smE7f9U23AMuLlkZZIwFHbUajwNTrODNiimB7giJTi8kVQL30if9p6X3xCcUZD2/6GBRl
JPB0Auofael1HnqDj0fQ+bGBWzf3JFkdrgUsr3eGlrKYFGxypXu2jgmmP9Rh69/2Psow9l8JWNC4
r91Nwn5czHwtSkMrImOXKGKv1UgVpGRicuew+1gWudcy8FOgkOKkYJ00Ec5nsjd7fKdl5A7u2617
3XG3LdJOV0RTgOFVYkKTxP8xd/RqALmXHRLV18ir2NFM3w8Ah4aRcQox6pABPxsV6n9CHlj7Y37A
QEx9N3sKLGfPwaJvOZpgxbL64PyxPUAe5QcpLrWvDIusVEkToQwx14P3AdA6/FaPJrqWnNvkYDkm
sS+HZzdLc+UEpZ/Akno14W/a9K3LRP9xiBybOYfyhv7pHdpMvPcpocq1O9KaZYYjOWu02KRihTxY
W6pf1DgJQTQkiTkvG5/ANRshbR/DqyBOabd5yB6sPNTu4bUkjplnlQEJV9SZGeunAqb6FbEhtSk9
m5UdEGUOkRsd3RqizuFifrJfEg9aRYmBNBCCBiAg6IRROIRGvmlHWyoPP64rgAOwf4UkdoZhbqDM
RqV1XpgsAfu+TC+dbEcsEn7953Oho8D7jF8Pp7LtoFDTfQ4bjCUmXYFFV7hF8qGsapbKuTH8e5Az
NYgYj+wltYXv402w0PagOFpuf2MJNjV7yQ708L0XBs7Ozz5+AjApE5Ppd8F+9RC9ykUcqQT6grwY
ELios97bhcCeWRZJin5JZj29WxWynYuwr66icPtfVZo3UDwNr9Y5RPbo/ZzvkFayEeO50KbOpNpL
4af6aDkyJCL/9p9D6vpWxUrtjdUbdEUvG1+8eQlKGIf8toa9Vf8gy2Q1t6GhHSJqfER/vMzQMyMw
un40Z7zI5f6eW6k5vXvvI3ileWKfNIGulrLVxaRo4CJcREbBGgaDbD51P11aaJZgru5HK3eW/4Iq
frLdo31qxbyKu7hZsiTNB2Bgxhh37Rdh8t0Oc9qpU+w5SW9SURqMfqSzHzAWwDXm6XbzlZs9y8HD
ws3uaReSuiWtGgUTunlNTvoVAMvlTTUPwxgyTAkWUdsQmnJHuEo2Ms71FMkDYgXx1UXOEGo6wxKx
xldIIWi4a2xVwCiOr0bTK31R/UKDCjtLbuPkBFlnuriGz50K1U0IlEOVR84xFQqRL7G2Gxfd2sN2
hDnLs32Mw2iiS4warJj2SD0UkpCAkBIIa8et1IHR5sOaFTEBBDHyuMluyQJUbFgKzMaVeVjq72Od
BzhKZls1EkrHTUEl26OjOEZl/sKwg6ehttCf0zfWfOJzZNNjm4+Iv8rxEnJK9sPrfCTeqTzVz/u5
yPIFY0yU97KeWUS97LClmx/pmKo9LJDRj6ZTPdmOKV5k4PxZyaO0Rw26aZEGNZoU5POglphIV/1q
qE40vuv5AhHyDjhRxcxLMdwRXCWYLJCRaSjoZizNNpxVdTCZMa2O/PSEJEgaJOBS3Q4XRC0hts3I
JLhsx/BrPXDXfoPoVcTsPmKK0EU9Zcb7vQB0CK+dggV2cUqCqDB2lIEmOGhedhVJCYWwQFdyuqkO
KtVSyXqbhJVisSCKkG7c1nv6tj/vfmCBmthUADvk1cZmnIYG5sasDi9FkJdt4jJevnvLYJMIo6ub
W2KgSv0UEm6d/FKpkxCwSoHPvnvPmpKfqQ04Mj5koyaYUTY3z8N5GlU6WyqOSRZ6oo7CJ6LtNWBc
5nL7YbUW0pSHRw6Z+5ifK5qQjnM7RGgZrhwG3rnaLKh6LdixJQgCFFryWPIL8RogxIGTK9cTWEXE
Jwr6sqObWWVqD9oKN4p9tFxaw9mw12DdntPEwgD2IitXg/ZD9gco5Nm8Yyk3LVrmsRnMQKVUgfmk
4tRXIgZ/Rj5Dqo7ajYLQh3RQ/5c3qBiUP1X0NQkM8qXv1aNj0gnGIP/Ln8Ou5oTxRdkGiRzmc2Mm
dlnZ0r4rKx6iWQlbaGLZSj/LXpKfCEjejxLf3izFV828DchVZm8P1YOrbkjrudGv1fY2yI75Tw0V
Pxwb6IkgAnBPw+uOzbbKoHvPjJDdHl/Ir/PCy/kf7fDZNdxDZ/LJ7G8k+aSYI8n8ur0vXuvASGY/
z1cPGxU+nC1Wk8BWmiwGB1wj6+R122rg3w3LU3T7Z4mHNGljhtClbSdgP/WnAm9RSgPJ+Yy4f8L4
cNKSXhKrAEEYtPKuLbSsyaI/sVObO5JGuXJg2CSjV9N7pr0WzGSpVH58u5DvrrhWvEr0mxvc0/gX
qxxCAtAUk4kbEJi8QF6nXSc72zmV5QS1EBcQTKN6ovIZwcGsCGID+jehIB2wgxebV8wmfAT/uItT
CpXSfT8WI1B1dxR30qB/n2PJaiCtQ5hXOURqPCO4XWVism/Hp4XxoFcpBBW/y+2+/4tzXe2ImktZ
iXndedIu/EeyxvSPaO9Ut44npMm1LAvB5nFlhAOooVA66FKUhrw3WjxXzNToKA82KEbrVJtYdpCD
gA1rCTTqQZyIRp8PRwLiVe5sK89kFisUGt6ALLgzlPD+SHLWOrOQCY0AXgv8d2IEXfpif5PoOj1o
ht7PwesKVL49blwsUC+PkcrQRv/QZ+7DLtP1bw1exmx4zlqC9z+sUmfpRpUDHMXARtpteaFBvdil
RCB9AGJF0EfEhgDgK725cJ2X/iAEiHbXcuxqEVFjMDRqiPIDfrx2kMCbcQF5WKKVSo2Zd71fV60G
xL1b5sXghCrjGVUcHjVSfnDwiTInm86TjTeL5lZK+OP72MLThDaIjvLD1DXtkVcSNYh8uHV3zpbd
nKwAQBIyTwfU5/9ItNnin9TP+oqb/p25yr3J29LBZ0pZUNbjjj6wHje7fcWPLt5mdthJnNqkvBXL
c+FQADXvoCsMfCeJTEqlh5OG0VNbPZj9izk3Lx3P16+s3flhrn5PyFV1b5eZngdqvWUxc0wCAQ09
HMJahdsPLndhGg3iBTrkW8xC/Xj5ZzaWDA51woZbEhQkHBXk/HLNDmU36giYTmO347V2UKg9D5Ri
u1+nUR6QZYZmHo57B2AREuernP32rJ//SYkTi7XIMlLmktj3GYu+wftEtYxLsXtzewhDT1brn4Dl
+9QedGKU+yKup0E7mScltNBJ/H19g69v9A9hBLhGNRe7w7zwZh2j0szuMG51oHDOpaCZM4un2sgJ
Jt+LcVpEqSQEf8wdAxbzfFqgnz01HbkUEygpHpW26JPsYlV3x1kyIBj7kwEk8rrb0dQEj5sG4wsC
mbapYrvjXW6g+Do6uRSEo0lf8dAef+wR8hj4a/4jxREOU2XXG0GXOUwDsHNeclq0+8cHj+z0P5jJ
+8iSNHvSh9cGE2mF5TW09PyOwXUvmhb9clLm0l+YKByakMVhiCkkQeLisx1rtTM0Tt9Wq6YvGfiZ
nCjpnzP9gwBEUpCfDnS7kHaAiQB0HCTCa6BsTR/ZPrHxOlclJ34RE9IqzoJFM/3UbjREn4jzO2vo
JlFmBH8+7QuPhOgb4kNV7YjhzMEknuM1I9p64fCQyseH2LA9l8YWuZy7v6ynoBH+GZMKNlGd6kHS
NLXWHFMCwbYQm3YopeQnO4VDLZcCEXVy2KWvhK01avCgsIcwxxGFfiGwfcjMzW3l7vBpc87cTB6+
W+he5WEJKlE+bRLxgE63D80T/6mv9Sn4kY+Q1BmzgkeUpd7OkW/73A+i0LVXKVK+DdXhO6YtK3wt
30KK+RzunUIGZu9gFPA1zfq/lX2t+wUrHW/DJ9oPvmXsKbh+WkyZJe+3gnx4oWm+8ITEGejkjINE
3myYzp45L2eKmd6rneF/r0IiF1mb6bAW9cpdUsoo/AM5TH/YDMvnzLeBFiPP6agYux0Pxp+YtA/q
57kFGUzr/XiVaafwfXrnPsGt5qz7pRq68FETaMPS4sjEe9v/zs266jZfWv6lIpUIxu1zshYzayHi
sc6SraKnF/s8kLXRdTtFIVik0Ez82dPirBgA9iyXxHVvfQumw31HFuJ128c02AzHbXUwTgWsW9XR
usaVR/5M0Qj+7VMyzm5vk95fbMBfXDVVmDcDvhYh7e0IEz9pUN7Za8BjoAVdFbs+gHsHIqmfQWOK
uMCau4rtd1LSF+l2oXVhMffCemNJo4ijTDkIpTD+RA4Ek0hRryGc1wELwvcSZP33tw4y8fee25Q4
A+5u8e6D0nFOkI4Q3CPe9iLPwJNN5vbE44EPTUV7znoQ1jaEXDU+2RTUuz/RXmiwgN+m7SokjxwJ
6vuOE93AFnr26Xngm8oEwG+W4sbkWwDBQui9YFpf4XlGrU8D7NmEBE848Mj0q4Q1TrYAnxwmKK6f
9h3oRrUy22hdmNOcRGxXgedjNa/C5cjGEPFMeT8qK6OFXAqV+BXt4qbhK0Wj0dTWoodozo/4ikaj
5uFSc8ivjgzLfgAY/UA4hpTJoiQfCkcfZ93o5DV1Ww3edydj5HyXMK/hl68X+QNI93Zz2xVSncrE
S7PsA/VrnwZR114gDIuN4mYJvivjmLeQdLAh86tZCQ0abmT2fNG9VzBHFaPj6s84Co2KP7evCoSv
igLrxgxVhBc+2lqJFUXPqGzyqnBnVhf8u0p7iWN3OuG9ktaTVaeET5XWpB4atgZEdx6H3EcWKo3z
4UDMgOM5d15EkcVUNwxxWCrFTb+fg0YZbx5nSMUcyk+rMX2rrykHfMQj874KhJzshZ7yLsh7+t5p
tj7crcOL1mmbLsJlVQfWwAuMwsPxMU/Q8NP+Ck6mE6o6+VEuKbvRWwLbZ2eJPRmzXQ/NXyXMo+HX
FtsmaGgOssF3VE07T+JC193hQagzUrMllyM6DYQ00yV5X7SHmRvN7WXQPzRgWC4SwRbI59S3pVMF
elUkKbbqP8JBsG2NLKh2C0qlmS3iLtMgQQQnmkLE+UNaDFTZKYj3yLneZDDTJ3lfJlJ+pkViJ3fW
2TZwMd8bvTLttsENOvjPD++XcwSuc5rZbBrKs9LWCXmoMqp6pI69bUmb0EQr06FILfqyzd8fDV2x
4U9fUByToSDUKNyEHmV9SYgIPDZy6zaV0Z+jeIBSw1hXyu2bQXpa4u1Ai39Aig0tDVDm9q8fHxYA
HB1EdXUqzUlQEcKJr7hVlhe72lbGYCv/bxBGRy7ExDK5X8zxxc4Cc6hLHin3nTmTyMJJyTcDUb/W
dNPggjEXErn2/CGbVXnw6VIxYsalm906SSIhMLzilvSfbqX4Ll9dqbWxgf/dlYy6SOjTpVupvQw0
8W1AKEovKOyqLuMPsG1l7LrgtX92Zd1xN+J8acQRHRxWj3VQEt5SWi1HmqPCjgR763r8GWnFlCMS
6cxDM4775sQxrjMC/L7t8uzjQ9melHl0qkWY+mZzRWNZk+bP7Ytw5yr1uQdE1x1oQlzTU3D3BfNw
gprwXgiC4blKRTV7CIxfdTKa03Y7sFll0zGfWeTg2A8YzyDEa0kZmVeo98Uc5yLCmsXubI61t0Aa
yIxQZg2HL7cZXbJwr5w9N6ChrUfDzOhOVeIMbJn6bLBS+ZoW259X0Dr33rHu0+aM3mTWg6FoQDFn
nmjtZOu8Wd94g/FVhhiruNYWp4OS+EwI7SZxoWpvjvhi5dEQVd1TmQZTivfGmztb4B37qIuPiq7f
JMQoD3lts+JaDpB6j3jWKmhi9JqH6OH004wPL36vN/2w5xH45d14etQinthHDpvqJiAsdgb9OqDO
bHOaT+ZHoE5W2kY08wqIMX8Vssixxn2fnLqIup6LkGo4JlhglGQKm2mOQOstkNj55lTnbgxufokh
niYzi0V6AqleR6r+Te8b7sIqgQTahvPwBDnmoLMOoQxfKeVxOMr6CaJgCdVrhi2Y3Bo0ukzSeoBa
jG0nqRh7jP8/LPLeP2pIiOhRny6x9z3RM1JNiQON/7JfVAXsiqRCEb/PPLNmBGGg+pIsu5pAFXKn
dA3Os1vLP3tAKO1GejTuGr+34pPFbD1mEGxvdh2bSTrXwfMY9+rXzm96SCYKc4laC+kAJCXfPSYQ
PApT0RXMJI0JYZsg4eC+dyjl6GdgyYZIfuKwC+X4Xcsz2eW8X+erCYwaSt4dLUyJslqfNGbXnzVx
d73sUWm8hvfYF/ocVpVr/k1lzbeLapEnr1phBYYr293SSRqd4W99ic4COWRrz3EBrbkHx++HCnoZ
UOTw377sZh8xiEDMJefJpZFZFPVkt2ZsEkIKBbqU904jpxHr0LRDPVSADSE1aTuV2WrYHPveZlLk
1xmIkkF7HsZ1pIVJZwhGxYZud97Q5bCglABMQtjM0xLpq2kFEhKarkaiucbbJU0c6ztMtDLUB+iJ
GBpII1JRdaNw5ptwo+EcczPFWPS7MhsgtmjJR6JPpmP4nQMMOFHV6cqHKy15rVLGI+gkHHklLJy7
hkVWNqcnDrGErXjfxNPyYJwvpG/SwUsrZrI/oJSWZfitFrxNzZcD7ElxxFjtCU7tjjwLUYHs6hrX
tJXD5TQI0fxNwgbEPqzPrAIx3lxF/4Y/+IdBR2MyK2bEMlbv9EFjj2kuJrgxZCp86C8IDFjUOdMs
MKoddGJHfxJpCli/y6us9fZi6nPD7g63aqdMxbLMwyXvMZwnWcdnPh++mPSRsSb7O0jeZOm3YOWC
09Uug1IYba+4R6GNyGdtjniKVJBANT88PYhWSlXgCRnhheOHGXHaUM0ZH5L94rm4MjZnX4YDp+Tp
coK2irm6GrplGpz7xkRG4RuVMSYHpCscUlQejmiIwqaRZrkU6iBDRPKtE4tLy1m6GJhzH6vx1Fuf
gPppI7Ib7RBAlICU8U8Nfuq2DAT3NWTZ1QvNMG0Nr+BQBhXPLGOdmBnee3iBxp7N6oq/jmDtOlD6
BF+fk65mM7Ufpm+halnoVhCGUTCovLr6y3qB6j4QFBZ3kD9mfFlE0Wp69dMfgSAPs1EJENwi2riQ
sBskvqTaB1fu7aQjB51PUd2wNOH4dWaw4GjiM7FwB9L1Ma8tKpztQfSYU+GNh3l3QVI3EI2LFi8f
ovBJNHKi0Rk+M/uv5dzD6U5WtVMKAplDZy1WcIjXbwfQdSA9mtp0Bt6IFqFX9O7nHPYOO5ffJ6Lx
7JEJH05sxzJxg6tnmom0+xxwBfyblWxAEGOQzK9BnsXvSFmiTkpmO+RdoKSME+rJbPv+jjOGq5Ni
vaTUa/D1j6Vpo/9QhUVKY98mZScK8hZ51RznR+eWcroU3VHqFvw/X+GD1Ap/7bBT3sY3HZryLnIm
/SB1bDuF3DdnYDRmqTZ7Q92zj1VYUoXy1cu4yNX4GxcveB4n6awuROWxy/hZnGMxUwf/iRUUEUqR
8zpSJU+g+jFOR9jLkHqjk9WU1bdGTO+BleLiuR0+LJVtyY4Y8HvZDUaIwAp1XH3iZ9DI7oA4nxCa
l7ujVtCkc/ba6SP/rIv2Fz2UyyyR0niv0y3tYPC+iWK/31abghRjXTD5gt4Uzw88UExmS8KuOLcI
ZjtmmY6YdXxIhTekd6uSCLuDQNNllIUwT0PLXj3iDGQx4HaLU+fu1BnN9FUqx2Wg9suItbmf82Xj
UHaYNVFzYQQXigPXcfRjEAQyrpH0FaCKM4m0irTVR4WuPun1M7QZfKiqK7kIt6dQtzMfOnMgmYJa
zqi5iw8EgOTnIx2tx+VxSIBjXmDVLfdK69mmx4Nm0qpvvoKSjd3nRPj6ofvybvwkDaIvuqX0GuI7
2sJQqfPGfMWWoonQve6IOmDV6jkQcJJnx2NPC4J1aeXZBqa8I8/LDaOt2QFpKSmMU8/FM9Dzrz/B
wFPBDvaiyeH7rHQmgKw5wWryuo4IFfwA773BkddAVaRvEzXNGyI2c0CyxaJIb1EjnY1XkNutedIj
qDUuVrObNAHcmbWBbdhWVb2TWlf/K+u7yeTG/1Qs0tfHm8baLXNvr3v/Nvbo/Hyb11+KyOw29p73
gNaQT/1hT8rpTJEJ42u2PCpMd0go/kaNVKl3+1PWu/6B3z82SaRYyZQEBP/jnRfadvEHn3F4bxlB
WllLCRrSPu9K4UzjBlweZj43xOsyWShcP0GYwj3dKtIR4LQD2eBlVZHaeuFyWJL36AkRkHA5xVJX
MyTza2RE2vMD4NHca/vZ0j+xbc2nQRrCc+7btrKQbiOhlk6RyPkX/tkLZ9PYgcXfsbOF97VMdoix
xWX8F56W8nD1DTjJ6o8GMOB6KJLniufkE6MZ7ozwQweCUVLRgme9Fklzd9bKCqn+qnvJy+N2o0HT
5uf4+h00dEwFJexBLeN6DPjirXWJxy74BvAxNspNUwTnW5NyCYCpxbfL3Pgw8lEWqtf702jgBOJK
dU4StvA8xDsSchOh1xhh6/arAt+Q4JU1cIEywFKyQrcLgBvDNWVJAP56SNyXFaqEg+RZHPa2+twR
peC3PQrHE+m7vq9FwnBUmVbx8QHJGCM+s8L9VMo4jzt5GVS6X6TIPX4quvnps0di1LY3Q0QRaM1u
WWSE7ay13efOlrdzTIfvj0D+J140xZa77qiupQ2WbGyskpkXQUlgowSxNKcE4qLnYAfnCbeZPhTC
asQ1jZ0H3o5pJGnvD7niHx3eIXAYylcuiXbN/uSerfbGKH7MqiMq0Xm/YkovP/FlXMAFsYpF/7f0
zes1RIwAnJv5Aiwf4dNPYWP5taK0O5ERjcOaAgUhbtVyHPPXyPzIkhth/SzV6qRJVLB0Ev7pxiUX
0+6nQZPfqYI/tLdUfvQX+48KdtEjIH3K4k2Z9YrkesUZDFejTc18wnsaisKfKaTEVJlB4uVfOZ36
qhi+RAEGaPiFc1wWYAzz9YZzEyCbVgaU8bnEoWPyFwtA9bVBXQ7oka19vj+P4eh3Mx0gRLqN69cV
HXuGhbMxQ3zdAjO7bqbqsp2Hm5avFEiGLqGI0S6+yuFeM2B8OEffC9MPTxCt/lr9uEEXNJ46nB7w
FQDaVb45iljh+6U/EZ7uTH3AvV0H/kPXUFWjokzTjcZsYnQSlbP4Xba1iLOLDsidq1Kp4IacHgla
4jg6/EhIVyWlDuL+idHAva4YvzmZ/V0clWhw9IpS1Zl4BEl/a+Sb0PJrEurEz8bUfJhqVZHrb4zw
ECdOnjkRq1UBGFsSmPQwDvlBOgyH4+PPtULtrGjY/9qS74Pe0Z2X02wrN+r/TyNq5h8Sp8bBL36D
0C/fObCEvcusO+Msb9W3cS8jAT/ZnDCr27Ftd/6Elu1+sGH1nAlSbr+EFyjDGZNcytM7cGxEX9y6
Z2HUrOQc3tiMn8T+XnIyZQCipPVGZvWcBFrx1WPJH4zlUwex2JCHQ6FfFYMbbwk/3b038QIMoz0Q
p9fgbRItjZ+9rzajEYHZ8Ldw4QwSwjNgOlzIy3C4nmOnF+nM2RLH4x+ZIy4zzrmo8StAyAcBzBYs
yHdpmos4VFTuqx/FU+4+Ap5L4+RF5yg3lSSVhQhiaPdqKhiT/wH4hb9BENfXMKmwkdsmso5Q4jOF
vniU1IC3udlbTpYaTp3piCgL02qypSAXyPZXvDKEf17Q1dtfVNNzLLxR3rg0wjZPHriHd/2E2pl3
v6jXD0cU3alcD1QCvcvSgeQ1SiZpNQgXwbs44LlHBpfDbQUVoIGXpjmNuLGJZU1RXtY+D2Ok8xqu
Ar1leADzuJlh5CetiXzucunu1A6a7b62sf61bKUyoGZEwdcmyMw7HA85UtvSCSNKglQyMulEexx0
MpPw6rRqlfqzmbCOKpUXuV0lInn8zGgXVOukcExTBzIRCy2aiw/Oym4LvXqaUoMHl2cirNI3YME5
zchGAmnBDiShraZJ7YBtlITPuNH4NLHRdA/UkD540tZnCKxQQnFy3g+0LYYAf78WYLr+63Qzgfr3
7jbay1hI1gpvZdQh/jvFwUV8egGTd7xtp+bH+78QIq4T1EZwYrh05x/5jIQLfIJDgSpr8RbG8zm6
8hON+mUiUyiXyXH7hCxLOOp/jqIAe0j3n9005DKsT5N7ncKbT4Mf49XsWZ1LHEwwoZZXVBwrfmoh
5OiCO5Ys2xmYrjLJCNED4zjW2EwEPdhiTpQyGCqmiskrKzxqkBYFAtjtTKiIoXDln9KN50stVC3U
RwJI8Ds+UyTZRXidgUbArH57mdCO7r4367SOvDpz1SfK6NuWgDcrzd14hs1qUhlGCqe17VcOXuhj
oTDvy+1+w3H4qPL3dZdY33T/whdSO9igsVLo1g0tZBHF2Alg0+OFnCBmOj9bYHdn+PGvv9K5u2Xw
8oKt/ZvB96ODdhYyOn5xAVbc5xJte17e7uWRDa3Nffuej+AYQ7q5Wh3YtsqNBdFW0G/w7nUB/Iwv
k/iALZWTiYgeAMK+nlG+tmVNuJtfKeoxUtQjGSrHkaY+FpkaET34jkEJ1BecuKMeEjcRXDtKQNwL
ySmwjEJLwNTyWCbaJXOzRIpgFCsaUX8ackKlHyZGv48QZ+9Dbwe6le/9IM6f+M2fO/R2GvbkHhuS
ffYdwyf9qacVPDRs0ppDag7KbjYSDAJy+/Hqa1YznhYiqVBv+ai/EKrNW16Dj2ZdtGquPTOV8b1Y
BfvhaPdbJ+bA1dnRh7gKG99xDfxuKc/hiB9vBdeLNUKkqVPByyHFW94M4Og30vyapp+jYseedviy
WMHLXLif5+pZ30B+sNWPGcpcVqIta3rWm9JXVqJVW9oEPX1Ss8B0LwNpYV2XIIOc3J6gRoYt1nKC
CUHXuzFqKyhVpF2fJZS+7dS2ANIqzLb1oKFeBCQjlchfLZYUmtqIEBnTRI0OjbrLdM9AeMxvyJUP
dNaaDnGagM68UIZ1Uv4VafUrYLpyHSSCVYLAdVj/IznomMm0p4Am0uTz+mbblia5G4Cr1fMyCPbY
Wd7NXH37dS/zBC3DYAS5xVItx/1tQf7yyqdkZhtMvcDJQcJCxXk+aKmJicXQJF/OqUEWUTgUBZ3o
D2kpSvhvXw6CnAg2qxvxab0cIrNXHnZDRxiuUhKHePfh6R/qoP7CAZkW1qEBN0fZEmuIoDRm4pNT
xDXK/VvfuSp9aTmru73Fhc6gz4yJVD40QUuC4yM40j6N7Jw1VrxGarCdM9dVG4kNQ3f7tT3+VenN
KkgymECn5FnhqGY71z9l4b/dchRUJfjXqKsCokX7T6/St4dROpcW/1EaQKiVzpM/R6pg9u9WpIhg
3iSZ9OyoGzw6bNR2SUYtIP8C2e6W/fZ6xa23BNL0ajxmlOhEoPIjUu44vJuGDP1NRG0HTWH3MASP
ER4+5X/sn7BpTrUKVSCzcG3Kp/C0nvDEEFkI7jzbj1CTn1HXFwb5BYh3cnTiEc0PdU5k7f2rx70n
/CGH4BFbVgKQs9WJvr7wsoWQDwFikbVEoqNc8VCBo8VrU3FVlKrcJzM7ohNuAiXItYocc93F7/BO
ueszi/ZmRA+UXo/vO4PuKYzte8Qx5QVMGrzJxzAF1Opb7ndZLuwpQcDtHTW1M7UX1EN2lb1Z7LS9
jxRfdWA3bdNGd4gM7UunISIVh1iXAuKVYcFIaGE8oAn0g554OK/tSQsIApE80FwdVwyE8EhgSgk2
ofXwvOx5IDA4QhjxFU8iklnMTTfQE0A7WxyGQa+QCOzW5/VdEQQjM4aECmCz3peIbdU98aoYDoMw
FpaGpusWYw/tZg/I21mJP24eZr1F0qwgSTTq6LIbwunPtutVH2C3Oam4dYMF8LORCEJ2XdJeozDD
rip+01/ygnPDWyFhbn8j8tLebLpenW7uRj6DX7MiQuDkBEb7dF7Bv76FUZw0XBXj8C4BEWgtNrrp
fBC/LVVeSgT03RgFzayJbhPmh00mEun8ENmdWYFGfwXtGubpaKPvNnvMcnAchrug0FH4IkMJznro
lIb+4fmuzsEWcxEjgsjfRtLngz/F+EV3YNMzGvsi1hjOrGVABZPSeNOs/dOKPzxheOt3iRVdwzym
LY4K3eMQupvH5fGV3nYP0Q5d9pgbVwnnRAk32apnVNm+93NFXgr37fT3HXcTgWd9USY3pKPxW+uF
LG3zDh1oU01JU9wNPRubp6SrUc3n+eLe7JaUXd/KRjtyayl4vU+7Zy//OcsCf3cju78xg7T9Ic4T
uLWBXALtDegD/tMLwblcU3SfbCWQTQBgCaEZtHGIXW/sOQMb8ACB8xK2GahfShm7nrXYBeopDuYK
g3dvAOJ5ey0kvKBjTGVepb1HPTxqPpl93T9bUrQpx5VqS7tN0AZv36FjdIDvY+MnBMExJhHnum2q
Ll2OBWP1NMR2h6O1vVWxdjPtcyIVcciyofyPXfSX56IWKpl6mPKdYFj2xCwKd7VSG0T0oxUCSinH
nUP1Gwv1L87Myyb61IryZt/56Z/Z/mxN/mLa0tqRNeuSd5oN3tWA+5/kpgr1vuwpgd37vboNDID7
n5qBKwi6bYlZyp7hLYA4qn7kjDN+28Ke81IA5iSv7UuXuLr/ThNv9PUFG+/YNlv5w4N69ZDMjybX
KfvHS55LsyMnkXsNHzU+PSJOOH8E7zHD0NJPtpS4Zl2JlOtDN8av7VfmYDuneU3MPoMRzp3w6v92
8ZVKVD1/vxXBaQfqyc1Dy65nuhOzHC59DsW4MFr1CVE/uL331bmqd2UTBKVXRqBDZHCb50YYHAcn
7I6luOsLSpJC6twYgweQH4v63MTCahvBu26sfnTbP3/Aa6dSaC5gto/7LwEGhXMjz/X2dIdHanp1
5w9KDDw25h92+21ScD/SDhomGFlfFzXo49Nso6wTaJIa+TxYcjLryGhFx8GdUK2vyoveCF5tV9lu
owtjO5z/S2vEMGINjEK26gGLSYk/jbaxmujgpS8DjCqYYC77q0hmdZcPDt9Q4Z6NGEM/9MKl/lua
tjEPoBTBPJtt4i/AFZo6ekBfpI/31rMrni4dkII1nes8Z3+MfgBRLCe73fVgTjFe2bLjNZP4BtQ1
C0CbkgZsCiKGAr0z5wpbuhgMohZ6Wpt8SVHRcKUHrE/uruR7C73CeUJ54XOLoj6PeHbZJdMthm/U
B056I2oASgzN0xfZoSnJz95+ID6AXHZWA+ld1PCiAAwhx00pKvGaBsYebJqhllKxibv9Hhh9YgZe
26koFdf4R6k2OsNY5bfGdxG+9vaOj++ZIUaU+5aB3OupCTKofzZkf9/2e1p/QP0PPs570qh1VjFV
Rkhh0HQ1y9/Tpzp4T0H6MvWMDrGJOZqKT4FT/W5bJ8pzfSRA/TTX4/FJAvGFl1Cn9XvnXMRDnU2W
ZPcyY7Qi5rxi7EPw/HYUN+/fOtIm132zfBiGNQUfmrxu/Cu11z0xUzolfQ5bAKjSsTsRamH7rEfM
Kqq3xGInA70OE2irpq1jiEtoNS+RJvDcq6WSJxVlXqSDhTHCzO/7Ndw4RVEioIGUw8T+Zmx7Re+O
NmdvKTaNov/uxW/xghn2BBXoQkBpp21vLa+W0jGzVDZgopO67g9XzliV9vWm8Y63bICn8zR+zl2E
N7qMmxzx1xUA5r0UKkavbKPG7ZRX9tlG9yLlDD6qV57ficE18z3Kz27kEEbhvJ5BLfgaJ2as4vr2
JbL59aWsWMf4oZRfsgstWlQg8Viyfwi0nUcdlQkVsOdYa5pTzJ/0ILW103Ko3aAjuHzSCtouk5oo
p7OPXgGPLGOKQSMlUKET285wZ7uzzJYk/8LBMlTgb4IVZalcFikta0S0MDrzaNPPC6uOUn6Bud0A
GzO8Ir1/XlbiJF1fxEzEii1W50gLgO1Ae1FyNUInXrr8oEro1y0HuN+hYQ/xa0vGRqZxUZAlVDIS
d5xHGfDQ3UffyVwHDskpX9KDZSfnQCiysd+1S6zDciOfAzs9YVAQnE0unQDxGJkyG8/ABEj9Lazm
+7Xx7E+z69/NuH2fJYXP09IvhjCYKxby05KYZmfxI/Y3FW03WbfRoo6t4eeDwjIBIM3wnqdTtlBr
l3JERmcHr7VDFDe+GiXAOju5DBxYgfBr5g7qRb61IfGpZT7N7+wKpEqiHoqknlB6XG85FfsE/PkY
XMLIJ0KoBFJzPmdEoF5/mC+GQYbuFvL9TzrUFb1LbZ8lCE8/ucVBTQ/zuHfhJuXEVNc8OGHGuc3l
JotofAnkGlyur4fFMqqbljWKaz3tYdydEfMIVPf5FwP7uRJL2uDDQy+rRCbyGD4jESK+GzlgYpOv
wopr6lS/FPKO/tSv4zYRCytIiFe5xr8BcOWUJZvG248QhNm97SNLfc2DfxKDTnhg2NPm6hSgACfM
OZ3H3VhpTqlW6V+z00+JE8BcLQdRN6ZsScjY5fR4nmfaeCAShJJ5uz6mGz0RcA7UqYjYvNkiiDFw
T6a6JKaD2yQ47cO8RkCLRT/B/w76QlNsA8HUv13IXx8wcX15FDQOein3tyR0XScvcel4inzUolXY
YA3zzW80NljwI56USM1V6KDXFXfty7nHoQY2C1NNE/M5Xlf3TeOiTTTQBNxBtHvE9ll2R62Eocg4
BcZt79/OXCDLp+uVpXPa/HQts8rU49Dth1QZGLztJ55cxFJopWSfIl7lPxCVpz/jGpzliwC//9EH
uIA7jMim0hbU0rqMjKWIg7sSyOjRckA2awGcTeqDfwyuhqZzKxZyCKe6DcXNVR2nO14XD5rn9oBb
8iIgxH2Kp/R8W3h5vozMVTsKpcLx/427HX55ytPP9Vb3A8JXnzORe7oZ526Nx1ngfPsmblOQPn8v
PnLmuDdSnuaLtiZ2GbPahPAuCEAhmhDERHgarMJpYVsotSvGEMPyyt6wxZn2KzFmDvMFd2wE354o
YvB4Zn4oLdwrY2ZSv3zyn4Ho6pXBqCJDrpqE+czo4Me2NLXBwRlJGsgt9giLgkoDJqc6atNNjxuE
QJm3V4+Wlf6Afzcfr7TrTtNPEChU6y1xgScE0/y2JLgBdHE6g6XC+CciExe2UPHY9IaIfnorbTAh
GSQufr8CB002r4W2isDdv/4XT2O119yxXZYWnp6AdDnR+o92oahUsiMhAuc6odoNvKrnE6x79vh3
vHckviaYUy87qzUR0FKsialq/HR4Wcr1b922LVzaYrMcDMA6WxVlE/croIHKZ09b3RNmV2eeV40T
ZvSV46CQHNj/L6C+D/a1XrBgYDC5A54VF0CQ13l01Xq7i+24IeZbUl3hbowzDPK9gy/e0C5lsbDs
VtHZFwuUmWNeyaamOUFn2ZTy5+SBYh/r5sQDHiqK8HMkZEvB+MuA1o163fVhH1Z91dfyAQhyaIm5
CgbP2RYg8YpTwNgyGUgrATEoKva+ryQ4aVXev6HAn2wimZsxzRJp4RteDVqnoORldLdiVol7OE/F
Tv3c7ZMhlo7QLdGpvqwXGk/pHVtMkYdzKiA/M8Z00fxr42nf2EToH9lDM94qIx82Alkqq0f+EJ/F
sh7jXDbq1Dd+y+SQO6pLoqOZr9QUNOzlSDlhJIQFfRscL6MrzgazOO04vhKbBJzUrVCyVcS956i8
AwXFSrRlqzlu1QkaYAu0WKcu5rL/iHH8QviIb3JE4pG9ymck5h5U6xDy/qgieNyVxVIcOAlBh6XB
7aULhhG7nugLapCT7j5u3j6JFFQZvmu3xep8KHibS9sreggcQgCFk2N3c5OfKOe1YJPNvSavIIGu
E5LID+lIpKWG5tdud6Wrquf7PkHAn9t4VMeTyHsB4N7TZG7RJXFCPBXrh1VuGHlhKhs6kPk5XeTj
Mlix/XPQNYTVi8QVOr5J9l5wlVGJ/3uB7fPEGGrFRRwzNoCvnAFezm4JXTSzXiTyPJw/lFsCAEI3
H1Xw5FavGGobcxszVpnJsp6EnfthaUtEIzuAvMtXVcT0wukzJYl7/E213IhvKtQSU0AyesTbL1eW
3cog8k0tGM1P+LkNESFG+/sBp651j3NKTaJYfp4ke1j8HTUwnNLysoJnfqh/iMBJgt89vlwl4rJQ
E736gHEWKCXWpEPlUAGho/KXztkvwLmNlfr7YdLJghHBa63O+k2fXOl8Ngn5gr9Gd7VF35DgAmXz
1/BZv5/U6e3CT/cpXA9jNbJ+pj1tm7hRBYEAmqIT0uSRCGZHvhD6ZdnZOg+gkcouoZsO1jk2WQnI
okjwftQ1BlHKBudFMIIvnznqZsEiL5ibBmpWaJCywpdOTFhmuQfq0PEPm6XbL9KsKa1qk02qxGam
PLhl8tdIFHetRrHYp8XmQwTaIQlL792CtpOS0d7iW/ZujGdENlaiOuJmVYIAH7+0aLXdgluxxio0
Igv1L92HuG1cKrjM3E6VdPBj/hIuv7B8UZ5I+h9wqCTY26qjTQZFjl2QICZdnbGsjfWRLF0Ge7RN
2i1DZXgjC/fneCTuuliUTyqHw8YArijOgmrRey6KWGLjRmb3DjxjPIHjj4M1VPvzOkUih9qC4h3g
PGIrTeFraExc5yJveR0bVrYQ4z+RWwa7GeAf5WwG3AGWNbNVCphCDIA47H2r6/uNonnEg5zklkJ0
w9asRQCxchthh1kQHP4HcJaKbiIxzgkuFgyjEHlacF8o2fE5F+3jwOWVTL/fY5Mh4CE1X0MsBKmt
clXtwfpq/QVP86+VLgq6XNjRk20qF9D2V4wYdnDKpG8aFBC6Sjc9thUeMwM+71fcvdnhaLv2c6wK
TqHBjy69I8V/GA3OXawwM8f1i+g9peFRIKTMzjnPWczJt2+ZGPAWzuUVqZLpd8zR3T1U65eCp8GI
p1mEHMHvinaYmX+HN0dxz3H2qUiX3IuRa3/bjztss4XKp1qoNddmDJLM9Or29RQ3zQi64XdWdQ5i
nvEtXXCZbH9Nzj593ORm/zVX/3nxUMXkvXnWVvfvHtuRq7XgQZUOXHW6s7znG1yYtaN+7lW3s41P
74kZm/pOEplb6o2Kk3a0Jb0BSEga13Uc8LwAusedPqD5bIMYggT9+2rUZLUxW72GAqF6Diy2ypj2
YIPmp0UymZSB9vpw4t7ORCczLZIF7soplhGKnkpGabkDxRvEqEaUuAasHPAO9A2IDaF4O7HULyrP
j7svr/ZZg50eoCoFE13WTKJHGznRlbUQvg31un7+ikoy3D6hF6oArK8WNdfFeuxCA1aLl+WWKbJi
ebKkWu0eGEcdbwrptZtxoiGZYBlZHS8CKRtqlY8EF9fbJh5kh8HEI6km16WpfROUFB/2TAVDN/WX
V/bmYCUhfpbNzXAwBkqFn7RFWQ8GCpCdxxrI9MZN3ubTO4Z0Tklbck9DQ5VofeA/k/kuFt5gPEX8
ZWwyYusD/sdbg5FhineUV0sC3sKbCxe9tq+ZP+PCRZR8OZsEZOCUCyB7qhWHpWdY1TjutGhZDdKw
R2CSOUxTAPB1PMYEX5Mtp9UbyASeC8U2wtfrrha9kHQb6Fpd8jrUmju7IbRUKphu277eUPou9J4/
wnQxE5zwFPGSahtVFD97Yc38hr52SPYz5ayNmbptPvFfNhQ0tvoyYfC9h7lz6YLE18w8QjeAcBXN
W0NstJ2b1T6kuY2z2EhWZZYQ9mqbWuXJ8aSsICgBKyzNNo0NT2ZxeQ2uzxzAZUU1NouY+tYPc68z
Km+S4ihx0wpi4WgV/4xa8vq7G889YPHtKvI5D0LvUxZN9YD97iLz0S3utCUmG0Cu5rHLb2l/TSr4
VrW0BfTGkGFudJOD+IGXpOLG/F6K1cuOIc6XMd/OfgqTyJVd3yeJQQ03SSjZgcNNbYcMm1fG2/Ep
ai1r61jQHsTrdBCodAsUvqg1lt1Xntw3xPrcmFPI1hsnz8JeXRlQ1zJuUA7IYk4EtE5gV/DtDiiy
AXRbJ6q7+AJz/CbqoKlo7fNqqDuytqZ7TigLfvXQumIhspTvD4YduQSyXmImsSePIH8afcqW3m5j
9ZBnUa6YRnemzObqQJC4SHzxDL1NsuWvqGVeBNy6daD1gePou+TAi8jAnirYfKB/pfideKIeKmdB
yPw4mGqfsBIyXikbM6slvPBi+tWuUrql6h8kYPc/V/B3DQ4h6FjpP32Xq7Ta5CLaCTXROq3foz2L
zZNjwdFfbKhaneLtDTnOK9u5KZhCznjwFgXEMNXF3WyqDU4bcJeOORXe/zPi0Q3EtaDqsVApWQbi
W0U7o2W1drJSE45s2YgA0croCgvMGoKyrZypJguAMVi615R+rdalOnz6XtCOkSTOTUfrZa5Pg23X
WQoKvbZfljqCbbyxHw0NTNrfw/kMEdo2N5ti4cR70XmCJmuMHG6jIcwRA2OzE0ZRJzvBzooyrexJ
Tl3AP8WgCcukMHKgEx9nq/wHRYXdznfkX8lYjlJnv62Ov5FvNFpgN6OnuztxW2fO7tMmaqu9Di1j
TLs0LxIM/Vm19xacxnYjTgZPNzNvMLjHZ7WjxuV/JwOGexgeBUre0tWZEMdI1FR7Fp0J6iQwRSnw
96aHSUUXK+xh5qIgMHjlrQ8I7DIvhLTUYsT2j7/2/iJu+nNHxAOdm84Zae0DcnXYQxV709x84ark
jHRqroWGLPhV2pCnMCAx4/tt/Ciz33+iwB4uMsVTQDiBsBDGiLtSJox1MSrewkkEvXtqcE7T6Aa3
qSt50OfJAOJPPyalk5dvQ5Y5+7X1w81VsMmes1fexacOq+Jl2fICBZ1Kmlu+nABdGcY2ywIo6kSi
JzV7CIxa1nteRiVSgRVFegICdM8ARxNqRRt939FwdUVoaIA0Lknv9nxQ0QndFvk/16Rc5bJo6jXM
mjQuWnnAIpudJlyzU3AR3RtSKASMqDHFP77seVSwEXdfTlWalVjFDheudkh57QDrAjqM4WyndO/b
U3reyA4bSW1hz7pluCKnGXNdL1eO122bPprDaPFGze4vTLIig7VfQMOUM40trc+EBZwHE2ZS7h2s
4+2DW52f5GrXCZggMbGEkhN1+0vZ5QuNeLQ2/do5ycFcDrs7QcSQnAjLwRj4WrQfRtjl+TUiZ0/T
NC8tjKQbf74XStRzaaejrobxAO6mOKubhnd8EWmSuVTcO1uMHWGCymXlfKZrSeE9eLlg+vi/dWrq
uRoW4Xn6mYMUnClusTq4z2egelXImJ6oeel3o7S60p9IWS5vElyQwiQlABADnq9vAxy4MsDRi+P6
pYxCxvZ5+vSS+q/OyNOeUwaxNxj890NQeYdpWZvlyl3tRCZzLma99GY5KfMG0Y0n6zyDu1wAT8nR
9CdOsLtrLciK33qTp5CX5xFtkHCtLvY7gCS5RlkdoVdQPDVAWl4jc/IRVYjvoWQn2qnyrs7spZpq
C9klt02K+W2G9NkRRx97OD0RAdL5Sd0E+FM1H+WU7H5GI0lzy2/cAPgB8i6kgbXuka/H8xiz1X0/
/IGgflE/i1/+NEMcoLXnqC0bKRIjRWF0iTk3loS+CrA44tbkNPTQ+7ouyr6A+FpYzKQfID/IHNTz
o+W42A929EjGwFdC72YTNlyh3DRMXefm8x6lpAtrgveEfOmi3vfB79/GtjTd7qqyr24trJDfD/UN
80Po6BD3T25o1JVKbvSARaey3RL9YaPNnIASUlbVXF5ppOeIVUChDuYP586CH+vZ6Y1wsDkn4Ioj
aNBX/yoqDztRfg02WFhw0L3INocqvCJ2iD5LFYxWhZKpLRsbTSXGXGhRc9mnSMq90nqW6zzIv2Ga
SnD/rANbjABJL9dnFnw7rYdw5bPEFz5fIlBfI7fzZQ9sFBc9tsVHt6vq0G3cm8fA8joQuQ5RDbnp
wH3nLNmwEq0WOP6bfvn7Ewe4/gW9tLEf3Hp/34ynKdtpkOjplr/xpfz6H4Q2Q0Uzd42BjTzpdw/6
OMiK/laGXkdkc1p8cxljMxpXbAnCcrPLYb31HiOrCQRIhadQ/9tmhJyIK3Mby5Sl4BCPpuJe854R
xr12ooipcc5g7hecF/jHh1wEuDfJ4QDN9bWTKT1juz29/bOFG7qI03bb6pHEX+n6qlQ2khwW8U/K
Z2dvOm4Ux9LP9vcO4xuVHFCODdptanGkIl7NFGHo8Z5Zw7E0aCdampKpAnRdqZSYfvzjeNTOIxKC
Lx0BGh0nvNqy+l4AxEWNdvt2RbGZkT++k0q4YPME/NtCEXLk15u7u1tZN8FpBECjJUZn9y2nLuwR
7zQklHW3PqADt0pbjC6bvzsKlx7dsg7zDFWpca5dLCH5Qx+wMuxR4ZoCy9fczuEz33QM1rxgvVPD
5yipd5UspB3NLJA8O7weMI/2rHWK0kQH6v+3oXolZaWR9OTpHxBxPL1kAnN+YSd6IN1Wtemld0eI
gnY0yrd9H0m0X5ScTDeNSMcz9/TvQtCZXy3A2jXsWM6R/uh5G+K2dzZz0Ux7XNhdnS5NBh8uMngc
gJgXsl9LdYDI7W0EgTbli9KmVFay0vgZaIKGWLbh2a8zxR3tmtGY3w33FAmdlB43E64w5tCI3wqf
Lf5+my8oeRWQjg11rPEIL6KMsgvE9B+/pZOeu5hdYCTtuubabWUdcTxw+lRjuLSSqesq4NRWQ3YA
CRSjM1AcI4zlwG2Kx+891Pn+TWt8dG0TZqLr49cCMfyGHy3LUJmS7EX/4bL9TzklmewoKZ0/vcbE
/AGKAaKLn/pyO6UbwLiQ4G/pXNJ57DhhUW3rkZzM6/V6rtutwCeWk57x+HtpezemxrCxnS1YK9T4
0DKJh6tT6e6ycLoDF5OtW2BDJQhTyRVs4ycqqEkMbHAKCarBNostO1/J31Q6VSaFha72O74vtGF4
Fb7C0BoC7WMoXFobsgjfhrsJna+XuufXuX5/gK4YBg4CorvE1EGU+Iw7U9dCVJ1gfmXJMdT78yKE
w3c2i9LjpRH9jKCTVod0KgHMnRPbMaPHhtEiegJhx51uzGS0mE7rPfZxBvDVIMTKTCsBYqnxSL2J
4o1c6Vdm2/NmLVB7odf+z3cag4D4V2X5Kv4hl5fgC8HsSrcEFsGj+GQHQf3iFTlK4ITWsNs3qogO
rCEbikYN230ZLoZkZA94DDKLk4IgYqgyYRiU73ZFR3236Fl8rE2O6xHNrdt8isd6Y6mDXbVA4ahT
mJav/XxEgFljt8Wjaky/jhVJl4k/4IAb5wlE2QhMrlY20qVtllNm6cuxUzUhUzFlV5FxZnGr6OM3
jXyp0YSa1MaUx7VHekJBOXbXv/14aXA51qY/jKOqxOc4BbxzFC3GGXu3tK1KF1E6d8jLSj66V/tv
wPkMMwb6gZIHocBWyOR4gCKk4zKarLYS9EGZehV2aFdkmh4CxRAiptzbOMsdXYC2GQideG9HU1yP
9guBF3Fsx2VPEVwXLqLO/rDvQwlNYb5dX2AnrS5tByhK5+OM10vQxa096vc3zTKZ4ayNeEqCZHti
n+MgaKrw36X9cPvQei+T4PQ9dKYgrT7xB0GyqNOKJeHvNvHYucEIS/9YsA0oHrPq9g9o5Egp5IDT
voyoQ4/y5RkizspcEVd0uXPp4yApVG23H6zTB9bDWEKaga7LkOanfK4HNajo2R4TXaQfbhUKNTdT
vZJjJ8t1I3QiL2/jeEDLJMqMqPnOw0BAIFA32j01Mb2xpn0LGvl7kjJfLYwvVOxPQOp0QttsNf38
uB2w2h1jHgDFApaFnn7yknQReO5IQ6ycsRFDElPE3ozax0Iodss6kO6KRpdrK68veKmRqblFIIRj
ZXTN3YnmwQPOSySRc/TnFJIw6sfZG6IShSmiOx1cFDa60dSl2307cz2lqgo8WLqGoLcAsR9iOoop
xHXu6qUiSXnGMWFtwmzs2MPiswLXkGqmJs8UpftPXcadkaKon/EXY+8D6LNQb6D18tOrWgJjHDwq
daBNcCjtylGydB30l/cBbjosyqAr/OYnWY/5ajbnNOGvwR41Hu9TrriaUyNlHCj2Ee5TJSDhJz59
xDSruCmNR9Ii6PRNK7WvxlQG68McQGStoZNCbvYx28WV7cdt9qdEfLEXqxlsyPYn0vWODbPOmoB0
JRk3s5YqCdB8wQhy1l111vH76eWvKTMQXb3vDG8CmLnoICp7EEroU7KUMt6zhNhsl9uIHkWcE8eM
WudnOz5XGq3wv2DstMPm6z4BBoMvEfXoXBeF32ghBvBpIi81DKvNYapB4oqD2WzPoXUltwlkHkNv
ToW8GIKSYxigHBL1C/1iTAOa/URPYKYLYgne2sNIs+5YYWbam1Y5RjowLja/x3i6upjRN3ThZQE7
G6h1RTiCz/Jy6p3EkawVcOAds9krWSa3cpQFvsIC9s1QlWJHOKZJS3zUKHmBdlGgzUxRy3Y6Nqpe
smQg3K1kS6SB6SkH2/ifH9vLtB7Din+LiT8AZ1ugiy8OT+Ncmla4H1NUpNC5vUar1eJBYKoP/dyu
93p0MVEOJyKT0a0Yy5iNg2AwsUaW+ZfFIIilZQ75VSjz+9ZBUjkfxrqLUZ9wrOwncaC3xpy2Zw56
b5U1MkERjYee+ulF1MuGmGtQOgZoNQMEe6SJAgYxSmhJirR0xAihdrVkfBwL5vG1/nbwvtjI91AS
LMtut1xo8m1FjsM1ZkukkF6QwG+F5aRwGL/QmcH9ciYrQ+ZZ9WaWad7/6CuTlZlj832o4hOE0iMh
FhyF5pVVjDo/Hq2pgMEUgADFkcWFSa5N7Vu43Su3zIHz7j8Ot1kP2XSGIOz5ygApNDee/JMUPrGL
T3vfugvnrm3iT5kN8m8NVaWja39QieWFl5g7G7C2sRpa+wXnRBHWeqU/rXnq6c0w3eWg5/uZvrdd
XEtYsvZgFAaw9rIkSjGcjgaaZj88/Y6VwKjRooH6XatOZujYOTsu/EyHdfYIg2JQqQAXpnvTQlYG
yt63V/rGwnl+11xb7WR0LFvnkELEN8ZQetV4b8QBIYJ0qwp76mb72oF+w4BHkefpEzmd2hrPE/IX
1Xh+8fg19/PSI9VnWuMdMjk9RqOvofKZ2AN4OenimpebGP85FzIHe69k0XoQOY3VJBdNS1RRcT1Q
bbDiujNHy35OEhXXRavr4MC0jTA+VGU8W2ztKZqCRPUkFeRvK7ZhXC2Rrv4DLzU5Oifa8IqEI1dP
sCaT9jRrBdFTn1SI1VtlnFB9cNv2Z95JiwTWgiS+FFfufubqN2Jzo+IS12BD3gpHvxiy1D1gVoBp
tg5Za5lFcJgztJFSvarNuUCZv8QSVldD7GMU2JMktp5epca6avRCAArQqWJWn/eRJfYzhPfhUGoE
el37+0oelU1eSyvDL15QNRQmbHYuhPcVUA35fn89Lg4esCuAgRZ5bV8+jJ4VwThlJIxhaarOHP9P
8nLcvMrg+pgajPJLeedigxETGXbKhPP/uIjEW0xFMyZ9iIqj03yZOpVS7JBKkql1gezjJbqZTZMm
rF0ZwbNfOxPhYIXBMGVEWVq0tp38i98qF2gj6J3w+7g4EBlWHVeD1nDKxw6yHrUG/59WjDF02eLm
uhnpoJxY2p6+DpIUBcxD4xm9k1bvQtcL1dcwRFGn6c/3UrciAhlVqT/Afl4JCHL9HKYwuI6+oPig
2/7d+O3UEYgvqafMv7VO733rdExUXNTFFFsd/CaF4m4l/m5F1aJJAwO8Rouql1OT/DlRKFMcu3So
mu9tYZy9/do0pkbI4lA+UHI76MQ7K0PbeJBCvVbVUT1KdSzt1i5IHdexEiaZyGZr0DdLoxPpMgf/
G1/ImI2hpwcXO60QA36nd4ordojRj4/r1zGzb8r/VD4R0W8qlwA/pdvIW6othfrArCjaUR/L1+07
b2iJFA5bgHU1Z38jEbf3YMbdnpV72PfIPp7aq3eGm+LXOXR1OHcdwsaKnt4uegPZos9XAYRvqUgP
mVr3C/1yd0Va3eBbpr3p4f1+5nIdYPwcWfb7DR8cInmDqWbZ0WHu5q7/1C6gdWPyvvGyWHNK/CCr
ivZkOToOW2GhmYiktexRjLxI2ZUMPl0HdmOwRpbKXdv1eT2Xrbrtca948sbZlacgTlxCyQpH96Hw
Csn0RUTQkUuKQkRwUBdpi1pDscgx65dh1qWhx1c2KLEIIcE5UX4Z6s09E+B3kKYD46S5b+Pd/4Vh
NeIAswvwX7JbBXvOYUm3Yn2IOm3ogtGHg2bxwSGOaHCMjBxuqz3U9rNgC9pElKFbTMAd0Plt/QIk
j4ev+1orXG34IIJuR7VI7VgEmrezCsLhyl6TqNCLMOEdviME4pm5dLc+L4j1CdKuZtcHsgetIVhw
iYWWd09mIDMwNwfIeoWlxviiFVE2M0PSsq06G+CE8UaBqZiSKbWwTzJHzhmU9Plzum9/+EBTFsKl
6Us3KguWBQjp6X+LCDP7NmdtOKIBi228uoubWK7EQfeJFajcuDzcBepRjaCEONcky07+ePg/qb/B
94yZIM/6Bpjb4F40BQp6FsVsbLjunZHa+CISlpNZ76GLUgckcOB5mNefud7lRiK99SCtv4VyNZ1e
ecGEYAXospEP9sIpLyMz3eSSZhuk1scRfVd7vSJgUpMBz0cuOCdMZxRTshQeUFiVPbTFS5ERngvw
5yQcyuEgsCU+RBNu+kRF52HbQ0+gw37ZZ+fGse4uvky/sKIsSmPONkiUDiMReoHeW6p/FIMUdXRQ
pGslQuMBeXjpitR/dEf0Zy4vP5IS7xlhZEy2GziMzjEHXLTMyxIdlAramdLY3C19bzE+gNwIds6l
bSlsm5JF42pthc8oELvUlRajv7yY69mMaXpv8StXM2rEuw7ptp0RPiA2Sa5JlRIrsTAQTN7E8OYa
rmL1LVLD2jNCw+3re2WlvbH/bqAURwqmaCC/jgdFGKsPNWGBfA6ZWYUmfG0hMou52tQdUcUz3nBi
LQQyjRjZI8dEpMoi/OFnbT/AW7x+f/05fsIjALGLC2gM9d1KUDaznFnLFiTgcoxvhAhq85peO1ab
VZbtYoRWLIw5ItqCDlRF7GCt6G35T5ItDInWqavThIGANSzhdnfExzaOSIqlBLlYp+CTU3/OaQuA
+8YwBHLkwjvUCbemclpeO5v7tcdVxMUNbrmuJBmWUcr/hZy7EjcjYTy5xKXrrVDj/Bqt1nUh6y35
c4OjGiIGE7wj+2Q8G2zElpijMNA/M6ONo+XnGsiZyqrnF9YpjpV1heDB1a2No7hrmSV5hg7SI+Gu
oESzWeWZCde7W7+jw3bdCdadfBAsWgHvKTVItlpd5VAIpfghXJiRW9XvRkFXuAzAVM5QQlfYSB/p
sPzJ8K/1DN7nK2zrsiyaZU8MDUG7k2urglqhMG2XyOsoB+Nl5aKkes6Ra4LkE0g9tcZ1B31tKSc3
aN+Rjnz/A75vSzoGg2TNwBvN7YV1OkNLGtmnaHbKw2JIOhkCT8XCns1swLHwiwueLG2BoXGn1Q8H
i2pQHFZCbh5VFb2WfauNTKp1sxEHUetbId084HSafzmTafcFuNnK0bJ5Fxo/EQy1JOl11wx+odoS
xxYWdLtgrEqwuUa2P9fEQ3HT3lIrOvIYHG3FaCTXzGeGsEMS0tRSDgTBsAEzmbqwaTGIhI0WBFSr
twub86p5bzH63BTkMoA4/5xK0L4lh12GSgeqgTpN1YSZ6UwzNMwlAQxycPRM1Nf1L2W2Xyi2cDWQ
YsG+v4ChBAkEVnAhiMsyHcIoBcViJKTWkNB2Tt/HBWVR7WLhdv+l5UX2G4EH2ntEhHWvfIt1g7x0
7oUQfGMp0Q00KV2n8a0xa0m8iPRsbP8dKLfJFmEC/gEVYXxiGmNpbFF77jhqYLnCdSlnNMhBzBnP
wur+QtPgLyzM0JeseHBPfFxZyFWLqxkqClOwY1OVPT8vD2ADqS+NQ1Xjw7Bqmnqf+QshvY2RpwWD
pE5yQhNxqu0g/yrM1pKFOHe+1vYMUC+HMYtVsXGz7QcpuPU+7l3ZsW6UiVt1mYCRwUN6Q+prRagY
k20CudRKzH6wHFUL35KYEnFeCjzODt8Gp28hCDyUJnoCm+GOwXk60U2vJrHFDyhNUXTsaWp2ITX9
UT/Uczl9O1+hALEx3qsHjPYAj74CjsZsD7xgTj68ugc0cvfHogg1U+MgdR+s9KSqbpRo8YtNdfiG
+bqhYF3COFFTpvdiu/21JNuFcq2sOsZ0pnn145icJuntLUnuHFX0eDj+Rc9rwtMyaaBXmClIdw6/
/a/Ho0AS5HSR0uPOHsviieIbRi+bs907f2CJytfWv5avuSTp5FvQNxif30FhwgJI1DIeHr0nvrXm
eGsCcjmP51kfZH5gvo5rHTlKoBj2L7y4wbS+wjAsgFtQ9IsJocxSeTh9c/X7ISfcceYEF1Ddyxso
uNM1hca9ArdPnXMoJSg3kppMzn+Q8R6cnKTCrmYygwi7cC13jurO9duk1y6nxWZGphJfWywdU40g
4yDB83ZnrAi9jam1LD4Btle3uTXJ+70eYee34EAZ5ze1MxldjsdGOC+rxb7ZVYeqXXpu9TLzmZI4
HyziNyizdUQozOCZSUFHVE5kWwa7fsHBBL0RyqYPInunMgmh27lmzwP8IKH0uKz+kFkMg94ZNawN
ytw7Kha4H55onzR/3fi1OdyoxbBYDLtRW7tPKv1fTLPTiOrKIeW4jhsdtT49HWuB3xY+QgCYJXQq
dRx5cfZZ1/HV10QGRNcgRklR4jTVh2a3QePOeE717XJTjI9ZWtL7/IA8lMgIzNX0qPi6ZDmLX1sL
/WC/0DjQRTgH6i+f/pnTKe+DtiooK0Uycl6DajK5G/6xIxy+AmUkaXsZVIRwicniBo0aNZ/hib5+
DfrM37S3kHOiNzQ2pQlWeaiOhpkRDqKsq2cSsAUqMzD9XHQCp4UC73T3H/YcWt84sgyU7vUttq3G
hGqWKA1KnvTrBQTYAiyyKPFlvrp+Ex57yCDwnmMXW7S20PnRtVjoQ02omkmvRmtdoNub2vpV7AcA
aqPNeuqnZFoyqjV/ZNQumYYXUah2XlKYahH8zyyEa9L5VZ849C6xzx9K4D3EdD9WPnAV52RbRiV4
BLnxo6op55Be6bEzmxDM8vJoUCM6jHFoxEW+BV/bEHt3Z2y2CNrBITRhl1zchDYPvqfYWn6Omh/H
3VVLGSpjT2q25gdo5qrxPIKPR75It5/cIy64dYL2vsbr+IZQwVqH3agdYXNWHTYaAS0yRFumGRkO
uSQM0Z+WoB5dM+kChQfU/6HJghVfyp96e+fD1DAGvl4s1FQTEd+tDozFqjlIXd4B+UCP5yMsO//e
SOZpldTq71mdOX06m2hzhBiK5SgmARQ4l02oh79CXi/8z+V95swK0NwOcHX0/+faq9polOsKHEch
pxPV/0nDTq+YFO9mL7tPw9F67l97Nx4T78yDwDvxOAtBrvIyR6PpxQyIk8YhykQ3a+3uOU/IVWZ5
HUrJc2lQojh+E6VYBQMT+c4bhXyrqwvMaxjOwZC1dQk7gEmSNpQ87V/TWAN/T5AF6HSn7QpQstIk
1jiIlCIIf5EdPB9spNriwNKcAyfy5QeXwToEEVNIej1HyLp8R8PJjuCrLA+TCDcTvuqC/l7Tvi9R
vBGVb8ArKfxXKSfAFyXJf3sLCJDckbuZ8W0O06czZgy/2Y7FGzpmLPOQjtfVZsRrwu+8JZjEf7sq
+3ijnp0kvSEDGe1/rESFr1VN9iL6Ujl93TEaKtmcNMVbz8oSny94qYZvyhQSPSnQmKichubXD431
n9PqFTZ6CwVtEIlXEwhJhR6qN7jCPOaArUS4tDzRLAXKG8fPMQftdujdBCTlLg6+HOjgUg8LTzFJ
kfAGGZ4813JMyPzB+TA5UZ2CgKJijmbef3qDqNlJIj5+eKbHxJa2QkBpz8N3Ef4iykfYdeiqxaEc
QcCmuVYUzfhFddJzvEw0iWmBsoktrwPq1KfV2UZX7Lc0b7Wgm9NwTYaQd3fv4ZMxj5UpSU4il6uM
xklEF8rwl0Yn1OjTQyr24ftNM4GA8o7H+pQflQW/pkKMX8ik6HVNmvooo/LR27R8kmgoSS9nhLtr
5LQpfjw0oreBlrm+72li3nESnKjXQpwgChqkacUzGuI+2exn1z2QOGa86aqzoSj4I0ahox95YUJH
FdCO9yAhMRUwLF5h/XIDNTlH6jjwiDiDWmRX9D7g5t9aDvJZuj9AqTUFB3P/LrZebBQzjRlz2jVb
UgnRkMwfSZXxFXSeMM62Mh036LmXrb8v+sAvzJAG2S5nZogdwTDeaL6w1pWPvvOZ8DxWBamcSFo9
v5u5jA3eIlLqydlj9oesGNVOf93Qv6VEAu+7sIHnfQkpl8sOyF8FkEmApXHuBwDpvpY9FWcX+GTs
IX00Ms0ZSfMp3UrSK7OP4AG/RZua/RqRfSzF0Ctwi2PG68LWIkzSYa8webAgPJJfLQRtQ9GN/L9l
jH7Zd1o1W/frhCeIa9HsPp0YbqwMcULtKRE85343bBKRGshfzm780qwJ9jXPO1pi/V5OC8Q4nyTQ
ih8Tpje9ngbN2wTK3r53LuxS3cqGPx3GBxMVC3OZZqee2lehNxnlAMGNXZkNF/Uj65Bu+NMM18rc
3jESQY4BJmqIZriS7FtkwyCzLollITCQwrQfHCPumx+CINbiX1H4dK2ySzrUzO8uRlLulRkIEJFj
1Bovixs9qRF9T69iolPEyTbWclKZWuMnHmztprsS1SErEi0+s1iWbfhhxqD1rjOPmszomOf6PEN3
jkox6ykgVONL7J0p7D0rDN+LT98qKiQDz77T47F965IvlwXq4n8LrpT7fxXRre11upgmqPsYsorw
6Y2Htn8hO/ID6nsD8hcTAjaJd8KRg605cSrMERlegEAROIfe/mjKAAitxXsZrnjB4u5cgqUA5O2D
Hsd3a0Dep0JbPJ1juh4eKtXjSrnBJ6rWt/TNgHf/UiW1VNzB2Z24AqKcch8MAG9o4h1XnV7Sht5A
TQZ9vuXxHW3cWwgQBvj/ErW8hVw382Xe8HL4spnjJbiQojOeI00pei4xz61Zk6ifOkugGsYMuZLY
Dxy6gsrmCAz/SUS+G/j3TgTLgodd3VL78DwyLd+yJxMvt7iOU1rWm6Z5/VIiw+Y/1szKqoObnF80
WVeigAf2lHff5oSQxNgsIIJktkijho/JEH/DUsp/CBVjF3hGH+aOnfW5WCn4IW0m79jDfPUVJqkF
l9S8Ic1s2OP9wGmvpgPXKs0sBeE537djlWNSeec13Z0GHbYnHKUUx2k9eqhhiQplAjqNZVDj1oMa
3qg4Y3hkrcEADboor4zWcRifkgrnwseagLPPkO1g5AW1QX8Ebsb/A9ZIoNSJmCrnjKIQ0SaOFD1u
pBHFP5lu0UB9c9eu9fpqUfPkBxONux/ykQendHodufntUBCvkIa+F9s8RKF9v/H/YnMD6DhUjXo4
HI34eNWqVP6C5PFAUWNnYkLUekYQqckkgUSp11nFSeaB81jBagZXK1crh93ov2FniQx6Ys73oWMc
LvegBQ98KU7zb0VobeOvpn9QUdos1NpQ91rmdKryT/l8D+y4Xzu3PbG4NhhMezgOJVO+daQd/F/Z
yYrfjxFaiiNbynPipWtc+bDdDBm5Wcvu41ncqpaePnbA7ceVqNRW4ivtgoscVmnKaeMO2SnZ+zsY
efT+gCyUzjTWs0UQ5sE0R/2XJn+3H7SRKz4K1bYkIJKf9KUtcPSOp3L3MTHhlOnLp/0jIMRAvmkN
Rzyob0B8XgkRgn5No2AxjlGQBVWdaWhs1IU0TQTk6wv99n2S/akMv3rm0R6JE3nqGzz8QakFdkQh
tr3b8CGM+PG7Q6NpZq8UQFUGMCcTpDl0V3vXs5EC0VEjwN7y5yJUHjIh3sDiCeXJugNw6H+BwVU/
sOj2yKLH/KIh7HEEc9qXJEebu0rAu2vGxjNhhD/wjWXlLR85S/iPC0s8tpoMoVXY58Fapc4Z5jWO
dALKIkQZsqyHsVuZlNkMpsmqNYwYPQCGaQ0yAf0mWBImu3bFjvbt46qlvOySFEV438MdKA3fCJzc
iVq4LOCvXD8ZKntZmOU+QuuvAkzvHetAZlE3oDqJcq8bW5S1K8Uhy9qHwneMqL/0XLf39GhIAEFA
6yLyqpfJEohrwRDWAcm7PvPLlNxx2Ys/HoECjrLmgdvNPTkQ3iONFWHKwDRPO+yrlqjEZUkXKRAB
yb8wtmsk8ls/nIRzcJcPrZgdWfiutBEPOP+5RM+A38JUYcSXDaWvbUSkp8uKVtEVNbVyTZbUHmKk
tRVIwVXbgVVjtHaLhkjNEV8K1Cwz8dDKl3CdhGwCNW8TtWS915J6WyMqk4ppVd7lTpk3/ItQpGNU
7PxUhoD40K9vttFM4cRqmQc+hYKAvHNhTQZJLGGdOrb2jAGIcec9yQKNOcjoq39+mFp0TE315mly
7rFadT8M+2YxJiO/jZEwbF39zVAVWZqEgfJtbZWEjR+tFqe8RBYI0R38X7khJhPCdqbwbLfVaddX
dBwvbqEUxN8b8awocGmxEUrWBOoh+eHMFYUOsXGd3NwDjapBb3M07944Tbykpn5Wbb/kOtTYaOAy
L1hUrND77CmUUH7RdrX4M+NbphrxyEDyetRgXt+VFLdxR6o2gn1Ww60/EGuisgBUXS2pQdnNctbg
Gol7G5p2haqBrC4xEExcW2uUFSGOHdHFkP3JDuBjMZCN35MUWZcuvzSCr0OrqvD9aYVMvUrmo2g2
OP+YqtDwmsMHLzCQxCnRJ/HrYfeN+4/oXMFULv4LxlQ7yuWLUPdmOj5nqvJH8cn4h2W2eiBvJGGw
jfK09JJgwSGcRXm+B+WSODFQPb7Q0w8b5Q68r1l7qdzs+vhh+n9QXSghgJHsRLQIBOXFvuHUWY2l
nP5U5CP+zm015VFhHcAgjeveOvDV8itZBl83Ssp5mEe+jY2YsVD19Hs4pIehXaT39NtzT/A+ckZN
pFUPYl6j+FCVZmtMmyrIPVS8HxlNSZmqcMd5jrUQvFM6ZEaHtogY5wEYkDFByeezA2RkZK15XfCX
lZI0Lr/hl6wNClBQkaO/5KGdPpPNdvcTMh6udXGq+5y74PTRK+JMKc7a9h6/iXNdm0Iz1OQH+bkd
bZU7kVGv/nfcLuY2zmVVslA+8goNfBoObSq0a54nqbVQe34vSEUC2N4c6XbCor2ojquyF+mYlXeu
K74zqzP0urmJaYezTblheh3wIrg4lHvbM/OsyUUkjXOJSPex/MDcEpsk0f8ctgmrDTpptDzsa+3Z
DL1QlSHyVDBbKEqXhDtVvU6wti4YfON3An4SR0iLH2mXaOJO/lEyAn7Fv6CeKd8tnrwoDDf1XosG
JoktWLIlAW64WPAuy//H1VRVg17wRM7HD8AubBbfZmscFNwjbXmvKg27iuA+f+kv5jGxNCLixt+b
jISPVyzXLqkBTGZIjrMbW5p8Aq6rWixuzKUfGUQ+ONhIjeMplpvG3p1OvJgZLkPgNsNglqyHt4w1
JjcLL/163UPswo3Ho0LjVYXD76kUWa+ddLteZXJIFtfTiF1sLh4zSqai56J8tEO8huOB0n3WbIAG
/Mfq0Lb8GiAPEjREMeXv62Fu8sMP/RzsyiUuMfMpsagOqZpZa9udN5H3Ez/WnEocVrV2IXukP02o
A1MPqdEnGoRnBAt5YdepiJ23BgLDP5yeB8hRt9S5uG8acTPXQ/be87oYy6kw1D4HlcrrKZ2/3Bwb
DSpJNoe6arrAmJMdN/AVN+TWPDGkPUkfipeO0hlxCs6VC34b7eEybp/pKTUAnCdP7blCiLPitBIF
121M6+BeSxbQxOl41QIaH3E9/pYSm+832UEQ+SceQrH5TvdkF9wO6IO/qzTXDy04GDLQJiJgmiKo
ExQwURPc37AQVkPHOZQGl7oT6aPAFidNLY6xvCwvnnuMxBu7b0hLX1LfkZZS5SozXJ5FKKPFlg4p
jtNOK+ePV9ZDQSF/9K2azeblSvMZoRPITmL7r6lRXpxUjjLrfW9P07xMCeNKSgTSQEeEvHa4LL4n
nrzGlxUX5hrDdn63fQ8KoNNhUx4l/hUA3Ptpkir+SnFP5r3uOnMQ76p9sny++9KkjAbI2ooAt0Bd
Ewxh7LKCJETDP6AOxXLWvi9YMURI6Ok/0LE0iSBz3Sp3voKGQ2/xNIvrapRt+HWkoGdtOrWSs9Pi
MdaGEq3ZLSar0OL5LcqopCVYdTwR+Shhv0u39R452a5HhhpJkCyuB2X6bONs+YgZ6Khqv2zKXrDk
rYCrf9xa061PpZNYgGCMhwCvVlBFPtws2E8Yd+Q4K+fEN+1nroJzo+DrrbTpMlYaOYZ8I6zB1lcb
TY5F//H5YZQqvbvKOWYkWGfEx3cxiWmBhy3vjivwvv0oXyQXZIMcmfRyjMai8LsLWnoyh18ajx4u
NiwHpCa+Hlth7WX9RDDa/xCR+0Hkbbp2RmgXt8TEZjDtyXSikCaTiDntxhFvdwhk5ZCDj3OhrTJG
BEQatmWvQpBDBAjc+rkqre7jBGW09izGcvteJs6UnS0zelrIPPiaEQUt4fg9HzWYQrxpUh7pv2kO
WXF/0WyJWoc5ujGmQDKUdPE7Q5Tc8ShJQN1Z+Ez8rgvWvdgSIejchdfknQa9wVhlwmbKBb4knzjt
VILo3ftCtttCSmywkyjbmXcoh4N39wZX28o3jz6TPFtgEKyGhrNyMm3DY1C0SKmqYH07rPmda1CG
Rav2Ln/OGHzrPsHDAEsY9lHyoZ8L09h0v9jGM9kCUZ04STcRBs21X150vT/dwW8+n2d0bEr+U5Dv
qWaWWiuZUO0khI/M6kMZWRB6NbXiFQ85fb9w6GaBZA+p3XJtJcppeAz+TCKyL877o9kfxIyWhGzB
g7Bd7oBefEx9oP8C16iJ5QvAL+/KWMJNzHpAinUoYyiIspbRLXtRfWawAZl0X3jbKkCN7cXYACeD
k/GNNBYfCveZlunLtw2bTOpE6g3p7x2q4EDKVIEG+Jk/zcSCpXntxfYJjRbdOx6oZuCXI8aIBrz+
N+pF5owlIB7I/h6bwF/zCfD3tSeHISkjrJxUOcw2n4TIhfWEdpyASUisRY3qqEZz6sig4JoFmEfZ
YJFIOfGODKi2Hky/lZVhHUC9X5YD7YfBhD8j1zXuHjF8069PpyUw1wim4DBt/UJiawz1fils8coO
KKHxeYDNzWjl59QqG4441DXkqrGpX5Uc4dv2zHl6/M3srCQjpTUgBxTewJZYk6mhHBzTTCyTRnPW
xo+/2ewOiEjLjRxAS+ahEUGQy0JullS5Qsovw8u7HwfW8RjafqUfbFq4ORl3KCKv+MlLScG6xYRH
/H7TirM+T8pPQ8JV9dN39/aJ1W440jOWb19Abyvt/Hxc3hpRcEhIem30+ns1tF9szBk8RwKgQGIH
TzL26RstuagzRszeMkVEH9TarWxfpMf9+UcJ5sLsdqCHAEiIloj0KuP17ye7PYVZYaa2UNXv7C1s
snheH+UPVjIml2XxLewxkA0fXRUdBl2Y11AAf87156MAX1f0/bKTvv8m+bdS7YIcDewS8Cc4+BD/
EVc3t797vOAjxGB52XjqJsfpwiBGw8S5o9BLv3qXW5Syih4BTF4KyLY6I+Rf3vQD57mtXZsY+zgL
4nFd7I47ifpoiKwAXCvmCx51F+uCU4HYFqRtuje93NUTwa+OcyJriIevMe0gPC1Oz/cQrwZ7MxTM
QSYR3XBtNVM2ZP0e3hPGbGhcGRDE5JjfRW1CUHvn1w37h2an8CKZ6jNQRwsbjwKihHVrsCPQWsPZ
tRcvz1QgEcAKJnnBQ/tYPiXvJlBhpNLRGbUTZraVR5Q1QEHf/Ju4tOpplYsUmvfeK1P0jxdp/46K
LVi08q20aRE6BUab2HQM5Ohpg4udhEhc6izdinbqLWS/GU02/Rdpf+YsWMNXq7u604hmEbt966VR
wvImorKsGTFjl45YwSjcxbViyM5gNnvu4rjSkH+iKkKFBvRrUaGoAt4Oi/5NNBElMeRG6ui78ZS6
0CmSyJgm6k8wVtD/ll6XQnysU0V5Zttdlvax0dmatqu89hOGVzw/kRyayKuoUol87+Wv4RrzKk2C
t5AMX4akxUZbMdJjZ0jiUJ+jmMR3Hi8l6Op+Mfn4tr5ksYTz8NDYilKFvtP3sXsb2vaLsF1eSf+u
tbAbycpARXxEIc1haok05FvUQqiyzFInS9NB1QL8EKoqdrTJyMRu0ZrSn5rI2c/GK1rcKCtsqUif
npvRaqaEQ4lbELCIv/RVK4qgPrQvrfyOJMwtrml8ql+WFaHTaDFz3hNvUYkjsk1biF6yF8O+YF7N
s8IZSRfKNij+QeYPyewwk+ZBQwoZ7crVlP3cW8B+nLergqRI4dKwkvVyTHIvS3P7GY9rMJwN1TLI
8yieYGcmEMiRFNB+GX+DGuURrkXHnYN1tEHs/0MUq+7OtAtTaxmPt5SHXrwDEkLIcgqsSQWH58JB
34nHg//qCSYRiEQAv3Pa3CKfwtMy8TZgUts42zD/NRS3NpsdAhCqZC/qGTOu7LKlKS+KkaHujJDM
ZDPaJfYy5Jh95oFQNRA5U7pmzGatgBPo0i19xdUuy+RkT6RG3fidDlKdX8W1hE4VM060kgQqb5JM
PKDN3/D3hw2ZSEhSLoo0JjPO02XLVLeG5oKJrDVmzAAVrwlzNUQ9szVqP7EbaRX1VEBKn/npy5KL
sTjok5n5mcSG6I9oCPczeAbxkw7ZxzWY5Nu8d92vnCBLPLdMY/o79V7e6fCByyOQ3rNNzCoTeDG3
6iFV+WjCQ4OcqK4Qp5QKo6PJIMilOIfpmW2b1fQH2tJOIwPbDAgOrPYCfb8IKAKHyw0I1ojVhDrx
RYjGZJx35oAe4FV4WMbtZuMe07qG5XBKvQEVqPYKJoxuxzgKGU2nUlQDpODg9ziHkVxu6KqJLhGc
GFl2cGr+jL+RVKdNALn8K5sc7fYcUdQL2e1Fl3ZMLjq9svRcmsM434ioccOBXhnofqB9ijvu7tvn
q6scKt9eCri60itqgy5OzrOY2E18EjfzIKGwTTxrGiny8cZJ7dxiT6c/ektVfwVTjMvrCzpw+S6O
DTjP6C24P5O+DiqC8UXAc9UMrPEOQsI+w1KyBgm0/lNWTgGSKQbwQeAgBedGm9xna7j+GO5tpGu6
EMhiOxtMX9/4Ty8DnsRlhe1FQXc355wTe+1CgeV52qxvS8oDmnV0BO0U8TB/Iok6RpsUOXGrJ+54
IkQcsofkjaZ3GmM//n8VE6eUvGJB/LIHf0xZJcET6C3PwtoSe6PZ302F0+Cmg7fX2W49XdRFVfVn
uar6rUSUeoxha+3m4HKkeVxV57qCxjOGGcnUS4zchL3y1yqX9jcqEHxsGbZ4pSYOILJBGv6lU32D
oyOMzvWWoDIlCNP6Ih6MVtX5c8Q62NhGdONeurOGU3lRvUouKUw+eLoZGu8iBoZhJWkZ2cZWM7GR
Igz9N9djBFoRILLIk1/8tdh2kzhDMQ1ywdSAtiNmWcTTwyHH1L7ue+8fqFV9c+NcrJGZdqCxt0KK
T6Rd+X2MUDewy4g89w0lo2XsCrAw88zfsOEXr47xVvky9470TrdWEaQO+1tC+AxETUJSZO/b0vQc
Twt7dt+jIQpLYgiLMR38YUI41IECTL0lNA5dDnVwCSoe1Ow4yu305kAqi7FXe9AI7RK8IijQRqcA
mK3bYps+v1rIsAK5I2OEVAy3TUsT5ObCwtulBP1qP5N7gtIGTDFtKFRPrynBPioBPEMU5fwvgDhz
UUIDWBogNGIjEWI3cYyR8FOeZzu32nq4hX+Rq3dFIzUOtKEzU57SZx0ACqexKSR4rPRZ/gBh/saS
7UPw8eCT9WuimxxdhGB2lU0rSMefopDTDBi/cG1ib4fuzfyHUGtSc8Rwvg2yK9ItureiIQc/iBDr
stvPyK6+XCqtvbmANRfiprIpqq6DOx/ubBJmApaswrzqovrOv5TNg7hWD5GQu7NRtN/TKp+0U92C
BBAkhan4XdZfd5D5k+h1+lF23RWTzV+sG0gx2ZJ70B/dH3Z+uLOSDC16P8AVCX1s7f6dF/C33B5j
j0bIWJ/PlU+3Xd+0fGF1OtIkXgzDGFNco+3XAtZrrN8ZSwj8AEvFAKqW6iYuWIVH6MJPM7rzu0UH
z+/j7k9h5cFaPGX5IzWRSOjaM3X5Dhd8b960Zdme0W2eudCpIU9Q8Rr3+N6Zv5vbImvk8cLFn66x
Crl+Bk4MxDiMtu1x4MMP9PqivQ+FaDNcblsPUA/8J2oUZHK/pQm3SdVjbh5Xdupc45Ip2+lQmnlw
sEdmIcWY+sYhRuRRcbGRjJCZ3JC7Ps0zgLQ5Q9NpkKtizPpYOJxPkfei9kRFjb4VCNve5+k4sRhn
ayJ067gpeVrTQbR2P8Wn1h7JMra00vS+8wIGu/rnhl9n1KzqqexZQv9GTDRt1FccoYl6AULvVSTL
3UE3bo8kgumMFwwb3bJ43UYC93Y66xjGW3SgbFFVikRob/rF71JdyqIyS6qV2CXp5FVGlJd4a1SX
tacr3ez0xenJJqny+/ppiRydWKe0FZRzgcTOydVBmk7vNJtYM3pb5K+8craHegm3ItKWeqEQw2Em
/8jGt2nOhCyyBUKUbjRzTmYwpgI89G+Fewt8h3LdT3vxpN/K41qEk9avHsgtKNuVr6RtrJlh6MxN
5QpAWzeln95Dn/oH/wJm3QdZ1GFU/8HwcOtqT0y1GETTP1WbHPbKaodSahJVEVAa/AeoxiMo7JhO
ncINyX6tnpeKc5VtJV5WfSkHyHyfx9YFHeklcqDfcKEJDuR5SizRv4qeGpW3Pbs09Fqf9OYd+udK
N3cfw8LQxO7fh73pZC3Q1Bv7lSsYAgDrllsIANbIFjoJgkz6UhbLnJrT3J6EeeYgh7FHYRrgiYGh
/pKYPaWT8ymR5+cQAl/3N3OlfR92HkUJpcPeZfap6rgKZMgdMwXpQhZXEHuqimlLoI8XH6bY2yeo
PwCKKQrKUxCVQLwPGwDv82qc3jCaoyGWMzxOPEfQRNrmlPt2cbwnGhclhEkyq6omuo9u6v8VUIL8
SoFWuW+833n+7NnRZf86J0cw+quSqhizS3yv3YaEUTTZLSNmtHaxJBFIG3VUCLBaHE2FMJWqLfXj
dB8J1klXApG4Iqb+a3AEqbyjECeN2XlaXmEqmdHT5e5cmt7hRVFGAx07JdrYQwEcrQErOfSuB+iX
dl8FPxNz9ropj/BXM8VQfcwHfaKQ87Dv9MwrpcgvkbHbMHlvE33Iv6oGCnPBggjm5RNIns/hwTPp
x/3Niq+EQ5+Au0W21o1ZQ3xxqkkl/PBG2yTtmqQGO6NGZZLEyu1OV4/EJOkNsrCjD0gyXZxm2APz
GdHjora0Xtc87rLkrTc6nIRL5bOB69sat/zKvSsbPXANRPhcqYUQX14s7rWZAnZ3HcAmbFrd+dbC
8z+87hbEZYTx9R63g7J34b5hEh0MKzRGtXKg7JEVokyppLEzsfE+I3hAj563tzKt6U2JievziiOw
07KEA/418yq1+wUo+18Lar06GEic69DKFJC7P2rFhIeTZfMmCq1yS2QoomE6X4gEA4HszxtCF/9X
eOb1PysifdJu+O2s5WCxcSLxHaeGHWlEeiDS36iSOogHovPlpO28MAKhrn6cLtdChLuLewZo+c3x
Xr2wY4o8otaHSPSld7V6ysfSL3GCH+n9rbtYR854PuBzTNCv+STOhOHPgh3tz/9EncqBnI6A2OWB
QMDKdp/uej0E0HQd9YuIiK4u3xO2oW2VPHa+pUmvzJrQKVU0b7Kf+NFMNmJfewgEfie7MILbd+CT
0IT//uIgwuL4klaGlEBJROauCbaji9kNP8bHr/q5/5jqGhYMe4CMpOvwH/PU4oN7qPJJJQxmDDbL
ANV/ryBP/6ExhBnRc7dmM0yiE5Z59v/vtuL0MOhOQECbHvnH9CXYTvFooy9q6wYV7woCoZZ3RRGW
bYNA/BoOOhs6dcFDwIWCue09DrOFCfezRdPvysesjE75kcdCPGf6qi0tmA8sOJ9UVunAkDEuCxjD
qQ52X35Spce/kgZ9HT84GRW/7qLCpj9OoBn64gsqSm3hK5HrT4fraMO3r6zAR9EFRnQ4n/N9xIdE
Boe2tup6AGbJfXdcCvOibiyL1AzDaIOzUORE9jvyAX2qa9j1rTmL5H2NWNQBFQaxrHsMdNNQ9n2x
LHAbp3aanveKn7zOCpi7Ube8vwGojNdHGF/cWv/k3kC9J2UblZ0y/8E7xoPnf58dqOm3M96KSCH4
RbmesLySkiD9o0BHL+/E7SlMr0PF+uZn/KHkU3k7hwEmWBXrh/dnRU97mXDkALIC4gcKAEvp+N19
Z5ss/copzyotA/O5rBmamR7UXLP5aqjB9GnbwCvmqOPAc9xWjW9RiyiWDoUTrNYjNWXF0lGZ8xJD
OStYbcKPJHstZDSZHMg4P0C83NxohLEYfZPFs5VcXKAieXB9nQUEGBg9iuKfS3o9094nU8tFxZfi
pAC05/5kh8J5A6WGlIzwRSKnSvii8AOfbHSbSB5/fXVuoKd3CVg/Dq+ZDM0nDyxKIsF5QLv6v6gQ
r7jeQPyLix1vpDIboLoJZtIOjnCzOh7sLWMKhonGq1iESEX2znJi90Qtv0tGxt2JP2ye+tOb6bty
8DLO0KcorPtkSAja+w2XBSoszpY44vxuHmXM6/Lebdxay9nLAxbsG1TbkEIvdX329vhiIlC84pBx
72B+aRbOexOWe0slN2dkdHgV4X2Bdm3zHlGTWH1J1ZfN+PSqnCFUbt9Zsvp3CbjCIht4IyUUAawV
WfPLOKl07SyhQPeylipnCQRcOHVmHZWFXhQI+1E9bwYooZCveqandI5hepLTEAL9LEYJYCBgPJsA
Xx5Ah8WBEBgXgOJveGpITMpcgq7lkhLzDYHSGZk6bJzyyDLWsKi0D3TUSX3oan3k4C/X1VjqtyKM
/Ur2XVcPrcJca3bNDLuRHe+3d+gzve+SU7sTInTC4WV8zgtaIPw2DKr9p+OuefHhvxZeSr/2J85R
LaABu1amRuLssBaSBA3OMcgSKX2EiKjVlsiPwTt1IZqvQnPY3tlTVdQfxB+Odfo3ajm4FyrJxSIe
YdzFVx2ytwL5jNzfP5vp8N5b4AjOE2OXC5gz5Yexa/Lw8Vv2h9TCNDpnKN6QOnPxISa7wLLabUqT
P8/b+ZtuQuwWV/y9ohzRmD+EXrddCUeMg0bvCw+3jwVV+9R3nqBmm7GQZEsgY/NtCnDMighmnaut
3fMUgJN+Cm2iWQZcUakgbTHZRrKG4JbnmZxUujo/LHs7c47ioWTX/1kAvjanz9nM2ei/YLzldHro
ngGw1KLHBhDHI0XZpBqOpUDUZ3uEL3OllFT497dnQnQxCDfj7YCsB6B8jy2fwqNHZotOH6Ey/kNp
OXS0hSSQSwP+PYbicyVXegz4SzLVLNIC/SEWVZsRxDX+EbUmdPaFS0tB5KI6qe9hiDfF5mcLNA6A
DmTEUvLJCqqAXO62ZeZdIrIYDhUkW/+ZMzpEOISLNODkFrnWT5lll7xfN2ZBCFjrIQKUqBKTR4Is
H8wRt0/t87zpqzIJMQQSxh3gqtMHOmSABHikopwIxRxvS36jOP5Vwadb69vn4wb+NqRwuJpHnsJC
TBY34JL8hLVcViJgyePeTtDiRptM5dsrvoWK2G41+MoMmykdvM8soCVgSxJhP+ssVg8XGF0f6/nY
2OquS+zJMiVTnSC6f85YKCHVkZUpqys9t+YeuVYPlHwHM10efiMwAo48rcwVhP3TlgFZnG6ac+Nj
NRFlda4h3V9gG1NjhU5L4IG+gJiVSxLQdu9+3KNNM9AwZjqzPyRKYId2oCo8uoqjzO6Xev40xvFK
dfpQUKGkgKIJRaRjW8oruOmzkle0FGB5AGIahc77k9Pak6xjJYpbQNguMcWVYr4Z8o1Aw7wHXmQY
2jAMRfefs/xD2/ZvW4m9t4BwJOqe0kggHysMoLndzwI0uL92VAw0owzv/9QNYpqOGy/6U3BU/Xhp
ldm8wG4D8xFa1T8iJdJmkuuKt9DaLBxDmn80KWrEDjl7HXwkRMWA8qEmnhVMziIzteR6V+SnP2AZ
3UnTndNoGvjtFvnTyKx6DEJBkEt7pfFVJYqwhfIzc5q2RyeFPpLtL0MWw1DnpG8Uu7S3uXduvkou
YccctkTtG58nC9fgfY3zIxZ57V3NfVVbrVWztBY7frqlhr+jw2ziJKq3l9AFQkbbAhmACFBUeY1H
4e6Nmo5sTpygLh1QU42/mNvUlrcdG/h6MZ6ybG8KRBhq4CzbIeiwnrCRkXwQNTxKaczKlyPMU1mb
3htD+PN4hbQhed0rlU5URd0YSQ6SQXeG2NMTOe46+5gDHd73YKHkFpN0LD/6EaoKl/pEFR7AYryg
4RyStwHrGrm7OA59vgX6dPwMvHNS05PWCFatkb0bT/ahnHuHh8Zg2gmtrMXuA7Pn2Lbmf6MwnBIE
0SN5wrcU5j9rChRYjwuseGhB7TK6JvVj0ijSjAWYUlvQcqDMya1i3S+7nDgX8usAwsNA8+KGBv0y
CU5o6r9pT9wcLuBa7nS5q7hnVaqwSCCHZ+j7lAY8sA8XBwwjCYv01PExPW0Hkwu4G7vsp3KraqjD
KVlwRi6T069EhhyDS7uFcuWM6uxpD8KNkUe8CyndeE0yVLOHSu9/QdxL3CAxYmTult+DFbRmgAzF
100XkDssBP6wOM2bWY3KE2n8rzy3/SLWXMZtbFjupsbrDfIfSgtUKsAB8tIVG/L22gHn88fUee/S
7HMDea4/2tQk4uMxKBnRpwrYYV69p5QgXLEmntRdV5ic6ScolUnjbYZYQYXwurmwjyl6TFQcWUvU
0ZthW+3zlr2NyOcPqdDR6EX7ocaczpiabpT46iOYFxEwkSA8Fvr1hcBZgldf/RsM4aXtbWNiCz5q
89BlxBSIpxi2abDWLaO6p08jLS+ZifmDWvADEQxaLOze98O6Lyez0a9r9uxdwpYNpQHLII/HS/8O
Pukl+sI4mlNtb1y2XK7TVy5+OfAKa0ZVl9/QgoWhOURFBrujrj+mg2iCB0rwM8sM7c5cpdcekxwk
WJL0XALPKLY41+s0Sh0SBvDIicNCPjxUGgf30KpPsNGZ11GQGmTBWXsD/kzp1ghoSEcKq04sfPAY
sKWtU2k0AH8+eg/AXMzhyrZcIHUZtxImMkKaxyTmgJkFM2pvz33Or6HxzBhb7j90GOukPU+pJFQ3
j6bX39LUEgO7kK9DWGT7ED4n/NESBAicSVPcKBX+6p9athZoS+K5/pepltoV1Aw124WP9yL8KMSK
q2a66JF03+5OcTlNW+Mbm/h7d6EY41JxA8qR4YeBBYc8yKJVO6w8CkG4MVGOVtORSlcGQ1v3MidU
Rc7JI59rxp0GIufg1cKFa0zSwWP5kIpq8+qtUFDQNpsPgMgdBCaBzoFUTq5uglXhztxVY3eKInoa
6zIq/vVTyJrU24QkVSDUbi1BkGTR9oRocy4nFjVW4NqwpJl4lsvq1QdJW1thENoxhOTWIZ/YOd35
IvLxsWDY6gJ/+ha6hNEKsINovvlVdmzViILnpJ4n2xaZ0aTTmiPlS7yQOF4YJlW8Uo1gRNA1rDqe
1ffkEyXw+fOibarHQfKhvkgPGgRBm3VzC1HfjSUtGpMKHyC1mjHzCgqOBv8/SmzwyQVxOeD6ONKD
y4/W7XcpJEArmNrdcq3O8uZh0QBK/duajg3GECcXL/i8QNgAoWqB221VEN+mD2ppZaUAaAVD73+8
ijMHUEI1BURcRwwdFJrk08oawbztOy7uh0yfUW3HJO9PEGXK7/X3NbHgUzvc2VAhQl+BGrzgq6b7
E2MajCgWO4KE9hQy4gwoZ3/hb6j0U4j9PmA2IWh2jI7J+tFZ6gFsR4ebDK4IBjdHKGVG/2/NggVQ
qddvuwp/mDBrzYbSu6ILJUGn8ROOvwKEdwdGk9OVrex0ovCxDWoa/mEQ1kdbYhK4Xse7LozPDoq1
dX1lp/YTBVnSm8RTs67Qdc9Nf6v8wK7UOvjYOAG0As4EXcVkeXsPD86hl4XVf4xxJx2RfLt+WjOZ
Bs2K5M7v4fiqWDnkjFhZJq3C+/n2H1AzXKlaqPgonnVm7zXA43xVjIFeMQyCTwSnlnkgBg4YrpJ1
14SCRNATE+/vSNiTynAWCx8wF9p4Oagj75Nm+Pc4VRT5R7j3ZKRaLbEmxai1upqFE3xSdz380u8R
cpa+ZzxLm1n0wOHcsTfT57oHJG60ZQOr0aauOi8owChfPjbrDlam2Il6kFteBI160WpkItylvrT/
quoFXcRS3yi9BaL6BiH5SFutvgLEPv4CaWrlR/05vVNV2rIArICF7jQULYx2nquF8G4Hv6aWcrfP
OeIb5Jlma2Zf/WatNfRH4oX5FEkIZtPTJcNvtU3wMZtMtBl85WvwDJpEPkB/3e19R/BQoK5xQkK2
KpjIVh27UGGMEeN8EfLIK5GWZ2o5uBQgNp539nnIHzvA8+nBQWWxvTqm2I8YJWaKn1Bh+R2LLdes
OcTKsW7Cb0LiAwoiTR9Q5IFMZRU70FWAFEViJawNrNApvrIixcwMSf4RmKZyV+ydob8OnsTs49dA
J/coyqSTZVOABAmiF1D3v86Hljk2FH1hDXjdymz7cs5pXsGK9b2Opb2zmWgKqfRsIF7yo4T5c3Ll
h4Ks9nvm6kO6I6UN/9aEuuCBNMZu7Ux40kEamQD5UjTXv5D8nmAguJa6C/0FWsHryDNoUC823JIo
rRW2B9MJcvR22ILnEhHBRdPpXy8hD66+2Rq3cpS5fkUDrvviTsUELjNVuyQQnAJyMWHyqpRrTL35
RDJidn5S35a8uBp96GVyMNrGMOvy9E7SCexDebQIv9MaUTs7mkS8Cv9BwmGF+/5XjeW55OIVz6dW
tK4Rr30VGo7kULbserEcURlU6raKS1EcPll2KlayF+n2wyYQS7inSRFlV1DSmFjLl5KVbE3qK8oB
pJ3p7GgU19hdmyPiV6uHpTAmqWHXBMdh8KwnQ8FNitrfqXulH21n+DyEiHdglSck5CgkDaMexc3M
c8aXTqsx8aOcLoBLddd3Mnh88+mI1A+4nwWeDmMSRRoJ4p6UzgXdX9M6lZEY17mrEvU4JLo0D0k+
Zb3xutDKAsRPcUqf015K7NrBjzPAvno5AekuXL1AWKkDxV1SiI/6xHh+ZU2Yzh4sMuiT/1EJlSXG
SPsEBXchDh4wXM8C4C38NVjxKIjL3ISIrJLYpZ22TumVqSPWZbTnkDdxKkhjFNN5F7GeKMVoi3PG
chihG47Ldj75UL2Kn2LaDAW33hkCMnw6256h1xsQElAyT3dfUvMguYMxEQsDWL/BGthbY5Ak3Jsk
YPPKfj8IL2ySABq64UlNGmiDg1f6/V717JeK8WFgIW4+mTMZ+FfPumFgvWky8n6NNYgiB30MVPwP
FGCLPm1EX3AsnB5OmsuCvbDWGh7yQQiocp087yjKBLtRjm1AEovhbqJRr60uJjZfNwOkBTNCImbV
vtPcbI4FpPcHxLrneqMvyciljpZMRF7n1JcjRMM2Pwiy6FvxR82yHnbgghVxpvnKjDdIZ4vuFinx
/kg6enrP/Bv3gPzdRLILsSw40KKf0ZGYXT0ITaPwF0rTlR+gA3Pa8QpLQqxhpZECMFSQvg3j53YU
mUM8Fe6922Y0y8ZJHZRyV0tArV8gqug/jZpwqpXez0BSv1NS4d+/GDTqaGjotceEvQOEVtqeTkW+
9jj+8d79Zhsugbab4KWFBzr925a+zjA91yzeDiHfgx/sZfOXxklkcoQNsBGMNHqbGOfiq2k09F3Y
MrurQ5ZLff/S5jNxf5bQ/FdFOCrLrU282lbUBgXCzaPanyszDQ6tRms66sNOIEW9sVryYtpqQv7y
wae+WndG6EwKvX2j4ARykY04rPdLuUBlm/TKW0CcnylIQZghb+6gg+vbKRJyylmsIxOQUgdJelBi
yRrU26P7AlRXWJej+YpVn4AtQx2f+jj/Hz9ITbsIR7QneCer0jkkJ4xz9QZtJ+64ntILwBhmGA7q
tdP8A/Rji747YlftAI2S0LJ3mtcGXdWQvPFUQ+FP2FVcQcYTrclSKafAchHX8x34uJAmvP4hvupB
5KgQMMCNQ9rSyh/Oh9glzVArM2Fh5JleZuEW9FSPqbFZc5LSORH7m8lhV6aem1fPLF1DwW39vwWa
iT5hoWho1xdGH8Jtv+YG80sGR6rzCVzuEczS0fZHmyVdUXzFrxm0DRQQhYYIpu/VU4rIDawB04h3
qtEYqbNBHgQOoIahXvjeKNh8mECPIcY7WhktaeQGNYaQlGVNcDDiquA5ayUF4vyf30DvC0LjgcJC
8Kl4H/jjU/Jg80zjEPKotaEEnO1FPQM3ZAJdV6ofTq7RtigFU1GLN/m0qz20CQ6p8UNU+cADA4rp
dQvdKFZZKn2mvoZoyB227FsSmhoURJUw9p8I18GT1GFoH9Tw8oW/4e1mKEIX7o4fI4r5mODAfV7Y
e1veVZIzumVG1W1ZGFOMrhrP+JNVRU0p7myYCzVFI7OsoRwENYy6gIahfbUw65RdUhAIRVN7T/B9
2mr4hyrmIOG3Cqi4pDIcmXo9Vw3W4Ng4WWPKtvEDbW1F7tkmOfBPJvkb/XpF6rgn5F8ukhNMCb8b
c1Udf7JOsEPOkAZ9I2sgswaJEcb2EE+BN1c3o5ExK03bENcX8dPDFs1K3lsdfyWVgFwc2E9yWTrm
73xmzex4OT0nO8kPGWYMwvAFVQBwK53qNhB79nMkDoImYCm9mpu286yHIfO+F6R6Kv5/sgPuSOq/
sBh1HvJPrqoYTR68B+nIqREiHH0tRjTPFbzjxmB3I65PI+QPA4hEzUmsrS8QsT1VAIKgGACtC1XH
4dMAgzoTSVFQ4BtLJXJ5Pqck2WD0IANn+HFVOiAK22ABTJ9O5SN0G680599eZQcxGCEMWm0Ln18X
69nA3AiHrv2LQB4wS16kq5Q2E0awBhCk/WuFppEdzSNPvD7mhghmL8L8IzIlNNjG+f38mFMNAmq6
17r2y8/EQAiHpCxsR0s6p8JwAjyvrYPoAx57ASywmNU7a6O+jeUfX8WHsS0THz71cMp6K6B9GOWW
ixF8yhE2z/qKABZldUp0hcyff7Sweq29lHPQREtOFneRLmHZJSoZjs4DuYzXZmXQ/0j5LX0qFfZH
t+nt+X8gfzinfDkQWiyqgvr/ECi9THAj7NzIIACMMg6NRJ2Qh8V3fZGfiIu+hL0Jt9xZt7mQA6am
CbEAmGZvz9oPVMcgUv70cw9yQ0JLxDaDIJIodatsqZ1is9kMvC32zLbSp/23mJq0kOBVR0fSGRxG
/B1GiRu6gW3SLRR6nhtRceN7uRvnrou7vZbIsLLmGOb4bNhXE0LNFf2shRERy7KdEQ3X4weN00g+
9urhaTVQVhmbO3ICSofOKMe1Kt1WLQt37SEBJ39fO0CiSG6fCjfyx2m/t/CcirUzURBkvIo1xItr
hVPDkwuu0j59+dw8N8nwrZ+2stWMmnoYzcihwCP2N5acinxpIXi59ki0a10/L74opjzeYGT1e6uK
Go2Jf1J/4+Y0tB9udtDe6Wz66TxTwjmvck7xRXxTOKMP/c1xiYcMaEkJ0VS13nYhKZxxc/P/lRX2
heIMyddVvLpypuH6X97yLsSyJXtyQha3X2kbgJbcz6kxQg9pOVNfv0wvr9ROFWWYk5xsNzaUm+7y
rlS8Ust0u5wNJYRZXcPn1IjVTvz4OJcF1F9rO4WkBLt0nqJQNPkD5S85N76Lo62eCUw1Gcw3vPxJ
HaUOmZu8JwTMC8bitLp80B92keq3NzYs+cAiMVctKcyDYIaYja+usJ9IZSwahZ69EAeEYhBU1CpO
ZlrVrnQvQll77sMZHfg6ZC9ZI73+kcc7q7apqB8LRYLWY4q18a0DMjvZGuUl1Avm9XfjBVdRFEXY
fAeiqelMQ2d600/A5lbLFgi+fs80WAa3y3RHBB9UV8ws+D8YV3O4CFf+ROgzrBKb79Ve4pWVp9tT
OoCWUgyUYydYgI13Oic2H2e00/lPpN0Zv2sx3EzNl2LtSRUpPy3mYGzrkTFY/ahygfccyZI6UnVZ
RFbTqsQTkXLfWq5reZgYXu125i5B4GrogYM9NbMPlOchxU/KbLdbS4+RWk52l9EwBfk4YCC71jLw
ZF8HzJ1A8bj9DpuBwmMxTM0u0UXbPfla/EvT+IS9sLuT3/vLVbluiyB3PWK4hRUe8EKRyNtSx69s
5vPensdA06IE/0ZlV7l2GuXQwxCYtpBxi1gtfBukx2V953dswT6kVzgngCl058iDmdi73+M/yPcy
xuLu9tyBKoGkwZci7BLJv6wvGJ5i7SiiZ3R5PA3LLxlhGt7RnKYQ/N/lDX7hO8Vtz3VMxmh0wv1s
cU8NqEPNAoyTQA2NI4gpRCRUlTY36KC9c9gHvuEJ29oW9bLqPCU+HeqhyCNAhB9DHGCSyDsyrH8D
4SR6jl8AcOsEcmnhtE7mKPNxrNrQ0okFLLb9S8v9AI1MmSe83Uq9WwNX0KTzwW3CfrKcbK2AGM8u
ZpCPLJrwrWP6ftSKzX9mr99au9dR92W4qb0qu7bXcCwpYM+o/s4I07Dym/fDprE+C/fTGuUf/GOI
N8UBwvdM7xo/vrH/3dflaKLKo74htlBIvwJsEVibnHuCQ9FCWxPOh89KBYlUh7KN1duShYXAtYFH
+Rt/KavrT3o4IUL1blF3U1ou1V/MR9p6cQfqfMQQQGS6uv6OEgWSsCikgL+2gLizAWRplGvRJrkC
roN3rLnZncltn30lt5paAneXvCMiXeOUGc7k/vUlMk8cjY2uNnRRVZ7fWNz/vfLfb5+doRLU9aTb
+PzdNB+P9cVJfcvd+7D4tPM+CWjJYpqU+3kU6Im3khpKLxNhbV0xGnnvo2vhiq+RiV0kP3fPzCXq
U7sjYSMc5C8j2senylvjquct6ZrYMekgywiurkCaT7Uibua+2h0Bvp+lMRBMiEpOzmDk8cGeHYxa
DWwniKyJI7/prQT93byANydgdrLnTirmMxSE8qcHemOaXa2RYkF+BWsPDKiROtMxkbm34M0XBZkr
JBZwq3C1qVA1Hj/Ty1rq7EFHiQC82qYp5IlrSUr0P2J2izFoLVzpgc24AvPkiZmss1iOWCEJOLJ+
oh5EpWdLW9aF8NjcrSSpZCuXZwjIVq3FTIckCkEdkzwiSwM4CU5jeaqEYYZATS4fp7fxXdYRLKwi
8lmKgW/BSRJpTJQyyW9kjfmuQFOuFS5cwNB9BIlK4nePhWaSt/E/OMp8erFES6HkBLzIG/dFGxnh
5L6/3pQzKwl6IZIxAqDjJ4OaFyH7jwXPFb14Kl9nH41qsOrzpdyf+HktDW9K84RtiqEAg6NijJRG
gvtRB9yUa4u4DZ2mzGCjxIr1LJI9VukCj/hehsiP2g2lNXkypm2LmFhLdjlDTax82f0CcEpKlibZ
MjZ9pgiJrDBiJM7cRh8oa4QTssxurKAUGXtdfVSiqkbjOnFXToClrRwX7dA2wHS1wxcZIhRxXZaA
xRLptBSQP7/opzeA1dX25202hiop0FNKgK7HaYdK6oQgnhxwgXjVvwMKOWyUg1KlowPECE6YsGUW
83azCBymrv8r7Sjbx/OUK0nTp1P8yqQKzYXmqRMUAoY3E30+4R71vxFmG0u1aTqFL2Fh24chnT2p
eRavdkUx/kmkn1gUPdN9Z3TJ1eSFqM459kqnwtODH6uTDaxEv1iQ5fO9wMogfjyziex9ff3KuMcq
ysb/XRKhmwIhxG1nuUGo/q1Zydbkgm7pPpkMAIe9LZre+2JzCgYDaFQv4JotCUbQVMf6ETtuf/Om
Ys1YlIsG+YmFIAAGVFTu9Pdc8mZSbhtsYKNpg9AU+rObo55Hw54lb8uxv+30q4/9iJgd1laIpd53
TVBwnpVRwknaJSdyyiHUL/hwybEiGMklhvDAYT5O88iB5Jcs5Qi4VHAe6p/gy5XhWi7/P6kDwNa7
Vj+v6/wvyy7gHkseW8em0osfYYPhx+Y8r5eMSCZNlF0Y2aI/edGOoCg4ZGePqIHnLdobNddMd5wM
w6CKVTiYVMT1cps7RdS1hIDt9B6EmfuovMknt2kg3vX5i75+grsDr6TzWkHwviOKWb+/ooK5Jte/
Oz0I8KMRSgpVwmBGKD1+4y/2P0ySmXHsIuRJuFKs2/piKP13cL8rb35RaHQMJo44QXBnqt+cYts+
0cfBR1fQSjhNdybpuRrgtMSukMfKEMgzVD4qBdo2sJ+yDNuUa+gfoYUQZ+PfHTa/2rGH2tHE5Kit
ZUccVJYneXG2Aad7e37no50KwHvF3CxTkQ675ncCfeZRiNRSZalOxyw5UV30WnUW8nJlBlCffwi8
cqRnGFzMIo3IHedyRFPyFDdF1hhZhc1GYSyFf/GwFPO8jrFlFaRgCf9lC7cyLg7ybpuuazUaI8z0
LjP7VahQ2+QjhRCAwmn8GOczQaz0xMP8rXu6+uX57txw3LnWyjTl+ibNusqc8ZbR/TFXXNV7rpFr
lwe+PP7MLi0XG923yiXaJa5o/3PnMorS0dH4By/87o4ulc3A9W/TNWczawDBi2jFKcCk3msG2+7i
UB4XHEYZKnE6nh1je6Sx70LbLfUQfAJ3GK0h4q1nmSh6BusxPXI+23zkDPGlLUSGKQAjn3J6RYVI
NejmEOJTdeUl70vEfohRQdYWjobhKvzTAv5Z0nKhGVehuCCQY/am3OA38A24s5/MtBdlM5hhtpH5
iXLvGduuybSfwoFGw48eSYo6wRX1tR4ZFZ95iqz0Ot2XhvEP1w+DeuVs21LAsBagy9XQWTX/BCdm
WBj9VdWV6sCA2PMZ7DoSBoYjgbWhDbHNY67iF49pDM1V0cUyWua3Z9KIToeRM5o+o6bd1BqQCspb
l+IQbU90FPbPJqwxZe13YOlGpfH+dKUbFAt8vribrwshsAJpnpN/eEgV15wBZKpALWcSK9UFwYJw
JAN78eu46/Dp0WchESAaa2J0n4UgxeNRTpO/bi4Vr6ZJbkKHYDElx8ZFikqZUpg8KCo7mtlxmJft
i/I42cFK3fXt5wvSh58BKZmi4M2EKJ2qx2wMX2GRmXAFjNn4hyuL4jtABGk2DoljMQaeCDr9g4p9
BjAN6dQ/eVIwpS9N8eDAJiTTKDioWeJvww48V8KfAlEjVfSq/zIQ7Isl1gW0tftZXhmEZd1C/DVz
VQnfGA0C7sDqNiCBnn6rNM6r0IvFHicYQsOXTC6C+HaGxpTuSLeEcYsm+vZa7wBqt8bYY10qQKAE
fOVxoaCsoVomeWT1B9gI95jaVBKLPqal31fE4F1qQN19UJrvuQ3lmVcbhd2//pSGIgKBh/q+Slc+
489K/Wv+uT7mCZNFGSDujcP6/fue9WHT39490ou0Bo9jqNMa8vRo0am1KCo5mBgEbPWXRsV3ePLC
HnPNU3V4uhbjqGubksuGDne6ANIIQA1X4whUYwKxGNWX/7Wy3142/Pd7dS7bpEwHjxQl0xVet4bQ
r6F5kCYPlbJIKeUBsl6Ostkpfes4Mq1YC1dU9wi1p2pHBBc3gkugq6MqoEBU3cgIk6w8x8McLvzs
b06S4CzLk1J3eXXBmhtCD5mW72LbIv8lgj6qYq7oeUQr4KrRx1ntgEIn6hMwPf/+M8EVimdQ8LQP
AuAIygP4WmlfDrKRX1G3uxUORJr7dRNrzOmmzPN+GFcVM3dYM+jNu2v5fupv+y5iaW5THgokmxyC
soGfvIVwySZ/WaCIN0Mv5PkX11ojOlJh4tfJOXnOhtXFqoVXgNHZG5K2upmH+ZGVxn24y4uWac1k
uoyMdjkbQmSq3+LL8X1kGVOhCMjsrmIsdb3hhMuA/FtaIEc8m0MndX3OfjAmIWKf/BgTL02AQbJq
xx9BBHTbG2zx/Gh2nBojprLqusnBLd7quF2/3hZ2K8ooZxYOr0dRI/gM0ImGRxMsdFf4h1ImHRTW
SQ8kntrdwdiiVypT39P952ej8AVXvtBsHKfAb7fCQP5QXPRanjniwzD1Whjs3KWDzPVQUshd9+KA
pIay40a7gZt6L7CKSvuVVc4VnC2sO1GnkTw28a0GzXSF85JaRc7XoFxSGNnyQnB9U06AoB1tFmxY
AUy7UWbNZGuvMef5bGKqTLNVqrYjVulPtWvh5MrnN83fwczALR/5l94k8tcChJj0W6StzyBQUsut
NJVutfxzbCFSeIZDyAFdiHZoD37kbkvKxBOfXaexUCJiSCDj+VriCBs5Feb988kwzdVz3CT1d5Lf
vUkVfJvjbOvp5VYfD0qFu26rdvYk359W5NKTY/bKhKpBGKvk868/BomwUGSptai/KfD/LXOTB/UB
mJ2jT59f+VKgMM8nrT42xX33G/Wg3VEdB9hJBcz0UTKpiVZYuMBzrgNsxrUG2gcQt3Uislod0AVo
Ft1OTLeaCnV3djpxxRU0XWX+PZ0mPzobXKo2/B8I4uvRIhxcAb9c/c8Oi44Wc2jBETg7HPwxggZ3
z4NbrUHA/GFT+V8QxgDVdNRVaZTaQGBGRGH0JFXvFHS8EUMzuY+cZv0b8A/gLt9Vkf1S51lEYP9y
MRbYVNzYzePZ5QdQIWFKDyqwnNmDg00CgsOXsVoWnMBB3mb5Ccn181KXcV21pCgluARHEuatMqXh
E1OkG1GuxpHB1O5U5X5s4Sx2eev+CrK2mPRG/ED6o24prm1OYOODsqZSVr5oAX5HTJXiXgoSaZPi
/2OwwJL0ANqVQHvL0kv55xVZP9keOcTyv7zPt1A5Ce4J6pPx7ixXKfddlhCJRlbt4FDo09zIotAX
ue5sI6Wx0To2EaOTNKnDkxd1lToeCkIx/X0g1mCCW18ro1cXiycjKZWjQmRmui5tc8PagyyHBpXF
2hX0C2n9Qm20BAXIgiafBHeLCh/SjHiFrbAYPc4osREwND/daKviSToRbR9CarfxzFhMP7KQASmP
oOPG7mq99/j2Jejq9fIc6lG/iCGTPOhQyVEzdYax2zEBokuWUCKVuwHF315NaqUpS59dTY0iu3qZ
caWhr5YrU243+bUxZPFN/3dAdllKuGx3Sm7softSvfLpVgli2JzL3Latz0cX31JHvjx59K+zaq/V
5fPyNxvjdV5EO9u/RAyiDJDJOBmIQv+l10cSqOgG0z8xwgVsOjUYbRd64SaP1VP7cF5MSyI4imo3
nrjHfF3NEgbGpVOmAUJz++NoljJqHN/EpPQGwDPVBMqIHuspJqDXIV7TZt5azO7yPsxZIxhkdwXh
RjmbFU2KokJhVs7WSkY4LlZ9gZ7nPJ27WNaHNzOlsEpz1nNgkcA2w6SVrAVaNeCk0iabM2zvgvBZ
+0Itw4/XRRRV92MGABqzm05RYH5X38HOWiR4TZQy69BmkA8nNHRw1UPRENBB/NgMggbjpbAxmA7g
+jqPCdjLXGMu/BLfu91bTumTTCSBNh60+Rc5iea5qGVSu8+VO6IhR+2VUs0Zf8Bdh3AZSU+69UR9
v/2VOFjyvlicCMRHRCSh0QTknFbxIdBQ/UgKrumMcLQQfAx1stEC13gvEw0halWE9MXPqPDA0UPX
fmMENWS4F0Mugk/dvu3srXo4tUee5P9tuxFb23+EFrvROk+XyjlDAjfvsgBT5i+WZYRpgLl2sODD
ByNN+S7p+8OCjrcY8sps5gtxLxLj/GgyeIqj7yjDFolJejQs+Zao4kqun+0mCGzCaKUfrZnY16Dr
DA4NlxGAiAOHM/hxwIwoGXexMw4rib+cJkW/XKHXjbaucWuwvr7BtV11gtYeGIjAL9+rQy4aZr91
cZq/ft3vLA75L9iBlIus1GMzXVK4klM5Dzd61+lJNzE+SsGOdmg+h6vt9tT1Q7QqtlBq1Y0OrWzT
8OfsaYwHPLK25SO3hbljJ0lDipyvnJPRrspRX0vZdBqmH0+fyvxIB8MjH3SD9ZwV6SbQymsupRlV
6L5Q06Gzww/0A778bK+OhzC75l73fB0udFVtvcREC6bqfAtHtEqXjWlM77/6CDuJDEQsQqu/DTiC
QOeYqVwBvgm+dCftqME8QoY7rEQR0I5h1PFa/jJepWrKdGvCXPBfakB0J76hIYK5qw4aYGUPWAYg
GiL4ofQ5vc7irEdXAXRqabMvooyf2MuTNsqutpGZ/agkbPyTdKJpeThtezRTKVqbgs/CDLw78zcW
2+P/oinYIdet0ko669Oglpw3BdiobyYHD9DsS7e0rcxobBOKEYTRdPZf0JyxLdt35+l4CZ9ibvPm
qEY3z6GvCvbdOJxxP37i8NR+ImtFOskoXEB0GrIQt6DGSCORHhb/NKZ4uxdX+y5dpnPd4uw7PCbC
/0g9WUvlaY73z9VhaM41skC28WW6QBx6hTUW+PDqIQiUO+unIf5ONtl6wpPzn/e78JA6E5a0kJI0
Rx5CV++WahIU18SsLk6nOeBeUdZDCfplflNjwuKLtyeU5tQGc7vgMUkyRDUCFyGQMYWyRIIHRV7v
YIPeFllFiXHUa8kNvLkcgJFE0lBHk3F0kRukG6ygP0n3wfEMmz+yRak9/d0e0yvbUy69OI5je++d
+x60qxlT1Clvxx3LO8TUuaiwLxhjPgFf06JvTRjzLAMKjb2kU02UCMoNMVVq+e9wbxKT1lLEYpXZ
bqruZ50CX68iP51Ox6A4KZ0sBQ3J3Lp6sM3sLwX3/VpSo4SD6132vGQRWGWurbkevOUsKjvRCiwj
Sa0EnSlJ+fsk67G9/GjCkMslAIatwWwt1nadO1MsLDbAO9DW7DA1c+0Qabmb9ZWOAvgmZgiYAp2s
PnjGe50thyaBZq8PDMD14II789V/1Mgn4fnIlE5xDh5nxkwNVmT5v9COsJucJp0IwVUds0raEpek
XKsAGizMTNGhoH+o63gwcyA1fV5+sB42dzzS50Xp3ZaUXq4E/wQ/QfTJ9uNP0s6qPxy16bh0y65I
8zbSF1FYo75Hwb7XHpUZCEcYkQk2nbaXeCs48S2BXkK0bjsYpybz0Y0cZZLSh2DVXvaaQl41Utlu
AeyxBsRJpzntAl2XIAyvmwGwR3yqK/Zd5AMP1m+xUbRdVs2tI+g5mS/qH9i4tmXWO4kTMo7CGdBx
VSCLVJtOWK9cRU7TjGrnW3/CRLVueAQfGBxkDMMHGqPTlBin0DMcG2y9HnNh1rY833YLUq7nOPEQ
9fMJJ/xHvVFER0z19+J24RyvIQz+maJKecRlawcrP46DiJeP/QbD+vEB3C/AfJ288D8D1ZGuW5XT
HAdyC/3pQcp46dXmum9/P/mCmi+VuhL7VP6zozz19sgnSCcpD62uKRqDIK2o0J54yF0UOFBMEJu9
bM5u9bTiqtmfs+7OX+2G0bGL3NG1Uds2OQPXgsViTqs11Rvak+grhzmYkWM97GMmRfp/paERrnVi
6XV0oet4ShsP2H73a6bY7K5lQ1m3WXpD91BjO2D/bvmBOTPr9g6yfjjIIBD0BCdtHKOPYnYQHIS9
OssfOz3muTXtAYNK74ht6Kdyt++tV7HfypPJzt0OPANhziRnS3PnnbUbgM4TzQg8T9WQ0NNvxbhy
Xds+QYKnJvwFVvlJgTLNxm+xFt+uIJr3x7jAJ2f+xLMTUSuogn+gy7d9JuI68En/eQN3kaE6L5Dw
59QAs4Jeuu72LORPfawXQhK8Yha63U34ajOE8DMyIoXW0QrL7CaBJz2lsjifUGps46IvUGYhWZNh
stjdvjz3vfIf4KxARJf/xZM4WaKPlO4Uf+0EHz+bP8N4QK5V5/BffSbUxu2BctnvfA6J8ky/n17d
ihMmct6wVt2hV1NyYekX8gqpj3lVltQ2Mupc4Mfhi2CKCmPIJNesC5cEGGLLLjmweVa6tcVHk0Y6
qdGc/sRHvGrH6doipx0B9ouAnuKbpjLHMs4WQ5dpEXvGwCaMibTslPnqQHC80hOZ4OIDM2RoAHnu
nDA6Gzv9ZCcpzUrVg5Jsi4w57phuU0JbXTQLKP1CLWnCFWkGFUa949bS/gYKf4VttgqHFdwrvGI4
lSnKewHAW2BSCxEt4EeV44SfQV/ia6HBAs9pJrkaV2AfMKCfVQ6XDLSVMjBeJGC0GfPqmnYjem+s
imNgAvux+Rb6mM+OWddM7zpak0oAcyGlItO6/g0JHRWELA3PhJ3Z2w07hrDo+34CdR+/H9uVxSiL
WSSY8ViZzOrPKoVY6nYgpNEKrOhWv5a7RkSaZ7u0xfTO6z25kXTBe8vHiKU25LY/raxG9IrY6olh
VaeUIGexKGgWdksphLkfdSrIhMkKJjx+BFIv+D96/2pf7scFPBSmHVVfqiQyI8wTBz+03buUo5s0
PpZLWG3hEnLIpcwGpPOigWGXsy3JFhm0PlWJ0IJTfKL43Aay3cidR8km6hIfcGEYUyNI0kYXKE5J
WprsUxXITsQSNme54nCPivm+aDSZXyY7wwSeeOh8fznRoOxtc6uSoolwceyvpDFZPR96gnfdG8ra
s18u8LnR1rNA34TB/ZjN4hwT8yrho3qCxSRBbLUyDWET1BUi2A/lUQFU33M6yWd6g2PFnRNQIMUu
rwq6i1G6dchXbfPaCaqLP3AK75fDNLoRoO/Axl5Vw6vu6BEmTAKEaOox/vWPvnJzs+xYPPwOq1o6
Inea80LWpsYwZ3ve4vRgfr/8F+MlaIomCgN5YZnghHevk3MNQoc+GW7nvQQyHVbeLRYAioaLIWDm
hT9n2wpjqvZXaMy66Cazz/q9PoAYfxD0tfCB4Z734XcrhlfFep40hpFJsOwQgj+H/KFoMRUAugX3
0TBftBg9AEbhHdGZXtKwnJGifPuGXPV8ufrVzZ4HJ1Ntzm/hJBBf6dzMhxDnypRXxs26KRXX6YYn
Zq3ioWn6wAYqEPloHtCdhEHj5hq2jCHqqNWu7sPNHjwIBLdLQJrBk7kJ9ks3YTn3/KV0QbWlKzwH
udzq+lzdhgEed9re8MeJ2CGLv5jIFVrR5Jgd4de9GQfWbkVP6LU5C9cruHtB95m9ultoLQtsDdgZ
SiI1s1h6YIarBXWZ6HU8yThysBWGq/0lcbWOT1uMCTvUaMRbw2VvwezZ/wuM2+AI4zp8SclmSHUp
n25GoF/66OvoDf0md8H8yxI/DH4Gy187KMp9JYA7TYSezIIaZeb4Ej1bhVM6wTvPe23xlEUH5Oeb
Kh9VEPZK5WYD4m7aXhEO/REWemV+cNCjkagqxyXhl0ElYTvpHvRQy719w10BNdcxjpN0ZjUQXoHs
22S3V5LtIv8K+wzROuK2eFPRGbzbhn8zJQHp+V5myucrrInW4Jj7yz+Ag759ugucADTUc1wj2Szf
3fJd4hyUjEWt4JTKdIuGwbzxzJHQZBHmErCcsI+lJYCXDBnew8w4o/bCii63nzSKEoRpju5Z0hUZ
Q+R0ZySIHdMTv8S/QA2Co1ZJsJG2mNTCEyT4V9If7OdSijdu2l9PtDC/IeR1j5tr3c4YkB3sba0i
w79JDt02A9/YG9IxeTjUxkc8QfIVFDF77rBHXE5nTvnKtE63VzHUccv7xdOLOrrAGTQzkze22pel
RaOucFjdxUWMaCsfCkRUZfFIQII9eVidSgS7ivRZHLdKmQfk959YGAH4KuBFHGvOkJs7mjwvR4XC
Wtt9QQfXjy/dWF1nXIPxhRDxTednFlk2WUxquike8LHZq13P9SlGcfTHYWcP7NBZ9FkXlyMHwmdL
SVMVbHI+Znzr0JPMM9jMkU1KBVFFpsmvSV+LagFXvx8dtNiAV2GcQ8XfJMGE/b0buQwdLWs7C7gj
JGw7IOLEDlUYYDWHBDPtprE9qPwmtfyC6W0yXBr2bKYGxuFofCFv9jPjEZRc1EZsGZjmadgFH9CF
vecPaxaQybk4XDJvEegKD9UXisNYJwtGklYFZSNF6OXvg4y01E146yB6RDIihYM5rU/eHWaPBrhw
iaqFCi4UgITVD9RFARZQrEPA0lT89dTVLoO1g/hZTiXftDw9nh3HSujTvE+pQO4ciyA8gDcdSdG9
1rjtX7zTN2c9VT3/CsBmPPpmHyNcJTXcUGhgCHfQWkcicZxE3CPvCoDJd9Qlr8noayALbXEizxt+
yuScJOYc2owpy3QPN7CmbWAOIubeJh61BUF/45Chv/m0NVHdGfyk8SlXYsEziXlFTm60rHGihnXC
OZ7SiRyQpcz+pu5TSfpObZk6/UJEBgZ3YDzAUbEIhTPhwC5um0d4Une2zG9loY33/6w28eY8qJqw
h0cDQCBKx/DAdqUu/muDNHM84nRNwmTlOIPmxRTrocoTvtT9eXFfi4n2BkyVthYS8hFb52oHSftZ
4ag8AejxUCTL8PrRIxtORfsKrpXCfazFh/UdwGc8aCM9bPxjh8aY8axCOI+Eg8W9dzrbDWjscMjK
MepwikvxVy/12Vkj9HRcmx22vkahwnnYgTYwU7HQwbvhLznxsfjEnKR2rkOQT3AxLtuiz/bIIJcF
xakSHu10EcZ52uOk02e+4EK7XWgJdC8l1jp9SZH6o/J5IeyL4RohmJBwG5cKakcGSD8BUCXvXv7W
O+lbPf2US1pY5lEo5oYQ2BI2Cdxxuaks2WdmRiMqFI40hLmCZfdBYVImP4ElxT0ocl6YTyCpxsSD
JSMlCnOD+/2SKZkU4fLazyRtG66bE2JWkZ0F/3KF/Kxc2YKARsKdBHGB1kBcF47+mwl8tkkvINlz
TXSiPcQU8DHqCpDsLuICEVUoESWI9O3753npF/Y0bPr00gWkrEWahf5gh82kSh20qWPkyGGisGOg
a3h6GC1UxheZ1s+JguwqogiYrSnS+rwUp/eoo/CUCvfDbl32ETZwu1CbamidyjfQd1Tn4RN/YolF
jbJFPH6khu8aWbZfWTh7QHATUaO5r6rgHMvWdah/fbv61BWRzvH9idaGcKSdqVXXYRul5+fSnv79
Qi1XotsC88ekLzm4UI487Xm4rMDIEdHFAhyP/osNRpjlnlXTXl+1a8R+mQVg43Ui9BLpVTq8cVYj
Y/+yebG1IVPC51oPNXcDZz6KJfHpvdiqglytESnl55k1DoKB7wi5/bVUDWg+Va0EMUlH7WKUrrye
UgRo7xMWH9G0TH+h3EVHLywsgB/vxc8jrlIPe8SVA5VWpPCyg/dzOaCYpa+V/SmIlD8rQBm79gge
LOu0+4/Rsg2W/aE4xxQ6qg16kLMBPfcJsNG5UdSFzFtP9rwHeqsEmFz9pDtnYsQUQFnGpBw6Yb95
UKbkvwOqv0cDZNpyeHImQxdz0naIB2lMihbHQpySBRtsvZnmxNS0ygYDb6KHXED3upU5grtwLU4g
X+ZsgRy9wE1Sy+kqXXKqN7f9U6AHzRlL0SYocWJ38rWvV8cM9S0F67zFWD9JNWF1IipVg+cprD7W
HdM4X/5c8JKkwQNfcRfXCmb98d2ppvc4zEXiG4eyWMrhf4Pk3t3NtATJKVrufxiKEvWHgLdCg9/I
SkQgBB+QDnLn4oZlAFqUtLFvNgsCHbTqPfLRXn49UCYmID1nt6dyubeJoqHsjmzp78XCR6vvYzwU
/uwpCLnLhQBYvzDjuVgfuji+GBR2MypkIhUFU9QJVFXypbtKrh1YvgN0e3iqZy37JkaZxHWeedDs
4OQSGTH4Ty2cC9TS8Pugmz9z1I1pJtFKDzA22O3LxdUJmWT8We1uP9s3iUTv9DQiHBnNhyJ4YGLm
gnDiCFnNBbPWOeIWiTiZs6gEF3372jUsZeRrEgh1BdqYm3oVFASRjioZGnWe9QFUSbUMYYBGlYr6
KeVbHJ+VgCcOzelIZ3Tc0ECg6m8HjM/rvKr2BRjqJ8TAeFO+3gVffRa/4NZ1Rpf/1GSl6YDO9CxY
AYIydsW2U+G0HjAvkfngl2Oh4WU0ef6fQDzXsDCIdBsavu8dCR/C6rMM3zAaCX/jJkGlWNlTLQS7
0qmb5ZtETEbjUyq3n0zTuSZLGqW9ECXokHDNhYnRd0Mvz+yf4AxkFA5r0AeaD1lPT7egwaiRbYe5
xU6KjeRBq7U9KQ9pspzB6JvjG9Sp7c6bqqEweRkZJE2OHEzST7VfkMDxVn43eu71knNmxSNjnZNL
Z3E+CeG+TwHsa86NQeT+xRkP3LtdEDFQvw2BjnUEzo3IrOUPqfF5hba9n+8Pr8RoI795BxRhChSy
uNH/++U3CTtpQtmB0d8jprWgaTuNgWMjjdqWEIkcxr3IWhArykaRPFQeG6J5FckRgKcYdGqdUg2W
jiqmKrkCd4uCn75aPDhFV2mupH3pQCQonlarASksOBzXhjp8B0FFdusQR9llKoallZVB1/9lDVhs
bxNV8xYff3Ylls/9CHj8w00Tu2J7kQ6lfDXQt4QVcyAgXOc1os7+Qg3LMoJiFBThVGqDfzNd9iwq
vH4v9lr3jhLK0GPZVbDkd+brBczDElmrJl+EaOprOML2hQNptOUaickyxVU5nq2vHCdPvnsiie5L
24WgBbWALLfEOzx5xq02+0ZpEmzUZ2dkjyROmip0wK1eWlE2xkKMnynZlEiileSGVaUcSREaKBlB
KD8aQyYEPDM8UQ7YbxgnspSh8mOVe6x9bzxK/Kaf3U6FEJxIDC6rVfwDtiQ/m0nUwWAk3cvzQ8nO
7M5Yg9cgtinBmOM6iUVh4Gc2bpjWW14+KPHX9V+F2V8LaBe2nNoZJkeUD6n1lnJ+wWswnY8A9IH9
kXHWZjLQXXTGcLtvLti9su+2GnP73/2mF7hf4lk4nrVajnnxZaS4gHUdjY1Bi/byGYWx0Sg+Ztme
3cWMNX7PCGBOTtt3BYhe68V+HLHu74gUuvGX3pFyi1zSl2hkaHSNaGOh2ioLglilHjUF7YyopMWB
xYg/KfzGpgHX/TYzjZbp9Y2CcwUIi8eNL/cbo96djPA063usBnjvjmpD42eXyX6BaaCjjO6FRY8/
e0I+kMlnzV/cvTAasBkrtz60FYhkv8jfdBGwTw2awY0s1dqzeuYPZmDEXj4hFS8j6cFyu1TecaDP
5lqo3z1cvAa5uiDcZF9kqAmmCwYpH3fTsB+8liNP5PrTsbD1MmAo0DYsGd6byfkXAgpntjZNhpnE
LO/birELZP2ukic3NiwCDbaQvkqDBRZmPP9Mq5LGjvDt8ncJJvcWWnDQQOXvUPmjeIeDxYazXSu/
h/xUbEbB+obdwM02VHinfSFAfJ/Sn5gWP4sTMPjiTbN1g5xqaUFFuCFpky1qyO6oZHFHkQl9pSPS
OSUmDi48ZGe33IkW9m8MnVydPrx0C8e+eF7cOvsZwiEE1XeX+AbEqS+h/V0w1E3AdkOvLHeB6/rC
mzDLMyPWyZ+FLV7KpAgkxgDgMTUw4eziKDgZ44cQmVOCk+Ee4KiWcWf6d1nsGM0OMa/9/fVjsyi9
3NP3TzDCogDE3eXnEke0jMuoU+Ys2088+bMWospMVE5gUuFgaUXq1G8s/40UP08yZGqh3kf+K272
ET9Uaa6zkTNrhcWOepeuk6u4rvHES5tkPi1TA7+kPkgXwtuF6XGKrLLYHiUDOexUG6HmGlkRyw+X
XV68F26ED6s8HQ43tXexmu40cOvnKvDm+Wu/hLT4DRBRpYMI6e9pDNVJolaxhB6BVR1ukPQWEMuU
Fk79SJGqAaxRjp5ZCw7l3m187uAIWK35Nx8YIwGlZsK+gjmw2uzHt3IOinD/y7TK6AwOven4Aesr
Mgkf/RD4v/r8YJP/Dt3yy3BlvIiQZuBfGCKDiYeSPGiLcZOl7NjKJ4hjVPVNoSLnDtZRra4MCw+P
+3hFOyyjSaSKAP9FHttj7SQuZvv8P46YBcIB1FtqRx1cg/A4jxVLgp9m8NjSr+2v+GNLEuMNzNEu
Q8EK8EiuaU0I58DoDwFNtT/3h3qol7bmDSrXnFdDeiBVfLcEAhSm0IdAaQmxWTCoM5mRbiIdw7xf
wqkYP8GmMymif1J51iWhVX/uKIFFQx1AxBzGM+hh4d/jKa1fnkahY2FMLgBVhZvUv4zK/1nNpNOv
la6Z//vpsDK6PBJ2ZwL3KbCcGQGAYlXwnxC15Y4oUOnUr1/90gJhK6yfRMBg5rhKIvIouVxADQ2p
sI6nPW5VNFOEPbeSEv3bX4ZOSpa5JFhRIX3fPt0DXOOzqBmImUJtv9ft87gojYM5iCCDUXA+r0Zu
yC6McG854jIiUsxgi4jbTgl9qJtfBiTGnZRfB5qUpzVlXOD7vw2a5I3VW527wGih/uvlB7e7doJB
fYV9N3CHSBH0Su9OS0XezFefNKXG4WuusIt45ksDTBRpzpWhxCZKO9hxa32UtaMI4j8VlXU0Y9Hf
qsDYAgQfkuMYDRb7uTLIpdXnJggkg8BTzCSRPfEcUgkBSDrwHkMy+AcCgb8skN3xPZaGyvpFtLnc
Rcabl2tlUCrWj8HgVHTItjQS1luMm0TSfD6+QZ481xAr6d8fBAAuaBVgaop8KcWvEn1aClK9A74l
EOh7Kx0X9bOHlyrtzq/Bab2uK4TaG7qNCB1Q1AuDF3Oo3fT5anbZQowfx/MeDY/t7ESM1jnhE2PM
vv4cgsh0tLI7uS+B6SjGGM6xWkvrSxSO2AHydFmSXUNn1/t5PnWGVo+gIuecv6q7jemiZcWOew+Q
DBUWMsNhTKhHbljQdQefy05OsSe8veDn1L82hzwoUYfBOJJPoDcUjrCPipw9Em7z731vilms1HoG
bzQ/MHG7KaRtE7jmy//z3yrNbdMje7opYhaORk3PLRY+dXZGccMVM2ANH61USRdXnzP0xcZ9GtJe
Cgb0dglpsThrfhQIf5WAyvTUCjpBsXsKX9ZOn0z+l6Yas743iihhZ6J+wUuWk0j4GTD0SDvDBtaD
fy6SF3UH7iuC3QOob4vx8dF0jUw9KSf9PYNBCmsZkluqpvrlSW7BG8DHzakknXrjvJwwx1zcHXgo
lturyGJFaYTFI5vbXnB9n8zfzH/BFBDBk2w2pMBjYxoKCdtX2mRpQ6eP/WRwgNKPnECZjt+mm09z
7HiEsFLeXFFDWARkP23Wi5A1lLyGicFQWPEDZ70nyHqAeTL77AMeLaRIs0UHnlBbYFccDsqYyTCo
L09RqtRSRy7nyHcZNi4LW7T3T+TXI0F+0s5IdBArNGO2wl/Obd5diruouyT5KdOE5WVIXLgic9eS
B9zGWA3IU2ykbYwEUCRwft9P6O0RgBWwvFWIjWaLsV+ZZ685Sxe3idXbUD0llpUrP1Fsd3atJZ6N
YIgL/NqzIf5cqLHfrBXF2oLcIT42QaN+hCWzjmL8APPZa+BbEf+4teBu3iKTvj6IC9WW//T2XXyR
8Fd89YCKgrnUmUeriDJbl15I+A5PdUz41RaMxB9FwGheT3DtjNcdUwyGs4Xf4xYfuqjRIQD/8idg
eUMLdvyszt9O00h99OwgFNdSqKbMCAD3nwLf+X6IxQDsMzzQcT4aRvvFqhToPjX1+4up+uumqqdW
g7+vLMj6Gi2Is1mCmlGBfebFirRgd9PiMk5SZf9R1Kdz538xRFRcWg18YrTtff4XZe0j7dCDDA7B
GavCgMrZGBsGziVxeszNyg52iBhcJAOJnJjEdGjUBark1aaK+4WdSOXyNdoZ39raS5Shr1yY1kyz
QkJosvzdu9AmxnlMGH6BfWl4JmDn8SO2KQSSHBszxSM1hqoENNJZlo+iGPLnZWO9M6+wYena1C42
k0s9Oyh7yyoMXe2eLr2pOTVcen9AVLViyyGvNkhWTNze7CCHp6tD5+fHOa2plWzvB7KKV1fq3KF1
QGGHHnZkmQKTTk2VUbYY2QGAvYDPeBdy3XLVUiFbog/6LccZPSuw4quuUPumq30c7yHFk3SLJ0y0
jR3ZJbRoCz8iQW2i/l4rRt3ANmNKS1G7wmy9HyWHvTofAKDVVy5YDQmqIqI/ngA8sRppwdUFcfuD
ETIABeX9o8nydIn0xO1UntOrhuMWtpjhQTHM/HCfPz4iBNbfdlYL7huSe1E2Yr0nNIu4+hNIraOS
3R5tdhUBaEZG5wmPe9PTgLV7ktaP9XxeTw5DUBBcuASJfCoAv3kq024r4PMYVhhr+kIz7fWdR/dp
mCdBshgzDG90sgHBxaYu6Sj+NAKdfo4cvFGl08+FleHcsvkPUowVYyjtuX8X0lLAscqfSYQG/Ckg
yTCzAqV+T2mBnXxa0pCi0qzItSJFqx1Q5UmCQxrIHrFzO2x4LbK3T1oxSST1IfuJRzdCZRg3WjfW
5TDJ0PfgPe/4wqCFv8OmVJLhwz0l03QmU308C7KSX3kVAXIGaOHZ7c7lgIWmVMK8shft/CgM1dwT
/k8aEiOTPhjDZTOE0zcXvdesvI74g0G+5/qDTrCFuEJj4qMLEyGnRQ7XPIynREzveMhnPS2T2z6D
xD96s2233nK2BJJzsnz2FteMmyC4oLopFiGyhOdiyWQMGy0qzXPvt524WGIQcTKYGkzrt4ouDs96
ezkOnwt5tmqHb2/CzwVsOq1fd9ypId+526L4eeMLOYsWGV6gr/p5Br3iDZdAch0kaT00oHO9eBod
k0LRWCPRya1YZSRygjW3C5U+keUIB70BSTaLfmAOHHzzNjiPHPbBow+ttL6+pxKvP/SWKUx3rBcF
X7lug/oILpEX3z+zmLLo5yd3AAvt//MY1LzixrDJBS2E7Pe9/CIdsGd4XzKqsQI6p4hS0Yf/YUm7
w6xrIqoTrDpNGs7Y7zN0GOTTl23BCbce9EHIUc9l7jVnJ7tT7MC0wkMRZadkpPvxMzWLZSaCiqTE
Fegl4CBGrMNwJA4/iIB7eeqNt2Mk+hbfoWdMdNlHIQlIyMOPlMUdZ/RmstIcqLiRcWhGwpM/nlHf
hF5ca332tgaNkLLOWX+ppUh1rzvdZNlHoaCWh4B9ASsik127g4zaaI0897FkkhPdIWqU1SYQMSfU
uW25kbd7tKQDX+LAy6CtDGP1d5qIGmAFyMFbtQKP/yN8GXNMKe81q5u9BWZjpXNuViAldieYuJuv
iG0llT4wnX9vYndC5xsGalkgIHe0yALoopIatwc4B3LDFz3ZXMMGcJiHNq96iiYI+BYXcG0PhtnR
JA5HQhCYfL2yCF1WedNHxSm0nKe4N1o/SGicTVmwKorocff8DJIstpENQrDzkpcy4JBwf8IXvjGj
LYCirLagciX6jYqvI8zAQAWjYhht9yC8M0sRhEAYrKM1xiUJChY+7uWy6pxJ+/bp6NsUsna3d4nM
H+n6v16volhRmfL9/5bxwufme3fBZAUCS9VRJnXpGctvO5XBeZ6vBkAHmP2WrsMdvU2tkiN91Q3j
7OCiHvnthHAEG3y/pC5yf5aTDwTY4SLt79B7YoOO8r2QFXYvAXbEBrFDcu8fd2pMorD+hwuE6YY2
uaI3BtyNeu09xDlC5UU5qfsDeSj4uRydy8E2EI3Pqxhv/l3SsgALy8kUoPlG6GdhvoyNxaZRAPME
ssMyszgl3fL+JLh3KCJHghPsUWGGcEW1+aZgXyWQT/BnRrHFAjmUMkhBsfiYgLctaZWbGGPWXWjS
VjykJgtQwHzHdgONfKy2pYAaOI6xeCx2mH0Ekz3pnLyGxRf+U05h8uvGuwo97l9Y0ECXx/+SXeO7
3+MGH7wNKMxCyW9XbCq68cLxEg+SYZpnV7T79LFRou5CHPMk04vYE9Ysh9vIjkkI1GjqT8vZFjfJ
R7NA7t+HB12qJJ50Iy8fcyd/CR4zb0ezCD4UX0TQufiaiw0XddHx4zBpcPVqHM6ZybKmasI72K/l
Ks5IkQfjFFFh7Lv4zDBkpIgU5v97DUX3mJQYP6ZHqirsw/GCzcCScFZLJtobLYRQLuYH+9B6a64E
gLhofVU82+UQilea0KgtKzmZewNK7ZA8gjngQ9SI6oX4/Gk9iim1OA2sHkAKA+PFcleiujpOF88n
OBTKqAkUiA1OH38Hk9Q/og251kQZWDuBXPvpTm9+bszQrQStIor5lh2kXx0VYYXwVJCji3IZA+YG
PQ+kh8cR4WAgOLsBXJe6si70eE4hrs8WDRQqZzdZa3AwlSZRn7wULIwI+AXZU2JC081rXFAZhkqv
cXcwQheVDZU48GqgQsvtZibzhzX5EbfAIqsrnomezsdQGbLJrv+n+B7Qtev/kk46Hg9KZPmSXhbA
5bA8c2eoV5ytXJk1kKn7PNVdUIyw2YNlRAzoB1tPK3d3YP9CVKJM96WLSnn/ZWLUtNA90r/VK2gT
348Q5kHmG2qxAqB9fe6AMCPZsh5tdyiZGPaodq+eWBZnkczfOfyNPHZMUycMSnEKlhKBBPMQCEhd
Ta52+S1Qyx37oQAz9nTCzNZWJ2UFltLNkX3RGZg/eCqtJiHOxCra5adxicbJZ/Qd/es2+ciMpeJ4
OK4gbhwgr4jV/HOfi6IzWS7vuVZGqpbqD32coEc2HmM6fTTgZPmhVfdd5+E40x43mDDNNtbwbP4l
4cOhXvkvc6xCFU0GRUziC1dlqxI0BK3dRzfjsD9k8cM5aWkHdrNtVaQ2aBzZ2zoho3mZilu7b6ym
sosm64Z8AkF0uZt8lEVg6G4nL032HuwvF5twenvcjlsbEYaGjuZkZ9p/OGEmPmWU7fW6B4Pwvfjx
H9Q4zNQs1UrFl5Xj8LK24BtGi3UFJ9+L/6xaIh3yZskS2q35UzxGllAqVTfDfdPsHSgI7/WrBuWl
wbz33H9I5fDX767hQsu+c8Zt/UjVIAPqTqkr6Aj6K6b5YGCUiWyEHKA5IEJgyQkVtvvUN2/jZvxl
Cpc8zT17+CXfXwjyue676B8mIYEFtNGOpI5cSME/jpeuKZ3TlJeo9p6lWCJWOOP+5hGFgK+WN6F4
1o8vG5LGR3vQD7GV4ctU+jrhF1EhsQuF40iY4H5kmr9km1rv2ABM0P/7DB2hqtRkw0rA/ewwNawd
4T9Eg7UFzKVF4qqcKe0wMmk2icHrEuE80s6uvr5M/+Mrt1olU3N46Fb/beIr1TNzyDhXMF4CWaHp
y85lnZGkXU4NJO2qg0PicPasCh/RWiRw+KkPecuyHN7VgpUmUqmmtYFmMooAYexaj/ZHy6TQYrcP
NfhWe9WasnclISvZ00jOJLTbMlupPIE7THk2gLNYfCmMrAvA5N5TwC6GEZWA1NL6jtHQhDLDIKpo
uAo6uujRgij4urHgVyovHJSZI08CnDZFf0aN916wivJApjxJgvBQkIkDAcS8oa3lLN2Fn+IivWS9
SWJEs6C/xyh2isZDaKRl5UJSm05sXj/62n5YkPfR7fPRyqZkJ4exq6d16RXET31w5qMAgO4JmvmJ
mzVl5WBp8HHk1PUU1iB2WKn4NFvbbN0vKlBtlrNDdxtlKYVmZINHZnicehQj38rmBCYh2u9KsiQG
ENPvUtKEp3z8ZmDLEKzbXQabGiHCwodNAFIVKUz1tB1tKQbJAcMUPPUrH9ua4nkAGMl8mzVfpPRo
3nMktmjZRu265EJK/48IaBZQAV6X4QXZXacSDkOI4Vw/FGv0ac1FTAs5GUUk/3/Tjapp9/Ys2Eo8
OVz2rtbXC1Dq1Fd0GWXK2CIosKivHfyX1qlczo0dK1tor/OWzA3xRT2wi6azyyjGq9TlNImVxIS0
OxizMynyx5DZShFS1K4H4Up17+IPrrYm3s1VOiIZGXKGCW4uTRtIwB/Vk7cDewZsMBs+rhuz8lOK
n5A7Xl4BFqpLXqPxUI1UrGLyr9BKmAdVfCEPFhqpERF3Ab/ofdV6Wto5roq2QxZZphb+A0Fd9GO3
FplHyLH3ca6nTXqagRZExxEjrByPWXtSFSskGwV6OQust/Sod/qPFrjRrORKfoebfoJayHkPjpkn
oQ+rZdE81srVH1OH/L5Re+jKqdZw90rdLwNtKoQdcpKJ7Z5SrLvCyuJoFmYOPE+XbolJJsmPN7pk
Pd4Sdnna8OshM1baX6s+M/uXb03YCi64AIt1we12FQ5Hy6dg5+CycJwtU9ZUME/mHcZdf8g0cw7D
jgnQszcxP1ZPVRKY/3eIAcYQcYZBmMLxJwxvObSBjxOu9hrkbM1NarrcWPcw5I7RyCPgRts+mhUk
3GquCJgSDdjHYWmLH/BXL+NdeTzMD7g8KLKXj/ous8eYgMzeQCDDOpZRW1db7ONT2/qUXyO4wU1z
0wCPTvTm8ZFY+NBVNQShMuX65xEIfsRKXpT0I0uBiOK2bXV5m3Cu0hoTu+ZjMzz+9eZoht/VwQJJ
jI4tsGHKUccluUZEsRD9AtTjTSwJzfCqsXNudCK4nHuIiqn73bnlNjVF2Cg1hSpB+lf7Mk9oXnbf
XbXI0mMrgPQwweuYztjPR4gLGVQjIte/IlrPArx2dgF0M0krZ3FnuA113nY5I/cFNoUy+DJLjaJw
qNcDPdX7j9hHu7Z1PO2UnZmC8M75WH2iouNLaBiuEc5RGsWZm/Yxf31a4jLDqaG1HSSO5YwK58xK
gO74nB8slCo4sZvRCO2Pk/RKPGDqoFwQWCLKJY3LpXphvRkZfVss0BT9NR42ymagiycEu86Bw2xR
pwTEzmbt17Smxj3lbeQz04N4vYN/B+pqOlXZuvA9opepA5uLfDBq51r6Ps8Ne9hFvVYYhK3lqTr7
XCIut1vYiimcVj3pqDwvsNr9ROg/jEMpT0HeYo/tC3YoegsZxJzDSrDfaKrdZbf6grgGZOzlAs3Q
ncyD9cT6qUc3Q3AOtk6ssPjrkhRjSfXnLMboqdOvfU6RssMi3fuNMWUrwsiPOfKwejN9WqGwZr/G
WspmXDylX7sxK4srtFP0ppX3wHvcBZXuPAhlZS4uGAMq3btfE7tNw6lScQNlazACdsFy3zfpIXiX
pshCuBjyC967/q9Vubefgsp1HjZIDsvCQQ6toTuwqoAdcrWsJ3qor80KeJzv0o1S/hwSzr+Php6h
FmEtOfe8e9ZbV9DdkImAN5lMfurQhcLr4INTXS7fJEP3k9LlZ+xDNoKDzSW5FGd11zIeQ8589ZSD
4+11m5dXUo/HxN8b2qKxHGNBVCAteJOvUHlQIRcdIeSnUKzm0TQnAaGF+lVBIosOh9vXLZFMKart
b36bQ+WDHlWoam3Rpyym8nSaJSt2uel/JcY/6pvfx2EeVqFS0s2uum64/vP+D+mnHnseOQ4DKEJu
43GpW3Yz9OJxjq72BBiPBjxfsNi8r6G3t2+8YPFdn/RVg6HIh7KYaGALvIaIrJ7ydKwRyJ0tD61H
cgZLsNduyU9CFWYe7qJEi/xeMSKZ3qvrxQYcsKIHMWi8XgI8RN9vBlJGuFnZg5qWRiODVFQmKGRH
xqIEq1i6jH/1xNXCLRmEShX7JQihu0hWJJJbKkargQ2ddxHXB2hpXP/7bGQ/HevanfotSd/Vfo77
TKyJOl4N7LhoZkt2frjWnHb6JX4STRUHDnk3Vfa7c68UWudDFSapFYAxd3RkXR4bR83O4257kmEQ
wobeigy8Keq6S/GwxdHNk6ghWaeBFkZlx4ktck3bxVezF7+9Y0eXTuEgtiV7yNlcJY4dux7JgYK8
JKaPgZSNEaMs0jVHQ88UIbj2DhQt7IxGkDp/Yltg2C3KUaVBTsJAMk/dZ+LrE61s0U7jjC8Uar3t
Fik1ryPvfRL4n2rsSq959WZj3TA/9DaI+/B/1T5Z6ph0BpKzT4SFpn1W9kvXc2oAlF676BhYIVd5
oolNFBQLjMU14hjBdSQkZ2S0SGAyadpaGI6L9VVV8O3ClzKxvtuyaakeY0avayj8zdRq/pnURS3H
BmsX22A8d/FqJKcJN9xL8ft12/lhKY20uRP0PEDI8ywhYlrtct1LHYMwhmtfFRpA9BLP6wHJcJE6
FGp+8KtmA/oFUdVIPdopCBbMA5w0t040zPjKOKkhnAEiRYXFuFtXECQe0Hs09UuVl6xHPISwqeSw
kzBAG9GZNTLk/vObdVp4STxo6Vq4TEOWCxEFyFjJvls5E8jD/kuJ1nUkC992SjsoNVF30grB1+ee
M5SHNNohmmmudik3TznGIvhYHxZX7JRSZydUWbvnWubSR2QiT3gEkjIlWrzDHVArly5Gg7LCLrPN
eGoQwXztkjfCZ/NMCcIGEyWSkYowfQLebT8fk2rGRLDzq3XyeWFxTD4/JjWyX4YLO0oPv6wi1hqI
Sc/0a/I2d8IBa6+9UajW+ZVCGgSCGi0BAV1VsvLskcAY4EFBpL2oXeKrxt8itZnUfuoMItrqF1dz
tYnD2x784O9DMPITw2q8jRBu1qAtm+t7rT+E33HX2AG0WzCrZKbnU+PfJy4HzNBXJ3L7Ba6gI8tJ
u+90Uc2WY36v4HihjDiKwyYwbltebc8LMcrlqh9DEKcQubS1qW5WZiPcLsR2CvGSyNwk6ywswJW2
xddPKim0ncVgxgJIZhoH24P2aiwrkT5zdSdUgeMD7xWxZWES/1TkzAdi7LD4TnVkVyq1PFkkQuYq
h7WcY3kjBy1A4d9D677wubyDD9/saJeqhIek5axIIHzTCjWeB1ahuby3qaXgHU17xCEqZ1zQEq4L
iu8xkbd4FdrOAe0jfM57v6nlL3fR2oTD6uTeWBFgntR9NcMDU2cugTDo6741ZhgPWVygyz2v9Kbb
PebcQ68dULpCHeONAG3gqHJyTm7Oqwu1faULWKssY4kuQDgK0MVAMAeax3bQd5UmsJd0WqOtXkTg
NKjnwalTKz2RS4rh3MgNl7aFLIjyNHi7oq4dHGmartdx2bChJo5BrhyVrk13jAf8GIIre0yj6BTy
4Asaok6JunegzmwwQS1jTaQ1ejy5ZnGM6DeeJYyFgbLC1O+83Er4FPRX08ok0UFqkUQ1i72dr/yH
0x9a0k8AQrkSp3g41IaiEmcjIeXZ1olsW/5EY0vJV6dufhllbcxPTBeo5h25ZCxuXSM8hUZlK9ZP
w2jRATf2I5Pbx4DHlM7nUK0k+lg+42N8+UYMqed5djJ1WU2NFkkU6VhY3Me7Mtcf+3XWEVphBPKk
2lNEmNH77zCMqeY4wXSoIzT9JK7lBfJtC9g1elZl+b9QgDuidtPmoYgq+st2AjRGPFhUxXom1Uln
HGy4cgDklga+yvL278SqasMCWlxPqxWu3WM+R3YR12ALqba66eiljWM4GZ6i1obQIsR8DZM9GHJZ
bB2L6bbUz+blhk9/bK+vNy4h8QhreUm7zLJzu61t8xDG6liyRlRCmuwdwiQej2UnT78rirMDmrfM
GUzT5W8fw7V0+W+gND94ttsZAV5rqOAi7gBBpPJ20KQx2jLN+G6cW6UvBjV2IZd6soUnmGZwEYPf
ypDWTMr/Fpy77TnUssWNmnhgfYDujXmCeOoewzJAEBWQQgcIMgUP/D4F9WgIlbRE9JCebl/VfYXf
WF8Uyra/Ir8rLEMHErtcLJRfZJhOdvQKTBHfGkZ0OGx68tt+tvPvz7xWGC+4SEY/mEJI5zg3ab/N
O3r2evDrFJwToqDaRsINb7oEeRJfxGS88XtqS/M3CjtTEhpJAkBn1h6A6DSaPF+Yeix9B7jP6uYu
aGoC6V4IsBQt3587LWyov05k85cnnqd7tnVLWgDciZRaGb8fZniCpDzypCoiWaO+lZ8ZN71/0ilb
4jc8EoTYahlUQG6H3bjgcZ8McDFkslEC5o50AccUaoSJeAcnFwJtJbuVI/ovQdduvMHNull0l5f9
UB1ZInqBX+wW6RSsuD/2c318nZcT0U+KcOdZ4KPA2KvgeqHYQBMEME4Fr0/PNeHqFoyOZP/utA5I
xbUGvJP07kH8o8O/jDV+SXKEDJsoVM5TOJp5kbBr1GnEzC3+6/6p2HDSfdrHzvhGkCif/vCIsONz
5N5D3pDoxyQVZvBcWsNxZwac8W9kbZvtNNBVB50X/WPY6qa9bG/zsJji/MO0HUnCWMi2nhOB5DJu
XN0lpkmsn88FW/po8maqI/qn78bywr6eO7MeiXgkkeP0kS39Tvwp4i/uGfptW9BBVrhH4oX9SbDO
SrOexkeuhNY2uH4YMqtx39kJc9w4vjsx6rQzHLJN9HXaOQWN57mO832fFbc6nxSgDcprsDfX5Fs8
4Cu7bmbXDlGwxRDFpT19tey/WmD3hZo5gwD/MH0HWdo2BoFGj/+MXcmvIJmpLA7CDqzL4HeVrYqe
Oz3s1fWuWW1yHcvmEAVtxm5wB1QqtgIUsfzhyvg6Bf235YJu92yRI4msm1VJYAI+Isa7AoPbeI+i
/8peCxgvwiMkJR41pGuWnMCK+KMt5RcRcaO4j1rLCuPUfcSPQq/k/wATuNbfngnQyyfGQ23JXlzW
cgWus4pTb7ICmYa7T8e537C3wBGFzbE9TfV7NoJB0r7sWE/DViKSKoklb3qJ+mQnP8RiWgO5znsj
o9QejI423S5l+Hz/zBn/8J+Qs0OukXAi+6Rv9rpjw5XVOn0h4GqNFzuL0yrCMJHGGKlOy6ZWjCs+
OSTnqiRdlLlW5NxapCUMY99Z5paWkKbIxScl1Clt0YgRUzPQWVGP4J27vyYLbikaR+CQGRhxyO/r
/UrGyHD0pbk1WML0gvEVpWtTKSQkteWRcggFzTAWvK7dJEnM/cWhKJ357j3PjOmV02Hz4aDF18k5
zp6v6yP/KuaXutJ+o3mHGQ1Z8v9ypCq6Usa+/ABJT+o7J+QV/6/i+K8m/zHglxDGpBQ0CuuSWhIQ
odLQ4UIXv0Qg8IIXOA8Gn7e289b9Ww31PXrfxkgW6KKVzM9HrHDxry0nRjXtCIcdWD3DrioPX4Jx
mKkRFnt3OcUXsLkTKS3M4e8G5jCW2gL8JM7wL+60/x9A9uxekez/Hh5uHz4RCBBSaHXCe9AXq9Rf
Nk6pY+zTBxD1DHtTTJEUrX0gSuYrmJAwlgWP1TDYib96GFZbQxY0VxOS09+cqE3NJHxGUsUp1qmo
+GMFGDepY4ux3uZWg3i7/4U5yA3LjdxG0fKPNuRIAdbuUspCKZ+XmiPTLl5TepWdPHKftVy1Lp91
e1nGfSrD7ZMp/bZB9JBySIga7Xr6t63r+c9bh4Fd0mLgBkHm4whfWlWRuRk2QyWQw/nJa4MS2Kaq
oziWOKlvuaZ8C5Qz1e71y+FtGycBe6tIZCyPzLOilgr91MTOvboM+EFJQtaXfMUiW7Sh5b/S/3Xl
2hGAR7RakoRz0Ey1R3+zmHyRPRKfcLN6UoS7WKL2NsmRQ1YV/oFWzhi52zP6N5CQFpriXn3mGlnp
7ef1KH0HhUTPq18VXu+/Cmzla0nehGTqaV99fzd2Hg2vNxCvUwcelTRZ+tt4yi2ZvYYb5AMRsJAl
r48vFrZxbm10pDtvcI2JpD6ql4wd/UM2OFEcLHerD8XOqUrGU/nfuPcCdJPXPjqUHDpmwJ+Ay0xY
VOL40eJ7FARkXrh72OK3dk6bMBmozWKioeaR6XmcDrSyhNW7kcw/X3NOVnXzt4t0viiTXP/mdO2N
pFesCGNkxCktc/d3ftBY08cPk8useSCUqNP0NQQBMfUJvS4wrKAPMQFAI4uaDThdDuX5nfVyUfZl
Ii6Y9SoN0ecNIdk7D7yU/5ooP/p4lKDoeysnmLzg1NIsFtVFntcLCrwcj9KjcQ1mtpSBDGoKP/OM
+vWsFgnarMXmDFrhNoWkOlIvJxxx+qoXWwgPBdoRTeiHbme/+rPSKvgmd3CwxWRLGf54mo3PXK51
3FTveaLJnd4E1JswDDnJFRoSnzRzeQwKOtmJW2ZPehommwu8CRk6XF1GS2OamD2MthXYLB7W93Z5
v3tmTH+/zbptCm9y9WXNdTZTwev7Iy2R0AXzHq4F+ISl8E1kOzHqSeSJ1Xl8SVIIlZOxa/+dqd28
d8YjScqE3WHpggaNbXbmEriRrdpf5IsFnr0D/IRQYT7C2qQIbWCgdkq8F4oWa2Wpqqoe+/1g981B
toMBkmovkG0hqdIHzCyxyb/bfKJ7B3dapCXsXjcxIsf1rI4NvKFQCAJ1iVKPVeJk4NbTtJ5aSRwo
CIcRq0MhZ26Hj9rdMNsIL8RiXorlfYPkydpKDGPQgtPNWdW3lO36S63TeD/wTejcnj4ghz5GBzgs
H3tgbexZaWO2+IVODH7zXUbNnLMLAr8ffJRfsS1tiXq1r7TuEAfcKuRgzGyHej+3v061eM0Qx021
2Yq9s6sqlIYNZpcpZEG8TxKwHU/YaG2siuZktht5CJuy+oechP2DauIldQrOkPp9Zb0l4oLTBug/
Mrs2iTSLbAq0MM6S7EJqQ9oIrhEVeIIgbhFjbFAw1n5M2KjTYtQ1O7WzSv5tzrXw1eNmj0kJE26A
4wZh2s7h2ABKRPTJH9SB952eRYzrjg9tX7wHMPD4fvYFycwWeSWlS1srpXj0KfOa8XeFJanGUL+1
X7Is1uD4lxCqmchexsVsK4G9iU4+IAYZPs0yzMXjz+GbqWmUuTFI2Ef8wD4q78a1WGq+q82VuG5G
mswB1CX2164tetRJS8fxpcQelgRb8/NHRUgGwKJGnF0s2hakVNAHJLEqLKLmBzD+d/EsReWMMS9k
iBim1caOA3SNfpUalgfA3Xhi+N2stcUFMgHnnUA5ayB24OEnAhdURGgG9uVMwpUp3K1Hd53FnzU9
rBXzXxaKP75Igx2dCKQz7UT7rPZYennCH0b7USHb2wZGeUSX4IYr6tY8F2L2QhAYnx3uJdD1zWvy
6InbgK4T2Ty8l/lUmdJeubsgE1BuEQKtx0izNdDT7r3u8HW4U13Ux7DdWP/SEGVA1zfgGCBA4P4b
UWkU6z6gxSdJDEOiyteE0A0ov2ga9a95ZPGph6gIC58j+4znG9Q0el6Fsh1YIH+dd10hOuARe9wv
Mh7qjS7VceVfsw/v1v+OlQ6Q2Ahs/IIH2lBmtBXdg8YcKUE8fAtrmMyv5BkzKbz11TuVERwKrGUG
K7MbDoGppdTypVOJqkcTDIhG5tCpjlm9IoD3p2Tq4JYfccpFxINm9ZA0Q3pWg4JEjOfGZ/ipZBIs
Q+ofAUitXaiazkLHZjQA1MBIYyDAHw+2jULoJbOOz74K22BsmQ49A7V8CbtixL4XpNcY342/2IJo
AFqUod2+0WbIZQLUDMYWcy9GMl7DffONm/a1Py7llPDDsXk7ijU4p3QS5ONzJ97lBR0vh5ULGjXs
KY5i4oUy8qH4RvA9cmGA1b/jDnadAohpLHRY0rdfneFsDjxvSgVIUMdEkW1e0CDJEYHeNZda0uow
uLNzI/e/dtfdH0C9y8F9+BE5e8E5s66QQnuZ2bmc+UE1DphdL2CZaup6kT/g1ncOu7Y43FT1WIRT
urJemuXuP/X6bjYXjZ2KwsCKRPvwflGBBN1hjSHaPVic6ifxj6c/jnypBkV28zdpY2dc9C1AgBR1
Opi9dk3zHYtgIQnOuQ0ZXG+gJYis38pRH0WcoU1TPuj0wJ55FvS08AZuXbXbTR7OU05tbWcIjUGC
AHY6YM1JYdWgTTka20y3ReecgkPQs4kS9LpGUqmgfIhoOZAHRnMXBLiuVsNGgYdiqHDJ8GXuCv7e
mKPWOzzZpbltXJrmAIoZ0Pv19zDSVwYAbHtUGT9ln+MP8v0xgzRsZVDnYF0QcGvM3/qt8dIAY2IS
IkZBrCU+KdmOxjbxygD28+SbtPzImotDzpFEevUCMHpJltF1YCfMf0JX73aslU8O/eI0PraDE8Nk
o6ok1mCr7+JChkfsQHGCVd5LEDw3Vwkqq5vpGPGRaxjoQiFbdhka5cn+EHzG3iTlExG4FqT81Gw4
nTkk2l7WIoJIit/JzqjVDUVMrdjdsjIGfzfcrkwINfZwTgcSwUwg3zCfQvJ8UpO/hXCM3oOQByPm
a2LujUvVLX43ndcIU5YYB+9j++1cYA2E7QEUen8EawxAgf9LGYZdUcyf5d4WoTCwws+lTEEAChqx
zjnTyTrDDJ4l8Wu8EF7NeTwOk8yih6a5MDiNX/FZWTDo93v0WAlhaDVZ8NqNZrFpSrNKYu1kzHD+
aJGPQkXrcogoFm6gK1myMY5uERZhn901DlEF1KqpofV1c93RqDV5DqCzgpH+eaU9tQRFyPML6U+0
0yK6uvaXkXK9lPTvweUrSHgik9gznDHTLt8TvtNUt2QE1Aopui7LZ+mW08dAQsZmsEVr0tbIbZwn
ITp8NktqTx58khrSj5Becjd/JOCyMre4Rs4EvldR5+HWTwhJjVC+cNLUl/MsAYPgpirlEF+K5rUc
CLTUxVb936VqybKMOpjGVuJo3tiMdPHAc6zoo5zcJ8vNineivOUOZy38T6wkrQejGZD4TgunOxBS
yLujjT0erew6+k0PgtKdvTGtN6Ngrqc68EoGA5jsUrmLrefI6/74uk/wiN7BnoBuBSr5cT+Lwy3m
QjYxbYIQi/Q+9k4WgkmxJIm+JTiJ/foVOr/FXvU9sqydVBRLpq2FZJ4uELuatQDwKEl+DIDv7ckD
xYnPLcUZCj5TdwEQItIKArk8sx+ozvmhWfuaJurIgS4flfsQZfj1l/RiB8x/+W4FADZ9ognq0gU/
kAhnJm7Eqyy18wcVjyfjhWf5agzUZRBwh6cY8a4Fe9oD+Uk8QaBCByOmUb6m5GOMm2HcHbZZycKZ
ShyeaVPZS2q3qsuH5Sd35nKsa/5Dkdg4PAqhCVOxlsn26bu4hmkN7F8AFJud6UJfAbQq6OmryMYA
PPDzkONw8FGA+ymqVxnkU1JqCMUAsz9Z/M9l2nH7yG+V66qFQDk8Ud/f/9uzL7+ldIFkRSHygbAl
L+ADC2q6WqSXZ8klKLKwCHJ9jk7ZSLlUySVIgcmtwCTSAPMq2uaQzWK7Usiy0H1lhcXChC8dEtUZ
gbB+oQ9DYwWKm6AzbTkMFRlJ+91iuPjM2pmwzvRuN4Ou7ibdwoSvez0MHugz2T6b/ug+LZx3ULwF
P4gJYzI3N7Z8XAp+4f+lPqnNAxb67Lm4+oASCKlrWSZEravI4XGO6huw9xxjAhiQijBj/LC9Rpf8
0WBXJcJi86KAwEQ/80V1kvcweKOBzYcXajiF7bigEf75Mve0S3Wn0nnyD8422dLG9P7SZwVwVaE4
xYtSatojEer4uxxp3YYzF6KImR0fvIWpFj8/8G3zqgmVr0xrQNQF8KJJGlnqI0++KQ3FBcoqiJyU
IaRSxn+vb8rreGEwd7oxoMmqwN/xpa7IEXwXGEHF4X72kAKrs1ENWV78qO1OOJppvxkanrWi+Ttk
orG4ckMj0L7VKsdlalq7jSq8setUS9ehyCJLG90odobsgnAj5fxs8MuWOBVfiFjP3LfPWsWgEKim
2OiiJcfGTwLqp1wnM9YsNmarqwtZrUZCNVGf8PX6wX59CtHG1VSu7zqxv7ncFiQZzsr/5QLyUt9i
Bqr8I2KlNpqRLQHVIOutsoYptFvrNVlIrOlbyGpu30nQLkvwluqt9ZaEwqPYnNH2WTtL8Cl3ZKrx
71D2zAezJox0cPyt/HiHiV2Ul5NQMuUk5BdghL37a1BFNgUcCJR3f5olJcSsTcvAjK+T8SirPhsH
yxBPIFGUUxc8QL+ptKIsLrswvyXdFcTxVSnTZPgEMsoxt+Hz1Yml5hnbsMcog9ltVpp8u29Kpmab
mJjLaTJP0209yDAfPbP6QDzgXxYhXaSCBYnyBCE7lofwtUJsF9qfQ4jQx3ZZ4rukWmciOA0+J/eF
olgrjBEc5qaq+XCNeIzJonw4RIfKJpTvVW2bjhRI/+XMH6WlhFq1PsFCTVCCBgeDN99b1IfLsbR+
yZpg8GL01EK7f0Eb/JZEq690US9WH6W32Nib2fBbmq68m0i47B2yxV6Nd39Ioj00eqSZPCUzOKFy
jkpe30S2Q3VqFzzQ6oRzZeoHwGZ60RohCElHIsvJ1OmToH0cx4iFDtNI2IkttTLn+95wjHIPTUVR
4aePZYsFWFmX20ZVmZWe06M6kLRTNpBdEdKJwLkc+QEtmpnYfW9/r5WeAKvaHpxf5kPDD3fD4jJT
CFJaOw4/7exJiQ5dRtzwB+MZyhvovDxvBhGeCwUofIn5xN2v1QDhQrWlmhfjdzX1ZDxUl2Qkkev+
v2zRH4cFu3uDHpoINdCvPwwkf/d7p7UIOC69GPplxTTTknlEeYoZPl6mVcAnPpNAbqbKyCfc81zW
doNMAEMkmiDrCl70MKh23fnzWtgIJaSWIp0oBts345+kECD+aJwTtbmiCiOCG3vWw6vhrg1udpwB
Im5OS+MJlwqCGgSyOzBdBlXV1UotgV6DNtJAEjWMUi7poloaOvM2TQM30c636vFHKjzu0ofpov8p
aBCt0H5DIkH76suCNlygPmEf9YbK49xnJ8pWx5qn2gQTSiMnVavthOIcx0nPnn6JNFAaUQVXOdqd
ate5ZGeVm60zyyVSs4H8T+6d0D9CQy3yiGgyPy+KqyetmZkX+ZenqDPLpw8O4xbxViRAo6tydOz3
Ah3bNRuaD/ByKddR5cyMZS+oh16NUtkmbUXE86uKUH6R3MUhvPjfX6ILhwQ/tQXeny/+Whaq1Nh9
3xnUvlrAZVd/yP2A1VrmNqAlE28nXCLIvt/CVyyy/TfQmtdlRAN3t4JKnm2URjM6S68B3YMpYWoL
VhhICq5PVF2R5bQMPUldmj7Ld07wfZR+FaJJKQL8+5958tt+O2dFG0my5PoVklDlAPBfJ/6Jv1LA
C+CDZHFySZ8UbUOuMaciAtzUiy5fe9zu1b2jE8UuzJKsj0TLwgqoKy6uO6O4UszTOqRYrvhiE1Vv
0Qait6TOpdR93XiTJvL/hcMax+sGDxAcXTeSXUzk7ry9UyM7IhRYVh2sQE6tURtYhZmOIBlmlYK2
eyUAeHq1wskBBwmT2xfIoZHgCEdI4jhwjDY8B5/8GCk4Z1ZUCAuVVCmCXX89TUAxRGoo/BbvpF3K
Al5JehF7e+mMfIQeHXIWSTNXGyrgUSko0IUXKdlu67p+GG3I5q20hYO7rqDymzeVNdGswnC3bolj
Ri442yyNvsZstMnEmKObbTi3yhlJ6oQfsXAJY+eC/g0JBwz1S6GlmqlXConjP3eccsKDafqrAthK
6iK0468eMEcy6CrPEa3JLr2HWww1rJmtSrjKiXny0u3mcYt/O9oSs0fK6VcX2fAp/oWJFoe9w6RX
tnizmzrfIEZkgAKA90inMfgKf0+UbRYR9PQy44qZcx64bB26wORW5YOTS116CrarIhr4xrDNIFVi
99rkVSzwQjbkqElLTSnPsvwQVFlBg/KNQYL4pgmG9fGcVN/6Y7QNLPAwn7pLeFLLeibLMzF/ZsGt
7aNjKnKJGDv6CUwBYbA6ftMlikB8YpCMVjMXB9S7D2QlHUaM1+1jk9Q44rsTN67QUK2yYIW1652e
QEwBMNmlPqa2YrHrjQ+XF8719CCCH1qoatdgm2K5bPsRnksCMotbBcvDm9VYoHs+BwPIGQjnCfYH
L3knzkQI5UebySP4Cra05lRtBuOAvBrsv6tFPkjJGDitR3D7cVrD1jZxX131cbohoi4dVdL48aG5
BqpVzxEz2s71rSx4sC8VC2Nnzr1ZHa6s2Hbrw4WB4A7tVOlYIBe2+MEbOynSwBR4zcqUrmMyPkcT
T9RyOtotbNCppWg9Xz2dEO2+xb0po6IdwZDQ0aGePJBl9vGPjFnuUP2LQ3VbnZ6mYIdMgTKWy1tS
TxzgIwbqa5Mkmn7xu/Vkf13GhrYePUCYh51nML6k3LzMgMONQYZfkcFC07/ytPqutJ/mfxeq2EBx
75trolHxoxxSLSZQSh3qGjn56rLLDQ6oJW67F69jnMTJG4TZ8QGjwAxfod6HbtwSXCCdx7DTWWmz
MOQvS3aLLSUcoi29X2jNZHhJTXMWL3bu/iodiY9TGSv8Gwdru88zL4E4MvhCb/eBgLpNdF9Sey0f
9F+Um9bDkCwhmMyKt9x8ALdEu3pvXXpLM84eRAvnMqkXoQfMyy9HqqyLMWovdzy5E9QCnAHdcjOc
uhGkauYdhinxmvTtB/vNx8JgNoTgV2yl83/hByMpFKHyZaH7TKEt9EqfAcMi6QmOsYSanRpD5VPg
2mNBfCqzHH81+8Wk4S+VDBZBBfb/XsQ9BHMVdiV6SRigewSb6LJYtZ5qwRohP4+YE2syIwUZCqFk
NK4EoJtkP85GmOcC6I/81u8Q5LEyLf5PzWctYfDgoy1jkGliAtVCoTvAYhkUn5ImllV3sbJgWsuo
Cz4Y8CM3xz99dmLtrL/c5x/21JSQ7JlXN/6C3k7Ley26uea5IfwPfNd683DVSlQUEDbkTi7Okkff
H75ru3fl8gAD7qcZ++1cyF5qOkT6FoKjk7rLHSDAeAvyhHJHor9rq8Z3+pzjBS/IEZu0LsvH+1Q6
sdGV0OzQCyEXxdRymoPPmdBgGJqlTv5htOUfh/eKxkPRJNOfz5v6fvmuW2q0ZNjPNfZl1EoxtJsG
hrPeuZhidUjeUFKSWdHlBoLxXTUALP4/UlfSI46Jg334jVy3hVOSScc2xSvCD1C0NSu7cigc5qWt
AJ9aJNwXSwl9e2IukdsO+LrNM0PErvxV3z5PDWM0agTmoEBceMa7WpdAMhCIi5+pnwM2n/3+AsGb
srzlzNqqomI85UGTojeuYSAK9Nruah5eZd8murEzRaBVxJCCR6dKB0St+lrxvE6zC+ZS9gjLujsS
CiowvIyM5pglgcu8gW7n5PsHhKIQAVnO5uGye6/BoLlf7GTnib8Q705hy2B4BZE+12pDy16SkRPo
XVGurHlYRaV0s2vjgKxf4qSOr15s2ENJzhMd5p794X0uUXHRGqfynNoFf4Lb3T6pP+LKWA16dbrt
A9xajZI+++KIdluq+D4HiR+bCW0YDByt4YXuBpD1ZCMYCwM929ulVURMgmBz3LioJQCBMrU/t/an
6Af82a88G7l5s+UbXWfHNG1ox2B75FcgBOlR3KmwI2Nub4qMGpktdWyBDd7zzdayfZOUIZ5yW8mE
hkCKpufl3r0QqHP2A3QTLwLWLi3XDSaAcA7dquGSDy4SY6e0+LZ1/5rk0E8Nl6mN5JBJM0pw082Z
Lh9JWFHUaw14G2l81ckXt93yxxnZ0uNUD2Oot2CSy5vaM8/IhA+uaKXPRFAlfmFBl4fVmpHBACQg
qw1DaIvxfrzroGYzmMe0bCeTq5UwhNEJguMBnGOUXUCuUUMHjsF1QKEKNs58gA3FDkpXqftqnSsT
yjRWcm8m8OLltme+D0aZi/GKtPeIFPT7AXlANg3ZBTzfgAYWKhL7mwk+jqtRJ3G4EwBFZlocgnmz
JjkitKw4EW1qWKaSivAhQDEfIyX7jNgD/LFHCKZhPR75nKEzUVOdCRxsIfsOG6mQ+1QabqqsWtha
poaq/xTVswWSMkN5pICSA4VvJXJ3qVpAjXvt+MOSWg/IhvBi2uowVdfTGzXMZW6nJbn6WSq/+az2
sL7o/6iXo+cqbHZdb25IcR8Lj27EIc7Vyzuzl0tq36OHVXOdur7pDrypNs3KvhFjavpHQHmeBxND
KQfD3PGKlGPs205EWlF1Sumax7hfg1YnzDTaOiiWkR+esQZY5KmOsGPc2UDwCPUm/qdeME04iLCs
xPgiY382Rwrme1MP8o+Iwnjyh0zbGF/SYfEI3LoUWXJBFaWAlYr4tPYscY1xJbuZuF38oagzQkJ+
132mCtUJ7qF/6QoDfv4LQh9rSHfkOZercTS+3SDw5xe3RxBgZ6HYJ9rDgtKewBXSsS4TI/D5g8HU
p6sjnxO/E9MGAi9EaS4C/Q9KZGTSCtOWWiI/N9fLkmFO5zuuLrXSzFb1kRzG/QJoliavTtkSxIQZ
JbF1dwga4hA8ww/muCCRQ1gwrA0Et60q4u5IxfY2OdtVmrom5YJUcR66mTKridnynSyorrsfSZ76
PEl5poW8oO7h0Uzlwvncpb4DJZfnQlATM0fF17643m80i2LN4I3p3KUSXahFdA5A+H+sfV8VT375
c91ngNRoc83vum7vo5t8vnZMoKWjH5xdtDaaF8k5vSpK6f97WkiW37Ut/kbes5zcwI3yEmQVHtOr
yLp8Ho0LEOrZ6mBQfFnIa0Hvuvy0fxiymcVlQ8Sf1BcPIJNgeKrQ2keU7LTshBYgHWeYh+vy2z2b
Z4i05IXB2X4QiEragA/QocTHxcABitspRtREQgqQDKw3chSJdXcQ4KDiP3SriBHf86Rn7Ti21Vzr
/9M5F8ev2sFGw107by93roB2HPtA/QneamOYRWHi3fFmzccR4gxITIU5PZm0nRGqB/iJXp3r+3nX
mUIh0fHATmxXsFKyRwlZC3qJ48A6if3pFBuHWQOn0M/+mrboqnjnGp1oon/1TGJx+efaRT5/qLtI
kjS4ytM12m9fmumfgkHT9ZSJFYFonpharajW8Hw+yGCnz6NxJ0XUaPK9YeubgDZdRW4iFG+cBPLq
NKZ8RiMbyXScs5iAJqMv4SqMTwfQPORFFo94/3RAOwTE3FH4ocP5cMEVyqD0YA/CL2blXUudMbfg
eCA1Pa6Z+iUb6z05kL4Sa1jLJFvD8WKVhNLKJjSt5J1qzM2ZPoZZAO7eMCyp6qOkvI+ctTBPcmcM
Nr9Pt8ZXLEpsWeW9OJ73iV0f1nnmThNPlvag73ylvd4GjqmzKELZQAZPxGSYaSv0W6VuKcZvDKZC
JCiTDxVKGPujCDJ4aEVfwf69YXjURpDFF0WCXQnJeOvSt4hR/D5nyDZ7EWMMSmFH+88cFu8T8TCc
SCk2WvNgMZLSFlxS4ImtEmJ52NaxzqzkRVKsIDyJVYuhOSc4yt6fykGeQPfZJ6tt+SuZNkItnHcM
/0xI1a7V9cruYDcNiI+GZ7oqGQRy6ag+D42KmnIb/e19MRkfhS/nCzzxSkgCthknEDBP7cnCTxSX
63c+31+Y//P6Z2lF8RazcFrI+OS+jNopokTMVcOWGUg0HlQ4oNCr9dRRanseNe7hsUl3HZQbPrxE
0F/kUB2gIAYIMKtplaGOcPV1OoiGLdi/OMePuU4zOGkH2jf9ktY/HY7yy4SBdFGKE9yj3cIO3p7A
uMyUlF6cfHLlRqQyfOwK6DfDUfaF48cUcTHcXvTarl5KVEtvbhpuCBHyOy1OIrxAbvLMSfVAzGOw
U2RUJCnYEpiL8dpCGc5w+2xpdKeSZjkPcnMeJRos5m7hubAWsgf0qLFP5avTAmX7/MUIwRAnLxgY
9PTb2IiENDka0xun2dpIb5WPemQLkHReuswItRJhG2YztdvsKbdiNefcDH8d2t0/IPD156u4tJ3G
N8ED7UwZ4/focQFvqTKhATnJT+xqtpnZX8BaErvCOsQNqBxm3nk8YEnWMFtNVeqfo1X2El6kdvdQ
RbcVp/o5t1HPyStwmxG1uAKdMiO4BvSHkaK9wC0XVxDnVH0Fzi0E7AEmR17NoJt+kj1G2OsDE5Jl
Hpu6CelMOjHznTv1HtwrS/76H5dDob10YEa6sERrEegrEme3D4JDA1BBZRDtEll5YSzbY8hMIK3r
Fa8P4KIm+S+uwX1i0dzqWUCuXrXONN+1NjVS8Zsxy9woWDhful7gEqBtZg6ug0RWxpip4842AXpH
G7KTfePtKcBKXtnfY0c/9S6/1/sMNdF8a8i8J+t2nKkwDk0CRHzIH/8IBED+eFD3oxUewwl7llTs
hPsw1gmD8NMdP/cIsHd9gUUhrmbYfwhi7IN165hv4gbPVM1lKBM1vl8sKC+LPOYOWnONSaeCOgw3
216bkoVgHXgVYOCk0mB1fMioXWzAslAtNKL/TCNVkMUuH9hEDmZmwD46NpB7ABgliBe/MHY3+3kS
piQTHyDDEi+FjCRGqdbUCJeAkcaLsPMUnkItOKPWEw8n8LXaqENH0I66sxQ2DNrfgHqKg6k4TpzM
z9kbPWHIf6MzSDJhxnFygBRqE8CaWVI/npkyqlT+HXx/06seD1ksEJQHrM5UaqEC7Eke4QtIkSkO
/bfEeb9htj/gVEqebQKc/jbzrdmg+nVmOsSG++Wp8K4X4MKgLrrj14cLhg1rmiv0VcYrKUMjEL0N
J+TWKDw3THhZbZapc8iSzxbbL67ILAEyMOAI2G/WtpbbtzLsqfLNuHzvv8hwdByNcJaBCeCofQdS
K6ImxzLZ953jHLL/THQA5fm+4rfVOiwUIaoTC75cuDXJAdGhy3YWpdu25WKCbCpwfQNsv4NysbIV
43p3/ZwbygTUwkQZ+AVPwz9Y7hy5VxYu3Syp3BOvOxyerZLsWrsh/nyp7uIpeA3pcZHcIEbAKLcP
HabZLxfVyB0f1ustUfZh5qqnYQKWFRW1mkdoozXG1xyIQk67bszKesiTUtLddpW52JuQNh5mHMcU
MQI0UoAQaJGKIlGBEk7Xutd9VZOTFgeOJ+l2yzfeh4CuW6Y7SPvcrjsqx8q03w7updpviQjszcHA
BIf3VKhiUDJX2cyulrErQFUWDPdZbefhI0UYzsjOEUwdTB24XZfY/iJOQMqWlRv+dzzw2N2OGBnI
Gxtub5qOLBHslxR/aujQMOctWghZyfBXWFjNXuUxd2XoAwpnz3zKB7DaCooEBbrrCEjO2woRFsJB
jlv3QLqzQvBAQeS+kuKUKE0eBQNpYhxZDzY891AfHGYWBfXW/96c3okd/WYeC2U18uRITBLGTRZy
MnkJLsddgfrO/7oDu6avXGO4a4qfu88u5N+8zx0G6b744bbwqrkDTZNMQSyZwUJIo/AjKGqAemU9
gxl+54OZUPr7dmM9XiNhP9eRWbj7ji85AVQlZ6pP2/RFGY7FoaVz1nbCWjmncQttVwp2FxwGXIYf
aYi03nSlPLfKM+zau5kRQvBUuQyNHQ6iAYVL4pQ1hjLiPfNihtPcPNTaX8UT4GUBfeGWjHI2nbrt
WGRDzyaDtUSiA0C9M8TMvYX8IIdJkUuzREb2za3inZnyXmd5Xw3B32kYjGXFs0sobfwXqxbOeylC
RMl5FPokwGoUSYmt1Vf7/UpbSnrbU+tIza2FtdVS+LGouFGAebhCeJKkjipNK2nrRQqN0/1J+cGi
C4p8Dnet3fU6LRIyJOwwqJjZsCBU8vLPpDM+uWQs26L3znbrEj2nn6fFiFXhDc+7sGZoHY93l4lp
ipdTKwMCh+EtXVFxkdB5TY+Pa9N/cxXtXKitid7NnzKetd7szTwB2TWJLeOZSNPDZbeMcfIAD3Ke
ZMGcf3pwtNK1WJfCXNDhPSJyu8vivbdrCZueDhMII4vy/Wgx7xAT0AdWyvrjkDi/JMceuggXcg/o
ES/BiP1+HlfCqzohOtu2FYyxV8676CB8hS4HSsKKdN0a0Oju+a3Iqkkc6HaRyHvu2ZYQwNoEp0As
ePq1qp8HuEksFJMRZQg2V/RsGjgLvGZJimiDZPUXpwTZhbn/Ri4c7lVVW8uvrWqr1zakDx6bzM7r
4PvdbxnUQtah18tB0PmfUeV33A+mqsJk+ZuuxKZrG/DVxfdVeVUln9Zs04/o60QgMlHzSGwmzUCz
axqlxRD7SJGL+qcTN4PSOaophAV62NaQsN9VvtZ5mGdK3RkrsHBmMS82YeyudAub6yXvOHWHeqqO
caKlBOFf0iDz+aMjcVKUS3OxdGE5Yfa9krOlT8J3oka5XNrbAiNKn2EXFHvqM1Kqpd/IwbGK7R78
Vq0kFLRidQCcXfaIOTmvgxqjxaZ//JvAPGLezWBNZXB27F8XnepIpQJ2yvFYvLRZ7u736rwc/zDa
akUDZCfl4VEAjTFFWkUIwmqdGyvSnYBh0vJHKjM/z1BppMfU8gZEBHagNGqAdDANGS6UK2kML+bE
v0RK5jWrHYS7S0nCpBim94hB6YRV6wjp+6WoJk018/VlJYBDInuR1bnRdpQ7eDH8oKEmOS9D5b+B
6dnTAUAWoMa579OC7JU0UrxOQmmqO1zYEbIWLkdfv1x/MIaI0Om6RWzW4NUxDIoYrSGKGHFccviq
cieuDUPT+TZ1LugizcWKTYRO1pCUzRQx1HULZ/jJ+D8+64miOyYp+bzfqx/v0kXyEHEpIKjGQCzO
t6KtFi21r5KagkqTo4+o/a63g/U9f+ObtckFm4bwExv4nMvgOl0A87ZpC035aV0Rx9mvskb6e3pi
LbKp0QD6HYue9R7sO6gg9kwJvtxuRsj0MK3MD2KbfgS01vGV0pAAoiWipC0XFl+yjMpHbxRPSw4I
hgAxAiw4Dq6q83Lx8cDR/STXqBK3/FIsXhPN+2nkpFAkZd75PuZTJQX5HxO2kp1nxfP+bMOPiqxn
8mkYuzxpomrXVnGevVLh5lJO5l+fGnDvECz64QaOs1RitdNFa/irIqcS1hjfqOZB4AlOcxXjHRb/
ZWZ9Kwdfup3D7Q1/lwAv7YifhpF2OaMfY8kmqMENnHrQZ8Zq2TC7ySbxFDzwDzeLw1VtAMFKv8cL
FdcAHB0ZMZuoSAFmPPR5JmegEBvCqCXXOVlJtUaWK6dnK/nOLKoWQ2KgknK+wjx4Ewrpsr+LPJkQ
CFqMKJpYTUywl4UgXxvybThKrpMqA9oM3N3zuobV8gSai8RYg6h+0kRriVaxgU71ivElFaaZdTSz
9oT4oxLF8p4x3WgWec+1f0k2PFqsernmsKO7U26qA3CqP6Vs22Of+hGmuC93ES4t+BYDsF7xpk87
tYebgMN8KwwBj1gAtGp2YT0ep/4n4Vxk0vS96jvUz/7aYJ31CVPc5cvbAJGUFCi/qIOha/x5aMQn
mjiqK/gKUZZPqzNVTCj9973RjQTsZ62PxpWKq+18K7vF3tLYMYeJJUqN/U5emtoyV5VnMF/UVCz6
bbCgEPYk6NlhkLCHGJ4+Ee+HFDEVnfbU+g+rxXC46tZB+C9HDtHOZ7+Rr+zzNRv4Eq1m24WrQV4c
gJI1XjjoQ7X7szxUe7gKTWtvRuRL5i3vCflLXQZRlzopUG6aBHlCImtNfyEo15dJ1v8O/PRs5rzj
SP9az3WV2HzAI47uh6SwKzS4T9GTSp4cAKiLql2XJawIt9uRsMYP5NhDFR278HM/d39EajpmmJQJ
/o9aCXaUpB7subRgO9i5mIAdck73drKUPodo3lWQs6S+U/rVIow0O9WPJVTHPKosLqNMb4CXT7ck
rfRL0FXHkFz5Rs5rIqu+50xF6LjGmdemMpxNOn4lehMl3EVWQTQL7lYUG7wOeBqCrEpgTmBUOzz3
1oTBlaFxUR3yQhKq+4iAz3Ei4tnITRVtY/T1vxmVro69ENAtN5eU0zQuNobRCTkSqAFvMSZ/67+E
aJFGp3gQU2BYavDpWYoRQwuMsIqc2eC8diIaWvIko1/L7I/RxNaULE60eSVAjLpt8M+rwep73iCs
svbrXbmqbLdG2OxraX8asICuIpea5ZAc10l19tLXijf3yll9j3DNvPS525Lqc0lxTD+Ywg9nTpqE
Ku0PnNYcq6Hdrn77/NhLv7oeUFGEQFAHvy7bs7IeccyRvQZjMOkBsBRfvdXZr7TFxmOY+AJGHZUp
3RAsuEWJ8Gp8zhmA2mBc+KibXMa0U8OZhQRNQzLXDiH2xhtM+HUX5cX2Y3NSBcaLE3vqMwvKxBrN
WkD0A/xNsWfAy82kFYYipSCP+1UgBAB2yBwCG0/hvZ18LvDjIwnrd/NqDIoX2pK4soD+wE/h3Cyu
EhvOcVQ1CNZDWB/nNxzHaNW787WpkXlkbFiG/zJuR3Qy2mULWR7ywzn4eKJShwa51TOwN8jsEoOs
n/5zPYOzSag5k4O0Y8blIWCAsgJlE0jgZ2rIu9VtBaatTIwmuH7hluE3vFiWdGqlipCAdYax/qfw
sritns8RwpDRFPw3q49EnLkZi9Wg1OIPcgsxQPc9ENRINNLu08FPSxMlxKfmlVXuDVdTC7LRISCj
RytCsHS4XCTV+9EJhzxgVh/+qN8sZeESxSU3PQeX0oA9G2niwcpbYA0XMvcP5B3spr2BUZN9AW3S
PGZ2yCYB44ljBqUUmd0qM94TT/6rkSb1RCVlX+DsjeE6pOZDufjBkyO5q+j0zZQ5swanxIdnZ4tz
8zBNQFTvufiLKp/uTIZNbOHK8+2zAOk6iPS3dskZUzCkVdygpws6ft8DrjTSPA+thjSOencTSv5M
UMx68DNGWWTYUCKRIlJaJErmbb2KE/rR22q4Mnur7hi4oMJOEK7I46LkvZXRiIXB65NTqIoMhJeP
vDjfQ2QktVtt8muiu0ZAQ5SuoPQmyqH25SOZHYS5KspPVSWc5FKeI+HNsCqlFLSguRs4jwtKL5+G
OJDewe7s/jqGZaLz6jlkGLEPYTWTJZ78zWF/wm3qASMMRVUlgvZnJtKi/aGZAJuQI27mrR22atMo
I/vKEWBfCsVhW+aIqeMMcgWMUUSrtso74bKHFZCGwLB0lQV9Jtc6LkS9dDoP6lUL0cn22uc5tlPf
9uv4v/ok0WIFb7rfbpIBMr2Ec1q8oJU/AEYyUIZt4dpdtbvNCeKCqqRGsQ695mpr3jgfRdtblI39
+UTxY307GvEuzMaXL5Flx0q3Cv+QYibhUTcb5ckVrbhLhToD5w8LpzBY+0yCVlDYBIWfEzOSti25
7Wo6P49exBaBY9l/E3+5sYaUDmXVsCVgIY6JXqoc5OhiBwuMFWoNjNpLUzk3T2myL3GdqV4pNkVJ
k4CI6//lmz7SNnzJOFTevz88pTo1XpEmAs5afdbmsCOuL6VBMMLDUHVO8rvdg5DZVgOMIg8mhTd3
ts/IxRJt3l+MZYyesjQOVTPn4nJlbnE7bOOm3ctT6llGfkPUcE75fY5aLN/3LldxwvTMNsY6p17w
hHtT2c3ZNVm10M2DnJCGQZa+5XV01omZHAlZarRjH8ym7C5wEQWkD9srH5uFdAlAw4iieupGrqxt
VnKMLTD1BXYDhLxQTim85klKDjOjY2kpy/mBPei+yUl63LFN1AhbUQdPtbNCVic067vvuaePEzCU
N1dnTswxDm87Vi4Y5aHzJOyx+QcDmckupLZ4fLZpoBIE3SX+rBxy3RxL3Q0gyUitY2JRbiQtfQv2
36ZOUn7yV0NS95lIRv/CWcKHgUmOMHfx6DzX66K5qwPY5bNjVRdv8Glk6uCr1ieNbVTJGL83tYkg
UexO8X1R0ESaY8Y+4HFrSQKGU3Y3eSUYuQo7g/xTXJNpvGuWR4CEB1IueZrVfPOjtTBKjp1NtjOQ
lGSUrZPwHF/sUpSYTrv3jEVHE5Hq0xHZLqvDqhcvKyqmwfnYVSNS9yTf+rlQhXnT8RU9nhJ5uyCA
eywRGXYMKMLqu6Uu99B72B/nSLO7OU/xhgc3Q1mj1jT3ZMo9cxKO3zB8ltZGDGdMM4qHAC+OvazB
BfV3Om3grGxoGcHpL3fIg+FpCbocrzosEO7LnvIYNGdo405abPaTLstOnRlyjO7TkPeo4/QUtLwY
MIQjxSnn5o7mtMJxGsQLt+2BTxR6pQgU+vZblvc5BcY2Q/Z9/h87/AO4epnMw67lqfTAu0VM3DQW
R7ZBF2M8nsRD3PSzuh07wyztBYFFI2132XEGsQgXv3Zd82x4vkN1ZCpQHu3lIEbPi0wq76vZ7p+H
3Wl/DxwtyDMOMlQW3dPVFCiuSKsEHqiUWAFY5qzVpQ/esjzwJR2BPlEYIzTY369VXy9vMhHgzR01
sztI6y7KaLqMqyXCKE0TJZbxO8KxNo1e93rPs9Q2UicVto1Kj0ny/J91zJeXTAN3UC0+kWQhiB6F
bHAC+x7zOstZkVfw+Y0oH5Z0gmG2U/yTOI+vqLcFoSj9bcy/6uUIgO9I+VSrKDaRqIMSi8R0sliP
ijbfOdgSNsqpk8a9zGxR1GqW4f78Wi/Yv7TSsRLp1G6ujqCp2RaMH7jhKBW21iRwZDuPhHs4kCl8
3Hig7/MOmUnqMzGRi30uuhM5j9GIxFDuGCD/cD7V11A4ecikj6j/F0na8Z+J0CBx8HjTbVA/FVxZ
1YMdTKqV+fdpx5vhCv8JPu6DVTvXHcjiCzxnmNsVt+VK3bLGfkQ50JjxjzZ18JpQGGhugOv5QSW5
DLZg+ycC+0dRvo6sBbfplyjzTk35Owg/aF0HQwmXcQ/Rdq/MSH5CSccOGUSvHf2qymEz495Uub+4
qdpkUVs84yka9XLY1IQ8gYYfmpF1edTvAVVAoKaevN3WfTdYn5HI5DVmaKe5a36OfMFMxsbHY0eh
GUOcgOD1XkhAUl06mJXOkFQ6GtQZo5D5aJlez5zuqcCIzw1aRRRWCWIt1chWBMjjZuol1hQl1PjB
EVDLpf0tZFfJuXAEF6G4c6GgY97gZMdntNKCx7V9YPCu0C9xnk0SuhpB3w0RakIbGGGK9ChyuR6B
IYXX62or6mWaTqaGVZ6dJby4WLViE/XzN89pSILCYxhTNRF8grKxEYPQtHDcwlvCIE7eyuvoSogP
tBoLo/6ZvW2NaVCPAZ0ibT1F0D6vmmi+v8WCe9keig/ICYDD6quiuWPf4nFCAao0BM55jCk8vYn8
KWVDum49JSyIRM6I46p9JtSR3QVQIHQS954uyoJ6MHb8Tj7VPcs2AhOj3MUT3zi1VVsEcFSx1Qx+
Ns2qGtAUMMYtv6L54/WUaObcGwCpSRfMZzmMDIpJJdXvP6J/E/+4wyfatLEb2Iq0HrYfztKQ+1/O
NI7xIUxdqLbSPTE5AUCU1VszilGhwTNg5GptXTyJuEonFG3GUCeEkmBLZ4tGjK9KKbQgSEzo1RK4
w+mOOH0litpnMYBhU66dB0CQ8T+QkEBDPDwvwd2scugSVlD8vWrywX2hdRXvhdVlNtp5+X84xXuD
Z/x8aJBxmjrs1VhYo5yn+c3Dhck+7d8Ji82TdG1USDM0z1PBdcd6C8gGEbPHZGN0muGtScCeISmm
YEa4nKE4tjLxXJcsLAwwkpGLAEqfhnEKJL79MqWPkhIxpsRtDjXoKJiEYx77glqLP4TX8v6YPk8r
4Fxq+JarQ4iji+TVUgtoINOpQgawD7wUuhpGkSqgoXsdiLmUGamwamImG1GR8tVgn20DuiGG9lCw
CvnLC9Smtx8CCewCiCeJDacWpUNAbVTErtXez159zu0QuBRP5YC1ZINYH7Vt4UHrPjO1PIyHGmND
WvdjV1Q12doXRSmMV33eWmRunOspM/ZIFn1KcFfLAyNNgDo61BeHcC74j6t1LM153vqEcmcYDznQ
aMcZbLfc4Z5LIXBU7/JMYutQnqUJlyi2/8nplXaJ0FdO/XgXmIPi/5VeRaDm4cfjHJt/tOPqnDO1
+ndhShi6He7JXfbbjeYlm3IKaHVGSDww2EaAJ/ruUSvlOejtyPp7iMpxSXDTjJqM9O7S2WVwqTqE
zE6af2GDn0SqCCYzyVYR0aCZCxGqFxTcfe0g6htD6HITXgz5klBBo6esBzItwrZJ7/mqciYQ57GC
yyhGgcqsVmO0sU+eJgx7gCW/taFggAey07Us2z5lFwO5B2JUv9StDy5mhjp8NPtDBaX3AssE7bWj
n7IdNwm3DtAb9a9QxsSOkLTrXBWor0MulqgG87TkjToDZZdHZBrF5pkVc/FG0/meU4RAiIFePY/P
qHfddU0yntaSyLcxf4D53OCEnhmXbtDRifzmZWdK/FjLC7I05d1H0Jm9ASQ7dSlIA9/f6ZRcJKxF
mghX7YWV8h8piM2kaQy7Jlusw0SF6TTXtjtnFpKW53Dh+woo171XROXLW71o5/M1boA8F+i6hLyw
8aQM/7QX81uNofWag4u60A264n1DIoH2+iGWYul3jNzK/C2YoddkJ0yxFzbkdyZk6f6oKQZZjo8B
i8cEabJrwebdmtPTh8MdZfp0QJ6+c1BMrHRxEfBqmIjAg5XcmwN1ErZmuBxNftUNv+2v0M3pBN+J
6FOeRt4J7JzXOZmTZ+ILFzhv+n4u0w+WZ4l5tVb3Vrf/HvgS4EqGgaX/vtV9fd0pU+k70UiRECXw
QwVOPzghI4NPvmDXi0mjxESZS4aTpo2W5nXYauhbpP8yLv1yAYxg14iHl/OHhrnxgDtpNGoCvCTn
yK2IOTC+Fcx5Z/j8SssfRQHEqnuRF/RoeGnLb2OsQmVf8uj+n/abrx9YSAPfQNTuU5W1L+Z7Cl4P
ZYXGedONthm+GgDoAcaisowdvsfRViXiYv/5KZiBaQ55DnelHIk+KPALW8zPDs9zVdHrAAP0wcCv
prNnsgR97H1VfkENvKnq85cwF4Rq1g0Rvsp65qHqmc2pnRph0CFMVHqvpo2Vg6BZj++Yfi6OxVF2
lDWCu6889JjA6hoo5yFBxmU4iTgTASC6EX0ao6Ad3baEYkc8JPbXt2Rna7H7m06GSLd0G9/tESYm
4M57JTNtMHN75V8Rtc2ba0F+o7NuQJdVgjd5F2nI4ZSq9IJmYWnINxGO08DZv7CrN6uoa4gmjvVj
o1BCRKclLPxf7segPsoq5TUSH3bTDUlQAoyfUHQvvxrODyXl5lTEAH7TFe//hgw8a+3KwI7Vt7pO
0othisa8Y+/HEd19CychL2tX4AezpvGcEm5G9XFLoY2j50wxTDEi2gzb4sTYSFQDK6cyDNFwhG3r
7L0cMXW+rVOX813S6M97KZzmvlTnJWEqV/9LtLkjG2+N264W+fM5F4Y8C8ehK2QIBlRr3VVIKiGo
swokkgr/JybZ/oJI5GXKiEFQzaqiNNGQRVfibnr+s5Z7DQ9Y1595gBcQvJkhiz7zlny3GJXLrjvy
lkPxBorJTCG34RCNF8sDaQwrLEzZ6OwiiS8Il1sqLnr1fh0pI0IV6bPkDQYL+3Q5IcitJFzfEb0/
XJFR/G3Muqzw84WpN9JMdoZZ8sXl3WsAz2Tguu2+8XFVigLyPob6JhWpWQcLkfSfXoa/Nff6+vvv
PySlLTQ5z8o64w01AnsLtX7kyV74ZwvuuHdEvUHCNY6O205eCLSVypXNRqLkfJXdR8AseI/GiuKS
OEpMkRJFklYmw62V03phe6qDIpPooJJB9uQ/N6l6zX+3MEm2kaqbBNzpqzzChOYUBb3Gwu3brPui
3rsw+No692ubWglcM5nCqKwyNWLyTDRK2PfxV4RXF8gS5HCyy9+EqeoejTERyn9iRCz1UIkzcxoM
vwabJDgtUheObr86RQ4BfdMCwgq8YmVRNgFJLviQUsDN23f51AqoMmA2SHFXx9ZevyT03ikowBj1
DBpnuAYyofP6QxDbyiuIyRd+a25YoObCyMLpDuspqcNclam5K1oZKbTTMU7Bb7mj2rIwnmzs3Cs2
5bQ8I6Hzz8KHlk4dCr3BZ9aaX174RGhBwqLU4cTIlIJvqJvFqfXfLcPxgCRdoeRgagucJ56GV8hu
6XhWPVExIPyC7GopxQPM/fjTEJno6SkS0bYPsUMhzjnzMkBrFFKFG6nZuXaK2FGBOsbT/D+r0vAH
I1BfmHHE8WzT7nvzkCwP9eZYCX9x6tafMXx8as4xYkEaVUzSvaNT1SYThbtoaH19QSGc6IL5TpCx
Zf/Q8BXhvEa/QTh18bCEv9W0nhjTcbQ6xc/pc8dSmvHr7gyFINf+ZZCHV+cc3Ff4qOvwh2JAh/NI
3ejzkM6I+9WjCfh6Mc/BgsxCdTlED1+ek5ScxrvfZFF48iEzsg5chMxsYZYhNGXy5r3n/7P46Fuw
4WDvbQd3JLJglv8ekewS2ysr7Lpa5DTSg5DEL4Gu8gL0oWfJqJV74RICTBDPYbnd9yB2zCFDjpPA
W4Xs4awgZmZBJvk+MbotGX3mof2rZidLjIszAjOLxAKQSwxmBD9336iA6iGFF/GCTyEdS1Q7eTaF
jAH1HzMXB4RT0pCbg+kfb3UbZ1sV/7NFnclsO3d0L0fnK/MNMcYaBXk3r1iQmToidkCj4DFvfFI1
bPER4THtPi8n49fWTmQgCrSe5A1tifeee30+aMWYPzfWNNYgJ3OjVzVj3q3SNa9bcQ4ZPSYujD/n
E1gGzi22X6O6z3LOEhmhJ1QFcXOIdHVdLiL6tvEqeHI/+GF5ZhyjSbRxjqa9LI8SS0yqCXkXG5sB
o08/YoAw7Db2DA4YNWGWKntYv5OKk2cp/3N+Dhp12jGhXisNxI8s1vr+r5xPOAwwa9uOXCTrbxXR
VVlVixrGHyroA7Us0xwgYh9IJoRhIdzpaoZYScE2lDmh0tVojgEy3OlrIUe/WcLIWhUgizvAAFNl
iFTKD+8afne661BKrmDZyF18V0dTzKCBtHK75FEaAQIaOuRhAaeRp/0n+t2ERQoLi9EZE37p8krF
9hfcOXGR1ly2XvqrPJQ+w9AWNMZgk94X9Jdnml4Hw4zWgyhX8G4yU+35LuiaY0R/LvOJc7VrYH+C
GSTMQcjEQQvDiKTk0VXzW4in6BSAoc56nuB8Wtxf4pfHzobbleu1v8/A7jVGvaTu8Sjo2ALM1A4r
UdCd4owauhWva2WFV3o4eCzvr7LFUB6X1DfH5r2/BifqcEyLSDLw96pYt/mZO8/25OnDQXciTMrw
c52z2lZy3kw0JcXmeYttCUT/StOA8QmoRZqhYwHJibXpZjQ2teT9nf1l7iHgJeX0cPup799Kbtgj
SfPz+MewDYfj4Np/F4/HI8xTsd+NsIvuKLxxLEtfTCsjhVAVw0QtcSQ9dxU/D6MtmTWm82NwPY77
jMkuuUWgQvXKsJcBI9twiOtnwudWm41DVhHznjkPhc/+y+OMO1FgCdtwXefFor/YZhIpafGCAu+7
+Xxw1EMr9/eaLyPFOJl/xx8pVBByi/nVnwtxqJtSJM8Ku4DTVWuseMFUle9Mm3MFEO9hR07aLnIu
lsGBhHqeB2iJmP9Bxktw2FsvNkcdch5InCqUP1sVEJvhCklukhxFwHs49Ovcg4B0GNCKDSUZ69ID
2PueLI2c2opM52yS97xB4obSGQW4PT07HXG50YplWTQwRECcyidMzeZad8xVFfra8b8pL3XcWbi9
ONqsljUDgDJJBe9gZ6oU374QKlW1mFNdaYJQGJeOMUt90pKN9gsXIoJVdk2lr+3EcuwGE0jDtBKe
RPqaFQOfQqyYR/e5LN3BibCDFQBSsNBrhjrOAEQdhjx+ED4N4Pa/TVhtb235vAJZPlY1m/ch7Ewp
1Lgp/qqdZRHR8Xy3+glXhwhG4ch3OVSHr85vCTmZ9Iqvgl7cCg//pFqAWgMAoq5QRj3L/fNh4T1N
YLuP85MPmIXn/NwTjmz/Oha/dzd/4eFy9l5DECEDL9qQca5uiJif/aJ6wrOGNW6mn6RO3TWUZq5a
74SKBxTcpUB8lzHuIfFEjoe5RyDKr6bBwGXbSXDEztAj/HR5i4m5lTlhTXtLsRK2kkdcG9OxHEdl
KxIwLsIl912pbh8ILOR+j5e+SHr1HU801WeBIfZ9GlgE5dcVqxFtdDuKnDBLzGAC737komwT3ue2
KAyjQXTQjJabWE00IIeXhyJPr/GcC0B9qtbbsF6FpFtC58raPg/4qXnQrr3Eey9D8F/EAQOymIWD
YBYjmGtRmBgxRDrOVw9i1zSDxWGKfV4n1s5yQ2ZrqUiprUSpK7ukjaVWWTctEAorsy6iQWqn1NDr
AukvIBz1HkE1Sn7BNUwGp3BAvVgqYMlopaSKbBTfRQQ56IerTH0VoFqWVzFRjv1i7PKh3BUbO1I6
DqsdusG+8O2yp9cdPttvVnzGmUvPV1JQua3aTaxiCOxQRzP7r3KkOrDxHqRsfqYqZ1lWaeqZnmwJ
SyVg7uSkq5k2sYrzD6YUWPqU9o3vwCcMDMWuAjoCUpFE4Iixd8BN+dXeem3m+JmII5b7oIa+Gtd8
2A8qvW/31SCGgBc42CxdJoXxN59pgKZdTSzcXnfmHsq2PFWDufOGtuBn5IW48aW5AHTOugRjqgZA
SInqv+V+KI1dDlhttPogMaUY03fUyew0a+fO3Du0FAwt1ztgYZ2Ps8Qy7MFtm6MBjiid51ig1gFj
RyNKcj8g89yJt9eb/wMyhYUS4Fi9c/Mb7sOWERQmhuMhg9Bz+ntGdRpk3O1gNVTFd1Lblw82D+xL
d91RCAl/v3AQ7T8haHa3ooEjqZPHUgtfSDF8fHzEm+yGpnjFkjaH6qn53Pkg4meUDPpBiwk5D23n
gIQ6zTKk1tHWOEwZwnv5DXx6qsLkjDfgfCFw4GyHotTeW5VO+VNyC07MEqNAEZfQ//NNCYO9n9uF
eqFvFvbHQ0ilk+N5QT3QGvpGG9fSQMJ6Tc7wQBAGURIav2VtZAZbj4kvhhdlvafWPTEA1aCu3HcO
iEGhNCvTKYkvtzVaHlxWDeFJ90YO7GsTy87BXT8SgAtHwjeU2HNOD5Tv/TSY6NwU0gCPzS1NwCRO
vXr55K6PDmIDEtQllopkrJ24ebvkXYQaWY9SiN+WOg2N3HqJ1VWHt8Rh8s2YlQutTXmMrbuHcrPW
Q/5kcs89IciOdEkxBA59EcQKB+W7fSXHRMdeTnsYXoN4BfVQvHgktRuvqlaG60X8fbi3rGks5jy7
I5UbpwmbLgvo0y+uA/FOfe/eoPQrS+7O5NRprQtGOC+0TBLriep7iIixunrQUZBWTfkBgmMwpsZu
jI1H++lS2qcSUX0dOXLcO9qEB4HU1ORieCxpcfbFcq9FgkMM+6OdRbt1ZREhl+kdUGgNnXwqIHi1
tMRJYK/jAqY11jGQEcxmejqrRXn2aBo3akkfXaGambLVykEiLGz6rsumdhi2TI8otJqdUDjU/caT
o5dnzJJYQafRHAmtU4p8rhWXsUfYLtVr3801zbsRidAWnzYU6OcWPhPaDmp7Ek5pIQdgukdjSWVs
fYSfOXm5QA2jkr3JSW5A9iag+xtjRDKlbWZ8eId7m9yg/xR+6/S5wqpkdTgknsILFnz+cAR9D4nN
DaG/6XXHAOUq9clk615TCrNuewvw+phqLq6Ukd0BdX1DVVgw6Vnou+dyJ8vMxMp0Uor+7mticVM2
Al1sMaNeMCA178h9G0jjqY0uqWV6ETjHhvvC1KqcsjGWlyP4yxwINILgXON4EUnirjBbbYzc7ayl
ijWFKF91F/1wowET0h2vcl8hOJ9oSGYJWaRKOKVJPkmxff8eDG9MTsXTXmDTKUZM/6Xuk6hJ+Gvo
FXnAr4j3NH89xg3ljJ82DfhVHC8Lyfh1n94O0xXwiU9/vyLzB4//Sbp/wt+6z5Qxk6l91eE9hQ/7
Ebwaw9S2bQ2h55rMifNy2CoNobEZOVpEm0QLA10mDazG49nlBo8YIL2/7UH6b+/4yT6QC1OA5af2
ra/iE61pjFBA+Yfqe7pSNKlUpxJagMGtCKu6fQLOdMc44NHxVLncTuV31VQSj9dKPpZFZvhbybjx
uzucxXxi7SSJliym40D2zqehPpI5OVRm+pbDJny5QQ8DPAsiw8TDIiHT4YXwTv1Ve4yJoiXP+LT0
QQy0+KD+ypkDZqQGJP1aznhM3VD7FF3wv78YwHgSU0lUsX86ZOvRZ1xAguze7DKVs4lMA1V5Pe88
zF0ZiaxkE7uw8HfIymRUMD+cEYDb0n+AFehtljqu8JPMsOwZtixaMOSZVE+ISf+wyt4mJxKEm/qU
3/+iU2c7BzTfjGyw7GkkqwSULZKbHeKVn+xwxoi+e8ISRdjQfKv2cR8hpv3VdPlQ2VZqwtmg9k88
oOFeW5NxXPUNtyV/yPsWK0GxW2g+Sr3zp9k/jdgrGHhNK9oBjbMLpwwIg42NkvkAlagb7dMg99bX
AhtPS2y01oh3mCCpAiWnrr4IPL3++vFUjCY5pRhkcO3MpZShCfhbV+PEBtDttP/XjmcensuhjQHz
1FXye7WOT2cqyRZeIikNps8119lizGJNCwoDyst4tlu6MgxpD4vlOhO22HaRnYcW61kcRFHGQ+gC
DluxxLFp9Pw/rJSm2k7eVVmEj3H5JL6n9GS4lyjQQM9sE3+ny27Zd/03/vIb8oGeEDIAOMV3kUKB
6BuMV6wZBzj8if0YSMwBPjaPjIaxV3Rgch0RV/XkVUz+UZC5F+ASBNExPSO7GB6sULBjX65vaI8n
wsYEz7YuVQCGeGq05gg2J5eJ9z+smL+TkghbDOZoFdpdpDttRkwpS3JM4ij4PQcLWvMUfGWpgk8R
CeSDBQ7GTNmxNk3p6Q6q03Sfm+2cnlmrH0mX9zR0vu9TvD/uPw/7BpQBJ3kx06U/0H4hC6wNHYNE
DNdoyFBdGaPj3jOee5LGt2PUjwpFnR24sl0JmGnuKWIQhngnp3tcI9tvP+h/Qaykl3wslpPjHCQF
e5KHYSIonUN6oWDKrW1so0Aw51Rd755sYaDFRuQhAQjPwxIz73Pd7OhTKQfpONSMdoaet2PGKtqL
J7kKTtJFVkYWRxy+86yfH64Aw9fkmPV6T3wTmIINl1n5Mwt3F2dwlRcCCQ1FDKPBXWfGc62aun3V
7f57XJLR4M2hZRpWyvL7taLjgzFG9EMwbEYUXzFwTXhnngPX0M7sHr2K1FflcHHm5BgFqOXwFSlJ
TINi4RGwToVXVlgsshTWKkzrLRvJYwNcJ/hDwxC0osO5sb/Hvas/QpzzMPt8/Pp1Ph+NdeMBqYeB
6FyN1ih+HWOzxYXLh9hplE8+zmcL8FS33KpS4sbCyLMHv4Mt0Wj+FpVLu3Hx7JslQtilr8F+iOLC
uWTWeFI7VJKJyHcg8FhyQK3t+CYZEIvzNBwNVKcw3Pz8d6Oe9UueefG5i9ZLuiO1mLm0jclfHlSQ
M5oRWPn2RH0mYNYiruMJULIoKnZMVEdI+nH5dn+9bALHVmBpBwjDHQroPSTQYOU6As3pYcLVn6VV
G0UPQVXqY+vwZSxsHiQb1FWpTObv1YchW59B+3ShQvcgJaQ+CcgpJ/MeGbmyYmZI2j64Wl3cA7zy
dS8qrVxMjm/Iir949gKXge76+SkWisJlim+BLZaSTX0mUifdsznVsyduW5naXkx6GgX/V1pGrZph
Oj8mSWFHMce7Y/hX1Ii6HLzgJ3kGCIVv/87lfC+16+n+vg6auwodV3wTip3uBvmvcV/M7iCkAqNE
tHellpVsL40IqXOqvqVBHIKrDU39UwaZKpa2GnpoDZrVIax7NjRQc78l2vpHkc11juGeblesIHGN
Fks0KMGmVbNloVeOcvGzRpfnBH20bMFcWByVXMJjH5WqTNV0a5TywWHmE65uixnCQ7g3SONrhfAC
b4s96G88bIe0N3RGHD8FGPLfPKtsLltruBLa/57qrmTWM8nWq1L63gYzAP2AuU0EXZvGAkqgzzaY
iedv2iPIl6dUfheli+Agcy6rVUYJKo8TLg/5fTKqydDM3XNAhBW6FGNnrYzxCf1ydReLqX/dKvOS
Fcgr2Qu3gVIT0mZvfXBrVxnFqri9U7BEOhuhR4751rdBczlR+BrekxHG3MPBcrohrUrXzScrG9r8
OdO9KdC5ybbeRMfxZuuVkYbslHnRIUyIkGq1+2FZqROa9VlBfLSHnB6T+Fl5liV1mSAoU6/m4Tgw
5ZwKkV11zApnfzYzY6N+wvNcbQ6+ilPhhyc3Bo8dxB3XQiopow/AFhi+ovMkDr33/6Hch0MDeKbC
A31bYvJYRxIBgDGOFVXwFBPc/qBHBjPlCGSZC6ZdVPFqWZMweZvPC79nj3qWQC5uSUFGDME3kWFW
g0TqQ4AAV8l4IREI2R7/utQOja+cAB2vLAv9v2OQkLTUB9xGT4Brz4yMbGi5SMRKsqVRXxX38aZe
4qX7M0NVTHqh58wKASF3soV8M2bZKVhYm/AvWMJoyVNnA0uM3VIj5W/0Xjf6Rlt9A978ZwvUpbUW
t7fEnq2gt9Kq2ceMbQTLQGImjNCORLQrmYq4aRa8oOKwuZlGpEfYte51h+ZPa2uYEWqHf6XileIY
cUZOI50Rw8YUderhwigOjW1OIy4CpasSenDgy+sZVwnsFE/T2yozZPzSiG2K9+tHe612sOweeZnL
CWmSY1tiUFTHTWywz7Bqx0TDrjUchGN2hT/bmW/CLiKQbGPfvHGOCsraTAgqAUrdJPtFTiLS1l2e
vLdxZMaEvlX2xYRByAg3DN8Hd7O0EHW6IfcULRZwCGrhYieJW2+Jb43RpH4pxhOGc8WsrxzlZFn4
/sqpXejaMYYCuN8To13DxE+T5+i9joE2NsjQccmOMa4hexbzx5cddVis4fd8OKKLXIFkp/K5MWtZ
hiO+fmhEp1XLtPPFgzc6oAHBDdqpIp4eDSeXQVq7K0rcxM+AzqhCnNUGiQztfuJkMyOk4dr5bANh
85ZneGDXz0jhUuxh6IJZOhNvmLYFt7QEnTftkkwXR2u1cqNILxGx9AeFeRycJ+vYf0Y3xZNBhey8
OjH1RcZQAhl/ua7MLGLXJuhgYnml/WCYIzK/ykxJCaldfkRbsS0w7PDQzeTMOqPkN5wRhqrXiEnX
6y+VTWfeLfyHSwEteNZXtoEJegDfxqq56rq6UA3Zq0xQXRK//H1lG9b6D/k8/m7q8kDa+6AaSWOa
h7MPj8vsD34SZn0b9gJzOmyVbVHQRYqDNDF3czd3qZZGzY9zBS4oey+mBFcuK7YtCLVGwFh59X6m
wg3KO05dhiC3rmiIqbtqvpXT6NFgjI459aGFsfrSI64d9gN5TCJTlocU91Ckpi72v8pfcAegNqNP
YKFbqbxhYduA54ay4VxhD/k/C3rue8BFoE7z3CZksTvLCoPQ8XS/vY8CYn2tNkCJ+1/gxrGsGufy
B+g3GiE3Y7TUtwDCTxequMdPqzU1WGkys61xb8JnNCtIpvGm9nW16+l192jvJ2iGrdXUYPBpI8Gr
jV49pfEEs+zlHpBj6Rr7kC3Ivm6lb2ykamwSYrbLJr/bbNMLyAZzHmj3fRi6afaBlTPGBG3gzPJh
IMJdBeAfjsqRjqXH14kfZL9HBK5pSCrc0mRENTInFblhZlUi/4K1SNbtk/1vYasRxIg9I7gIib8K
mK2xcnM168nre5jYhRiPNDSdRAZl/rDQ1/6URtixM6X0pdTRoVca24lFzBhfjokf1E2VttssCD81
kfqgOWBFO+xHXXof0PtfCL84aK5spRhMKW7SzBG1LKDLmjVYxd44Q2U1H6SUxZ3pdfPHHGmQhYoy
tODAoQuAn7ZuqwShn6tmQ2Rbmuy/HTrmwp6PcmaFfsaOd4JWXGt/zTfCQik8sP2kuQwNxVXdJs2B
u4tX5D6oPTCKOMWNDcDcKsyS3eQePqOiTU3F83ff2D0TZQ+0EAx5vFPV7ZM/gxhIKQOo/lTr7lzk
TljGELIUd5+ZIHU1PZIKkTcnj/tjY9fWaegY8nIzOZQVc8xm0StiWWSZwRZnIJ4R1JNqRlvAAYmP
sqPwtAX3lV/9tZdJJHnGrO2vj/Z32N6wl/rN8O/s5JOb07uIK9F3W4f8eMYw/ww4P0vE4sFTNrdO
IQc7k0JPebROvOtO5CWcWwesMherA/Iv7QvTuONY3OhhyiXIL8cx0uAko/KesDf+tRngWgLY/Vf/
OIHkQZhfMxR1DKnd4IUgpNxtmFGNIbW/k0ClbXolUqV8pwSyz4gk0PLOPx1cjOqVD8wV4kpqM/wi
o27jsPYQrocYrSYY3/I40ck5OowB2lTRNKQwBYoFFeiarN7FkJIdfK/RU0A3SDbu1Kp+THUvCtXm
ktgwMipld5vdT/oJax3MjG/htF3l6mdEbPc+QsRu7kjbFYDB1ixfREpTxchLJIj5KGSLPOhpAtl2
qIXEqpHnetalpJE0GtrDowCrmaK94HDtwR5aQS5HYo85ngRyz4t6p7bVGwFbZ9E3CEoecFMFXPcu
q67HahWiVf5Qtjp3G1Tzo4MOE6zMuP5D2HuUpnNAMCOZ2bvdaRqOcmL6dH1uloa5MZ1PJnomIBU+
l5prIix4bFm52iTgKVSoDaLG56vs9GPbA7aZBdlNHDAhNvKE8Nesbh2ZLHd9Us2Q1dUB5RTBNOEF
r8sst+qSd9K9EqatfshxeGAvwoGjLS5H3M3y2PXsNXxC9Rd7IXj9J6HDa6SNKghGk7lUApjxnUpz
XuhlX+nLW4sBUy9wky2hGHUYg5LpIaXhkuV170kEHVQWQJcycluH+wg+HwEfGo+kwqGABTgnRdoq
fCIRjwyiM7Y/F/GLLajSgvUYPQvuXzPQaiiMfNkW0k16ddVcVBcxkwJxEi9+L/f5NP/fO0gOjQK/
zyXF8wzBgO8nqo3vLNdj44kTDGtjXgkgn8S/s6r8N0uraFfAjD/r3Qth1fdEfhDALIOajNANR39g
B1KCG1QwOHaVjLfBuCkg7PbTedl5+EloZ1q6anRkj5jCG/uV2JXMPn9WrK8v6RT4sUixrMF4Zn0j
Eo+scKTFpKuK+ldAnqqhcksT2rR4dKoqcp26+GWFyqwDclXpvwqs4NeSekvcDf6D8uUMFJVyvdx7
06w4NLXpw30ML96BDm47rcPGlcKQqRmHjqznXk/t6pU6knlueQSi92/YkS61N8KhlJViqYHM/VC0
xtUXGmmA2hAqO5jUPDIHlERMS05iwI+t5RPzObzDkF6sT0+uyAg91NdN6aT3savx7QQ+lTCHYYZ9
sg2nm3uLfWjcbS166SRHFhs0nXXu2nqjbh9OCBnsZ+wOsRX2n+cOJ81VAjAMtporgGy/vi/Idc6R
ks8nyke2A0vYQ2N1Wz6DpLugJY9MX4mSrjzl2A/hByHGciTAZlDkEm6kjuf7xitt3YpRoN864wVS
aDDPn+rYFk5IYWIl0dyJvyuZxtH+lDnRICvpWK6bLdN2NK6/cXeHUTVkZl+XhXEEsoZuzLYISSAv
KFEqNABcI30fpUgPTfwk0DeIMqe/Jvv/vMUyCxm2xMRF7vaCocm2YP2vGtkznCWiBp3SnG5YGLHh
SCGtsos2saOQO+vrCsCXiC0zb1Fm2e8tIEC/jTCtvWojnD8Rbvwc9kNg1lmsKhuVyzhDCke2EQey
+kh2RH3/I47sxLbkWE8EZYW0srfzZOaFRg4C6Rz1Jg0vJlbfFdV4hLIrT2KHXS/3kVrPF7NwPs0T
rNmBnMwEf/JfUIzu3jIqLnfvIlXVO5PKEMEpIdY/XTOKUi1TJvY70+lw1ftEUurD7p9Ia5eMcWPY
t1JfpqBRhZIC/Mn0NRgRcEWcshM/5SHbqzQLxid/8nhcd2SNMvLqiIaXxM3OLcHCHFUeANqfkK53
31QkjV3mjj1ZQFsMnZW/otWdf3oeIlO1+quOdpjBEVlDhZ6nM5pwGm2uhfF4rRlqZSs5H512DGRn
Ydh8W/8V5jSz4Ni71P46ViH2Q5qAO+LHT8U7OWUx3vqSvioCDBplt7EoVkBoGHiwE0DoY/JMlZxP
NapJMuzuE8vGoiFFajKar53P2z8U/a7m3SpnK7AQtpQa7dnEIOQvpZpjeVeLz7l55mTeINVU2md2
2yAM2utsJig02223FvdwzWBO0pZjhofMGfKjqya4S1PxAmRGn9XhzaAJ3/S601f/czz5SXAtBr0k
lwwMiXWwj5Qs/IGwcDUOS1zqrrfV62CYX098gkiggP+8uXS6naeIQD1tO6oA3aWvvgh7txT+rVND
fMhM3RCrQGyufCecGE2UZls1eJVIaSsFd2WhAyIABN4PhdVWsI/kFVsLt6vuvkGM0wvP6hgY5YKS
8KebVeD8rVnlCKy8wohgwMaW3Yd9Z9m1vUyqx7VKddqYXnehin/7Q5cXEjjXoT2jc+bRd314H9+h
55J5zVLQr1Wk/IJhp8HfF8siiFUoGPR42fAlCyn7lOWpdDWb+Wwhyc7HVIqC7mGPihuO0a3Q4e/t
Lr82l9YMKwhx6ujRAB1ctTmXkEsDcc7/4i4UQKcmpXU2nrly3mpbItYek1Dro7+/wMGCI3MQV96d
ycpZOiKWiZ804or4L866j/I2Wid/53W07r4v7ToQqxUiu8vLM4BopZ6aE/fNwY0Du3fLNVV9Hegq
gLzEwUpBpVl2lwuIvc/TApXhW1ECMn3VAltfP+S1zZhZnyHCyrLBqvbrIrP2xMQlVW8P52aQ5OFU
4Bb/LIrZ2exYKosv/hCmOf5dAj3w9qWBX/k6AkRPdWI3BNvEA5eX36kRlanc7a+pY+wI5N+rWrb9
UeMqk63wEAiAQF9GCkaeG48iQepQGgIo6C6SZBjP9uDpZGTc4QXjB706szZb5fcTDUI3D7N6zFQP
PZANIgp+FlO8CAooVnLyoYKerOFpCgkPK7eEaXLsrvub/Gai9A7hAM4y4G0pt4WQSEzPNJwFlhuS
NQEA5fokH2+hUHYSwluLlsAWs1xTnPnMKNwS6pFxKff2cP58q5up4S66ngpLFIn3pxqxWPGU6Ecz
K6Mr0SezKV8j3sRDIiQVPFO9It+9Xkxp6dEHWArwhGXA31b//kkwfSR0UwQmOWuCQoWMvcuGIcHE
cSip9QazXaH4Xm0WrOdVUZMovJ4/ELluy4hBNpYm0OgBwGt9k7wmx/pd3uWfexmVGMbfzKLStTtO
MgKiuKFSMsxleV834a9udSieXE5pjfoYzWbHS4gkc/qNHUFtCtTT6iMlpp2052N25n9WDzOSTHow
/6Psriq0c+7YVaiPwRyZ/Zk0ubvNVbnggKLlHGVFhaTj9kGUBaCuWaFEtCqhENgoMRjZm1bwAQZp
TlQLXqUPbkMEx29k0TPDOV9x7FtOdTr8jeHU0bcB8ZDRHQ2LN1GjQ4yZFdLyqxRN8+C58dRv8Huy
8AG45utJiubX2aC8FyEVqRrHzadTPGyNFQDsqekdZhKQ8QYvFCOO4YrmvfOuMMx9/hGx7o3o4wGd
0SoIBHlM5TJAaZ1UeYxD+jMRQqP6zMUfv9ahdvGEdHDSGUj2no3Wordpq3qlg4C5sfaKs2iNqT58
ldmYi2C6fCXF2nU+CkHiQsZPOpY9qq5iZAhQzxpFcmizdD3ZXnQFTI5g4d+7xxweD9YSdsEX9ZNl
rVmui8yr76mzK/07aTXGRYzTZdAawfpwKSI8ZPI8Gkw818U/L/RZZno4+RdF7MAk5sY60WtH66dr
zGYw6Ulkgmjw80fqNY4vUyW018ItUdTH5euaAlKtuGtir+CvhdD62LtE1CScPpVAaXFoHE4z8H/3
X7QChdtTvLETGiY9EA7k5wpQHEfkCCPsGVdBORPsKaGsYeDVnofsLqcOKvECoXTPxo2otTSkXW4H
l3DxNrMCpFITmIl6rznB7YUao1hdcumbmQ4NM/jUQJ1LtexZGVTG7aTIxZFUWc4VzDuKqyx45Far
p9I7MoeSzHnMzl8/CgUVLvAbbTJdRTsSn0S35SAEsHL4HzfJz7XLzu+LBUOdqAXFrlNI3W2JOSsP
fcZjkGjvrdhiRlu4oiK7CGPwPj/VwZkpnOQ1E7NPE2nmEngpcfJ8ZBfcto5FgmQ98gUQ0b5nfsKX
wTQSgf0HthAaYyeSs2SIwTomSxhwY6CvafZT75xAzy7fjY/WpuGr4LTyC2t7NsLhyMGEj17NEOao
BqkHjcs22BJ0aGArWcvKYuuOU8nyKh1XVFI+JoRk6GFviK0Y84P9ETbY1KAUDJlCT6ukF/1E4MlU
+gzu5FKuEC/xr5LcTaNroxXr0w9IMiqqOiU6FNkumuCiaYoX4SBQ8ESXz+2T/bHtqwyDBimV7UyG
XMd6jLB1jcPiO99Z53AwTAtxvgiN1hQPwgvvOYiCUOmqc7Tg4V2Ih9PxK6foMSqR3I74f/zegvMU
gaeyYiXHFZpQrx9Cz/CqOyFL/v80D7jWRIaDgSWHkQ9OaA8tA9x42YmFyBkjvE3dfGP9xbM51Do6
GI0AqixXHBttgGr2kk3fJsd8aCze5wcev9fqpxvYh9smxd0gUncfQwi5B9RuIvAxcby0gRH74JxB
r8EQIib/ZEBzNmGUzZDStuMCMj3vT9VilSJzLmmiKq3owEFWCdNhFXDVNBdPH4WZlNa3AphR3lrZ
1wQRwoZL/Aj066Cvk26d/oiadNzhtN8EN2dADnXCp48cMsTkMHjO+sDbZH6UuJRJLGxhH0Dgro6P
xS0HNZZHsQuLZg9gv5Hq0fw4fzTmTThTi4WSVsSWguJ/8W41MZw6oeQi52fmxgk8I/387T1GsC5r
M7XiL7Erb3FZthCUJHbnnb7k00ok05vsqktkUVKQuB/vJSggbkOMbY9Nu+oKOhVlL7uKR4umGz7b
h5j0Zj48SFFRKo8ih3O6o6kkZ4lf7e+s9nIe84wW8Fy6vl9CBSi/NLWuhGB+nkGa6s1Tm6aAiC9t
CfnUt80RvpWgLdM5e9jnU50WDJtUyNPL7oUdtpfUWtQ/O+I3zsELADe/n1ZnkaClwUDqEFv25p9o
FIzBiSCWC1NDd4bmmR+poBk+x0UMKSHVHLlj8PDHQSJM22DzPTyps0P1LedEp+t2VzaSEg40t0nC
Wsrq7DF8E7lqg5G9/TX4mQvj5Y36r32PQ+eDs2pRzbHTi3fo+K+imhBvuSD+73IOObXIVZ7JDUBb
t87sNyXiiNOvf2gJnLSesV0y/8FLUborfkNBXQSQENL2qkyqgUrEyBQddjRBoPsKNqZ1PJ/ys7hk
Ok6izbHf3YmVL3RFyL6+93Tai0rF0SE5xf5PXOCI0zqQnQMMxGfviww3RCGnQlrkoz6YCyNnj34r
ouUG24oL4WTseLO4/CVtnHG4JtSQZlm4Wzanwg+MgK3lTGjz7MXkkjx+wB8neyT9l+s6qQFvxwkf
o5o4gfPwWiSBGyiEGvO09RLUlJP6R/Ifbrv/MluRxEJu8DuR8OZzfR9VXkldVckWhBj5NfiFl0kQ
9Bcpl1CnbmZ/NifRE7EZZS30PQywsVDuZHozhiIqz/JX4eg5GjQXFjRk7l83j3Gk78s4fPEB5CP/
CR6dL3xjM8FS22xC8QgHoVlzz1qt1AK2k3LYL5sdJqOlEOJJoYzBj6O3AXtzIXhhabCuCQ22qX85
9jj6AgXX9Hn2sTuugtAeygz19EetFa623ZLi4G8YM66MCBDjBSym0euAimWVR/4m2CLGgj0sOboW
yVLqorgl7jsj68n5Fxz6LgKW+mELpRcSEYmohEzbd/HESLqfNpzlYvk1DEIN6KM2lfTaW/6nHWA9
RWZQeqztoAcuT8KOmNwiqNN5oZvA7v+mRgkzLOsjvJVNZzCXBOjaC3edZ64/ooEHlZBSWkWL/QPq
iJs81v+cuJsqNYq73V6aUXLx0JH61lbmZcweR4EYgLAwwrP8N1+VFnfPb1Ipm+uh0JvKrLcVLs4l
71FOub1VAzSRTnOsZpsdqlQp6WqKMy9Tu8Mqm1C8rizaRjgC3R8ng9uLeKmRUK0JzdC5CL4bJrvi
KmZWTvjh4gxay9O9VkIKHnxTbBGR81s5hAuznkOKsM5emomMHJVzlLdfFcvlAHNkQNwV0V3d7Fv0
kblOYrTROXbbKQg5PxxDk7Q7eT24agnwlcGgNdH/Xbvyh7pCVsG7I+cWcCW6Hga8vizOs9m/zdZu
WPFUW3K8zSMe5Lze9P1EGsJxw6YIjZcUXYleurKYwLIQ0hQi3B/TSbDhzuhR9M113X4usAhw6KxB
s3Rm0fNxGBKp4ciCxnElbGD0FIsYrKQ2i+d196hbxhrYlsEEYqG9Bm2lKQWeqaqqaj2DzjvzquVF
630LwcbXH89xQ1K5DxPqfviL9IuXir6J1PY1r8TaRJhQQybEUVwkyZ4i3iu4myp81B+1tEdNXyiE
QuxsHCFsJoJH6bcNaInjXhEhiEraip+0n9/lmEqB0othNgPcTdgYo7BjItNQol5pxwsTMDAoFCpg
ItWOwM2292Eo1Hs07gWokRfdw4F8wGLi5Q9KqTxHVHKdtnONFoRsD6cvgHtK286WZJ9sDE49+Qep
hDiqQjPBfv3hdapHXjgC2aJw+PGXIwxzMVZpC1H1VnekrWdEQni4LUVlM+WMPxLAaRHlzSiC1eQS
AeF6mIhjakBtgUvNXvl3h2xHn1sswDMK6acVL47cX+sH7NukjQan4/gTsqSAV0BmnwnfAAOhslvY
5poL+RmmcPaHnlKiUtY+eR7mQ0yMZ9mI24gzYnTyd9sLUA8zjzJpa8Qt6EsXVRgPW0dA5c9IMsRR
5xMQYnQppqKLfsOOBiuejl1TmGqfAJuVUBRend5hTy9VvdMIEEJpZfo3nkD1tlF4e9cNA+8oRPDK
bMIf9G3IQLu6KhZXVaVZwkuh4PqM0ddl8vP1MFqR34uYGK+lRMJW3yR6AFWDb0K8RNoa0q9TvRRD
eZWAE1PFbk8TzBhGhoi3rQM9S4G7vDSpTJLNtOMiM+a/0F8UUMlX2F+m2vGby2KV7vKkb8IH/Hj9
e8veuefls0MTk7O/cYCdKhKywiiv8NrRI4NSUNo6+z5dLmaab+RR/rCXHU9z+05T8SBo8Ix+QxBo
LL+UnEe4sdWXUGiHDSv39c87UL5y/sJOwbAhgkWiTQPgYThlmTyJBf5POiPLCZuSa/jz970Ll/59
td53150A2usKbJvdLGNwpK4jDOpPuQImg8GHhVtxZJctbxxFxv3fUvDzv3vBAPK1uB9wPDuZtlP8
gyThGfUqiu6kYXMZG/kDoB2jSBW7/UcDxrHBnzTvr2KGY9m2TuFrOX2JZwApe3sgTt4rL+NHZ2pS
yFmdm7xeMCTJfpPehdvBA/myaZ9C1c2TMgBhswUiZYx6j4hPj0CZ8V4ldApoQMgNVKOWHf8OAMoE
jAGZYFqYX7woWI+wyO/58nb0q8R6Ry05/aEPKgcE8Rrjao+O8y7I/KuY3IK8ktG8CldyQa7mRZa5
gBm6A3Ucds88PK9NaaCv79IMoLCQBtRcmb947FdB5MiGulYv1jLUbwcUeUQDPxS+LHw1MUS7ksVk
3B9fAQMywub81O5sTxd7Jn3dHW/6lcFAlNRLXYML000xF++bC5kjNeMxb8MAxyKTcCC5pWPL+FD7
W2kmG8tjOdqRdXpgCai/caThT90fCxd8OBFathtgoBSZZwKFMMokdkETkuATJIWNLjn9HTZ1/FyW
WG6GL89q6lA1P6aOzzzOnU9YXm9ewvFzhTo7SJXrKsliEdUhW1t5vOkBGom4/F4bLrsAtF4ryEOJ
3auywh40SsX3FsfEUYtCqW7ev9chN48TvPX8SBB0VmQhS3LOY622xaVtOPh0dJtyVEJSgfyMjH7S
XJjHNmf29QSLq8m/EpMf4i90p0oMg4Oj08RXACijOReDURkRtp3Tizu+ARjXhOSpVZJnLBJX7FQ6
cezCKMAiFaF/iDsTQjd1mnxnCBVd91qejIMpGyrhMCCJ6LT2r/7c/76o+Dpf6E8Zmvu9PlqQBBQk
NDLi2/o3jaSXU+f1YbGBQpbdZUQWh2Hpsxa0dfLioFQnciFZ2X231ldEX3JXDgJp4PS1bfVJIMJm
JodgTmx0yk4vy0xMVi3n/F5jD1voL6oXj1RH0XvsAoyiF4mMXlz+nQBejZXA649Xfp3vnc4CPhiO
dhQno+Y7Mh/Evsv5ipeNkhXDXsG0Cb9UvXZLAKH/ZwgVXGkiPZHKC/Er0M8wAxWrkps96iE/q11h
c+6BUt6tj7sTpublRrUHPY1v6daz12u5yVFEBxxLHEb0BF5sCqGI2K2oOdEbC0HGuahBrPkfVDei
nzMPi0O0BhCnzQV9Bz3bt1z1RwsGiWe+q8uCgM6AgzxqTOB56+GPGX9aStBiyY9p7Ab2VbIHwrBG
B8W4Oc2ITo3IJuyRVlnO9Vsy4s8mqjEW2gqVpIOP3k3J2XXjEKVP/rpgxso8bbQ91IqY94DWBpZi
JqM1Y/yF3XkDPGBW0cZCBHwRfBh/TAuihxG/YJpOCYPyRFXginx0udkjK2UIBKPoHY6ydxKgWLrr
LzS8o5NmPYih8augOmmokG6DId9QMVvZDtg7GwDwNws+Pp40I4MmhAGLTUujmo80PBeo1WNiJbHD
1In3ENVABKL+vDnRUQn820INzm1I0zwvpZT1OD9dnpGp4PFtqDoh6wilvyMIGUOWkZYsk+iiW1Pz
JwUxp81QvkiKPXV7omK8xGpE1Nigl55VvVT0iuNIj2fREVMRtnq2Of3KOrx1bKzSUpyjf3xTCjow
2USFgMovWTi1G0dUCdM8jVif4fwf617YrXL18CTz21fD15anEzdbY0hcCL6DDvlA1co+puYCgo5B
1xUQSmPpm9ZqDL8KfwKUXrP+GzHdF5f+QvyP/3ucMVZSxmvoJo9KnCb8r8LqXwg6g+AWxFJOjIDN
M36II28APd5q/jFvtTOjOybCtBsQ9AwKBW4o0Il/QyUPVndqjCui0Kq5HUpbHVYmwMiBqUmLuQ/R
OVTYtp2AdjtwGLOgPaydURO6FIy9H0f+hbbu7EGO2gyLBYHmraVBx8+1nlxi8/hXcaV5TU8zgxsH
eI0F1iJ0bCCl5jcfU2uy2gGP9V92u4HqP00ikbFyA5n+1PaobkXn+1PtWXvwT7zSB3I496rHXP4Q
mKpW3a3uzWKmN2jXgLmYoof46razfzefPvZYm6w/ESp4mkhcd15qYA4iqyej+tS53fG/gaCi2JI1
XaDOfT2Oc8Bn1qUSnFq7BCGl7P2BfIkm7otfCX3lB3v7j/TEhEPRJqp3q3RQoulNsvHvYZ0HaOwn
4r0MwfOGKgnmJarGux/4cDFbnQweqfnOQcEQyp8QtTXgKG0zTGXhfVF2l1UUQq0bt6avztly5jz3
uu5kOesX/jsLGt24IZn+ylRKFiduofokiOu4+P3rZVcAzIksG//pLnZ/eXjX5uxonxykDfRjnQga
PttRWgxl7uZy9AByqiljJdlyA+TNvt0n2S9GKHUH9WlJGSbeNCpo7fG4Lof80LTMaotorVWoIiRc
acAaya/9KJN4oDnD2VYvmxUpubh2JBy6qC2ZoMLvq5uCPcvSS6V/+I2VzkDfDc3/71pSGVj/KuGU
L1dVYSSSmAOIbS/Fkl05CXzn4mmwl/MCbZDdlsQJhslHQjPGJC/yr/XsIe3/vkJy6iClw7t8OpJP
ICiZscGupCbhfjIPS1wHeIKFesxM3QHcr7SGkLas/FnI2Sfh4RTd2iTb1z2tmOw/oDGd9odJPJmj
A7ACo2Xt2TPanGpcJviJ05owSX8Tv5XYIXNebw5teQnaBOwBZ0bqy2qh3Ky8ihylxKr5eTaBWhsh
6cvJGTCQ+Z0avVA6ssWzISscQhQLytINIrvo6F6fHMMzNhT3pvr0LqhU9y28rTpwrmGYB9wV8TX/
sZBrlNfaSDQhoc5qe7g7PVaHQSM1+0AONf8jJVl8gI1BrU+ARUSlntSTO3K9yDQnc5mAlJECMN1t
xgoi/Bf1o/gtK/U6qUIrtdO3aWjbMa64uEPa0WhTE55sGjPteSLPatn8Vqh+ewxuyiSJjL0nFb9o
b8EEJiDxViTqeDIRUo5j0EBrEMuk7ZmR+cSjx0oazgvaBDRvM5B4EupSEFvHjC8L4RT5k5ISM4Sn
hoaUVklLfFTKFI00qccBuu3zeyJ9Q25DMQqOta2fGH5BueMVCbOEsbKjyc6cyHSwcDjLK9zHSVVD
IKyIIKoKuA31q1W6SmIw2kMI+S2sYCcOaXtcSu1xtnkhKPCG6lRtcZ54a4d8tWzx0nbxMszUSqc0
opsuszSuDC/hMOUU5xHJ0/UVT2Kqt7vG9+rVo+cJVUe1LLRhoqLrzPa5go6Lrb1aUJxE6DCaI1NN
6cW+wov8AH0Cn9wY88prNmba/kciR3knAOyp5cW8k239kolsoJvQEX0XnB+cvcgHguH3L4+phoRr
SwrntNhqoq6dV7nWqiljD8NKoSePlb5/A/P2Ha/PHx+sH1xt4YGAwc9jiwPnt8Tkok5qTKh/01Ed
ouA1U/g+r9zL0nknRsEuoRBE0a/24pkFxx30073+H8iBSESOuX2wCQQjl1lflTCVV/QF3OTKJRke
DC5+EfvMLz3LUye7hRXXvcxf0KTrzxtyMvsWjHqJT/ZInhoePhb9P06zlfnig7e2ziugPdR/UfeJ
/nbP69K2Ri8W0lqnza/vJnQyzZjT023PWlk1c4b95ytHU8rbF2BFSqESsyGVjKap6WvbWfenp4Ev
zmHmbB+fNyYA51GZOSo4Ki2xrdvA6M1lHjL3xvLYGchQ9M3Z2asGJweMJDBH+E1ctTbYcNxS62tp
r0JbejSZXHgmcxL6VbEAkFSFrVT+FubtbhE5sdJ3w8ui8DhphwOZm0z9smUdApWPBIzVfwVi05Nq
KVMDr2QuUMrDSD5ZIWqWB9jZcmG+M3sPGiLEzroh/QXRb7CChJnjIV9zndUsM5x53+P/qqTKhWF/
LYMcrBUw8JGM5o1L3ekzSctyVuP/MQsDWWAACKNft3+tqCyhn7l2Y718wbGHMYNKkASUo82MFJ1S
GqcZ+tfBFc4dqPSZz0DaRj/VnVYI39GHAPMPj7DLFaYit4piK/BCH1S4e0UkyC4Heu0FwvNoau+w
rnTGOVYyEQ0I6oFg+vDgfB8Kc6BMd/sX2YYQRfouRojfAHhrgXZ1e4THMQDa1EOq8S+egy4a50/p
WS12Y2sIywnrKAH2MFQFVzxWPYtUXTQ4QaA5cxt7wYxTuBjCIGHb54rg2T+VIgHsdHcgbocM6/6L
g+ZVogP4pWb8lHvNQKeBPl+KM5J5Mj0gk+c6lLB4ImpPiQRTcYCXHw4SbjgI19OPWDdGh7j56z3c
Jw+whF+XNrZ4DkJKLGcm5xR1D4IMr9MU2U059f8fWR53q7/CCB2IOnWCbPfZVl/yGTsOYfN0a0og
7MCHMjvQZ7CeOeRdVlDrexHmLnNeCNqqlnxw7cqjzSEeAt3lJPMJJfS2G1up3TVpqhE0tkKeYZPx
T6jkTlQd6n1y+v/lePe4yf73QQwMJApsA7FMskrnkYqDBp+LPeuJAC9w4es1AsWlTu2XqA73mtLd
LybAYjHcZzOncECtFzDsrRn9T+ajBJMUmG5j2w+Inshw/d6RCct5/ABnAJMaxw8YGDZz4WMxLAUR
LL64dkB+qooqIGES+XrU0VJ56+9pPpYeUpfxgcZb9Xjva532sfgBVuV1gwQm+O7vdC/DOYSEZSJw
k+gf/2qfP72dUvriIV7A8Q3TWJ9r8Xe5RyHac/ZNx5hSFne5RlqMB9E/6yIyytbpNRRQFTq3MPMi
3Zz5F2cz5x+Oz+2iidCOZcAy2WcrafBnGgr9uCyoq0YTb7uJUH/7HSO/+LCTjTe2tUl0PtaMwEUh
IMNaZ1mOUTKc8eCAgKSE9l357/6Yg+RFq+NW2eu/C17H+tsWdno6nW7/M8EWsB1V2tFkAjKCSsGO
n+P1YgjszGkeH+7+3TzcaTL2O+fOtfFAFqiVv4Fk8hOYgjxnwKoeCedfZiGTaHPEEOHdnTTWW02l
xpiM9kh/rPvdGJdVBoC6RMzHK0ebEFJAHA//Ylzm8BJqEChTXHpPvQCIveyMfXvxS/X5CqJ2wvYY
2ZENl/pRRW9xbt3+sm2G3Sj197z9+uDuoMz0X3FKGvNb6jq3iQpB5I6adHofRR137h+xt/iMmmeQ
ny0wqk/DAyKNzrpYnd5s41AYWSVkZ03wkLBG2AKQ7QUnasG0gRlQED50ZMYzPGL3s6YANvuR1B3y
JcUxVaEubIuPMRTE5DYiuw/0SmVaEbD+l0NOxvf+kMb9rzrlFql0WAP1MeGn/DrF5sNavqTU17FX
Iz1kQBRPOzizDHdy8DUNAlc5R56dkR10durM4b5KbegCrOOo3bF0ynsBig4jW62M9B+mHWrvDnKc
wzy4JLROfGNU2e1EWUVnFKU790YttxbgmUNkLbbzLZRpmOsPuZOxzNnzvPIdIgIF0tggdR4I48zt
RXFblpygUoGfjo1nHjTKU9KYVp98neS957NRrah7zul2uI0kqgdWGiBOnLO6zs+xAx0N/Js8XgXS
4k521SaJFHz7TCdsiRWXRdQrPT9c2yR7IG/BivfyyatrkvdKVvDGGBrIM6Pid7MS+CAOWtG+EN7C
ERvGHsrHd6pUXsfutgAZNE1EAM7hLAK/FxVCxnoBKAYrUiPDBMm4ghsERpap2aCvyIa+IpV9AkyF
GOHJMFkAKTEABi9QqUB0IygxoejagHVetPRxDfyvEnZNfZGBkjLwV56UAndVMos8t1oUUXZyMmvr
D37V2MdoG+RHrksx3ZS81SC7XgE6YdilyysHriW/0W6Pk9FndtfY+p9AqgEw7QQDjv4ZDfV2y/rM
Uyp1oZJBZKhATiQWBnCgYLK5JwL2IFuNpKekRLfc0OK4rgae2Wg5vhVaV6j64eBLhUCuXHtAtyBx
z7YXrps4KMor7+K3RgC5/ekDoyQsc/BrwexZWpU1oXNRu01fccfvyLI2P+fZtLEqhuaZsquEXc17
glJ861sL53ZmAPANNo56lM7rHYi8Tdp/cR26WqVpW/PjYtkERnSNRPjFETZy/tPBOHNxuW0YJaWJ
f0bL3WqEPivxxGDa8/1pOe0BxHPB5VEOVkp91Uz6srBt030ysypRofSKnEqKvjEvzRICkOW8mMBI
iX2Z3iZhPxmwP8jAiUkWfqB6US8Db9GM45+2E48w1+TN3JB2Z0JwsQYnt1Y38jTKq4Ccgaq0sj8B
KUv0C2gLMGJRBAucQzgl9JK5JZJOEB2HdajJj5owtPOx1/6Zt8tbs1qGt32EHlIusRAInb6fgtog
/XaEQjEDtnbagNtClPnuED63WTpGUXXMDxyoE6MAzOCeUeuESh6Z8f1knPmZTLPW3+i/IitpqvDL
X7NItLy2ebA/HAwtvf3NX9Tsi/r1QC/qD+qK6uB7+r5Xmh8oH8qm7wSRPzDPVhWZK+1SUU8eu5Zc
i88XJykSbasquujg65TCUBMz+6/QaYYRbkib0fT+g8IfUi67344r+7w5+pYpWojh4h4vDbVAMne4
rWVkv5VgJEClYFufTToSK7DYcjShqJvOMWHuFG2gY2z0Lji4aWVio4x2Vd9VmGSW29b3eQI7BIH2
xnvfqZ79jFwOykgbsq7ycXCCw+povaiBkmyJqf02sJsymddtI6zpBLxiARlAFjWfn2AxvhypGENZ
e5pSo/dcmu10PXJRyA+oo4j3BOhBBcI2L8KzT85anf0ljfx36zL9aKRkl0eMqQhkGihKKWqL8IvE
1YlmfiB7Tywz/+jvJjE5qsFKnI7rqmELsTqv35g1xATyTVPn6F6uZL1CSrySqCEQWd0LxL87sn+o
MkUhOPnW9x4yzud3KhpEKoVbwJF/HU8481ypIWlS0yErZ12InIUs9RKH/3ITN1R6u2BOvJCiLyMy
lJvVtu8jPYYUcRemPjfRZejI/ealhU6u7WQZY/0IyiBgKPmohjSL9nSaEKJIoqT5Ga9AWwCd0TUw
32eEqy5EpVK8ZWmIJSoYEz6tEBvl2Qmks9jk80mf56a5Pr9FBfX+vDvG899HRrNTLSsVx7W3Gifh
nP+M8sfkl1YsTJ45BjjBhCym3Gtm+XJBFQnjGXCY1oyzGfIJr9OCZAI3iiXSpcO4CRCHnBYhvDN7
7PECaHSZolEdOzrI8rD/wcUIgL8j/z4h0zH5/+kgPfZcHyT9ki3o6+7Z7fSP4BbmhwQCTA/5YTvz
1Us5JH/g9l1GTGHpoi+jtTxA6DZaLzfao1Jmzs3Ae/r0Q4cf0KSTV5LdPVqc8xF6BgJDL0cDX5ck
6WEUFqDb32HkgjGZj88viGFp4llozjgKlZqUgXVb6K9RKs4fjAX4CORfHQZK3mZ0wIjpbyoPhVbm
2826iJT8OMdLDcBQOGEvqA7c0+YIgdLHIKoYwShnKSU4fnz1aHOjkpHsAhg6OgYj3SoeJZ54itAo
K0PZynuttRvieXdSIqjCRiL224g80r1K6iyWSDCSF1N/bDnYSd/TVdmMgcsON61fkQr3oOXJIR+a
+9VvPGNsYzQbhB+r4aprdinl88Acv+FBIb/jLHGWTzG6h35l8eTvced3IqPF9k6psScvKIGLA1ls
cvbiadajBH+zdJj1h7Ep/2sfRU9uprzoQdAB3AsYCq6X4el5rb8p2W19ddzNAuq61dzfeoStXUaj
Pmrv3/6MjSwIbZ2PAtMZk4SIKsWkl1VruTh9ljZfNSsvqjIS8rLkssoO5GptKObtcpi9eerONUqh
On4J6kD55HTDJqDIyof27xrKEj7ZRFLHotee55J1s90uU04zfuBmCtF4P0k5SGrX/AgUzPWTrRyw
JCn4byAF6aSWUo9Q0OJ7Ov7qP1Y4/bQhQ3CP8gTYtc27NrZ1hE/xkMkou/ruDkhfuiLPb6/OnLH1
Jj0o3tXHm3pEf204OV/D7Gy/FG8MRv7rcKwqyfRjDhDdwrFbhRNT4AtYL7yjPe4/GBweGEwFvVur
x2AcpeL4TNtzVrigc5vNuriO+x4m+kcrUOoXt1nSeHtl01eUSbZv5zl5f5sM19lIA/rII1UIJbGq
Rt5aWA1PyOppRcM3DJ3Rhzj7UU9YeZNSFHc4lsmJbPZPz4ktt/YBb5fIeHBAKQO4j0utL8AL3wJg
5z/GWVjpVboHTkIQgRVAZUkckF1QViwjI0IVG9JRImYInFSrJvO4+d9PQp6KYI9sUluLheS2YOEk
/98iA1wyvvxSyXAUMcz/X8BElg4dKF/WknHSNGjsDf1LTVTzqCYlI0QwMzKwowQW4/WvE/um9y5c
hUx5U6+6FNluydzinc6UaYiYhnEGWBfazqDKB8X8jsNxLFiJPlCeSY6yt/tYaTW/i7lz1vcqB9fG
9ofr1BDdAY1PaYKC1W3li9/+UXRbOLYyFZ1n4LuqHTlB1bY3S6gWr986x0ZCys8zBFU8XeD5+dO4
Dt3vwU7pNnBfRaqW5qTjrffdfEeORNKiM+/tNUgxD/2RPxSETVJq91Txx3qaM07WNM1P0HhmlHJA
aPVMd2HGiLvmpIM82lgYJXH9IGkvYgimvESgIHHn4/9MGxUWVMP7Y0BDPlICRPVClz3d8G9+5Qv5
TDVAwEPVrfOFRPhG8cVzVWiKHqJs1JOTb3S5tfJmX9RIN2qfhd4Bfnw/53yCXo32vm3RjWttR0eY
z0s66gqe9l7zEL1bV/FeDoix4WP3iEVztg1CWuaWcawwumHnPXzbGaSwFoIvDLc6qe58lnObTS6u
j4WsrdLlSBsPg7YkCL0O91LxJUrSKAuV90nOO/Y6eEFBKaQY56hJH0k1DpzDkd7x0ApBrR0hzTcL
e/zIjRCG+hSD1EEob0YNC5RgkxFt/c5/MY5Mjp8s2BbaLqoi28bp9uRMDRsXFV8V97p5014JA6rY
oSpfEvSQoYIhhMt905MirU9zq5+/Fg+c4MTdfo+fIKXAcEyqX0fZXGbyfh3weW4gdKNiYcfKsFsv
9P7c5iXmHb9UfSPF0fn0pP+sLJpqGmy8HwZwlW/fcPnSKIOIBfRt761B4O5aKiHcaPNIerzQNWVv
3zt7ajHDYDrVrZmvjPoZnLqa734/2ZPAt9XEICM++wsUyeou46PSpbMeQYEg7u3eU2vStYEoM/YV
P7nqgSYasrMxT3UyhmR+V9QU7V2kXqyNVw3dkizULU7fzduE9Vc1lbQdKqyGTw15vHL8OwKKl9Qf
rNt5fBGhR7wqGbDutuptVIytM82Z4p9tRJVlmmDNnO9Z+RQ1zcbvyCXGsKq5Iuczih2x8Jz75QW/
xmm9KAojZaUyhWloZAaA6g1TvZ5seD0o0id38AvKvaijYZxIZN74f1sVZLfHQ+756L/NmK3ZNq/4
pec7Cu0Tezb6ESLLo3lHC/ECCS4s6m9MePWXAKVsBsiSZ8zJmKEe7Bl4q0guv3NiVqIJCiUlkUhj
Udwv6ljcgkzylXtEcslpVIqmddW1ZT6deUDTy7hG+OTDyBBt/pgpuX7pvUW1l/pCStIyQraME9F6
KK9S3n2cla9MHr9z0EmDUoxuBNXcDfGxaci6PO4NqT0MfRSoOA85Q9iWPtNdJP5UDyMmwxDxMsx1
JhA7F4g4TceT+U4kRoK+obuc7+OUamMiGUjHs2CEnDSJhhTNT8qD93YDOK7jozoafn/Im7JDK96y
4cnrSeCHdykx71Mswbtu0SdbaILc7918aiuS7oMjTSm9gGwz+7PMykmDjQQ/Fj1Ilvb/4WxiyiUn
kd4GiFXu9WFR0SAQIBTNMyT91Q9v1465S/eH8ENv/zE/AFFWNoS/y/gti2YicFqWlqER4REM0WFa
vdj+Wd1QmFjnShSA55lu3hA9b9U+8RpKrENH8G+SHZSpPFn8xP+V0SYNbSC2PuKUeaelU4jQqxe0
HHlVTy0wnWUaU4mN5LsRjPTIwJRCWmzRQ7pjH2+9Fz4uLnqWdJ2+uRfGkMXJ7ii7FqNxJpGrQLTo
lWpvG+dFunMMUPpTWWjdO+ge8htvKOUM8Qtq6NMxs9RZZ2OWkE9aFj7fVHeta+zelQYFVAvrqZOX
iYHeku3fLUujObpOcDLLynAP4rMvbiqFQX0fLTnGSm4ROuYjYbVo0NSP3bXVBHPffn1S3O27RubQ
uRzDuGCLAUILDvE9O3kyfNkSPWRr4urykcRpgvlYKgqeirTtUTPb4R2n7PCn2UNSKILR6OQIfL9k
+wzBdgM92RxnlAgfMtNtdC9cCUZ3k3LmMduLgJ/N7gkTfqOLvImUGV4jXWGY18p+9Tsc/6bIEszk
gcCxUwJdwsjvbaNHPc9IrIKEGU6/9Y/6msH1+uQimgkjJfPgOD1kRD6atVyUXuZ47n3bw8OmeBpF
pRGUD9o+INq2JHPrQXDx3fcuEvnCXvMMzSA8gafMCSffOi0bFQlK/Qs0m22/BpTLLL2kfvmkUbea
OoPkUPZkNmv0FQGg3S1i77vM+WPHob95+r/WQTJg3GeQSos4fMqwxFIl/rgShu8D1bGFf2ULeG4b
Z6+mMtnmJdwYnfHFefaV3c7DoFrxgn7umY/tO3gUu/Fg8l8PzoXRs7eB4Ay08f2gW573dbpR+vOH
A8dSMVISSniKwrUw1cV+pfH7Lmo+dyH4Kq11izgsltU2PeWQ+Ks9ZauYkl3oWe2MusotgYhHExv/
PSSWUoTBAWy26oDiOuZ0eZXIft6NMhS784YbJtZ8XeyUWN6khwKz5uSTknBpB3/Hb55tH6H5U0Qw
iuByVEN6lvI898yd2Ex/36pM+ndfbggvZrFML1jgWZw2cbrG8WHGBasTikkO/QztxtwFSiuVK+Fi
D7d4kKCsfxZroGneNgwdJPqbYMPXXUarjB1iOrZe1Oz+gcoMrSTrAZl4blYNl9Z0kXFg1kf/HqfA
oy1BdATLPBzKOO3nzdUa1vrqP4qoa0hSEqxi80n66+JadPcoy5IyvkSfdzCd9QT5aeRTgLvzUGeA
7MqvxN3GgEr2BYdXIdM3rTzniyZHfh/JdU/T1vX3nT9N75gqsxQ+pufoF9JwxnEKyWXdxNkKnvH1
xT2JFqcXs+f3nj7/HYan7euM3usX41YLgelsFpov8rBRcPMH+TJd8/sHH63EO+QcXaLWLtGHwyVN
Nh9TSqoJ/BJ9N3ELWiOg3mgbtQd3wJyk5/yO7o7E0cF79Qp2wDZgIv6nRK12bWMrCFviZGmM4JvU
9NeG3diC5vWH8443J/xp9KYLZ12T3GVXQPkd8rb+7RFBbLZX1dtza2Ia+A3xX15PBh2isCWIpEiX
DfgVtkhdFlJdhBdgUQFkqA4lXG57VVfWngyF8N10PybQypIk3Ogor4t+A52nS3cEYCF4dEht2nvF
U+1lI+hddCoJUVlp5Q9GGM533pxx0BC2E+j02u+IVdtSdIXTHAeaAseCCKRKQZgtHxdM6pD8ZOJR
QfjaN05URH9AmcMqk0Il9oSMBMqtC09HmZIfcGtTE2oVJErfQJX8O6ABmImCaGTR3jOitCufjVPv
A4caL1VoizZ8pzuxQOm0gKSeF1YSUSxOeGicOuEJI3D/czYV02TRCDO+VM1Yk+tvp3nV5gieLsSf
zIr5d0w4OheX+vh28V7DFJ4igo891FyX1T83Kgx3z/76gUpDdSJiV6hrJ55iZl2jhqdAOJElCh9L
2Lj3ADnuOEXBK7TvfzaIBoNWdzwjZuxN29jMA+qFz6P33hZNOEXzWZ+DTvhbpVehtRTjV9Eb7Nd/
xIq3CL+zy+EPbwVTPa5Juz3o6Ky+EgEsthfbXiyF7tJ+LtNOH9TM9aEhIRTQkZVnIAsaufsReiiq
OuDMFufM0TVdU4HTTU4X5xYY3/lXlO3dbqZeRwLvCRs1srxakvXmFs9Q/+RnLsF7AQMykdj4d5UT
xWJ0/gEOdAft9Vp+Q3iHOmpDuLMIcGD3F5Huf3Ku2Z4MXMzR0A1Jm8C+nAWs+p3uTbVvqRX4HzCQ
DekeUWpQNAN2xfPqWWhaVPLe6NXvGq53r2UdiLSHEuepQVsWnUvL0UWSi7YZcYGDgL+dm1XOfUbp
K7qcHxTl95M0KlRMAWbzzjZIrfa5XCYn2sMa/0LzpgX3ODh/l9CFt3mv1CYKAHSDrYAB0yHslQX4
EYYK7DAAYztrzu1v91skBahBDP+X+zTm55YKh3osiSkPz4zcR5zBvhSdzdK4F1n7U/gMkMDMIniG
BwP3oI//Z5AY+PP5daQLTGUhZMs2mbD+tQgx6moEJRUiN6bfz2zvZcIGO19bfbySXnP1+gFBF/vG
sp2BtIRVlksXlmsZFN2NyfOLCaPw+3lYno2B0LNNp4PLdzgaRJy4JbJzD0V/Zyle8tB7tPemugoL
jND8FTqEg+jCa8fvmjoOYrEmxsD41O9avi+L04N4t9OllcQZqyfw2D7JPf7+AdLTvGfrY8rD72uJ
9wkeOcoBjFlo15R9UdlX53wcOteqUG/1M5aDMfm+JuKtjaJZRPGsHDUhALEtMBCm6awAXpzmj67Q
nnhm0NZW1hZnJEht3tEwdxFUBCCVyKzQUYFDO/iyWPQMGsotBp2s3mG4IOpnYiKzc5FEn4AuTXH0
aYYIJkoj2781rTeL0hmw7Q63QGptDSA0qeqvYzAFKMuglGLL52hmDAkxKDTTwsLsJFd26aWBbb8k
PdxSBYJAYEetfNsM2unWH+MJGDbvAE6AyLqUdTD4RFBY9W2rxcuO9BKx1w5VZyXZjo5wy7r/cowR
Vg1x/0ZG8LAo/cGkatHXMiZLuT24tXF8hh+ySPcCZotOmoopTfF4eg/VjP03j01EQdTqCSBARoem
wLpSHu3fu3eGxZ/EaGyNdEpy6bWYIiI2+7vWbJDwcZjjz+kl6TyCb52CFAR+X1yRZqo76uqdLxaw
Q11fwwr4EBj5A2F+WstzGdJ/bpGKDpF0h01IVC14un1xNIS/J2gYJL6qP1gVU4eQAgXUp02owQoP
QYHjWtSnQB2JSKgwXV1vE3EFzd3w2jmwZI69Qx1xYwy25Pms74/jo/10jZroLBiVlkBzwKEOhC0t
HP3+m+2tLyoj0IqPbZdn2g7Xky2YVzqXikRw1fgVRCiK27g584UE3ISKU4kJC7cYcv6PXvYAf5AN
50Ki9MHrdVFpiE5PG1OEVJrkb22TXTz5RSXmeIxYP+AN4nigRPY0Vxd9UH61wvgJnF6mjoCI3ytS
VQ1bST7pdi4gxHegq2yB4HSsgSG/PwSyIchhWyo/jPxXt8xKDr9xOM/flGJQzal40lHSnM6iZzuz
oTsGIQpOczboIsR1MhDI4kd08Hrk0A0nvFPQPZ0Cao/wHMfcS+N6MGL0byLXb1Z0GNUnWLUpxSB/
eFoAmBI0r30sQcg57ZqzUm6mnQbcr36L534Vw1DgBtw2SnicghymBazn6dsoSJnFdLfWWF8GTTex
ZPQ2aMtWVnuFnGIKFy4XunZKcPhRUVyj2CVdAy4c50STRyXzwXaQDQHVkJ7o21/ro2tcSSQFCfiL
8kmDSjDM6c+wxUQ6H4SdyGu9C5QtQI5QNwiQ15m17nFR3Pa5LIYKxhxhcE8mzI2cLLukZ8sSX2Ui
rjM+Wab2jkd6eFKKN56Pc6wILVSmj94inOP72ZA63hFaGXTsfWKld4huyMPMNYR7AMpMWJssV8Gp
Zq7QQovo6LN5+DVCTl783QImtAMU6zM/4h/mS97f7H1otcZnQFbk6GdH+ruRyAcLTIoLeXKpUwC3
tif+bv72BPj4cuPk6l1Dp0H9HAMWKd5x7KcOO0D1WGvIS0rCNSq/UnKc1vQc0mslrdJ1zUImF3oS
L0M3xaj65HTdRxxdGbC+iJStTWQDC8HEUDI6KKJGnypMUV5pOvSD+VMs+fIwrHjQKPbTG0N79RNq
qXQ6EQRUYOGEC2IFDPRO23G7f0DtK7qOjKeUNsT1qFYItbqovw8HSioPPx2iGu9881XdSRL/BZ+X
rkbRra4KwW9p5neSvceIAmyYiTFwIKVvgJlgCrT2Hw8aVVPz5t+9RnukNg5chqHi0MUK/W+Z8UUr
gsUmW0+ObHomxkTsLEImfTkwbqappFurQPialLDNqZob8FeeLEP5/aUvB2GYXmeHrVUv2s9kenzX
+zMnNHS0VRmf1spv9GCwhPtfzbHoJ17VYxA3lccCEBCdFh+9N01ZPrLpHEHJdFxJjdLTY4OemEd4
2YMxhf0h8P2JoFutnXJFoM7J/o2+lhRrSShpZAFIzaQ3MhJvmOTzYZ9DAXEuVXKXPl3ysnjIgGH2
9DZqr0hFZb62KVxDb2Xm0FuacF/aXNuGHH6S4yrrJxGfjvaMRylw1pX+k4Cf6iSciXCQLkbtCTHW
mt3XnF+15WXknrla9vyL2PZcDbTKBeac2YFXxCnkH6jQJMYEMHZxrJ1MQNWztGVJm8Oml5CxKTTR
Bz5LzCl1yPRIwy9S6ouPcXYUGgkH6XSw2rB6GAMCeB5XtwZ8YeSDk7bXC2yA66gjLBy7Te5fe8mm
55XjBBJ9jkK0facZTuBjjS3JklPN9CrY3GHcrCYXHbOs6fhBbRn+1laln0h5OlS66LZOP2JbmxHI
IJUkZH6OfmjnJqo2pizOpcp/hpW6fnDCnG4KvK4MeYdi04GGTZiN212tNnhDMzTBub43NYikj13F
34bK7dKXjFBkcDAFh43p439QiJGxUIzZnoHIkzVbq2IpeITZUi96K87LFESqDaUnckKx/CkxaUA0
FyhgMHMMWBjkveIjO4u6qs/w10Xrl9qccgwV9g6ad5m8G5dv3E9wRf3waZyZvpcxM6WboT6xhkuT
8gbLEtCYkKeoP7Zqr2GqeTS4uLvwTFufC9TxKLDVHdbqix+cFJjZb1KyRhzomWI4ptKyJqMMJjUe
JCMG2ru5dqzMKSpEK6ZgoyZHlkSFGA6KX4PDmErTjhwD4M2qSe3c1KgZI5pIzEU+wUzq5mbRZlr5
dqpDiXvoBRRJF21T9uYJt3zFBTg1roRtvzGBclmOuolPwSbOWcagbbIMIrbpD1ZqQXyLLkHbNRnn
qZQMLVy3gj62pK+M/w/9WZk9Pp4YBQDGON/Xr/3xQMIn+XV8Y7sB6alRKqk6IC/iVcmCx2vEN3rq
fq7z8MMC2qVafyFVAfnEUOHwj/QwS6bB1AdK58O1MrKN4GcrHcgF5Q7qFhQIZllz/ExDVwbp7eWT
vuBQczx0OjNVZH5Vx4e6hzz6gDB/Cj09sA0TNUx+SKurecuiACjy4Fu6Idk/DCdAhvLtm9oVE1xd
dcfapE5QYF0xCqYkV/G2/JFXYuhq/Ol10xZtUGbWKq/vh9WxHgI+NsoA3UtDPaK0Lb0EYHD04af7
bP86T2aHDBHNA9ROtVyip6BRWa1kpBH4+YXlmX362y1ajISRK2+S4VAv1kgU/czfqx9NVsQvTm7u
ztoBrH1y25B9HzNUzWjMFbeG/EQmL6ytb+04ayb+y+G7mYSoTsuFtt6U+izhb8JBhTtmBzJ5hx20
kEjnwJDrOpZ0/HO/vKUFWpaK1URPb9jAp2aatOysKH+lOM/zL6WbEKwcAL4otb/EYhZWdCRhF5Bs
Nt5bBpeioF2xjrrAYqPyg21sx435y7j3hDwyDd2dtR3/WS8qDPu3oX5wGa+6FaiJ1Vl89U2Gv/Gw
D2q9ahz2XYYDHFthHrA+8kzP0VrJ4BwQN5E9kVFLVhLvoHzsC9pIBWBcHoyEi2pZElMHdqaxF2TA
w7fj5mvp9qVZRpnxISjtEPwd63Pr2ZZ0om0Fx7TT7hEPA3Wuqrt4KOut+13Kg3GE7jeFt4ue/j64
brIjKlWkWaCj98MjbY1DFbiiBGYGCQCfkRZhwdVH/T9ygwAJBHtYShUxApboLr7N8jIApMFqIAr2
fsS52yCQmGyLh3/AiG8u+FraWV3Y6OhkR+zRKQIRxFIroGTBSpAMTgO/v9LEnVbJHsW/bDaXIJOu
JtMien78/S4TiQiz15zFv+1nbooczdhVoHRJldZozuxpQKb5emC9S7hFFhFJM+okgyCSVzlmOSam
rrCt6fO3+QiFvj5nBPXxlQ/btsAqdX8sxu9GN1DiG1y7JUO5P6hwpw6cOYsjw7ALJAWgyXs6mhoW
FcGFDDo7+E+EGlzMrptUFbnan+kGk2ETLIao2TuUCtmSpXcrr6c0d6Op8MmrweTEQuHInxnuGA6G
a8aGiwNrzRiefJane41pOTT6Zhfm7rfwe3ToCemtwBXpOLDZmv3JqfTvR+zVKZWLqi9o1H+7uIH7
Lqf9Yb9tQloxl3cgw9utghaHnJYpGtd7rKTSu19hh1Ls9nYfujfAtZAGe8VsAxKwSHxK26Ix55xq
gAfXyYJsz6k6S5qHHVx09GJeOsMYxOvlD/h4lE4KY98fH+rhh6l9NI1dkKyyp6z9k/IZLA9dBqBm
gGrkwJDTx8GcnIR8Yy60GU5CyjHR8btkOXudW2Th2t2vVPp9KNISZq/Oeh8j5HQW3qP4SaiqHeMd
USV/oJ4majWQn9ksqU2J+H3hyah7onyZsall1a/aiDSVMErUwjpGJ2AuShDvoEqM5kmg6mAQ1oek
0VWxUBg0tnG30hUfj+0X0zbMqAjfkFu7sOP8Z7CznkZ547AKfIkScyNXDxd4y7eyFDWvmtBVC6VY
6iIfs8ODrRRKpEDIhaay/9lSfGFgR+1xRhUi7uaEAWJI2XWmKOZOt8LQRWFQV6IGjmp58WcbuTvI
edJQSmt3quV+RkfAk3SQjOq+k0yXRCBXzPed8Dt21CkAWdg9bwzj4S9+rkYirYR4D6r04uOSbPer
Lkit7QZIqfq5cuXLQXkblQpaRz4Cauw9jkKhhdUE5JRK+3TQzcprBYLxsaXWxc1xPNImBWqKehSK
f2XDBlqY9F0ZsVN1cfPrBHc56iGWbS2sKh9Z0svhmekrWbRG7eOzMSD+NXJS3dX7jNgUYMn+OE9J
NZGrpukyeUEHUQTvU3+6PTymDUfZWBupi6iouHWf/2XfjQVj6ueJ6wlmq2VphAv9rG6BThFANBZu
f37w1D4QBPqGcynpEaEWvqervs/qi5JsQenxC5WJ1x7iB9prxAFRQz7UzHRV3i1cuPQ+k9XERL0u
aQCKSBshpj2jtgOtf7I5xd12Y1pwlMxXo/2rfMgBIgVq5xAmI4+yqleLH5VBTtMA+LNrvOY/p5ir
NOv5IjbO8QB8pQv0CImOnWbVa7pphZ4UZjWpxTIGI5SBksScmLgAX8l6PKEsoY49E2glDPHO+Wum
1YI0UYghpEyLPSP+7lW8lW1dsnjy+KbiVS4Bdv9DVm88IgEul5svtxoYyJM912vRbR9hYPtlfrwk
zG6B25WAQg7n13vvKT0ZLL0UGbAZX0oeTUxGQJ9zug+PESnRO6AQErobn6brgw1elEpkuxMAVDqW
tynWANK5er5ZQPIBEE6GN8mZlNJJwwUtqDf0ZOWMpAKk//x0jXdTi8IAwQsBXkrQcBCE3k1RYelf
4loP/wvnJFGVHAHkkXQZ8JYj2SqvR+19eO+T7Ccu+M4zgHRkLm6P7trkn9r4AGG65ekmuUpntaLW
x8g76h+W4L6Dg4imJKNsyGrRJpvunyazOnjch2dCNpgUT5FhLdJjbkIBieKpGM2p9T95js01BYPO
ddDqQK0QkbeKyBXQGkUMzAEa1td2255x3w0gB4IpQYDRwZ+r3ld4VkCCvlLQx/ojQjIoGjP6svAp
NjA+qJt6FYDK2xeUC8IxejVEkA7/KjRIZHzAlfWdO8wtlZ/unmetL6igjPP38NujfAis49QpDsNW
JY6T6HSiwljanpnU3UdGFXykVX6FJ+ZvKgBxZauJpF+VIz27cjh2xXxj288jjQrnV47ev4YF95cq
8AyJwmwu0Ow50fndA5YMt317/1tNiA0FJiyn9D6sA2dVOgW0a9kN3B2XCxZaF+QiourEHL+mh+mF
Ma2GbXeSK5obITqJtTl95W8a6OJFs53wkXafYAlEdh0SP8uUAZxUkR/1rBJUQn9hKXcHDN7dnJxc
n2q6Z9v+p+p2ZtSF7HiJrPZ8UoeUrSlBwoCmmLAJQdxw1370OAnF3vc08MUmdQ1QOfyJGUbhQjqK
9lIENmLwYu20eiq6GaAr3TRXmsk79JlwWWSpzT0iOvBxE0x/y8s9/auxbHkRRurZY9ZolBSXM7Oq
/1KS5trx/iZJrHakuAnX/Buz2LspQT0DqifWZ2+v0AIkwI8P9IJft1Iex2+MwNjIZid+uMh2eSoW
sv6ygMzW2ziUYmptZhfn50rWArMZX0MeRiyyjNSYXg5dy1Pd/uBD2mLjZNOypZMqum5G7nDBHJQ0
ncc8egQtcOMDVjnPSn2/EnhEhEA/RRQp+c3iYrv9op9rflG5E5c7ztUa/hVXxDdgGu/vwolzLbvq
jDKt6s3N6ZxJwDNwX8740N3IvTxk5HF5cUHu9miAWahr/7F7uj1J5scUsXtCBHHS7nOPksK9efgr
Cp/xD0STJJLOhr0yPovVHvcVtld3CCjmff5hPZuGv5PxGAYk1irKCeYi82OFPuQpv5dMpAl2e9Pj
0gt8Rc41GX7OCDqTFT5SKIr55JHOIwayeG5b1n2YcbHjvwrCE+SRlLE+SCzv5PM8Wf5SGmNyciGs
5vr6tvKWsoH29KEa6KtDviinIiyOKA+2djwyntLo1GePZlRl0cdx95dz5Rsr+/cKgHjyCHadWWNg
7hn1Il6oCVk4PE0IwnuK/F43HJrL38Ul2vyagYc2xzpRd6u6ekP3VolZvRkkwomz1mja9OESw4ve
jUxHptCilrcwcBqDialV6IHPPVrWkqNxv/0PKDgxMe+BkwPMy2xgrNIshU9+NK8C6yYAcEiYnSY7
V/rQn6MkFkFd/gjmSHzUgkGAFqvAZ3zz+lxlXLMhlMhEHIRl3pzWFbL+315a2EJmxUjqDcZBT9rO
5c0UnueBiewPPxlIeh9WlfH6DRtVBJaC54hikHnTR63ENCYgG9Vd07r7KiBL6pYkAPuhCrHcqPO1
auyZC3nYZYBDRvumSjChzoT8XdKFozInmCCw6/KSaRz8WDGiwpm9MIQ997xbX4n26RS6C9z4ODMa
K6ruCIJkqoDqIEwcV+CBxXUfNFAbBxIzbE3iz3CLfRuBuejRygVXNnWD7z8gj5Mcpuao7swGgo3P
tfGdZLGRtSlA9RJX+RPHoaYmGfhfyAbOojrX/lUsGcr+Ssiklji7FIDDiyB/S7AYWkVOjHyxgSE+
S9d+yavLq6ryMrj55yIilG9Is103yNoOu9atpzYglfsH+nOsbzYpbLcDoSDrFvUX7tyYu8YCKwhu
qsJZbDcF1sG7IeON4QpNxR16TYDofSVTEKjHgNoBqcpRtTcNtclNrvP9K0Dvm5POKw+k3B09Tzh9
fwfLdMoShU29NvsX/19NG982z8d/ZICNyDg1K3vuJDBYHwg/YRJEwTc8RJwUKHRm4DHkLg+8cWTB
eziwVoAQUJ9D8dqoLdgHqSolwwK3kw8hTQWh81fBrThvoZh5VnO2RphmJg6C2MA8nwlMb5ZfCkKp
uxG0kvVciurvS6RzJW1IAtSsB/p10odI1a1lIx1O4ypghlzwE+MNAGUJrOnWN5E4yhhIDjxGHJ0b
aTX3Ke0uy0oUyAOk3Bw9FCJOAHuWANwS9GiDY6puHv+6dUnhK7ADti9TAhYuB7DUGQXDrJtX0e+y
cWZavUyR4+5NUV5O+hq1UCC3TPhgAqMYoDHRS46CtEmFdUYjdptxKcRHmNVd4r9cx5la90v2Gi1J
YDbuwCAGecKH5szq/Ff0MNNR4/bWGO9f03690eJLiThSegZx7I3q7Fy0HH22XN7z05I4Cd01ZODx
KVOwe0i7el0MZppKD57dhSwBBZdvY8kcIfeusYyRz8aHF5Tk0857dlIB4KmpYHlAU1z+ALB0CTSV
bvp9WvmnwY2wRVelABaHtq+4a85anoGXh1p8NPD71p9GQHBGGgskzK9AtwscyKaktllvLLALex3k
wKW8T+NMJ2EYeruYYBSixfQu/0SXyvZyPxsu83aA0g0iACjTuDr9yg3nIV0JwY3LgGAAyVpKDvya
eGZ9367OrtAP+jpNffiQE0h9WCeKlFDuMPzgaFBofexuQEmHfo6CJWeaLxfoxgLtdgdGnkoNl/eI
Ds64eSmRx1C6lkbvk9GR70jZ2JbdgXAWJ7kG6pVlW14aOxYRVzhdpPl6SnXg+0/snjoF4N+S+Qei
HK4HOX5XOAPbQjRjCp032Tu8OKjD9YdyXpfSkoTn1f4CEuEa+BG0npdE9KG19TzzlHN0H1K5IO9e
dv2+lrgGGEFE5KkDB6J81xkDYVAzWz45r6+KrStyiEpSCwiRvRa03nRDentTo0lBqvK5y2oynggE
j8HkrmNun6A0V7UXRQXUV3Nwhxoddk9OT+FtR8MYcASHqBYuTLBvDeUXZZmTtSeesNsreCqBZV2h
Q2ZPJWmhzTpedbcBtiW0yidvwZGSzq2x36awAaSYCwamc2LBJ3W/c7O22v1idu4H3LHXu1v7xLVQ
JHtTngA8Nlj3DhNyPon81+F4BUTB1nFWBeZmQXKl+HK7EtmKMKZwBvrp4cLIQpt7WQAGgVC6jgq/
Undiz0Vo6zzJTohz6n09FC7vTuyVFpq7UbBVQaN2O623m6Bwiy+y1XRfoGnRPIZMDqXSwPwRY+kA
7+uqnjFQZArGV1VRcw8FUsSx5cyf2mJg7OKMgG2SLL4cJDVLBvZzM8JDXv0BbI40CmKGmE1tNZaL
VJHELlBbwqRMwFSYq+23iu9/GUL+4NeP1j6Osh6CjNMIm/wIeu8chPvYUzXzQ3Sf5iTwLbo30/Vo
+ntgOoBO91+Is7TYpAGBg+BA5TaTcLZgPynagR6682Zwq7kqmtWUy9b92C5nz1AomUcFc9Yb38Vu
IOPpFms/IKEGiS/aEDQTLwS3Px+fhAx2AO9VF5fV8IS5yURTjmnX1oeP68BCfD5NxEA/eQ01Hom4
rNoI+sWgLLyHoP3EOzIYPARyx7BU7Vg4FXrJdZuIrWjOFUlzt1HGHR1hfccuWDLYITulQ72aw/Zq
GwQWxq4cpItHr5yVxsXZsqXJ3lR24ggePQDc++6UyWPsC1oYsB/UEkJkSnjehPumfU8tQeJcI3ui
ggRShxvir3p/aqFvyUOgKez9Xo6FYJEKR9NydA+CcWwWFBgzvQoiO3lrs7eqvRoo/Qhrh7XbkwLF
/7xOyt9/t/G6Va1HXJ7KedSO0v16a1itzC4YQxu6x8w2fFff8ShDU73eQ7ohz+V/eg3MtfyVqRbT
Loqt+R8DWLNNYm8Zok3bt4BO5oNaFM6Y/h8kyNB5liDhkDA/+A65xLqiI6lCiCRPezuTXPtyPe35
y0C4hDyJrWbEPWM6uf2Uaq7haBqgAJHQmfvtA6AR6rUuXmd1y6iS+y18CzH5tkgiGBQyQhyKSGmn
KkKCLwtxQos/+Nh1bDTaOm++4tS2lQ15rdsdnuYtIJY79Nf5uC3JV+P23s0nklwujjNGijoJ6qSH
jiz85hx6EMjVz/Yhv18zMNIIo9PNEamWozj2CkclW2H35q3tRbsgjm5v47dP2phGcQMZyW6K5fua
uM6bNeW5l0N/APdf90Nk/zjvvVQYiMC+FPHJW+p4+B+nskSbrcmfdw6Z/itPeDK5H97zmDOovtdy
1hUAe47Aqv/klW5amBHK2KrVqL+NhOXiLy45tOwwPqwAEsccvYI/Yt4fSyDylNN7pFiMvs3W9sZu
1rRs9l2zpIuUnODyx2GlPaogZkh/yGUnQ/kMVWKX8F3/sKGkHRFTzti8MQ5HczSRj4QgFN2rLizd
7VMWz+kALibcTAdC5lTiAL2DA9MYleupRogT3tgWbqlYoxzz24FaddyVo5RlwEM2watqatRAQ83Z
CQddM2pLDkRy4GkLKo85bjmXEWrU/hY+gBdaAnVylcDpGk5ThbyBTyAy70trbnYEJaIumEY42/En
HJbSHS0Eh+hTCSbM2bjrR8MqRZ6P/Os8vrhkEuTFq9N9lBdC20pB/Yf1eVpqW0tj/G9q3aR8DwoR
v/lUEkyjS22vNdv0P9JvnRwu06sH0FtZZCM9thBXg+CHvupxvEM7Hc4dZyktlm0fgoSy21g9+gEG
BDar2CQb94CCsu2DEZJrEWQsd+lhB0vQ+pIK/lz3/I3PNIbB2q292F9w9KPcfPVzCDO+vofBV9B8
GhoIHRoGJbivSaSIp37s9wsCw08lPT3M53MyaNsYs1TFOfYO5kPN98Kappkn94gmzMF7CqqOvrmj
X+gEsAqKGR3PKYBHZkByHyMYSoqtAAgIitUkxYEK6Pg/XaO+ueYTQBwnBWswPYImmIuHn60WYisz
i/UCljZa16zgnonpWoh0PJ+sdn7DE24/YOcEwKqjetDFDryEB7kEXh1OOOeT6+BoGL/yLRSa/IjK
8lWIArXsKrrMsqY3Ze8L9PB9n+JZovUbkUrLbuOpFnDZRilEqu7vSs3oPpxqYhE0/h7cLlqOQiRi
Fo8qpQ28u4/ZlFG2zuECLNuXIF2yc7eSC5Z0OZ4WLW6s4eAjM6l39YA1MQy0/zmg2TDgc9Wc4onY
p/reKGTGbrFab9VX0fXJUDJJMHppamFOpJxAA1LDFlInFwKh9iC6Dy5eqtLuzVf9/f6cETF1bWvb
xC+mDL3jduKdgArT/42wJUYOAYWKiio7aZ5emb1DncBSjTnariUi/CpdhzohbW6wm61MqRMlGAQr
om5ucVdCtmDeUrHAfArken339RvhRmFjvREZCri8FgI36PrNooIQOQuithew+cuHEoSfS6SqwAVh
9RqJfHl4MpCpzkkA+UYYim9ttQ1WzW0yXvPgv40REs8toeBfwKTFYRy0OiRzv8p6rZ3y8nH/XORm
gX34Q73576jf5PwtQHUlRBrNs4jIco+nJLN41f+dI0rhLdlTJSEm1r1XgAi/nSlh5OCd0xJJq520
Athb7Mr+k0i2rhUx6FZedYTSd8OWGtmBpl8CvF9We70wWZxHeqdGcNFpEk3vi1g2SLQbR4m91Ssd
//IMXgy2rzTDCBj6MLX3JN7fp0h3dE52e6dhlfcB4qPj4oZVg5W9pUMX5M3LxCmrZVsYKRZIVxS7
mshR3v3a3gkrSjs+Psn7o1q/TZGnV7/8OE/1hbJxzOoe1THcL4HmDCKtI6yZUhu3iyhvwD45umuN
fjF6VeQ7dnr8DcgJ9cXMcChzOYw6ZuNW2qj0W7wsuDgAzKFApOoY6NY+HX3oCfRsO4+y97XQ7wZW
Wztq4fGkRweNzc/2DgfEuTcBJoMa1Fuua9Z+c4ziAeldNuPTjAUvG4snwElsFTqLVUTcBmTGg8zs
WcUEsUHMSXP/NJVh/1gAbq+VliHgOns7G9K9m4oycaNcDBG9bsGKY3+Qfc4YsRUcogD5eZDlN/RU
yKcSl0i6XJRmRoFOg/45MtApFzcGu7pZhIhTG7tn/suMC5rE0n1sb6yndUC4J4TTxGhgxdkCJs/X
nFOp9xrpmQLElyStvh/GTLBk56npNTxFnGVNEASCXTETNV8EUbKtizl04i+5JDs7HOrKkJkVmpH5
mRf5r1cUGW4DY0uKPwsNEHzRX8VEPHCYUFK8uXj0flmejEmKHRWJDYvXG38iUvkLfIqcC94VjDJq
jkKg9zzSislEB0wiOz7wbFnXOUBDFBaxFJ6VI6bGu7sNdkxv4ek/O66D4rqrPz4G/d2bmVk7nvLm
qlNeJ4UhieEehqqF3T6A/rTbB2MpckEM/OCn4RFyQ7JxAWQqJMfGL8fRy370wAclhciDhGDvwpiS
5aZvFgDg5AMLeKLp9WULBAux9xWXxFzr+PGInBcUQseQe5YRFBDd9tCLWQKIInYuH5fv2IHTcjOD
eN/R8lSa7+m9yO3AWrOSXJtXC//Ren/BSZpwUjdlOcuyQJsYhvZD+ZYzwBCw2+RmFB2CGIKcqDu+
2HKNIe+i+I9JcI6njKVq3QAS3d+gVdVi0sd27o/67NOmiLoe3Je68yDWqlFBC3krqh+4BAySrvuq
92BPFBCwrEuChx8wwS+Xm5IwoLVEqxVueFfOki3nJsYMJk3fWKM0hLKjeyO1L34vtZXh7sfJGFGg
yxSB9jYLohlTI13tnh2dw1jPrbcF7/eyzqCFhtdwGBlR+9aNQmbG5ojy26EuNMDvLRRuJFjEd7PH
GiWKOvYf7bAm07U2MCk3a7VSv1k1gAMVuwxvvnusr+s+t75BGdQFp46Xvt+F8vGuV+LSACCJ/jqH
oAv4A0U1gJCeCo2e3bq2wIP48lrGeAFhy5I7YZen8gFjJSdr5+kKyJXvN1XvVC1grDW02JhaImHc
j+EHDPxF4KcSbHA15b448e8/LhHwl4Z9fakFP1HsurZ7yDonVdiNejNFfpIFk8wC/gtfLTyJSiDq
EGF30mFVS78eNwpVLQe+Y3rtvMS9Opohb3kzPIYSsLALhwbzyul84hqfjDA/T8mTf6svP26Qr8zZ
N0AvpgQBfrk/cFpfQLQ0rXOsv7KBJ/pbdlftNW59vHV4zaUkXXE3uIDbALe/5E7N0zz+U9Giuqvi
JGLEm60upNPNBbDoh6tbw4hChtOaKF4UsFK1o03BLucQDhEMWmMLWrY6AoYys3B7Ag1krLDFR9Xn
wstbmWawezCaOwd3k/rsS3AzZQhGngJbjYXrQjeLdZLCnOwFZbqp8A5rGQ+7oqNGGc8y90QjCvhY
M3ZPipgTCunYC30eupEpYQ3nWk89p1bsbchbajLNL57UsmRpX5497QE2gDOHObvWnvv62+S8JXpv
xyv1wQ5aMdU/gOn8H1erYpmSqjv0eSr6bGIW292RwSZc0hXu4jaftkhw1gzRdL21PK6ZhEfxf+/N
P0GdJ9MHNq3Pe+uWghGpphjximp7e59ut2J2/xRtglxghD2S023A5kzHlL+/+iPxyqhC7qHn+X1e
y9e2PV5MKjLUctQCV1PcTjy6O3EBZYoc8EkRrGGluH8/mP1dohiU/CpRTlfBOxrxol2g3QIJ2ZRW
bEkvcZ10SgvOsy4rc2DabwjqV04Mjxsnjj4wbk9UguvTH4iO73bNVm64itMVglWo2Yw6kHeXAWtg
J7ZguLOUDsdumPhi5PvFLM0Fw9ZBHoFg6Bif5bcCugOUnDZscmIUptA1DHJrFB3R5f3Ao0cjXrRJ
KktjKedK17Txu4ESZW7ZWW3x1uylvjIIPxxl35anDy9b6GiQIYpGOXObNQt+6VBUZfZhcxpfS9tI
4qwVha1gmSjxnbBjw7gFBZMhwr5bMm0gYJJllRodK//kf43k151RAJTqiklauxMvnjOd0I9Uqrqh
QQ5jaap3ENWR59Al9RusAflCVYNlLDxkN2oBnHhtRkCRk8X7p5Jz9RZjFS7v8owncsxJbCClcICn
8Wu37sN6L2eA6g5loJh3v6+C22/NgqGSAnYxyhqL8iUzFHliSOW4nAlnNCbvtwVhD3I3agvzzJCM
TVwPEJYBW5eZNWWBuPtrw/NMjs0ywQkDmDgQjMa17iYiy39Dn6m/PinJ3k1CwtHbywnkyNEjaKwN
1H+5QhfBJNKrXScTWR2ENueGnRlpSasbBtg9j+NyOO1IFjfIKQLAE0Re+/aYwGvDK7w6B6kiJ5O4
yF/4e8+hc2OlnJ82QrE17bQNlZ+D8AHnsP1QkMzEj4q2ZPF9+/EfOg824vUZMXGC5W/w/M3TpgSG
FaWSJmeLdIKZlHGP4k/QvGl9CWG4Skn2speSFRF4sOpeEqLxje6X6f2myYyg2Q2ZNgmj7N3880dH
gUpIGqdfco6jc++oR3zaUe6JlEYO7nFhQwpCyQy+8JGVYW3tzHHF+YEmzK+ZlDPaLrHFJhgBqOxh
bu1qXbmlcT50qLC2sS8Wb0UlxCsvFAh8BG6L6teNzuNA6vje6GPtGbiJKzh6ptbi+jYQGfOhz1kj
D+adBTs35pOYvzDHoYZHU0n1lje2rl+phWgvaHn/kyz8pWEQc3JY1CbWN0RvceaFnqSHW/iiv7QY
UXdzDcYgA95Hwx+kymoBNm/rlgIXm4nsf+x0h7HxnXWYJO4A4nBebWJ+fCZT17tb0DUfAEgIAQz5
uQg0BaFZEJeHKQe10LKMGAteWmb0Xk+rG4FjlQdNArARZYL0wnVlM7uuCFznRC8xQRmlmWnjwp3M
qAtpuO6uglUhNrleG5kLOKeQF5GW0l7YZNwgWEayX2pB/oCbfWyA2dNxDq7rXeyw3pcouLD0/zVD
VpXfcLSVsKqUOIDob7sv4mNOo5eXNqoRP78fqNcCK8m2MM9E/AMv6pBM/R+731EEiukJi9mSxhc1
pPYSzymOI1RmCeSoRnf3EwEUv/rOe6wxVSjbVb6yE36O8cleR61WtKs/2tn3yYWkNt5hGZActRnp
Qrj1UbKGIrRg+J7ronnxd2JH7XjOHfbFVvQxf8j9oddYMowi9Qlcs3fs2/uxgl3V8Sk0bwm5EWEa
3ZgMadhwuG4z1Gucbm0DIHjN+tlXt3gKwBXCUOYNVFQFK61DZlJQLaELlayDEj7RZQPtKRkW1l5W
f1RSlhnWwCG9Hf4cXlNOCoywTM2BIUKo/pMNMKf3hgW5oYxd6AZvAA+dezBF7vic+0qK3gB1nm+O
YjQSxTbn8xmJMveT6QbHNI8Ji2LcNpyiFAcxJawUsOxAW42yK2NSlBZBOw+SUuh87K+qVWqV3WZ2
uARMk1oLbWYE3v28o93r6Su3554Cjo9XNqinyxynZu327WxpY+CjWgKFi6qjYe1LXZ0KHkG266pc
YcNF5/U+ykHHxQWwkFP+MBKkxaIqydX2XUgXMnZWC36clgGREeqgOsdGJPdw4O8cNwYbsOLykjRf
sT3Kz1YKpjtB+Ra3odb1/PUlvfjuy4PCbQsMbUopnxAmPu58G8SAt7uxwjspG8sJ4exxsPCEw5et
R/8Sfz5Bm0yrmeQnQYupZp+6OCOYscqXUKHggoDM1eD8wH3ZIM0FlUo/2HubROsRXEZg/4C2RBIY
IEZuRN9rXd4f5VlCS+CHmI2hKVBsix+2lJSX+TQU8QlaWZIL3nI93MehLwsRexMurLqnFVMNHxci
8yL6/orf5rmNR0kP5CFS5HmlqCr4KP9WEg4QhkNvB1eDOPWLPlDQEl2aLT5WQUgEplmmAPMtLtEm
NA3DtBeynNrawiaXPi3SmTV7eti+sjlAxtRBTQt4AeSz0iL72lnpv5+AJEyOWmucMd/A20+nMnZs
WdC/EyH+JpIAm0yDob4vixHlLSBQf6yzz1ZiW5Il2zQ97haeWh1PPE5yukxG8LpXYSKeBLwq3jD+
5i6vB4pgpNwEcdXWbjMD6zMP+uammO1EDN3hmrg0dRiRGDfCbFSFYuWBakAt5np8/mDNHuMvwuFh
B8OJyNE7+4h+jiEJtSHIdMB6kELTaC0JT7vN4QhKB6OX1G+RJcRoTtVCrldpJS9xmrrYrfrqTK3K
6KjDVJX1MAvA5wAM61RrpV64rUbOkF/AotpDizCAax1mL1K7CDWvrUfp2sxN05ipLC6LKs5KXt/0
NU0J2KC1zOxzeQSXsSepcWGQzp2rUjkfsEVuO5+5y8mF1YF7Ginx4udOQDo1vLGl6qmTUZ9rxXyg
pQHLrvaN3axTo6ocTrarqJsF1IG//3Cknu1wTho97b4+Cgsggy6pofetLJJXDdif8l9qE8LeWfu3
WwDuQy/6oUB80mVLM47UACBjFvVV3be+zfD4GioLytHesBrK9RbGGlEw0sbPsC61Uk2QvJOlLhm/
Ng79+jOFmkyFOpXQKd+RE+k4mgkA+OtIwiOiB6mK6LlRnY29C/1lV1CSPzdZuUvYS1wctvSBcnt8
pXYizY+UwY3NgS89WxFTYhcPgxdUjfg2EGdiWZ3UkNTJDJenRt4/k53NmvisAlM3nupeNIAVZ5BA
UoI9BFrgNn4DbQ1v+fH+KOyV5yVejeoOCA7nPKowtu6hxa2VS0idKN/WRYeGkjHI0BPIWDuzfyIS
RdAg/iBdA2/hN4MOvG9uhQNXUlrjKrO3/xSrJiaNXdI4mu2eyHpFkfvtqgjVqix1oiWr3xJWD5+P
w31kKWhLvScii6bb8uFcGGgxHL3TFr5ZmKYFJB1QLp5EgTkW7f7eW0o2Le0m3rqFhzAfzxb4PSQ7
3SRFXbeiK1dI/hR5F7sjLtibTI4MSyNw9w7Nca5ZkCYGeJZU9IyEAijx/XFxWd4G1tKMe2tLQXiq
FyAE8RZ8CqNR4oLIPCOcPfcCxLz8Uxpmb6t+h4Zm3juY3rjrdBy6L/9rMWtk1JLi4/XfV85rkIp9
wX8HfYMcX8HQOyo7ZFus5b0PWCER86hRwkdnsEo+tJAZriLw37B9uT6YgjoptY/TCw89nShCoJOh
1ObMhmWLiWZ8nGnglnaH76CrUp8ayV9dRHaLJkmgPBrrx6sSKKpBH3foKsIG0OEd9hvjmv2/Q1Kq
UOzR5f05WrQW8m5qAnkOjiPnGcWPpOnK8/HaD05ejviI4GRQGgn9DZdEXcloDv7orORykXcr1pHM
d9ko6Ay1uFfRGMFj64CxIdkbLr5v1rUlZ9rCyWyhYhsOy2MsdTHu//q6mq8B88ThvVNPbGC00rI+
Ht8/eGr0W0mFNVclTuAKzczgxvbXeE8ymHK0r1G6gdv150nTdUvcQ71nW7CLkmpAC1YTipYJwK18
0NIr2hzpBJQXoRsewbyPaKYs+rg4/eNRioeEAeSu+/TwkZvucxCzW3HL6IYmsAFELScmNdimd4a1
mdumoryJAkaZlnuUEuM0lgjhhLqkqPjqQauC+rmYmP2AVhdgsWbscb986l411YVL4b33QQhhGGVh
c41m2LMR9ncjV29GS/22ScJDw9pPk+RdTRD0N+e+hhWFR3w7vqfnsJbSXOtDR8utxhQMmRtGu38D
fcao1owwEo4VLi6tahsMjcp9MWzm3tcX/6EducDdZhg37FFxkKh4f1ij1Rny2bIhQBsO33qmewL2
khYYyB9lLOPQCIfApNS3Sh63qizidPvouQVonqI7N9f1wCQUAim2Vogwph90+nYSN56wIuubQy92
siOdNywKOe+qtlrwA6I8fvTOcYjka6N2J+oAR/hwwlvlkww5DPLO3FCzgLuvNcqMCYCZCzj6Hl22
Y//FZ1vfbfKkILgeocBRMkEN0oxGxN8uKoYSekEyDs/AS/8k67UzCRwqi4u5JhmCFPNdwfkbaALR
qtmRAPSJCXieX5YS0+8q80uM8JepKeL7To2VuWYJgUx0UIcII95ZJb03HL6cMVIDKpT+Awe1/vHX
c6Y9NouKsMed7jeXoYi5WBmZOPYkFhTTu7MvC98mmGG//N/Z1pANShUY1Q9EgYp8+agUcWjj2Gub
de4DsB+Mj7PhTMjC7O6cLwukvd218vd6/4rh3WwF2hToU9YVHAy98Jwi0SsWSGpJy2EMFopDGINp
AT1t8d29H6wVrwdzA3FtZpUD3ABKgXP8U1rrrdzyPkoFvBRgpJNXtSSBauAqu1eSPxCEODcXIdLP
lDkwM2HqVA+oQx3LlMRHM/TJeBlbWqJbuAE1Eg3+FRvVbnSeSHhWvxbrKQoYfSdclQy0GJscIDb7
96839pOCunetC2RxoxrQAnpB8GkHnY89o8F+XciuOg+yETeYalc3cS3itY/FXQvxeIwiHAbsu2wr
g+DF0dQeETpVL1Jriiv3gELUjumjHXQIftgla7dT0QvPBQfwxwOZLCGoRLm1borHvYf3rmtgU3ML
ARxySr3CQf5Rh6ZMF+CA1+cb9cDzIuDzZQLOQsMMVGRo7jtqDLsbuwHq5NGqvhdP0p5XOaXVkujS
p56b3PevQhfkODBhiiW0XCAJCsef7Tm1Ux364rYeu7iDSxcOuhDZ7XH5YTtU3PYCrx/487Hc1yrE
gxy/9hVqwAXTrtDUNkOgbqw/dCVVRrS7lGk0EWiNB/3bluEFL7wOHEleSPeaLAa6DaTWFK2ZOf/k
pkd//L/AEFh/L7naXL8PG46IVvDSW3JoU2wZVliw2mPzAKX3DoT3Kng+yDZPIBVyoU/BvJttkAzi
ue/8GGr9O7IESGAmB8yDFAd+gPC6scx4vYGSjxqMd+dYT9nRKYvMujniBTC9GE3s1y/cnL6SKM7q
yrtl8o5k9ugqtJzR9OM9FbPVNLr2KoWqYiySa/gucffNVw/ICjSqgJ7UKV3TMxp3KDuefDEg2uHX
mXKOwUFcVzMYJOCfwSYNcLnZgFZTy0mwHaLE/8FJZmftOw1miJpziVIATjOJkkRPpeYAxhrBAipA
onCxWLLkpKsPTP2NWTfXcj66N8tTTChnWL2iwTotoUY1GlfV+bm65iWuVj6FdCTkF+fAV8XyxICr
l5+GKgKFRNHBRAZ0idJW1wF1JBmJ599OuG/4Q1pq+XaSORWyRq2CXXeo7fGeQkrK19U6bi3j4pNj
FoXv4nIRuZN+nTJtvwT1gdy7HYCIIHFeseXaXieu/zt8eINWRDsRuByJINxjw/v2B4IzLEvab1Dm
OavN8q+lB8l07V+qR4UHekuYylgrgNYxp8PI1UFiGmeuVs0Spuv8vXH48L+gHU6V4WXNMZtjtBIB
TkNHIo3Bt8+/0ffwIkdLANjW8J027eO5QM2L3Mye26HHNd19Yr9SocchXHLVMkZh+PKKb/KEtZv/
nUxQHfJlpJD8WpNXAvpo3PNEH5a0F9svRekEF5OaAnmdTr+CwRnZZ9c7DX8VuWLewViMQXUxHXSO
VvaRZZuxH8BaoCTBE+zHUwPUiE/AK3G0/US1XvZvrHmc+WqyvqAAF3nlZ2SKaxdpYK6V3DBzK4dB
t+mPZT0cqzYyiXG5D5T1Et4ZU9l7q9JwAV39mYTLvBUFq6N6tAMIcieI1luvlsFAZ37khp/yVhKK
IfTwgbRvWyoD5219ZZTWkj6xaP/x6wr3t/IV10Y2E5ByCQvtaYO6T4z3QWTNUEglZBZMb3oVYSfe
6ERB/LoJvaMAk0g1h1f8Wj6eEK+Iw6KKIFZ+49iC4dkKd0p6xibvdu3VK4gsoaJCWU2duTh6L4vF
tFV0W6iLzFXz/KsmlW/0mOwNRWb4d3U27E+3KSICApZWH1K/o2+VkCqtHNcuDi8LwPIzATw5U033
yHWYf4+1EMXvqZ1U7QaYElot4MtDli4O4XN6wHNrkyEqljAx1vBJqIMQCxHHcrqD/xNMOLR18ASX
6ik4EqNtm56CVZSSr6mXc4kMiYtCuhngLs77K2IOTvCDXLAJ60aj1cgYuCBa1KlPllnLZz5QclNB
x8gkMnoRFwabQclEOeG2LzCnKFRgvkTv6s5hsCaQWHpsnlhoMvkWEPVPkFGmqKmMYwSrURyWRdkG
D35Wl5hjcd+cN//14UPD80cEk1r3y3/KXtdRFiPvlIs0NGM4KNvj2YXJN9QPwWz5DmyGB4bfQrF+
HrxocAsxEbEh6sbICb73GgsjeB+CXKMO74VbSQ3GwagUtbS/y7bKY4c7i2O8j7SnKg545dCE9DGV
NyYGRngL6/bbKeojVmGhyw6tDZUWnST18U1cStx0niBEyq5wRddV0g37+TDCPV6cm3ojCvZonM+v
PkH4B1h/U9Kb6vxhnrbxMXB9lT/1oI0grS97pvHR4Ur1MVyaRV2GDDxJXm/wlCyHqCdNCJMyWKjO
FZBvN+zfbKJKgm8P9CK9OS8DFPl8ZlXj2WcIY+p5y5M1i3cZxcthEAyuxb9Hwi1XV9nhbHuqPg3F
6LYMehmbwG7v9rnjHw2c2Kyv4w31p0non+MOeYIOnmT+sDo9oT1wGzpvbpDcn5okhAvfkPb+SGjn
jpfIrGd+Q9R0l4h4gjWOnWT0F0HCb7fxmtQ+c3lKom5AG3rguwBvPy9I7/xvlGe4uxL0g/1EOSRV
GaVKQUjU9N0YLHkNjeVtofNX4ohJwi2D+ES/3LGoNbXemkSWqyiN23wVT7KxlZWE9zxCklRuWrsi
cnGZCpOBOuoHYafzAQsa2AztoczeEAuEreWIIw6zmohC/r+IY856iorXGlvLvy8uZ6A0vMOC4emo
onymtAk3Vl4oIHwjuts8DYTkljz1XGOewqsN9S4YWb3ufXxtasZXunz/6/x+nk8+4l3rceKJWPDQ
aWI9kpxhEuzil3cIYpgEHA74i6fa+T1VfLdOaAtb9yD3JcQuwvaz0BZj35j1c0UNnoz9tSk+AYiL
TnKkdus+fyNdGUgsWu2EVy81zU5Jdowq25RusnLwT2rTc6DdWXvQtBxj04qSD+idxgGTRiMw1Cgu
nu/34mcl1u0ubyX5mN9QSRYL21Yn+6/MY6CyoRD7tdyyok56EHqeW82M3IGepAktz+LneuMePFIb
Odav0smrVV+ZkngapjIuprIMlJy/1GUv8aGg9PVbCMi5JEqlFi4fwHsspBpycVBFx65J2V2Yc7Ym
RWjaQnPEqzAGswkRV6bPwoMSeYVxhYPGxA6pE6x9FB6UtHonZYHgf6h/r+U/5DozjFfzoCrL4ntV
U7Ges0izacTHVnJGARebgxFaqqRg6Cg64xcsSiF/hxE8iKsvX8s10vtjoNOzemjFoqFYZzAVhMAq
XAbBhVLlScjRvYbYrSFNtQB/QDGUqaM6xJj0rVSS2jlJn2hbNG1wSAAzAoNtkwO4WW8hAGetyGW5
mNHYV5zNRkSWn5byzhmOLzf868XS4619lZKQJD0EPw7gOvsVH45J5S1BVRdxeMjudftU3gY43JlA
mW5kzBP1dMuwE+f5xxy2OnW/uyvSMBdShgcjF0EoPSgXYaa5htkS59zM5kvZ7ypSbx1SDilkzbs6
l0vtdd5yJ1GHXGssFgf4wBFP0/Cppx6nLzLg04QXaz81C4ECYrquDx/A6cXrHEIPafKUfe4OI5hL
G5GlgfByVNa8iYsqE7rt1jSL3GlXlOIRmz1CvDWwUl+3E7sVONZSkWGHGuUTxY398loya+8XZQbN
pwlNnql5Xhy2uAvaHX+M2fl6WTHCFoumZI3a3PevwfomBX2GTT6mF7dIs5AiWtG3+9NUmr4IZMQ8
p/1MKS273ovpjy/Or2uYHio/txcXvZwgFXJ3goOG1QcGgAPL9w9oEG+WWg1PaKjR/HbsFsCz3vz6
3t2zo8nnjT+/ucdhgGGHYYzvyB0YbAZ9ezgN2jgxvLAKw/NUKngyaGwzCjcxIx5mpUFGO33RqGLl
VxllymHVGSCLvxirjeUYTVMzydHSO8yzT1ZZkwHbJHUH14qqH4z4TuRBC4x0zrvA0y7wuoKmVYyD
fF3++p33aHYHa5VCwlqBhI4pP8MNH6aPHGQp4C5j/3S6GwHhjxTSlghx0xPOhqMBw53P6J0YgDoz
vWtkc0vtWKL4vf4NbLSPjSDFQ4Z82vdRKmmwg3gjDPZ5c5mSDHs0RWk+PAdpB3z6PSE2lBz0I9m7
h6bAlacr0AGX2QTsyMd3x0QSKmn3x1mncpEihlnDWikDtA4EZaiWUv8aduMn4pxs20HHUxlPEQlm
Y/GdQzsU4voZpNL8g85iBLc13zOnp+0uKE5Sc0jgIwmtRYpgFPI/GV3hdA0iLxLl7Epl7D2hNkwK
5XUIqBzOEQCwKpwRU1pcBzs+GuhzQRbH/o0a/ozjE+5QUMeFY2vvcVIMDifvXzj2W+GvJ2bB9E2Z
qoOETajkfxE1zEeZb6B5oN4/jJ+OmlNy9l0ML3DnOBBet0FRL4HE+8LJakK7725V2sV7bx0xjpQU
pwJ0/yMrKFTXAtJYmkr5kASugL4ULrHPy0E/mbeab2skynBCxro4QZxi5CnzrO9i/YYFQURs2vn6
wVXoRprXHWRWmxwEcWbnSMcsUqelsM6Fl7uBLWdMq1lxPBLzzyUusxbXEN6aOkFkjkg0fpr/D0/r
jfmr0mLUcnsxLTuwLP6GhnKFYHe3Czt7Owb+8I/zZznEx5JPGas04A61/b+6raZ9bztk0qmaDx7P
Vxu85M8RLF2468WXTJh5SgDUBaGGZdFJ5Chp7hDBSl9QO4dw3k/7YkRdiNiCKTacvhoNLLMsYeUg
mgVxXvsnIvy4ajuOe1haKeeRHwJYJTfkDBg4y/IswMo7FUPsGr/t9O5JGM+nb345ujG0f9J4Pv16
GS4FtZCmXejY3zbx+ntDby/h9HWg16j2/r/dkc/LJNj8wuFubxf06kS/bizbOoMbiA73B8ZihIko
n80bYJPo67yTEEbDjWS6RzbNMU/OjqOHMXOkfFKXo40BSevMdGHaU3ZfK+r/f6l7Bj0roU5yzcPL
5hCRdW4LpZwyhD0vcQaW2bk3br2GTzULVQxw3qUNHQMcGuEUaohE4oHzqbK/Tqc8hDQZvEcMTB1J
y1g53bKSZs+Ex/vV58QxjwpqHuW0B57oSvbS3+y5/JcRQcX0OSVqQyziBAiETyk+l2UfFjVbT7qh
7KaxbdudPQYCQIEWQ068ijJL4DcEoE+B9mOYMnVK8u5hlCFGDHa1EVco3SCmdiGKwxg2OxcpCClG
zHYFEBMayJozrLFg12mSRuzFdiZtfWXI+283ziQ5PCV7beM+BLQlAx+CkSxq/JvTAGC4Kc6kra8x
U4KRBJC1mJkjXolqkiD3A05s0jv2t1RretJ0Y0ncH6/MmeAvXgsN3bL097mKa5Aagd4x47s+6tyi
/EvXT2PprjJHKKY4co/VLQyckRdnXFrBnEufusj2HEtPGZoNKl3Ro4z2A34vU1Cnob+EHQ3iFudx
xOd3XXfCzh83j6MNc9cODGvCEgSf5ElFPvp4iMZr0vR3VX3Q3JZpVW92CSJN4Rz4gNFs1dt3GPsG
MbEeCgWs0fZmFY2sgLi26JPVgcE71Iz+++xQEBXcMSStHugTkbfUzEegrw1LxXNeOaeawvqIPGYP
99Md9kllkxFy484vvz+6z1CSGGEwPzy2yQ2yfZGgQvX881Bhwd5PjoQ/hPTe5Ah2N0frnG4TxCZ0
aRtYxBZuiEp4yLexKVfN5nleANy6U7Uk2D5r0ExfDkvExmSSGlv7d1ufwBgWthKyoIYX5RoGX7QW
UDFL2VaMMQNa4rQiA2zrQbLME78Bk5zP4inlJHra1NSw1DHky1Nk6ggeeJGwAck9NI2VfJDMpRwi
bn9HCNq2B1o3C75dT8c6ybWvp/X4ju/VruHsA8/+MEU2WPf1v2aPNjZiDXK334p7c2C5v8Ty60m8
OgVrhKp+MJmPJkoAcxqbQn/Ls/dg3BafGAWAKZBoywPaISHpasZdTabAlDMBn/1Tp582BHbL4bY3
qVmexS2igs3cthUCIAkBTrGH5WPl98dXQESmVB5VEsVf/K1s78DGwlMMoUoUGU18/p+ypsCZmSub
OeXp5xQnbHSu3QbnUC1Dhaw6KzYr3JTVWK/Pt/mUUSByutjk0K3KtAlze6FtH45Hw3QG7ap2fzOY
poWEHQXgKaVnQAmzH2Il42yFLe7vPeD/MAqNNhOQRlGcNSj7euqkRkXIe9/Z8i0x3Yd2uAFgkEov
7K58ca5YIDbB6BnY4gn4MwuNnlgxC9CkSj2FzHfZPqKBaJ/1w0zgX4vLvepELHFIAB0XrTfndRWA
jDheRwKvdU3NtyTn0IDc1V63Z7a6e+hMwtelc7z1qtOgKNKQzgGaiIqigxFiFaaVFbibcANSfEvO
SJAg+gOg3XnZhd9Uv4kfyoYgRAcOYSx6PvpT43eed6IbgaJbz6UP/4ehy7HJssuUrCA4M66gI2ob
bHCHhe/rIGucPaGkVir5LiPJML4Y9Nl3hWtq/b4rGzxHWH9cQwk7GJmrhrqfEfKwNQ2LjOzb5c4z
kU0jM/vEdBtwx8LAC4D7BnX3/7sBak13KdkNsydDr//uQoPkgKychqbGqaDVuWO40pJ252k8vFKi
yQLUY5AQNd2m1EvlxbGZNy7IxfOxNH6GrsW4EKQL605J3EsCIqB79o4FtgJEMeJ5cY6DwJvFZmMT
dcQngTXMt4iex6MyUOkNFrhsVeOjQqzAoyg/SeafaMgUuDRiau/ai8OkqJrR2ZYlArjcpiraxK26
MZqbQhsnLIbleBnlt9ym4XiIzZJ/E4W3qmnVZJ2aH317jrDf6gxuoSjn7vdZl+sWimFdZ6k9v+hf
ctBk+ftVjJg519iDidPhcnUE/H0Cc064PuK62wm3eOBq/0v0X4+sjRWh+sN4AeAGYtHRHLo0spMw
IY2KupOsaN1j4TNGDw9WlikoVlRi5pvq6cif979zM7OR+SV4PUpdr6e4crl/VRfcEnpZe8FJodxE
su4uHwNcWb4kW4mvEcZQhDAW8oiVJ6g2oZkXIhY1r1J8a1LA5eKdF4QFY8X1ogawfZfCxbS/H/tX
cnOuqiYNV7F01u6JE4qhhLGX201EfTXf1ee7SaDf8K5o493kTqQJbvN/c3IJMRlbHk2Z6Bp44Oax
dQyTRsGumdPl67p1//59FCoFD5tw4X6ipAXXg3FOnEBAZ+fMfXx35EDsODApcSJl86CteR4Fng7j
W5uRLmt+hWY94/CtjC2NwKEoasiKcJzaeFWlfCuOoMRfhE2APHhNyCoJwdcQoF2OsLK4CIQ3rKQs
TH5/cSDCLce8A9I1k1BLkIgxDmy4w38ie8tiu60yq8b0OXlmkmRTx+lHo4Ak1wGj+jRyCzkOXnRV
Q2Xx2qxeo6moHrHAcBTzodO/SWdniiCmmyYEIS9HPCxkCmcWwveE6OPOqP9OtLT4k14nDXrD83/W
yY9vJrpRmlWzXqmL5drrTfD0FFqTuYufagIb6RFEaTSFc8061sV9wi0wxNiaxp++6bVFQWXCy4My
J2trlkbgJ3zkPuQS7FZ2FShPdNEuJVabY2Stiur582FRIQn9DWFzSkrs0PdoIZF2TCi86XJeuqp4
Y0qfrpb+L60ybhMyeZ9dmRIK+tmITPB4i2N5qeRm9x1IhM0NFHC+IUDw/TsH+Dt4TcD4zF+Amz77
cT1gpNW2bNyfR8SYUBBT3xh++RXLfOR4RszwmLLJOeRflZHQiaY2wq8gi5Z0ydPQJyG8YodAIhY2
whwwwAmC34ZWsDx4Vqzte4ijZACJh2LFBUDn0Lzrg9JHBDBAxAfdWj0P03e+S+lIB+IQmEcCUfLy
qX8RL0Ar9MBY0PVFZExxmAveGqp7x96STAdklaQJ3gtt10Qjika4KG83+m0qpjloPTedIMVNsVLX
+2TK7IwVc1DavCB0gW6U9NdIZX0O2ieg2RJZ0UpOO1Tyu0lEmJffYTFV7CsEn8YTAdK65YVaYhlO
j7x/ruR7WVw6S9k4X1cUJrsXZDw4yaPXsC07XsWMryvxOn9xF6/imcQgxyXPIKJCQY5A12LZFcV3
kxri+hHHexdWfK5qYcOhc7rvv2iAWR38QkYDkf5cFxKTCwm/jEzx5Dt41IFYxhpNRV6K6R+R62vX
sknd92ydXIfCff9HH3c9PPWzVrN0ynXBXizfmVv12c19o3Cuoo4eD7ATYZx5jO24Rihs3fP5Zu26
1Cr8xP9ShxbvW+othdcuKa1lQFWGaD0S8p9kABo5LQiXadU2LmJq8hsEM2vPFp+lrizn9odu8V5J
w1rda0ImxZs7aMq8AnowmVs0cyScrvI84rJr9MkJfYJY7GCqXfwMcorTPVzX0yxUV7gMUIczyUqL
fRxeTbnc+IKcT/SP9h+HAzerdC4vB+mrZUbEWnhVXozCi+cBll9EtRFxVtKG7YjvoIU/7NP1QxdI
1iSqTM8GBP6cGfwZ9Vfc85xaZUsNyd8B4gqtfkjHNMnRDC3EIssQ6U+e8vwG7JlCIxsiQZclMNj3
Prv5SMjezA3mSLLYtWITMdSwcYyaSAZ0ERtwhxhw3bx0bHB+R4GsL7ALtAOpVoHxpSM/qRgOD5Dt
UByqSEaiTAWDrQ2JtMAolRfB2ZYgDxQUKEmYpYScQtSoQlisyYkHuIJJ+SPAIDappVMY8YyvNYbR
9+3SII4Tf04dEcUsQXPGnrWqcqOi2QiGSBTVwN4IziRx99I3ITzwfYoz2LmNf9FrWj7WX6NTAKgZ
Mr+QDrnO7u3cSeNFnWkwg9TaS3Df9BdtU+/iRZy0JGOiAHpoQROaGoNEXSKWy2EJJ8FZpOOLE3he
ItOz2t7T44LHnYlKxEcFqJzn4MHvmVA5l/9CQPXpq9TxTRFPPkVm1lHHj2yMkIxVLvZy5CZh94i2
ZjjENujEfKtZxIHDDYJFxfoW69uFUthvy8Ce7P3X5W67g0OqisR0uMJdbIDYq6SrPNU7DvhL4FE1
ZB891XToSAxoxCthYl7rIJ+d+95Uxx7HzopJY7tMadMHPLMg1bs2tQd/vgowInV7dyIYvV9kgrNr
zEE9Y7nf3+cs3jvuYyhENM+VjDttIPdF3wO1DZWJLRd3o/4c4WlsifzNM4w2fwlpMrtc+YT2WQ39
lXD64JkYaVqOM+D/AOBGun4CCMsE5BCtf9xlufE/Zw0hmSeuMq1Z+foy89o7FQeZpLOUtdQoCCRc
BH7J7n4R5sWizW63BLbpj2Jl9aWi1rQVu/gI1SddryYYd9xL32eza0EJv5IRu43HsTTxgAWJx0+L
PqDxXPACWj4TxW1uwpGKWSr6Ua+Ak8y8fIPU8ZOeUvQuUK+0fPPUn6bSEEBTFvzzL/FJPV1Jnzps
/sJWJzHvSPvcQ65JIpk1oJ2pfIs2ijoOZSM48l320krM2PeIhG2mpGHjdlDCPEDOj76QNuc8Hap/
G1DCNsiss5tSnq5kxM4zUw8/+QngOZxwbExFjYslJ+foLngZ9J586nT/+kSMuCyfVZmr0y1ki/t9
ijDSDDv0mNiRtjUlJ/27ahxSvps1UlxNd3zUke/sUrCGYohQoLzz1LyolyxUVPhUMGPut8tC/nHy
Tp6Zq81xAeegipdncOG+ehvD0TijoUBz0qm9N2HCcbQHVnuyH9VNLES+FLZdftCWyg1VuqN31hQP
SWYIpYu9gbLXcuk0MnXe8iKXeQHcE+YX0ZpG7/YN1h/EBuYMn4dF50tnX1vwDNgePYal3xgbs+Lx
3Fif2NCbRNo5QoFFBcK8K839laQVW5TLU/zbjazyzZy70Z+XldoA8dkzb81E7cJVhAyQro/KbYTy
v12DgmvsUWxOEn74ZWLadHIKCOidL76CFI7BTkR8bsp1WH1cx0zYQR5OBt40KRw4Zolb3TbBXy/u
2YXUzMZ+HxxhkJ9MBlWhGXb/bQgonYlryZob3IXdvpICI947YiReUlsNbK5+SBhzpWIonioq9Vjo
NhLJ4aKGpdPBxJldy3LxR0nchQE5w9qdznGZnBcLKHUYtyIzKMeHTulDVHMIiovVN1c3953/NPzd
Kcq4wjdDwR1OKM7dEncu4C72ZGWeCp8m4dseJgBLFXhTI/KCNqV+895rZpwuXp7OLKjw3opz55Fj
AnMxx8vu9qBfmXGruO6VXm+XQtuJB0P3G0otfLZyyWv1dGlxWVGh9e++e8IBkWJIT/YyCOtAl2wg
r+Vwx6qeB1/dMUe1ADPgursZhgN6SfvNk8cHQOF2Vn/U65cvA4XOWF6B64yqgqLNuxaTHl7ova9B
cr2Gw9VAjlUDpOx1fm859IglXqW/NJBK5K/V5BsFcxXto1clINw4/L4fK7/gRQyH7Za1dpvuEj9v
GQ35jQv0AQJGpBgYVuiebh/oGQzynsXG45ivU7+OiEGp92jPQrERarsgtCjv8h0cEh08Nt326j4o
8gbuNp/s2RjCWEUOajwHuVPme7mIWiGT7ZAJa2NYfQEVEztNmhHH/MeLMNqH98Y9SxgjvlhaOQ6E
orOPgCZiDVCpI5w1TG5SCkmyacHym/TDyLM71gMMIcSbjdErSOKmp6Yx76ecdMFVWy4cyXdCZaC4
M+SGKLMu4lIvcvg61mICqRq2P1avxExNdFRuyqZ0S4yeL5WtZHxtptYSg98cVfZtfXtQO9gNnef2
CXwWFPEKZUamPygnTyikRlWb2Ls8PUPbLzvKs0BQX5YqIS5poIwdZs5LqDXzN6AMQksvb2d9qfhR
W+8J1p1ckXPi54bTIilPosvonTsHnC1LDXcDhyd7SxSDbunU1TMUlFXi5kJV9MWDBuh7CUZZFsy4
SSMu//J7nbKy4Fp30aRzTa0sX//vZhJlD9HrlvqHSMTCt4CDI+pryOQFlnrtKg03OgNWRR+0Kpax
Zlsl9vTavjj4Vd2MI4V/LyXwSzqc6FwzjPycAca3H+3ODOaOtSElJME7UjDqNR0ou0z7g7gYjcO7
1FY7eZA3ojb6cxZsS612WUOwtBfs63fYdWFd7KejcLd+Omsmp1sig3k7yF5eFSYP862J9XfNbSgl
B+uu0t0+g0YIQssaanCkURe+7jz/dYW0Glflcg5z5p8eCGzLCJTptZMydyviwPqaMKcYwyEKB0vU
ZOA8npqHpwXwHjkGeUmin2OpCeAAMGDvZdNC72RaEKhf4P49cUcvQQyIfYPaF7OAI7wJzlvk5zh/
fX4fFZpjDzgeGkH6G4Z61KC6HyIAxcN8N3QL3WRSnMTFNOASKRXG6Db5dYuTFMSne9DjUu66Jp1r
+0pTMlTbQ6L2nlwZlSSh2QxLpGaO2jWbj7+Erzi+gtjIHncWUNYEdDxM1BBQCE+rj1v0wSPtUaWF
QBKwc7EO/MwW8v9u7XkE55bXiaMz8qSabcsC64yLKNehN0kiZnKdKrUhSxd09Qfh7BGYQ7EorBik
rWDAajF43ZBlemuGLx+t1BNi6CjfMOXGyYYxB2fdw22+QBGQkECCgZcrWJIpka4T4gRPibrac5Vm
i/fr4YW3HzzlT5WIax6p6lwOtgToRGWZjZTYbVZw124hokKSA6aj5Ssl0llEu+Em3RyuCCxucDtZ
0NCcL/pDtjTOZbzqM+FD7JBehw95pv5oeHjjS0ADqj6+DPPCFTZNe5yXEn/jki3ZdnhHQVtnp0OS
2E1OnVs3dJlIi2hLUj/O+OP15qKEev1k2J6s3uoGmGv5LFaooMXdIqqiKvjXWY+WnNMSx1E/VFuf
pVgQPImxxb/l42Ec0Dl0ljKn5nHOgpox86tQB6L05mfuFDS7FJwfLuRodtxm2q5viJUYgv5ohAI+
0w6bNOTKr5niY+DEn9ts/su9RUbmagAdQZiUEAOMt/K7h979HBGEXhXiqwVlihcGGzaxNUceLq3D
Vt2gYpgQoWBiRjwtfWpDXxJqmbR7zP3mK1SlLMEObmrCsg3/0OTcaoSJwtZuKIGJ3YsgjUqKGNdC
LwbK4LsAuSoIz4H4hgRUtJ1FVcQdoKJqv1zEG+P9L19pza41GcGYA3O6siXLl/0k8JcF6pXMVSdX
jCW506goDqU7/gr68eqhMFYJLdQuKe+McDb1JupCulgUdqHpSLZM1yfor4ini1asACWnulBdp+tF
ZBDqIkfmw+6TPzm8F5ugqTIqEbX3zqo3CoQkN81ZmFEK5KMMr5Zp4p0ragBqGclX8ESwmTdCgTOQ
bQcsqWC//ifwgXrKk/d9muBkNuWx37uNm5UpghKAcCI2ssgO6Ps9TWcA7pWI9f0RTV7W8B72oZZL
xzTZtJ17+HxuIS8hhPEroS8LlarOG+/IUClEbC3FO2/xp/5yvwxKQ5WaZecxRLhY9MTs9MY/nR7p
IqX3dvUWNfoVAztri6xVMLhdhkIrHmzo3fIavh27hYL6jnCehNepfieCRSdKwxIR6xwZREQCZ8OX
r4AoQUO6e4SJjULk05U3/KrxR0J9qcxpCMukseXCejUF9G8gdTvzeHgp7ONnfRGEzrh3/Sz8NtHR
5L8lpm/F4OZYngMvkbYW/vf+c5Fje0P78tY4vOj3zT6s3rDCcqShATbWXPSRGGqgT1qBwiwdSvRv
u8U3PXKB/JHHxgFQ1HZ63ok69PfiaFpIe7sFmPbEYns7wMkUL5MPm1G8FlQ6/eDu9z+x5sUFvqTe
rmbA9Dhaz2+oUSXUMmjgTR1nfQlmzWRib3xU2uOVYabrLqRFpv2VoQ9QEZW2UsK7LPUtPjolVjrp
EFx92xJhF8t3+lQ/HLgRvGjwZ8BslLHPhC/v6ALP+Q76O42OnEiWIe9FqBxEAiRLok9zeOK+XwlP
hak6oUndjgfx3mzT7IL2m7YiArW2WzOUh4c9W/PKTfzAttmy73vMxozim20ikVfZE+oZGbF95SYb
sFMPqndZ1S0rlbtObbFNMGPVd5ed5ZYdtx8hz9r/jJ855CUiEHNDFRx0OvcslE/r7WH1aimzzaH0
74/0VjwWN7DMrBb1TIrG6C9cdE9CsGZxG+ptu8RNMu1vQn0Mn7+n+tFyWT6OhPGR6vkFNfJMZrx+
9MAeDpYRfjqy9numNg2n8MK3/ph04ib0ILi+RovcFH7XutvhDfSfLekOcKU6ltq289jIYIU6Ri/8
olJymTGjxDajR1nkxxG+UOMT0I5zLdNCVe4J4o8Oox0n7klSzOr4KHAVY4Due1lmiJzpgFanC2Sl
6pHpN+TS8CYRFXOhpTxcdVqiyhQ+xB1WnNgT9yPsB8nydPXN+7fFrupca4iCtTuF/q1m7sez5qcA
9EpYpJwLg3TJNvPYoz8QPzUanl6hBk15ooPMr2TvrXwGAW+MoiPPLjrPkV9Vm8UmOxfQ/jBJVQ08
2E+hE0pFvzd8RPyGzE+Qelod8+Qf5SKIc+r3mM6ohoZBbjMuJuEUn8sEQw/QNRrKn5kagHEp1oPk
KmmKrRbdejbgYoWPYrJHqMlwkGMX6K2j9Td2YM2kZpRZsXhKZVrM3nb8q8nKWxgZyr7jnJ9p5SjX
NRr1fpOjyOektvVyKMAiD5z877YTbxVL0kXg+gvuFpylF+UjykGLdT3+9ribX5tA80oPsxIAQZjy
HkoYCh98UWJ9HtWMjOkQqr9awKEbNFEMLgr+t3Jgk/7vsfE6Mrs50gOzVMcpET6pKrIa+tATZ1Qm
HbgCN+wAum/5vjBQp6Eq/tGrb0mDjmfor1Kzm4h1l3t6wfBIyV1O6qTElXovOWjP7YDPbGzGNWT3
SISZKiq+8H5gSE6ZItoQI4nUe91J31S5G580eops51VEP809t+FokUkMss0nXWh9Cau+werK5Cw9
ZkXe+fFYzMJZZps+NVi0Wz7MCkKkTSoXtBQ0jdmTZgaMT8jk6ofurIpJYi8m0BRu5ojXRAoTMMEk
+fSGHTYhDQjaVUUs5nU65g09Vgz7LBZPfkWBGEOfCXZo8dXUi67ll2gkCpG6Achb37oZEL3GdN7m
eCB7hIQO9ZPDq22bZgFRP0jRwxLyxt2hHEbx2OadFZKlOIvFhGaRLnfL1S4zEI2ie4n5s92+zG0y
C3kQ0+PfNYEuhI20ldnY5NMzscKCpmbblwuzSMRCBD4vyu8bx62VZByd71MOH0NSZa0DXkVhxbBa
JZbub8q8dZdwC5rdcZHvbZEMSzQ2V+b9Q3V6szu1qrmksTOO11oS007q0OV2J6jZpSCgXKsxdHG7
YKmRaHWVfVqMjqqfX8L3rOjQwt3vuXguwSpINvYbaTCk5NW7jnKfTRNlQvamqT9Nde0BPyKDGy3g
YP3WTD9ehuj0obUmn+pgn9KQfSCYZBgqAvjfsHn1rCO+AvEH4mQROAN9hImmGkjKHGuTOpWxE9XB
TSdyQ5Zwrf7qvIH1a9UZK9zBn5MsEM9zo/fc5Fz9SGC2rvmKEGNs/f1935bZWWMY0JFjPksI43ig
l0OJDGWTP9LyLeG+MILHKxuLyPraehgxgXQ3JoNZj0n7lXISciKJsV1E4rfYg/J4j6hofo1z8zVJ
T/KLe4iVAryDFDNLuyOsqft7LIka3h3PxirwwTC2T3A25vXycesj+QKOo2XP+bKWrWoGLu9rqRdR
thD2DVXnqNVsK1MKRid7rjc8A43kBRG95V6zWYogUxuQeIg4sViazhODfy6qdXQggEZlD8HVc6xs
EpEBSGlo5H6GXBp6ygpvSwu4DIrybXbRZ+vNlJhZ4M8glJARJGNzQNQF34Jv2Mz+Rnqg+4el50CY
on4ZSe72v5q2Ght8oJ44/uUJTK0SAWzB9L3LurJeQk3B9oEhc8Ou5efU2yJH6YMDW1HSVlTtxWEI
A7/RZkk2CDV+D2/cI2Fb4sNRxP0quK9A6moTeiAdW8P7XUAc8N5IyqxEOKOveMtTU5JjzE9Tu+ZE
lgqKV+86TRnOrtFliDKhFw7GltCczX5lq1Aoga7gcqbl5Ug3iYhH56BtMcyEb7DgfIuwqdh6plMO
a4u77wImIlyHN70P71UyjibCGXF3XoQp6os3ZRHTCLTjJuMvIYfndNfhw7sWYN0n5KB/wtakpQWH
FXRyGAz1+jCvPT2AWdy2gwoY+FQ8q2jGDuuJQboGB/KH7o4hdtr/3LHHFJbZidXBJIzxYGbceemJ
krE51m4gv2QDDaAlVXXPt63XkmJr9nO2D2aBc59He4Sz9BdohZhPh3alcR8GTGjlsrWGangkQtdL
Br5B9KEslaGOcPnPVVx2ME2G47U2ziJBp4RRRCrW3H5z8rPG2eHKdjaaB5g8HU0uRqZlxopm/10S
UPuXUdZWq15rOhQGD/ekJHp+D0lTSqFUTSbOhyitQLJXL46PFVWsdr+hsoP4fqMlY3FXsSLvQWx9
Zv5UfSnifG/fhkpY1ik7zu15FX7K2MeyUfH8b2bPXurp3VfnoVd3aDcajl61H8bF9BbrapNsogOk
YB9OAqfqQOBp1oK/YyA7ordVohVC3ccOohLkUYga6Lo5wb08x4vUdOp6WMQwddYsHp7vhuo3mX7n
RP7jJRwLeYlc7VTDb8RiOz8tTA+M8+bdO9ydOmwz/9ZetAIQTUEy0p15Hc7Dsx8cm2Uikel+Z5b7
F3AMRbT1nBhDWZUT75ddIA6TaRkbKw+XM63YowsBfq5MN2fi95pr08+hpolsdH0YWE1gYqhFHjba
tkqlP99TGSDT0GtXAr/Ansug4MyzZbUJhefCHlOV+HGJdxyZ3Xl9EdX7t6NcaK8LfE4OYxXQE5fQ
vRXOz9wMyT9YYAmZtAdFi9QN/TJAHTakL/K1eoLIyHzZRmjNWW0DZWVjTh/5qSFE/2kFdjS+2Bbz
aC8Eg8HLm4cupysGshUUQTqllKPQIvrFjjVaw+XHyURiXSNsKpvgQompyFbFdwP4F4clCzVORqWS
zTQcEFCFwfR4FjdVHaT2hfcUDr2qRaZxvA98Wxn2IG493KMQmSMqIUf3LELLLzHDNGahRIgEP2+0
au+nXRQOpzFysKqJG0UPTU+4T8+qk4HPbWJg8/LTY7Sufuw50xFAapkZJMEXOoe7/LVzYPotA/LQ
DRYbzQp6ioVoR0BrLcTKe20sDgMpcfohWg5YHCAMUGZn37/v0ZbD754bfn4eZLEcBRWj3pU4I5y5
YUzxIHGfd48bmq+CVEtiazuzOHQJPSSmTmlRqAmknAVwTx3aJmQqKkvPdtcxL0b4/VbUBrQq0Ksr
Lt3DvgSCY/HcM+FjC1c1qH09BDWjNTuKTqSXip2YcIPoJPJs7e2BJOtqA4boe3VXQYorVKUq8vsA
TFlzF1u0gid7ofa3PY+v3ouFIzU6Bgsm+D90afnz0XVS7wVXXeect8emTSUJxHBBdWquu9EQGGuB
ZHjqLRLqZuomcE7fKj7UQQL65LUElJJI5qp3J9j28g7eOuzScYzblERx4PP5082dgDiFAaYyT/EJ
xkVlhd/VLJ8gjFb8huN/N4DTWftV5y9WXmGGKmytUkaddkfNbS5rPyQF8ImxMS9J2NJpoyMINoBZ
rYlry3bwCXvKnR52npYnOx9Myh7u19oOmybH3Ag9k2S8cqFtW5vsoUzAa1mmEH/BLmFfGiLg6pjH
m4xCvdY/cYdtlMzLCS3UH+ZA1vjIw7/IXbxao1bc+6kRbePxRlYvgZENPkcuF+TRmXGvLz9+qVQM
MR6CwcEh8rOiAY5rOO5dXu/7n81WZfaWNgh/y6YZzZSIMKyDlFM2gGzjWuQCKQEo4vcbo/ZzZW2n
dfRWYBlCeAK3uAg+hpy3MYl9VhfS1UH3Gm+7nfrPTrW2mXXZxZSSMMfMLdUKkjp2IU0Bsodashm6
JmRew4+4955s+aj7q2swThn3tPyfmjbwRoWx5tEZdT4vwnvUYgZzJghVcbRvuyI+xskeRzExEcAz
ORIoUXiqPBtApH1rzhPyotPTxH1TjbaliprtToXRkiBenhYMrdabnrx2oJdZHl670Ai8Ii69gO3O
HSHFRnXMd96HJX7a7YCpcj8mWCJOln6q40Wi9AQXui5RtI3Ra4Yhm5mrs9SGwPW2Amw5uh7s/cSq
n3kO9wtWE9lSe+ycbOI4+iT6+kdEYXH0b9n4pFkQeZH7zmyGeSS+9q/0XMfk7KpHafEDF45jmytl
sWnnQ3sVsL4lGltxvDqFE3vLkHwvIRhE8RaQC7dCNbJ8tJ97rXa186qRZSIeDTmav7Bf1OAPfd6G
qf7eOMPk2FOHszWn1S8N23E/NTrIKxu1WMpUty4pYpJH/iQiF/FUnz5Qw9hWIusgQNJkyBViAenm
0OYewY+dKllznPyrrM2deNLFENgfS0YwuZ96C7mhvf0gIhJxO12qbDw+EX1RjoqOY9eR/Hp66OPp
wgFURMrX+e9yso4J98d0YpoQbvAvTQ+nJT2f/Xlfij644vXPCB+QkhnMpQUwmwBZBpSSnpDg/wMI
9bY7fh2cc8jQJeOTQI661Fp7AkUpDxUX42q/UJQVfsmeo4M/3C4x17zDW53VJH8mkBjpf2kc9TIe
lygEW/c1y2+Cypegwjrm/MF9Jc8w0dt1mswtINBNPzgyf8n2gc9vLv7xfNVjMLkACd4bFuovwopQ
INJeRs7Tk3FO8X/+unNEzYD1R2yqICmjhdJYAI1NHvryKKEq/E44kQtbnHv+FQmDl1t+IaW8OVH7
Wwxa+Kj8X0f/wmQb98gi3b/OdNv7NpOHZUIX9ZdElgtm3Cx2ByHruU/jZdd9S2XBSkV6CoeKWcZ9
5tg6nFezkKumafyw+ENyPmBpm8br9NQOqtVSZ8u6o5l4dQUqzDVgDXp9SiUvWHDnF5UGPI5+uLto
5jzIOvQOt0q9qfoAYxrBQCzaOMrfSNnwCIPy5lA0rs47OGdrOmttTsYB52Kct6ZDbSEwkhxCJP2e
m73gniK+iCjHiDB1LOYSKQs14xsXnUJeE4HQpEaMfj7vE65MMgHzBvnfzItJESvxlSidoQ5vjG/N
MvYkfmSGyaZeRT6pytDM6nRMSpbBBTDQouokVPxbCbpooDueGYnLatMoJHaM5L3o/kkp/YAnJE/V
AOFffuFtYebx5RCxqi8zcvvz4Y6f08NjgBDrdBBcT7+bDbkqCF+1wgF65YqHXbYjqZeDHsmk5mjK
gXZtbNAuCwSH9z0ZXVpINAfNB3wjtBSI+FAmEtUFJlGKY2JbbEjSyYdQBW+aoXuQkG3Pb/KQxRMe
7rIn1btIlH5P1N3lb7JryXuUiBf5EhQROrzg76nuXeHl1oMtjAofn8VjaibFq/flJE4W17INku1H
WH0hIwVRz+wvifKLY30zQw3btyeY/svP+9OFxHPERt659w3Klce0Oq1UFoRwiB5ZAc3dwIYZ28tj
78BhtsKyRpLzfzMysi/3I6+UwNkWpuPYAulvvEsUd0ihZw6cH31lh6vCHpjJ7PJfD4y6iMB3qWpN
7NXSeL2K1lOmFJcrPfrtYsWHcT/r0snxW5rkjvwnt5Cauj85ebIrQBvIpSYc+r9kFdq6RgjAjD0o
qw1CoRRybmO005xSPUSh0eZo/6ZSHwO8U4tl5L3bXd0GNTqU6QSRWuKmwxLoHrR0M1maNlj5/dUF
NigLR9CbKqgOXRDOdaAvOUGPY9zK7tXAiqccnQuFUXoZ+cf5dKVcTCcygBYYZmD4rTKmveTV4AhV
8rFSvmVgBYmq+Us20GtCwVTwuAMFlwRCz3dNOThJ8agTFtTsCihtjzO4NiyGTeYT+4pLTSjUl+hT
qMFU0wrUH/Nxyp/Bnk7ZRcFfabWYwRkkzkc6LEi1pJNfbbxLM/XVAlNoeZrKzvX1awMrB6AdB6Zx
Jvru2F9sdWhBk0Gy6NyBmLaLr3jfAy2wRuhAe/T86kkmigA/GUEdwceKEKtR5YjQhb5EcdWVP/sd
CYR+pB9pNFaUX0srJvxTKx08I98Di9CAbKXFp+HcqNf0lnO++MbeL+aqCKDiE9GqjzQtIVb5C/wB
tNlR5neaVRZZ8eAQO36IOhtdDYA+9wjVlBIQEqm6LPwzs8lNcLzrW54yczm15MwU1Z8Ngj+WJXvW
MkOzyBHjCuThEIRsosBGmDlARTxbkxoJFG0KIbfmJnEfyQ01yDM9X/zm7SY6Oq7m80vhCBPZBmyr
7Hogosc8WxY/NvchiTVDbWcALifI5m9jX0fiSA5QrWirggfwl9mZrFI6JbiUxQFgxJQCuN3KSVSF
6w9QYmnUZroErnKjXH30lX5AU3HlTFVDteigyN1ZNca3KAadr4c7waMyWRh1Hm5flKycnks8ULJg
kKdRJvWjcmP9Su/c1jAKSdJ0+c7NH24503vk45UoJ+eYTs5J12wX9z7ttj3XXpeu9JVzT2R7DMx/
1a051htsh0Xp5Q+BjftMMt1S8rZI9uVqB23x2UgPdT8SC1/Nia/qw42zsdHhqVC+G2J45Czwv1Pq
PitpiHuOm5B67uo+k2cysbgOSU1jELuDyIjz4RMg+ieI4EnTpeP2BcLic2DxqTA5BT28dLaqIdB5
dAx5TkgfVpHNiQ5UZ7SgJ4x8Zm3ntdtGP0j/f2sThJ7BX1H3hoPyOaaXzwgFngUzii2gROXRzmZd
HujT4C9wEFZKt/+PHxioy6M3GI7wWrWJqc0CV8eGWIoGrGx2w9Ys+clmPC6oy3hYDzf8DJ6FGvjA
83fODwOAtm2q9aCVHT3UbYDHyV6Q7us21I5AZda0nxqlPxaaGFhKhobxug6ThX/b4wM2jzCGdRUA
QctikjtHC/Hs0Vgx5LCNHlNbU7s0Sp/UTiReCqxsIT5HKC4AprRBJVg7jLhYuPUKBR+4wk6TNUP3
2RW+OpdypE87ylTlfKxYpRBEGinb5wGlF5/pVTMsArlzy4OQcNAKIFDEpB/Ob18zZ8s02p966Oas
dpmox4Zhb8MtwuTbvCuGqYaJ5CUNgx4us6mcxaNWtsbSUhUpT2bkd/8gQbqyqfcqUtWt9qrFPN2e
Mr6r6QwHY5P1xaO4WhsnXDBXeumrYxyqxqHqVJpryduBqShvZLwP0CAMjBfcAv1AEs2Bsb/nr6mt
q7SinwTgnDW91JclyozsF63KVoSIO50ozrxT1DNIluTq19J9gED8J+pb18c3VzlR6WAe8HuNuhkb
s6CD1I+ykWl2BtwzSS0ebRpjWyTMcggsH4Gw7FD+jTu7ArZGOZyTiV6pB541bnG7lc6VVJ7AEuXd
NRUB0byOH3rq97h+kAnNfYKnPeSiSZoIgN4IbqjYHUXDz2Obz1fQjFncq5cbouY2+Lh3u7GwXtLM
JHYwa8VftdZN/8sj3G+GKfV/8c5udTaRuk54zhfV5tlN++ET2Id47bsqG0dNYZe4r6DunykRPDy7
LzGkt8iiDXucijibpUHWPshuQGdPCZ3GzMku4QoKtj3/qwa6AmSVh4l+zGnHC97bm9BuC4rbkQbY
nY+zW5Ra+jvOQRtnY4DIEX5b/NP/l+Rha3McwPhbYt5qqhGLF6n8vQPgqDVqv7rYXp9ZjzxCqe20
aqE6Ge/2P2DLWqNKOU4WNnqjOokovBcaBfDintQD2lBoTqsTMAv71sK28FHAZCCeG9DdJxW+9BFV
dApcWBccv8/ntZWlAqQ1gizDi/JeIG2ichIZyPeDQ+zzlW6NJWSoY1hoER+87SHSI4NXg251ko2Z
vq9oo53nEunNqIg/w9ZYhVkVikRBdGb84zY8mzMfrp3F+t587GdHbaiJ5QGWGmuNMCC40BjD07v/
LapANBm+yoh7V45z/uI6QuWUtBDLTLwKh+ydMwcvQ3ByHTbbW2kl8L7mYi/xbHoV7WeCspFyfyoF
5qc9IsI0/v3B973fCv9W1ChRKWUSWKk7c1Qm83CsDnKXpeR9Wow4K0YS+0pWpug8OlzC8EAKD99E
Ufi12ETR7rx6ev/4M6fT3NAG0ZGgLnMrvRhVrUE4CqNndN4G13UjR/mJDpKLyUrtKat+Rqrlgdve
XSGMsm9G7WeJhA1p1z7cTIDDiFq20WIugsqct/QB5NwmvvYTSoga5cZK3rvBw2T8uUlKOxACbO0n
aR3n/KiTC7+R8vfgNjgY7zLE1RQgV83BdDXOPVdjT8ixQej21xx1j/dXMmGrlO2nHPwWZJiU1EpP
0JFg/OhC7YNQoT6PCybe+3EsotqDcd0kgdse7F3JWkUQfDlunV59s1SD3a6i5EmIZJ5M6xT9sSRi
xl4RVVvhClPKuwbNSsZtQyPDu9wtnPDoOQ4sKW2nlij5IbMX2jU18ealo32KvEd7GZ1vRABiyq1M
pgPDis2SBoNNEXJepRPSti/IQbvnmDR1OSxIDWkqeNADNdwF4PBSxmTVJ/AqB/BWTuTf3suWqEr9
yF2hX76WuwDd+wPqGio42jyzVA793e3JMvOGxhbPL7TrXsbW8gT5sQO6vjUUhStFRtXuFDGfXEqh
fRFEg3jt5bcFpSz6Yx4G+s7gm0JzIitUGREmDGej0KMDMYu7jzTDYDRxkCM61cy5GncQxAozCjg6
kCPG0ku8eQIpXjWNUdhx+YYj3j0hdQetnG91GdJzUjX+SJsHJkC09g8jOQ8wMXvt2Pe3PVjhLS9+
FofoMDA8gLOMlHz/zb+vTxQXtEu1ap5Ojo273IEYZYQJSMY6spifz8P8yW+8e43URPClSdgr0wyo
SRYVNe/RuqEA1w+V+zLWyP5Dky3Cp242pNZEodFZ1uDP3HvtEWPyrPoSt/y90uyzlNGBzMxT6Nu0
80aqjX8kF3DVEBJAlJDvWt8F5bvS88Gzt6hUhilZTd9wv5S9p70g8P8pv/pQOwELqnQPoj8irHdm
oTNlbnyRRJutyzi74xly0qE4L/fPUta1sTmpZakohGax5futs3XI0HyDvqH5LpbW4OhR3F67CFHM
TxJAuBOKWyFZUjq2vwbHrjSg8oFoF9jnElNewN3jXeJttmubtphwHt4B1iJnHFoKt+MWwMiBPIl7
W5x5zDCLqokpM3hl1iZn0kb+tiOcwE3Aj4uZA3TxYabdBUkiRaeR7fLQuyl3xzvqdCJhvEzRseK1
RW42+mUAwOQCG0WU55trty1KOjRlpijNKBhpPFY16xTp/odotqNPUYED+imwhoh/BHprJjIB+jz6
kOsge5yrESivd3Wlcwo11OaXqbjHjRHiKlaeRWOT01ywbNCNnRDtFEpPCqLRPKXTEqWTVg8tutgV
7jK7nYaizOlkIDNUoAum37W9r8X/PCtYRg6M8l8y93Euw734Rn0kkQBgu9HVe5pQ+gX9wFQDEVzB
cSRCvtgZKW1CdwxYsA+Yd+SnvCe0OaqoQN4z8Q+zBCC39EPB2WXJnIpZEfsxFHDi8SXEY+5h2N2r
Au8YrnnZcoddBStObKZ9vpX9kk7TT2hctLB2NsKT+Iu79oJLqpjOT61nu5jgGJuBqW5SpuptPB4N
Yia4O2b0V6jaaUMxHI38uYQaGy1qgZkFXXDwl2YME6MUTsPHDD7bTOry4gXBL1MCWzWYXElWplBG
uGCjcqDdPZ7YPt+y5fzDvEmlvZxBwng2qGI3MrPAJ/GfycmhUqBogV8Z2wdYoq2imm3XNs3aRslP
/tVmpN3mTYUWXxXI6rUJC1YCrkQE5BVDAPqcRRCFpHFB1z+Xn1zOrFT227mG9zbVUpQEhMysRcAo
MDKwc8ZRIhqc9O/myuFhna9sYHuj08yHDSGIToTySpmPTSD7976bB1/Erzjkx4yi7EKrYUBNUp/f
J+hM8NlDQbIp0zFnc3FJCS9k+WIR4Mw4bp3SXTamFkTVVPIumFwmWVCT811kUs/pp3WeLIxgKVbR
SwtNHmsePVhNC2q6aKHaiR8lcLx8eT4nlmzOERY3HOt+gl1Hp7u9oK9q+aCpvMbHca38lTvQLP9o
iBDzoGKiqwdAnzx6i8NXoBieSYdZy5sAO52v4omGQuzTuHy8eMl+kZGgIKeSWwznmPA4r9Kuo0e/
3A0fu3l2sY3n3izp22vQt4vkJsFV+smBNs9nBbAUhAjRQWblGZptGrPmP8b9pF6MnLeJSviUhHOb
rCJlqiwZLUh2L7VHMVMfhBBTNLpSDtUGM0PUCgOkQJEIFRW0VPzHW9rEq6BIB6Jhv/QaDOeNyFHY
1Jnk66MEZ9v971BUzkVlSUWKhgvvHY2Dh7oSzwmGdMcGNL30Gjqu0376z1RpslORaicDw1QCKOrM
rnOKsVRnrnXbiKc/D+3Tk6s8+/NyCK6Jn/4/3JsqAt7DmyWFpSE3UP7qvV1uOSdUuKEc4YZYSSUy
bxX7FqT5oTFDZtcb4WoUbirf1OVQ4Qd24SlnDsRRnjfiGIx/o1l1hKW2nmbs9hrNmXUfx02iYnqB
/zZvciaZ2XWoltXmj+BBp3747PlmqCBm2AtylKmimXuLPxWImHnkHc1/NHvi3mwT8buHd1Kj/K/g
WHsONTBk0nyTv9hIoxbCwD/YheZSqeIovmJQ7a4z2D3QLxe574z5/gPJ+Zu1JtBA9voxpewde5vT
p0BgEtml9ZxFNS1MsSOOLEh2t/szd+tOmt54XfVFBcJQd8lMBf6O3IcVHMLU28w4znOqS0EROpYw
OdsCdzVBbsRR6LJosPjrx71pNglPCEsjNNLl3utcr2lBGXAyNYim24xM90OWcNIue13EMmQgTzal
9UYzX+Hvvs8y9tG9eWsgQ4smtUWRT8F8KILqs5+zTKMC/G62o0UefbDronaVq7PY8NdFdqPZLX+3
J5ZLfnfYtaEcuS13vIynsXPEZcm10I7BDoMkLK5WfRMW1q76Gb1bA1FAn8CTCMf+eHe8F7ft7OI5
pSJ4/5M0F17lYe+vvhejREGOy93C3C5VNsfgu2dmg97ytVnDYcrh6oP2tXYCiLM3l1iDQyVTJldq
nUcp6rwcRXeJsP68lZVSJSnAMRG7oyrzh43rHTy4BwfazU1qmXXzdshyqev+D0EcsGStrEgj3m9O
EJ+zp2uW8Dh2z0kiazEz6DSqyjcYTK3hZuK/YQyEnAtEiMMzso+TfT/Mq9dUeLxxlvnyfstag9Pt
ca++GGQwvpWouNS+i8fKsUNXyZipQmjK3SfJAMbG2A1PrOA1SPUWVWZpXIEn/nP8JmbhglibRUlk
W4ZReiCZsbC6HYLGk+aK69aOnBeaIKEdKyXlFAR0ixKC9TWhwIJNkvItoMxSkaDeJyG2dXsyZIu9
67FBpkk6Uux0vP6qaR7GMf1oJ/mKXrX8kJO9nZiKis1QNUsdIoogrGVkRZ7Mx2nklNIarbBmgvx7
5olosU/lexTLhUD0lFhS8Lz4kSLce7O2/nlf6aIgsHNd80ZrbiulvJQTJ2osy8FbzQY9C5KvVJtG
k93H2NmfRNTIvYDo7bpHZ7xDh8pQ7MSTRj/cEFxfPNxUWE4lXZWmmOv61OBfEaykWK3Onm1n6aST
dz/hQcL4MW5RAfi7lSLrMpZT1JBBHsh6LWie9Bt/jZ4CCP74RkHDbfHiRGufnlgdl6dU8PjX99V5
Po51wlDtEzLyyXnQOvzM+nCib1Iq4azMmcvQGDwdVQ2WbiTJCoXrkbeyN/93zGoGTFvoAun6fUI9
3/xNn764zjt+AnPErGA1QUd0B5aolxN5PHnd8YnXFahIAH1UrHqbK7yCwW5JrIvb3o0M+KLZFBUa
dWnaVf1ycryVw6+0kHsBMHUFs3ycUbd4QJKjfzIx7uRy8HtmhKqpl6hhH8e9E7dX3/sEP8XYmBcZ
rDhhR6ogCWUfQsGSUhJjMGOtSPeV+JWpg4usJIPA6bgfJwgKnfD55PA8XpFk4rmdOjTPHTc3xLzl
Z4kpXWQJrG3JAUNrQ86kTU2RaL21yblgzgScqKccV3dUmr7F/F7XIrumN67l/NYZykQUyMKcrSUY
L0TQVUM/UQqq/yOxIbaWzxUqla2gcKMWwhQjYsrZ38KY4dVyEh3CwWwvET1np5pWo4YBJ2ceSo7e
78hWAnCvplj3k23DLFXXw7IKgLSR2WzzB45/i3Ys4wxk9FcZkfmUPz6g1iAvBuhQA5mCecOtP1FT
IkUq/xt9Htfh6Ddtt791gQ4EyqY0oM2U2wHl9VWMMzO5Xy9bS3qGLJkdP//lH/Jv9RZWgMgTKTNB
VKJrkG6MIJACCU2ktJPWCFi9itnIGc5vlldnmAtVSnktCbEZUs9VTINfa41Fw2k3C0VwYXL4p8MM
WQzswAapB28Dorg2T2jxPWd4OytP8oY9L26tIDNcOov2K/KHkb3Ik+hhMnboaCOwZFFutUq73XKB
/Z/gAnxN7iky3hARPZhffQ8KsJBhih3koTrJdpJsC82Sy90dPJ5AUWyPFJCEfCeQx3WUG5sHaFsx
MnhVCTcUQQyKNKwr3CnFv37vn8Dwn3wRtlh4QQp+9CvBZE0voSub85sh1gFDZzF2HQ68i9lYjp7w
uhVTDIpHPlVxUakyY3DbKeNT2d1GMJTC1/NKsjsTtxwgXyKGWni1VGPtOajbp7oPUwx5XvIuZaS8
SUxQSYrQ5REwvPX3H/bn72LKRzwUqMS1bg3rGBLt7gWQBVkrZbj6uyXwsNqzkM0wg0ze8GFWrJTv
C2VNR/hlYiLnVviNpaXNwxKquwfUSd15oiGhiPNuSJyctB+sA2rZkFsJQGgBAOq0J3bWdyXPsJlX
v4EWtzIgEAQ8bdZhj5KztUT0zE2wLIotKun9J1mBx3Ra6bQC4YqF6XxoUnBL1zirD/5dPqbvkqtm
+WXRozHo+B0D9qbRQJKQY3GYXZEZ6sKmAa56vjiI1i1bzjg5VjQVrm8bNYL7TNkTfpRRfI+b6eNI
l0N+kf9T9mmaUKxgucc9lswYT2GKyguH/jdNEegeRJRJFVXv2JO4i20wR8K2H1e/meCtfnHRCD5L
RZDtN6r9Vl11yJBcCokfepvQ6JVv26iTiYwIWw1vCns+mzb1Mrmu/WH/Y2DE9r7gsH4QG/4OWtG3
f2SK/YhLrTO4wkpIkcuTnPxdGGzOcTtDw+xMHXNtiammY8UgWHOpCn53FN+hDRk7hClw5so3gt2m
pj/1Q0mhnRnwcZb4NSowodywHbRKSWqrCzeC9JDbnPhZ/t5wTDIoX74wj6p9RtFAwry2Z/RlNb22
boJautvaaNK+mw5XL34SkOyQIcX1uijNveGotkTYOw/0rCbm0yCw0Muwc5NmFg5fjX/ryEUvn+4F
HqfapJINWQZpuWTcI0kEse2uYDE/2LEjTqU9fcPbrBFwq2brABJnRrN9U9BlQIwD8Xd5XIl1txrU
naDLYMpWl0/nH9x1uOpQ1PRM1O8+dFKEj/MHRrWzetl74aX6dXTOQMJtP5HSMidY4YVam/GMfEkw
3nZmtEtO5ST9iRiWNzpU1uY0hf8gHP6er5mzblyPP0Z/riEE7MDRNsw6f3Abd27UTNyGc2a5P6La
cLUMPkr0Gdx5j/GmtUJMPpEbiKxrnfwq3U2gCpIc8MnDOlx6rvNm9DAOraFyJcqnCWxpZDdmBfG9
JFO7X9tMDyx2mV4v9CICD1chZVXpCd08ruWTGL8cC/mITk3BZ+h1lWOfqP5ZtYel/Y71k8gspVg+
wcY4+D5j5G1UbG11YQdaFdH+Ax2gsaFKp0mFP6zo4Oy9p4li9wJm3nrv8k7O6nyUnQIih/Adi3qU
LBdW6F1kEUgv5yWy1ADdzBfW3eCtyibB4vH0D/42aJLmfNEuvOIzpyTbkhMoBWIBN/jVkd0kUCZP
r80qWVQ+XLODrpB9LguVtffkpovSo0sN4E9lv7AhuHbEX6YtmiK7tTikcRqf74E5AU//rDJsf1j4
OQ2vaUQuK8d5BkRX6mecrwaJJ57scHIeZ+zp4VB4b4zx62j0ROsNH8DOeSCZER8ofQfgRdqjGLRU
36yxUmV2yKghSNYqyhkIHagja4A5pTL4q9LQzbFQ75aHFWskOr/jZfJnnDoDlUBmymmaN8qcXuSe
TkgMltxl384NOeJNksMPavsLU0fgnBX9mfP/8I5t33UPuOQLm77VBxL5satxbApyJD5G9N3AsFfB
1bGgZ7xofD5E4gvK6/oKRiKkhc6Yv9+SBZXyfTQvDzTjZuGsBTditzSWVVDlmYR1uEodAmxyzLnm
E87rZboHq2aqHD74sgOL5gPi3Oj/P1t1hDbv2AcJdyCEnCIsw2d/O/vkUWZPtpL+xafCuB7IFoCo
KAwVUkqci1XSuX5fbavbp8aFDGm5sfbNvSlOjAA5uTKMQflfdBaQQff5LN8vgAKl51Ic1X54CLar
Z6cJhJ+IBv4+8MYqjAT253vzME+sj4uyETb3SoV/5RUHrtSyreqP+L18WQCiw2YGlOMJB8L6B7PJ
eWIdn+KVb3B9JEmqrENSpXCa3WHpsfcQd1WqDFMd5mhiwGS44C8Wriq5itItRUvMDKO5NCRK6GpB
YYGYMycWvqr4iVPGiM+HHoB2/BSwuQiUH12fH3bDcL/1vi0B2tpOi/dqvhoFUSrERijqwfVzd/1S
a/VDXxIYevdNkF4pYF4/3tlmtoJe5jkpgchi6Ut+G0FwrqIrIw+VOdCF9km0SwjMcHBF/Fgui+fE
YjOvy3lAwUKjVxUxBS5Kef9QZf4hmKSnFwiP5N3cfhDLxCWNStYA0yMZBm/0bf06m96/ksJbadB7
xEDVaDy9LPYwb3G6eBJWuqK8BYxPbTuQYa4GSg1X+qw0je6hqqRz5SoNqhGxzBuUFBojaKpyPNDl
jBj3XNl11FlI1jKFqkN/VK+765wsWih5Jm1yu6a/eIxmoSwgrsTVwsrRi2Zz7oEwouYTh2iKQ30X
ZgOIFSRJIoRB8WdnkQf0VYmGOywub1oquGnkP3biI5QILrc59LxFnpm/X/7VUXgCHMBOPuxemIJ4
c6JKiTwcf+phJOJsWCaMrAjYMVKdMF+yRYhSUAmu3n4AsqbdR8uZAEkakDC3hiSzY0VMgIauNYLl
8GW2eieu8UP2tg8rLZjJxI9lqPAxQDOqGKUNt0evJ5mcWEBeDGgle6LZmXQMEr5iwnk4ZMPOTsV4
I0aqedPsqxRFVqtZsVITzTkEFeGX7XojFWxEOOGFgb3A17IB7PscQyhcNZg9LP74roMeARceCaj9
Ra6L6HV286RPmYFLmSPgint20UUSH0R7SO3Zmh3wJmaWaSvSg5Fy5mKFeEnoRUg5FpgvAux2YdPe
zZcjWMvLj8P5TIZmzxdN8qXPoRXaC8zKgjePWN6bC0eGjKWGrSqf5sQf4s1XeIobZejfEEBvBiQm
1CIkGcvV8Fctl+6ic1UiAC9HU9qDcZugogSG0N/XIw26vnhSGzKgTaYtddM/Nk51I7m986TmNcW1
tG5Hy5o5faktNGOItDDeneuWLKa+a8iwGpyQrDLF4tx7IGzYABe9UWT4V+e5r14v5pDblo8qgoIX
VQCxC6YaNLOcVgKPskJOEkbzhghLCuv8dFuA8rRoF/mmEVRVJ3I0IeSQ+pM/U9OzwtB2tLPvoMX4
8dMhPCDtdZrOIyxIIhFMV0YVYZApw74UQW0SUyC0Ct+Spg6wiFboqfazyJpIM0HhJ4Xg9DahsLHA
s1DV0dhNamI1nvFDt5Yy1aEwz8Dm5AnwESABk5q3orJiiUJ4J1HFmEPxSkShvVO9rBJExYsInbL/
aFmUr/y7RbE1hajbWdXuoHmC0I75/nYRM/J8kKw0/IAYbKiFKsIfP7Ki55s/Imrgdx75jT8inkOC
3XBBaNiJWszo8X0b4rsnnum8xzZVTDlR3j2prd+JWWq1iaTDNMzy0QAeNZTUnZENSI+M2YngKDEp
hAlGDYPOipKoZRuEs5qtbyLwif7CAJci+6+cagai8TDbYvAdPEUs+LjTYSbTODQ4c/cM75ePV+aL
1fDcKESK9NNipYN2flJCHPskuvcW4PJi6goaROoFjoiT0hyrwqciezSrZdnLl0IUnP5eF17rwSuF
SpElr20rGUjN5DBNBjVgUmau0RbZVc5Zb7V0j2agGQ4ny0NX0GiJ/gmaJTr3RyGF+Y6SmY6w202e
IxRwcGJee9MVboYeZ4u62RecVYOEwZFkoR4dM+EA7UeDDEi2FUb218Fqob3eE5LaIAZBc3+bK05K
q7zPGvAbHsxU95rSogqZc01eXLBgCd5kg2SSt+LyLLj1GUwkwSm9tMbj2BXEeczd/5GnPwVBvfgg
kwurEN+xNF/OBjV6hEAvqLoY1V4QjibL4KYbhvtIvLP104RqMb70GLSKbn5B72kjCnCyOiEAQQRM
KdxbiDqeGF5zMYnXVE3AFAWSVAOZzsBex7xm0h+TEAAz9ysVy9KBGoXmjSsEDCldcdZ7pE4eqiMx
ilDxTcllG7ywLJ0t5QOY8WhB/TdBmUSJq2Edsvr/2HfJM1Gsuw5iJ8CfJDwchX3CZrMk6UN4LNOE
fg2mvTb9FQNEBzFkZ14rAzkPcYSifrmxDi/447wTUKCy1fbrlzDULnGgAiT3c4CvWsm1ihjj2119
a5iwAQT8BmsdOChPV1vOQHgUDfQh0iX9HzKK9IaM0njjo6XDaeh9IZJnF6aJsWf7r9jU0UYVszZ7
TrBqbU9nKhHZIPjUVdRouBZSPpxcCWe42v+MauQE5TfZZTqToNaqRH5shXFye3BguCK2feCdK0sT
8wsQoR85kdogJT1vtlZm3Ko133xcQGjZir0BhVEZFqfb14FMqc5XIxjtkSZQhYrHfaFB6D/xJZnc
zIE0bU2IsDdQwwyUi02x0Tkxkg2Kr3ghMGUKP589pUQNoG0KYwzHqXwDBdfN4t+gVTVgkmlw0Y09
MXkZrKzgFH8hk8poVlXFw+noMX6jHm69YtFNrTad3EhVZ7vH/e2nYbQ+1wpKBwf8NYbqws2MLyDM
B9NOVo8MuM25HGSAZ6azvJeUjNQQYhezZR1DCJJiLZzo5YJ83mMJ6ULlfxwSqrowoE2YFV7IAaXQ
Kzdh9ct/9WbthJj7Vo+zGAy32q+9RUXNCgUO12Q8cbxQzMSkWq2R7dPhTMHAWV6t1u/gObZ9x/Dv
/hkEEtixOmjWwiCQkibKIHid/ezjO5OYGC+Oq0W3zflErTKmw09psy1GszE7F36whmxUl6uv4tjX
TqJvEwAm/UjUb+l3xWqd+nQNJ4oDvEDl0qCzOX7yyi9l0QSVygDuUf+GWmkKiXeJ9GqHrE41TbmY
0764sW8akuDq9t10i76JTOTkpLxsm8yegkp9LIAdS6wSweaShX/At+J+jm743CLHNarQbZwsEpNp
GGo4wmCJiNQM9JxZLKva81pxmwM1LoRkWASZR/WSg6mGr8v4FxtlbkcPzdCp71QNWoxJB2gZ5BVK
41OMt6s2su3iNr4mGtYaEe3ugusUNHw9C3G1mFWFFcR9A0PocVnA6zEbW6TDV7N+nXDVcDHv9U/Y
3XRQnKFpntFarYVGb4xO/lCK6W8ZF+4w/+CxtZwkFVO/17YusfBhCcy+eQirYZ/rHcZwgNiXO/A8
OHRGrQgz9NhBZOm5s5z36TyHExpuYx1C2LM9N4JDjB3HHD+T8ngBTm9BDySLzbBeW0G3+b7Xk+5c
FmFe8hwuLGvdnuijW9v3MAFpR/I3l5Ju6rf2IzXPeoykmp5tQnRw2mivBe2Hp7Vjr0elzROdu6g5
5d2JgjmJV0OZRDVO4KOzyP7wWTHs77YQLTKg73ldhhAvi+c3kkJei/3EQ2N/9hqGVku23BZ7n/ZV
ViS14XHRtFW94ToURubYrV+nq5DvZiXQAWiJ2DKNuSCmJfkH9lucUNq2wpNnVRvbOyq+7oBYAPiP
0E9kIF8DrNX+HPcNdX6uvxT0aY1ZuwhdQd6GNQSHWJwLu+06jBDyrK0cElJsSe2WbkDqFu7a+oz/
tqqjfzmH+GIMyJAQW4/tSyG17JeyXsBdX9odrs//bWwa3w00++ZPws9I6Oxe1/zp8rm/BB0a0gxo
lo1NnZDJoTqnyE6KdIanWxvqsDOGBp3Wj2DwUlw6nbt1ptsdnKZRQF7hHu0q3Bf0MCgvlGLTpxu8
ve6xs4YDq+obH4ha1vvTQ4OW4NWK8aZM+s/eUTVQmYpWVF9rfn4CFF+Z1yZY+BWG/ErKnyizPMi/
OTPoashLmPyktJpgxIt/1vvuyYLZqrnjtr3TXIN4DDakkXXxQaBYdLXAkRAyw/bM6C0ViHXpYG4u
44JgYbhgSIVvdvOoiEWI7IeKxqxdx98JCU+eHk1ZJDIe6wXOOjqYMxHac5z7anJ5V1yfeja8Gm3V
oj0tOSeNAtY77dF/kHcadsALEB8H5802Ge0Ez5f1vWsWqVaAbbXdYvsZFEO58wuiAGHR1ivTOxO6
8iHDAFVmJFcrvOGUd08qd9m5GI/Y69pS/VKRKS9arU5DJVTIogPlWqSRvhPlvoh+LVSQjh+ptNA6
iRh8KuVd5CQNDez28ZkLAAIX6vpZxcsk4KHCNJHm3hLA+NqvN8jzyR/tLlc2Loo2VlFMHBSRaz+K
cDdFaAbi6QYWcYY9CkhMrddkZtd5Pcx1Wglqf0AEQrKW+YRTfhSxVFzuA+byDDeLs2rbzeTk1tBc
yMTBmY1C/8aFxmNDxHeMpvKzrZ5bbfAKwGTRu9xYg+A6cx8PSaYjjOfiMlTbmi7xai4a43SiWSwD
jxBlZ+T5iZuP48qeJ25m2Lr4ANxp/+TFZiJ98tCf/Icl7/ryoxL1KlhW1VYdTPYFmBtFld6+vZij
zof4EXcony4QdNOqoonFxR+B06qdkaOdNBG9RZo2OdTICyLklJkI7eSa+IOo/v5bdxAxb/YwoEns
vGO716yhkgggSCAIv9q6eeo7aqtamxAB8471HwluVXfXgXZJ5Cgx7HuwK/Qwlu6pLV3e8io8/OtT
tt/DcnVBTB1DmLfxnttuW2SsGwT9LyxUyzRXNvS/ZEjmpv7410nLGU+oUEhKez02jyc9LA0hvoNG
c0dGJ0Tg1HqPXHlK+5R1fHuqA9Q01JQWRjHQXpz05isLHDiS3F+ZXPEFe91pWy23T71VjdSsiYbu
grCpy0isY6HaFRu2oxaGO0vBfO6FxZqA9zykQwXV2dJ8R1Gl7NpnJTTZKgBJoKKGYb1aWm3wYMFi
mBKtPu6PPdgVVoENWAUHFrFYrMWnImG1vjHf8iJ8u0rpzgXl4lfpjtObLBLVRqkvKUSUwQ/27yFx
mdGpKL9oiOA7+PJLFMbKMiZWHBbUqp3DqcB3R4t6pXQ4ChgTDth2rnKJPPWUIAWbMiz0Wl2E3KeN
EOzJUnWfcEmp51Y/Qu+teXB3XalrIyoF8YjPjW+m33Pf73aJ8x8IzQCRbvX4sV+0SuGGhvdXzBBb
cuAfrVuQ6j/ZbAgVuU+WcEgd8A5WHqVmBCeLb31PGIzI4Ocf/sooMYGNtoFM0/1WY4Nsl4FSIFFQ
yUW2kc0iDd8QAg8bQ6IymPNrSQDDSrT1W/xsUvDM+bZQvkslOuu9XDnQzl7si45JaczHUU6I8KnP
54MY3jckDU2YWD+DBdK14CzI+Jk1baoFRrVG1L32U450AMRM9CIOJN1j2fRdF91uz3g+TCylWWp+
r03Q8EE39VRnKPFiGuB/7FWUPDIvrc6cOfEW6p8FQ/daHuvvRJbKHqyU8Z73a8c9nAN1FzkKimnG
4ndMBnIawzm9fXwOfPgaFU4s8R/TPPflXZJHG/lVLABOLtFlqGJwVSuoN0l7UcHpDyvJrLoCLjL8
yoCTRMKyGyyLjGdwrJ5xpQKlvJzIgZnFlJXJ0qtYq/ga1/vtHKwXkT/EvuAB+q2K58XQmTjvDnPG
QKAxDvJWm9LttvXcxNVmufOqdJCqM3Imvlk+TV+D/stbZU2miKM35ZTzb6bHOxZoS82AJoje0PH4
MM2HR+WOWvTIhW3qbnqYkZfaPKxCM57IX89xolIuixj2SNLh/FQ6tg8qR74rf4eN4uz++kvuowgO
0BsLbmZgPhOb1O9YsjAeDhCPN8qlnSuVAnGOsZa1XvgbnxP7VZG5ATn0A+bEOEWF+7FxpK7X2YvX
iYV4tiOv3l4XXg69znb9GXfxRKFg+VvEA9frtpOgs6cYTuGdYgP09Qca974XD6FqI+eclHLibPBI
4M3Np+j6Ma/CV5NKkH+Q8CtYWmTx6IB0BUjPAILmNcmujGBqd56vA4SMQoycOJlkzcBrjgzY28CU
MdXadWoBN7FxJnkmA2apYGq/YOt4XPkZMISoS649R3Skk1dFjEnAHarZ0H76gzBY+FrDcGX1Wbu6
C3PyShkgB/aaBGjPqt/XvO2BgIve/UxUFb2YN97AoCnjGfXIprxG/iguYyjkv322DbsPOziOq4pF
Mpt7V0WS0HmWQKtdHj8kzWmyFLDS23MbIhWsvC0YB2D4sqTpVBxbPQJ/3gIrq8vehF6Dmr70fDfx
UjDnTDL2YFd8fqjhltm1yVnaGTdHP99dOfoZ4Y72tmkNd+kPeidHmNXabScCpSCmNyDuo18AMSo1
HC6y6nkcZS1W5UsJqA6M9msjZCbW3DHD5nkwWeVHz5rOgS8gQexrAR7vdlZHXzdM/y+01sPiYHFb
tm4L2wNTChu4xv389FRwRsaGnSiqxAkHAFUqz84giyLRNo3eQfeDds9tfia0NEqD7iDwiS6gn1/J
s5CYerIQtSMtsAhOBlH1VU6BgVbAW099xnkZ5wuahBbq77yFNgwdA7z916Y3ftKCrS1mcq7pyNWv
9uKm43m+aM3zu53a/1U7sG23x33dJpc6ulyRsFcGr2PPgCfpPktWRRRHMD+Wcg7VzAZljb5di02M
0YBTxLHg2rwRhg8Tu/fkNF/V5hBcpIYJdxRO8A4Sy7wcjBLAmojq62KOsYmgn7Jqov/UBP/hZooa
n+imf3wP56s3yiDxjK5IBulVMAcj6VBVj532K1wOY+rBGWnFoujpyKPOP2ImlYxARogheYH1HB34
eJlW3uAga44EPZFF/+/fZk6Q5NugYfiCfMrstUp3eT1BBJmCPB2DU+Zh71lW7YqmRZ4sS+HrizCA
tdndGKF4zzQG9VSsRksi92oY6xLksTizlFk4iXQv5WVTvXDoqUUu+yqO5KRfNWTYhigDie4f3scB
XZgH81QGEYz/ud588XxEwl/lj2p660Yf7ktL8gdAxMEF3vt9LeHgPcHcZKgSMN+VsqxIDk3x/up1
nQ1QD84trK5Hhs9wgRnF5oV4YvskV2aBYlqGAL0EEAoTwKoAbdFjSNwBFRGJzLCZOJpUPlzl3c0e
mRu0QBd5ijdMJnmU4+/ixg4nrjs7Kl1H/sbxHs3aIktFVoiBPrdXK/PfA136ol//5dMgwchthe2M
4qgyUXlxH+uVaZWiGwUTmt5p+0WUzPx6wG657qitmrhJio4AckO0e3nJcVu0JgpRBUIGlYNv1fXp
Syu+IGgiYuMQQcr5PclO41f4QCZAAQjoBpwzfWE5VJshRqrB4aSXCEBClMMEiHYNZ39mhBAxWX2l
zLqrWmoBGbO/UmvACuTOuZ05lbOmeCYESaP1PWSE2PByWQycqBcQA+eNXVlkKiZq67Y1PBfBMYyz
mILT1Vzk5SelFxUOcVpViqTMX/HsBFHfeT7JpVcHitLDHXRWOnKpMELlvpEW3ki/xEHTPjhctp6w
NjE5IAZY37Sl5rNjLohb1+5Qjf43N2OvX2p85tXqZ9/3f32Q2vZjQAoWQ7z4yVvz3E4g2Vj6Lm7H
o0Osk6OpF7osM8JncHDpKuLsv3Gb43QB04iS3vXEdO1ASyxmiHDvmOWFMEzEGP/Tbu0tpVUc0zSZ
OAnHc9x3S1PZGB0AE5gSNkXKOEo0vowDPdRRs3Sj+kliqHpsNOhdjZQb2ePvtidownebA+9Ztriz
ff8kE3mjlV7M5WcHhQ24L8Pjp0gmkpfVCT987QjYYpD7g8eHt/YLuQ+abFm33JbE7vc41+ZUch1O
6i6K6L6FEClYxrC5dGxloUxHv38BQUCqeMDY9h0U7YT0k+XWVt4KpcYRvz//mCgmgKI9NBVzPeVp
VPlFx1YaaWJFAI0sSajBvJuB5zbAEEYCpYmWfnolqmAu8xXZhRiDcoYbLfT9V0fLdpF0xTxudbSZ
wVlV/X5YeGZu2fYBcHwVxMy/ci+VM+3dXX6r6l3wAQyC+SDl18V74usGU4rTNauvYznbtqvnSki6
faB12jViql50LFBB8UT70GmDwWGdy748jnHZvj11/lOELmLlnqYGxRUEOEchdXmco2ogbN/L695w
wdFibudoRTiYPKxbNdedU+OAtgGCJZeUZIR8NkzdOTQW9SCMN2cWNmZ8Rc2UA97Czvdel4dagW1k
T49qBO5FFD4BPK5eGEkNZ/tQbvg40F8TPzD8vWmcDOYFAm40/nRHc1wfJcLnG9F/OnJxaGt9ZN/d
KqTyq9dS01loJt8xAiZR5K7kLqvWw6M0RPAgzc5KjZ9M6amuEIDCCN8Rlz5dV81tJSSBRYA5Ppmu
12jjEtaSe7C07P0oI33a9RClyRDrXx+ZTs67jAkqaBiwvsws80sY6250HRoBmkXGEgmTJnVOS6Ol
o7ZY7FMycvPyXcZV2aJAV0YJ41MeoQ5r6ZrB74TezgBod/ep4FfdwhPLVFy5HqCZWvIshH6A900a
cVXIj8Ky7JBK9dF7s1WKxpH0Z5q4q1x+tSP/AhdJcQDKlvbyqOX7MNEOXPYYc8MbVs1zXrtMGFj/
GFSDr8+JWdqazNS8el7LsvyXEeUerSYo6jgNdm3fsKZk0LMD6XatcNS1pWqVMmO9v5hUomnGUwel
kWoR5oZfhJKTjZX5JvsVNsVzMjnOo0WeVC6jneHe5kgamxM1WWT8hNdHVrIBC2yxmIBZH7cdjZQs
9ICFtIg6fZ4rCxqJDJNW9P213o/aIe9Q3JipCcakQLSZKHoYE5oVUWjSXZPKbS51+1VMeGk0xxSa
HUZTHKqf26KBTjsI+VCnlgz/dt3ZTnuqBcGEV7EHJL4c+GXPpVeDXwlnWasDEy6laWkoHe1m1vbZ
n3Ip6F9gDmG2reyH0fLuNohshtBAuicLlNCvcJleVA93u5JFIDunp5fH9AS1AS6NqzMQC6W+qi5r
Gekt+oFkkxXslnWbHFlwh06O/Jl8q/LILPqgK62OsoNWamd3VWa42gMQd30LkUPMuk2FC0IbIVuC
SGERJgcAqumBqBBB7UO6IKO/bO9bbnBBqSu++cVWBWDhVhT9d6O14lRozflGbfdT5SLrEzjO5JT4
yTsVFH1EIPJKHrrngbQq/OFD1BkCiBBw7RyMg31Qso8ozG4KNBq8hR2mavlMAw6WvbnFljYX1Mz7
vvBGy4EazUrJn/3Wq0LexS8+7xA+xXq3xNrx36RNbsvyHtWPw5FVvsupS4GnH/ATQKWgsDiJ6/IR
HgtXNJJWf2Rfv4s1/wLNzGwVMo+e/9cljwSCKIzuwrPAG2WsPjvDxrK92aABqFNrh1QROmLT+/oz
aY9kgfLNoRowU9JrSEeOSUwD2uAwCXvOt8QL8rBJBt2VKhmQROqnmAG2w+HOj/UiQcywC9r+KZ6K
DTkhsQLg36ie4mezaKRI05Nbivaio/sxKwvtX6vAUyfjtDSXhlSO0MophBZulnR9jlUTmPVR/Bbr
5lu9ELnsgNGg4KvgW5rp5YRnjQNrHLeRXjgqCj9epGzkL4NIkK9kymf+8uH+2WtaGF/xqYErJ4Xf
4f2l6YCbVmUKKqPPxvTqCUuLUUPIkyJau5wC7OqtpUUmgYQsMRxzXgM7gUrGxOE7pBzt08r74Ww8
dVJ8t05kRA6NWsKwie9WDsxF2wS0Ko8uPBq7IjMCe2umVA7lAyM//KS+lDiDi9EeiGNXA+QXVd2i
nv6oNqcqtU2RhTJwFGs/65CNCzUC0kTs5hJPD8k7rLqjGjbKLDVWBefO/lDGG06i0opryYccjWmh
aAQsDosdeCTGNhPbBaKzfeRukDaKV7WsQnXc18f/rgvqXNEXNGVO/3AtcmkrfrzhnRzu25vlKnmp
jgNBbPkXq79D/VFgD67wemT8uHaRb2oIZ28QcgHKaea2U+cBP+zGI/NMKz4HdxLiTx+fUBdBZYxp
8MB4wfPdMDD41VcTkXfAhzHcIpWiEl5kAn8jr0IsfyIdcmL5+eSS7rl9/TRxczbfdaf9j6ReXXdK
Ncru6iRj4MCGR9j708pk7XGI9aybvHYTID3dQwoy3naJQtPsluYgNQWXvMzUHK6HwYYogTkOLe/z
uAelTqbn5CoxWhfJL3g9boDYKhGOF3MGR0ccawpm86vQYJmAh/fNx7cFYTaDEEfYV53+mvKg6yGF
seEcBAvGD/JJU6Dgfv1t3lxv450yWwNNyNG5Fwuj8jcho4NbfHRDQHdqyClPnVahcdgwfRQ5XURV
uwvEhuA8b5/mGHqS6ItmGv3B8WLGrPkZN4ymrSxqZbALzj46SYKVnE0hWQeMKk5yJFWvk2TkW3JO
VhKR6RNYw1GzMeYMuNB2pbT1Y9wSWa9dAmfYeSjKAWrSmLcGt4RuZAGPbDjVgz4N4y8PdNgaA9v3
+RiwxQU0HkVBgPZmV+dCqW52DpU148JRNIlKCvtGTJWO/x07gvRGtKOgy/ZPZCl5vZNBkhobqvNy
yVk5S4rUvHMeYaKCo3OicJCC5DLmcDOJ5szD8fRikkv+D05P7SzGBZ3yAKJW8V67HRXv2wsiFl/j
x/4/vHZeT+eha/7NtFPNDte1HJ3gb0CWwzI+jwKahQPZVG433L4wedqs3x4O2eSPsN8LyC91TJpA
TvFrbvkXslmixIqV+in27EqfN7CXdFckcKDwVvDV3gefwy96XCZYa7kNfOVJ2vaiSX3wjY9mVYyc
Yqod1vrYcxXkEHEvV/XWM2ZjQXRjpy7+IjQH5PqEtRrIas5icpKNnkmids7ye06GyHYWv11oOZlQ
jvbZf8c8I8ebuJTsDVlgRSA2pYho4S6egbJxd5ru5iOuu67VP24Kxm2BoGMQDFb96VmdGGtY65IQ
9fdumKyZ2aFPjzjQre8nrzH/bAwufxaa3JVU05OLRTbUuM8cWgS0w7Lk3YSTNoONQk9oM+yuhMeK
tJ9mbtz/GOOQhlV2p9hXqRnRv7AEdxiCKChLSRtl9QZ1YorffPwxc/0/56ataPgzTvkivtNKwP6a
JBDA+CqAc4eNwUOD2202S5/2hsbjGBzqFm1eDMv0DNF2hVm8fdx+o1n/gTFG1cAShrgSUqZBsOsh
f16EpsWIxWNqRmZIXrUvdtqCaLbjBo77h1i8Ms93qJ4Szx2Sl7L0OSXlBE2z41AErGZ+Hym/0nYZ
yxkjRk1bQ9ZchhyBTCYTb2o/nbo1O/bXKm3O2DBSpwjuvLJ9yUGdUspBF6RTJsAYleW26t8W/UbJ
NaJHfczKpkQTMN0Aos0I7tOs+rLeR1ErF6rhnGPQqtNOk6LN3zmJI9Kax4jQ0WTvr0Psik67PeyY
v+VsuYGTINx2ICvmGmXppPyRwy16OrecMBmvRqc6NyQOj2+cuqB6VV1OwSNe2ZBcPeQa3Hkm9tKw
lCu7dTdODBMsW6yXEjjc7dcOOBJHacYxnJi4qHNAV2JZvYkIHIchqMP1/z1V/yhsOTL23ooFhza9
EAhxVPtc9jQg2WKuVrgVoFipi5BTUYGBk3NfZjXqMehm7sWc252w4T5NNyXfaInqPhdlzDPnFS/6
7/D8i0PYltSU0cg9FCJZp6aM9/tinCEeZZi4loufK0fE/F5q8S5vR6IPfIN9rw6kQ9UTyAERl+PW
RP6DAiZbfbzXHupEBbJq0YOnWEOm5vT/xRnqbP4ftOzTqvNUn4yJt/PGUfa7wAVmCJq+I3NRq/op
KMemIe2GKngmbCeYYZn5VP8+uylDhhpY9po5BAGCmzVu6dIyK2KOTd4PI4pJ1ozgPmYJ/Vak7kas
cFJ/xI/XjYdT9qWFRLi1LN3lyfARte4iO0xx2mCbhAmAqYEyF6RM+GWGTvr0kBRh/kmlq2VktCv/
utzQlUcrob0YBaMll+suUm1hp0Go0RtO7BAw2bLZ0YC3qSBmeomH87Rej+17o2izHfWSOoIlHw3E
boA/dMUez7jFKxuUvREkQ3QGICJIq2RKvCxHeI0sDIQX5rOhDlXL2wIfX+NdVPy0huOXiNImyCQt
hluNGz9vpbCiEGFRsZPCZ5a+fJG3NAA2DXlT5R+dwhpwoTVRzMu5JK0ZaZ8EmZjj5lBzTxzDQCCI
ONIJiLpPK3YIQ+Tuo4faI5DL/eQBh0CTVOJK3gckUDvyBbW2kE9+AG3Ojwce9CfkKfxbsMUKm+bS
2Na680cT3rf8IzxfXdn0XJnWPl02uvRlMjxvkXi11pEoBF0RPmq8aFhPW8OVKac4wOvbNis4rMOq
wn8xhDc6ptwmngJj6D5q+8uJFUaZDAu21F9sM71V1Ypl0GMfKhNM814Bd8aP3F+sIybDInlpV8Xw
vY9TmRYFNSSPkqjkRrWILow3uSSAiRsam5vDvEseN4IZF0GFdu9uzt3Ik0ujKpVepMNutqtmFbvq
xfv4LbFcuiPOihQ47a+gcyCdUgkVwjyNvRtEpZffwtgr+oub+n5dVkbD5t2iGX8gNSpAWSCGL5I+
b9QCVUNH5DzRYfX2uuIuWYG1VwWIuVcjEhTsGWOfTb8TIPUOKXi3pGs2WYL7rzcg1XAOhXD7A1JE
Bc2gXpydl6/OTEp8PCePw23Kr50p3Gi9pm2jB0rIDWWWic1UQ063rAxQRY8OdkIFB8ARNSqBaCDD
lV1Bf4GxWwbGK8i9Q85K+/0mkh6JZ4c6q75FspMZIYSd23zMaL0cevXXX3/AixMaJ6z3qpXxltVH
mbrInLdMBB7MbTIXrL2Pn+oeYaxyvfcirAUXgOzwhi5ZjTKNLAex7/44lQMDTaEaZ+aAGVtQDWTp
HKm7qxYDzMxBQjGjzEwZwcyGzrtWoymkESS+VgTVNWN+NLtC771b0812pbhQv3wDOVqn8ArRWfgf
WC+DKA+hU593tRu8EkzHwfxCyoFSZYnVJ3M1TCPjjyDzehyVUOiGDi5aDG53N0uOCWgDbo2IRVDM
QWP8AiAdw01icucnT0vWQpWaypu3Sb8H4vKzkz29/BiV/Aahz7gEbR0PbHFjQdb1u6nq7JhH0yXQ
MutQqTbQodhHr5qxvMZcxjFF0+cQ5y8ZmNglSk0IBVdZSevRtwcikrIgPJqw0uRNm2gwTSUkIDzN
xuZm1qfkPLiKkOrQiIqeNooh51ALZ4FeXPwoKxEOkGn61fkoOIXgTn7cLQ84ptBU2mGeyKIMWPCh
sgvSQPfSRwF/b08k66FL8e+xf8KR30bqpjsie4Ju+1QVzpfoxVT9PUuveUB8UIKoD2tb8rvHqv6v
6CuYfu+2AL7nk6rNC0MW7f49BWO6qAYkeMvVDw+Ui5V6DrTawshP2v7tgmhfUxHJMpHubCquIdA9
ZxU/hfTRHYcKaC5ZMnUKPBbpWOyPKZZI0Mw1/2lKIMSxSYS9NuMAsNXvyqRBwqv/6iIIEBWe/BAZ
N1EI1EU8dqSLpcN63DhUuvzn5W1D7nc3zJObkzdbZMYvRbkvsgoUVAh3QBg3rVrgxrIMXNzcvMpY
u3Yu+QLUv3qAQq5/jmHx3sNzOGyRHV7O31WBBvqnNx868N0QH5OwBUqSVVUZPlbUPXWQrmWLNNRt
MbMU5QDm0JKMYIpgRaNiqiG8ZKZHGKkyLV/wmbavr7PmK4nJw5yV+rfkBA4HigbJNg7xzMsD8eKU
HHSBLqgvlgs/V5uvcMIofSKHo1zltrvzAKMV69gWs2m3C30S8GIynfq2ij4fs9o26wWHA8+0AxXO
jM6pAjUDGlDFrZCvpB+d1bNHNm0h10puUb07oxQz9s6fUe9ar04Y/DjWIU1LhX+TJewQNAbQobTs
c+VUvCUV1Lk/zoi7ZUFsksFx8NV+Vy4DpsSDpEuzJ0qL4ozUU4HEjJ/ShOM5uKAij1l3Zck85hul
BT05DDREh6NquadtZutp51JKMQgIoZ/R2eGssus6l1uRvzYAJdp9JranbmJ8Fe7cvD7Bz1zJx0vx
j88klHAiFAf1AxA1m0DTjPWfNs65k1g385+AQ7+HekhGKT8yDj4YcugAILEomgARaX/pEN0NZgX9
VXNvGnPLWBq1EpruWOBWPfRK76dG4QIdN0TsJV7UMoYpJLqO877PdjatGAgz9MiPpV6JyevpRqdg
gHeemHy7f3qdkH4fEfqMo/6QitHxjL70n0GpHcPK9M+5tV5nqzJcE0SWKrOHyEQene/mK427FA15
LnVGbKyUrnqLRaV1I/xhVRmSr9E/wmF2cGKBdnk7R7V0LSi9C6I2shswZktDN7nXvdGOyBHP7HEr
+SQvPeus/bGa9BGxaE8lQ2AE1ifgFJ4okWlrc/iBT0juFcSNXGpxlhhOezqIkG8RMBUEMj7mvYX2
QmAAnbtnyF/dn5jqWdEYHGncGnp0YIFmNctYyY8kT7/2HOLKiz2H7Z6ckDRcZayRMiOaK18OEb//
mO86Plr3JlZppEv0/E4PvYmPTOnGQuX3rX1zH4CQ6XCzW16ktcXUD3rN1zLqD7gynJIwJ6ZmAQBI
rqi1q9KL64xDup7yYFIu3I63OoGj/Pi4bqiNnZc5q0kPe8jBNRA4Zqn0xFZveyb393LaOWtqQ3Jv
1DxxAKnv2/BAg/SL9HscxwtnmfBiwwplVK+pN+f2D+WMgATGjeOwUO4Z2AniRNR81uoKnaC+zAKt
a1O91j+CeU5f4Agbfv/QRoNUPu3kFoNlLCCAHBpt16fyUHBJu4EqkxGoROo+f895QSVwWPkSWPEq
0TfdolZyTSzzU0Cl7ALrPxYSycXO4nAaOazQPGvn//t9tmZtqvMpC/+ppiaRUUhidhB3VhsbE0y1
hyYfi1QfgZpURwyxqcjGmt2PvI7vXmCpJGTivV8B0gQEW636VCAl9VYXR8vg/HysUFDfik1ttwm/
IOG8sXclpdG59jfBLkqYYbji6xcspUzcL8cMoDBXTzURdqxYwDsUewZGw21F8qAvPfDpwwkey0Hm
9fYENcaSMPNTyTTN+AkPUOjsphKBlA2FvpWl1Ezuo/C3wn7zHVBmHuBsfgq+j80O0LPfpgsFzlXM
4+ifuqJ3+Ic0Ikq0eUivcvlAJ+e1BoJ09LGGWJul5eyrJmTA2xwQQf0Q8P+YoXRfK3ZkDh3wQeet
29Mzo83AyxZYzG4kMZN3vTOW+SZO9avl7dKPvqs6pojUCSnVm6tggGKRmccvHgEothhhW+vREDta
r55FqICPNRWsNfr3EJvNgL6NS+6+WZgVJHgAXV+SJO7rvULJ1n9CgIM4OUn59VQmV9tsGKUyPqc5
3iU794fTzLq7pdVrk5s83kRkHikobA/Uhsl43dipqWmZJHy6WNlhjaE6IPtVAUBYmRZ39zlQ8ehI
SEM9nuSNKkKTaUy8g88r9pufM8EJg7Ed485tvi0lGeeYQO1wCjAI2+VGH4dvsmfXsmvLcyU5qfSC
HviFiqV2t1hmZ5jMevK9wJfmhpBzW2j/cD+d45fPSKfATlZSVwSs6nq6pM3HTVPF/MHirKU5+fYT
pYFM0/xSDe+SvqZmsG1C9R/Nsnstki8MUbKtSaA0WyGhXeBZuwAbJqya6fkK0gpsToKHP40WoDZ2
2PEAHuEm8d1etZLCywUVdS9N3J2hhNnk9xVjfBgZmNCLcezpyQ2nM+4LhVYrsdD5YDvqi+qLLSac
rfR0JZCOcXd+qK2X/w1QAJxDwytpU3clRbXw42zsZTAlsgg916713qC01YH26vw3zoZCioXM2F3v
9s2KKQKs3SMUhu0FljFEBIOOXSlj+5FbcDGiRO06nUaE8pSvwA1pDsiF7Fo9+vNZcLDQ5KOyo9dX
BciMQil7/DUGyXZSgtHT6bpeYM1IOWU00ieUtbB9mXWJIK78jcq+FZ4EJ/K3hmuY+jN6MQC6Ss09
N6pFn8H+m0/mdJe3pr1aW5dd/PzjS3zNC7UNUCx41M7SDE2fvbLVhI0gVZZuuHPBvP3her0gpYH9
Dstv/hwfOcgJTWSBoEFxicRXj4U8he/LqqlTRW2egexdEcFpIg7XWyWTF5eNBo1iE1bvQtdqZKW8
FcA2tSujfSMPAdfsoEMIyFVWVqxFybjP5wJRGTCWdKuYywu+iVesUwlnPGCeiAbROMkBevdSBK0c
AsCUwLI6DIlc/zO7KP48zZktrht90ZxBUrYZK+RVcRt2gPr2lK1XV2k4oXojixEIdaDjljPls4Y7
tUV3P9RZUq7JSuFjSjPYaUF9mZo0ujk1Z7yA9mxB5M0pbKtuVxFzIRsUB+ZE9JagJDKwso+3tcnb
ACp/nAJnhONKOHZUEJwc76CFGhV4HcNRt84B6dmDB5bPT9xrSqa96F/l9OlPqHjUCPnWx8ApAUMn
ilSTOFo2g4vhD9mhaGOVUz1RUgdCoeQG6iBoY5HDN1w5UQ0J8dWIpEQZdflZFyNXyqKUO+wSAhLm
9cejJQvMpfCBvN6hc8MT7WW/raABvUvJQPYVrjI9pi5K+Cnwqkgp7V6mRB2QPUsFE1p4FIEnZnQN
mqEL0/Q/6J5jYkrTZL6GVuFf4oiOi+eDiC+QyVr5rGj3lN+jt25PAJYMVTvnIK/lfQmFOwUO1zYW
muJt8Rgkilnu8maHY3ENWNg2ba/vetx0yceliY3CMEgc2O8SgirWDl4WsMd8UgH/JSW4TCPjaJFk
mJviDw6DYverrfM5dFfAdd1dYoSJvyniB3tMTakaimmA6z3vHE8Mj+iuvO7G0UMBx6SBSR1dSp1m
KZhWWfiL+Ay3+ncYkg+XFXQs1b+nouvAtHdpRiSwjoTHVg8rrIGEnyC3xUeC2DCtaX3qd9uZIEyH
9OMDizuyACmDd0t0BTT+zP5Im/SySeeIwHV8MfUIwe3En5eZqhNdr+NtekBzD7+7PxseJLy5oZcs
vvvkw/4IKikC7f1vOi1S9iLpX/g6D2Xbfc93Ck4NXcYief3xRj4YvH0+eeNUhhNivt3Z4rXCAJVk
6QH+XWsEmIy4JIRcq0Uv1tTVcSAQB9Jfa9qg+3RICGkoh1nfqgKGMA7su8LuhiPyD6bp/fluqzsO
fnnXsqZ5oOACX9mdabLqo5LoL4OlrOVmhJji4BqLtiafG1kXi2xjVN3G7HJlQYwLt4f9WdIPpTDa
a/cu13cTwKsKWYq3BoGqzLnPB9eeWfdkYslUFPtxHVbr5XqPmKAFWAbi/37XfRQgnLiQhDEWSgFF
U/L/6JaKa6fRIn1N13jMhcx1VXgk3dVk8zk5fut5KePFkMVTGvoBhRmGvp5CdZLXWg7R2kg+8Abh
QjyiObJmW2iVQ+MCxDfPkOXiJxhjcLAUDIVvBKUgI0pNlOuvvBMgoId6sa0Qqxhay5mfjjljvcBy
QewZLAB8rLrH+MiqCQRdAEvz/e8Qt8Tzq63oOQE2/jP5nYLsGgbYK70xjGboQjNFDKKu02ixMQaD
0hbggraCUKrARnqZsO85yLLT+lNdNgmTBfQUj0kgBS9MD4srPU9AjmyHIT7aUvepR7BpWIBKoNdo
CfwQmBs/cnq9QkLr1ZZdvJ0FcoOjUwzjkg27LRuhBKNKA3CIsOL4bZwbrul1YS0O3jtIiJM3mQ70
9fChsg9TWbt7bcd1AcU7eTW5meI6pvZgcC8iH4IS+3pqBgJPOK2KjKoTu8nvPWXopFqjhpLXvjqo
YcwOUHQ/kQqcO70lD4zJ3i1TJke5dj2L/YmkdjSkhboGEMleropgMc1w0qzovDDAoQZQDPUcWQzh
xofO6+37ETWKRwXjxqSU9lW0RYhBYcqzU0XfSk9D1VL8tHzAoldMjpRzE+Y63ydmfH7kIGh4fomI
TIDLSqjv6Tk8ES0YnBVwGX6vnonSLayLkT7F5XXBeUQ8u8nY/P2/gr2ZSLIn9IRok0Y6GMnQD6FQ
6pwyKea4FXwVC0dKVxIVl2Ajan1HCfneM3KOAK32b4mNssx4JnYeg3WxQ30BBaiGMQ2gH14BN1uC
I/EZtLRgKuzxpkE3Voz5OB33TI8+la83cdXqGF/U6d1z2P9YcQckEaHZ0C1McM0vgebwcX1pIbKy
puQ3zHrkELNlrXAjQf9V2tuVJpGifn6+pTRXAq7XwlXCAcK1sIzNzmQuNpIOhlUVbUSLpoFiaQ75
/Sb8TgBgUexpFioS1QPqTCkJYq9BtA2rBmGjk+6TIiqQ67rfUBDdDd4EatQX7CbdAa2lzkfZeKiv
lzYIe69w2Fd0nUKmUKFAoOFYvnjOCM/LRy2piC73Ggswl7BzzKyqbN61pDPERSGUylCU5s2N4QlX
Gv+gMXcr4BGgnej9mFukGydcsHusZEE9IhteVOPzUN0vVWWPm3uDEDrQRGo4DhV5vXM1kyoE9/Tx
D6YtHa8aRdOr5uHeegvAl1L1Gyup2slAL+zZR01xkqQn8Yv17arcJ6orp3IGteS1ViC3HU9njiZo
k/SRm72HVDF0VUWA11IWwVwcApbWhxDeBj1+FWntaQRSLF1DrIo+7Ry4sKNtzLjRWFLLYNFQSxAh
HFfUgFV7O8XGCIweLSeZZbTN4cZNTVf/7OWuXqXzE5tGR9J50fNIM/AtqTzolRwck62iu8LgcJjh
81r4oioTfKtNYuI627Z4UqLNEeI1qJfuTY7AAWeofZt9IIA+L2ZC/0zHUpKvCkiIyLN+t79neFqo
K3UvzV9tgVpMY+eNwJpfca4GaJksDkgS73Mlli4ZJggk6FuzbvoRJUY6LNJTEhim0SDnWNkJ3my5
VJbUFgsbeyr1U7DDFVmtb+ydJ9guktEjYunDQN96VqGA42tse7RBzSPaFWZ2gWTzS8bpZrmI4Qjs
PVt20bDfL9z1vi/AF3XIXvsStkc/I9kuBFMeDEjiZdUceaM00Z1uZPaflTdnrEMInWODem53zVnR
aQMdP3A/0dgSR7F/qfiRUHJsEiiFWWdiSUnsI8HPp//IH1zZgEtYWL4insGEolww5vnVGkqAO/TC
woTqVI3smkQ+f9Cq7xL71gYX/IcuFSKCiNg5bEBXxnWAFIa0BPTu+sLX47zk9m69FpEW5fnGfvf3
Vkgtm5JNhKJ0TMGx9E0EvAbFYkHrfXfmSFiIIXeNCZnPmHeAi/+uVJfxLjZ58Z9GoGMlUffspvPW
GsIr0zUeDe3tNrM66zjyag+JEtBOi6DdoV8mTuctEr2LGMjNTkM2Do9n05M8/S2imnPi/szOJyxM
dC9LYncxDX/yVadt3s/c1nsAd9cvDrfOgPityol3SeVkFx115iZYyTJhXc3QMcnYIBYGfbD0LUwA
geS6/AqyUEkpVpBoMUZCLOuzvnxiHj5P0bje/J9CLUpydk9TFAhPBJb3gv7zPuIU+4c3zU8qxbsZ
ePjlfO5ew1fjmWsrTM/r57LI0WfArW0PK2Lj+BklwGeM/8YNUmPOXtFD/uC9ayj9GGtgdtTfjY0B
yg27bB/yLbMhUuI+3ErhnpBXaOFCOJtE+JzeHlZWL0jDgRcY4c7f6v0CQuFxPWSo0yYqUljZ2bEB
2Mm/xgg7cZ3oKVvde0reJ79rdVBaQMRkdze0Enpc/nmH+qCrgYOWg4oDKs4PreC9XPse3wqUfOkr
+/g6qEfbqR5+hKwGBH2PyGcrpvKk1scUCsUTprJCXdF/hV+Kzk9XEEr+CWjMgMIdONy86XHyxDT0
Yxj5DxNzy6K+LN//J6Gn+DoSjDMfitDSDI1aSV08AuSYgPASqoAobMRWHwImcSN5uwqbEepVdwTh
6VRjrvd5+ZeclV1qJoIGYHREkRe6cyG0co5tMFtCOumImH5TDOegLwFqEPi8LvVdUhK9yBuDp/3b
b3Vx2KMQ5A94vsui7cNWUq/pOQztVIupa64dFn/RwCWV/x5ncY+/Zw2TTCGn5j/XjlzzgWcFPh5l
1nkTwFSoM7g17k/pdHlIMBbULB723a3NCR8mYL2zfUD7utbnyl8+NENlbWCgF8xo0Knku/BiQxVM
XnJCsjCh4kcKLQHtrskwozidFTHnBnyojR8RfWc+DvVcRPpQylf53ri2QXKUfFq2AWCwFU/lOwq7
JsSQ99vIEbQXDEl0xsHueMvARA7cd6FqAi9XkcehgfpH5yz9d8HGboUDPV51yhBhado8woxONmHV
wTtngzyKwLURpgcd/dzWVAKdubvkcjMXUne9ZC0JgdlP2M/XTaMIIPyAQhsqbK1RZtyi5Be0Rkau
WlR2WqD93TcwABHC+mwK11ZirrVklxLqxBCm3JyysxN/XtjAbCkYHVi52yWbzOHvm0gPha0DSRr/
OixHijFyix6s0A2yF01JEiVt97/Rg2o1YI1zoEYHOlWxVIJ03Z6XDfKJuGaB5TvLqv+dfxNYS9H4
W79z8FzE1OgjqHGLf1fEYDJofs9EhLPF9K1PynEgYRJW/LzIAM2/xqbBiZ0p4z8kYcjkbJ2X4kaa
lT/kcT2bQ4fEDegcj6seIJ3Zvv/TYg61uhdG4WIDrt4dvzPIv95GaoZjuIe9zQFJGuCPlhTDO5IQ
rbZNxcMPEi7md0O22Ymh2OHe+gHI5q9JhBIQPixJ9XGYcnVL1wwgcKqk40gKeFwZX8gg98oAaZIl
BLp9TRphl2xrT7ehVggfQDqY18HDq7fFmKumkpZ4Lfcuf89SLaqwh/3QSkoZLKn2DgtD50mLjObe
+i2iolIhi11vJM0f65wvakrl9IXxiQu5gd48a4qFNT6JcDj6+gkZdzd4Xa/9cgn3r/f/MJrksuGG
xf7jUDFFkkkWfv9zu7Bp+NdBgRRV5UZFsuUCTgkUBrTIifbS61RFk3y7eObiOWU4ytKXrHHn9k0v
ujHdRqjhFRJbeGcg3WP+/wBNVbHw0T+Xk26jEAnqi1w6oKymOoMUzVb2uqG/OjYuprtQEniZH3x1
GPKKeOtQaJYwrp0kE2C9/Qh4bdYSXOfNyK1dpw6owE2pmluTaXPvPddiOTltjKFNd0PY+sEeWwe1
Wb5HFtRmRtKxPY90q6jQGwtFd2sAmzcm2hMbAG8FuFDHQQlo6fhhstnxtShTwnKR2X0AgmJyMxMF
hZ0Kuu6aj3kmKziFFFFKTLI2ywu/Ke6pGvQUBJQM+V5keyT6moPcQa+CTtLEDUB3Y6djLkGz7yxZ
iO7gGt+JnFRkc+Pvcu72pnPT3TGhms36VhuWbp5Klm5lY1cllPhoUKZkeNXo/JDZ1pp9fG4qc+9g
1cZcPa4Zoh2RzWCmhujao2stVsHB3Pz2U0BuchrfOD7KIeRqF9B9EYkYuAN4N40zan5ZwRgCkRK5
8DXaMxOFbxPccsas1B2FBGetaBXcDxbtTFCqRm1HH5+HciXQC7NHmAuGw4UVRRRoqGy7c5Dc5Wwc
FLzHCZDHvrh01RLYDiFc5cBPOedU/a/T5UOiZ4uFG98Vx3Enwg5LBsTLZQKsBMK3rQwxxfJGuZrM
z+XCUU6g/1TvuEox8zhSmV13f7XHpw7qPN/D53MT2JaRR44bo/6M/5Zs6DFKjOwNhjpNr0gORgFv
ihwWBFW8zr6CbZaA/n7JwMVos7upbPRJAJ/cvRS+XgATqXK+WU4LH0qHHmvrJ8Sru1/h595klDwz
9m9C2Cns9jHLYjmBIrMcGwpQFTKODDKxab0JrzNvGpTLPgIX00ib1tHiQzyaY8XZFNagVJj2dnmm
CBurzxm3Btk3pP1Mu9s24G462IS8oz301c0lXS89PDB5sujuErL1Td+uAJd9rWOOGGcQZEM66eC9
epegtKIB4BW/CXAxK6+lKSPuIYD6G9TCxLsCAQrIOnWS0ZpVnAqL9NbxqWRs7IOYXA7GjqN5NkYO
wqnKz2tF214xUgIQnpb3ZsMw2MwzUR6JZXzc7o8YlyFTbI2nna8xOBn1jw7eMby2Ix77OLFSYjCG
MPR4eRS3Z7gFyTxKQNBe36884WmBgYLmXXgWXCzTi+SDD0g6zQpFKVWC6DwHbK8/BaOF3Eer8p37
k+aDetco/22tnmVZKYomZcP1ha141AobUAPL0bX8PHpH2st+i2IVr64X5FG0mP5d+W7nmUPpgK0L
wOEM1ToMPsnOSV6VTK58fDzusXPKqCAStOq4xyhd+x6P606p+CQwb7kGnVYF4hLtimnQLGuY8iV0
EWM8DC8b4HewhKcgkzpoW50CIQd26y0fRIFD+mTtELy3DPR9bAGbNVgcQZrluUW9V2plABYlWZ3G
IJQWB0ez3uF0vXEJha7X56coRbRk+l2CXZZ5QW6AcxQeqe7JTJ0UnnmoXlHQe048YIb7ePBRY2+/
Co4uW+ynhfBhxRdAuqnNlRvgAvovYkDWsVfFbQ+aYDtc8u1r3KlI/LdbTYb0JF/nNYjaJ3QISiUW
oqpifwYiHVeGOVnYoBUVA4VnCKG61tJxI4qCsZ41qMp8eSD6U8+vDuW1USOZlN6HFuLwbPe33k3g
Tjpn1ibM+9z69T0aZ7orrYDLTlp/j9MJ7aXDZyim2hVB4ebTnaMhleQzGVkc1ohImOXkHPdFf/iI
ZFGOpWKqYaQwnyGCa9jCfdD9Mdh10Q9Ve8JWXfo8Pxqa6RfL89kpACpyON+Iup4V0zWTMbmRzGw5
XQTa3wSGk7b+JEOrwQgsqb+lOOkcgg2fQGjThkOVbTlAFkHjWmNUEz+lUjfoUAEgmS2UFXNROgyV
WT+wniw0/DqoXPTeL2yzX6vu95/5JCrZhL5fPqJZkGXuVo2ZWex5KgwAAld3aKtbUTdr4+nNN/H8
H3vjYJs77c6HCcRcy8HiLOTN/twCrbjzpIVLyYx6z2UidaHv9OOb6cbdRXl9LL1tmbXNH2qPQvwJ
RsSiea6+fmait657UiJhBlUqtu8UDt6laV9y139evrph0jozbuPrj02ZNFx638kJdrZP8n95rYEr
lIOOgFEZWnQYr5Xq2phsMijm0zbe4+AiFdErveq5Bnde81Nz/pOGVlzv8+8IWDihEapEFVhOitDG
w0aFg/mzp1abV49VCXb4ow/MisRQHQ++V6Mzq9bvybBSgexEm7Gdoj+fj1Xm47eh/1rsI9Ve3emP
kTGc6g3uO3QraZdeKT6JICEYYbRLbXLjwLrPz5n25IzRzc8uCl1IeSYs8ZYdBJKu2eslFiYi7Gtd
pTTS2k+OnrJnKG6pii7CN6//1ZemQ2LPguQAAfFEQWCQBn1n9iGAsy70yE3zBWr4aIgsHgZTmGqs
XJf0MGo5uEyjunPMFGw3kcQ0qbQHt7MQDbiYz9+VywcSLq+SYBpbbNtc6zu8IKcAYq5cEZaQfLpK
ZBUjaGpi96+l5Vg56r56ZZ6ovmXGGIFL53Fe5N4p48+kVQ/PkNp8Yalrtv2SM3zMrw/SAjIKvrMV
y+FVELoZJdXWwAP6YON4zCJ8BPX0iws5m/EmF8nfVAZIpJPY/jSHSM9SW25/FywnGum0krhCh7x3
O91I1RZflKQmg0Ip+a3jYCsHWecq0eHXf82tuxX85w/6QcU6QURK2BViHyJxGUsv4Z99JxjuKarr
KzQAr+rH0D6VW0//Q8KzN/vHKg83+0tewphsYRAJWDLliDYyNzDt0E3UJyxxnVVCL98GZPoG8nOA
nGVzcz+QPtnz6knUvuX+WOPHVp9vOS1qUIk6yvitZE/lC5DB3op5MpWkBxClcY/wFrBV4QEQI9ve
hl4YaWq7JeNcZluRGD/LI2KZcac6+AKQiMiFI49ND3OKDDVOKjwf1qWrA0Z+727H8hTgesbzSerp
dT1WrFjdUnxoQmO83h6zgbCmgelMkNt48GMCAERgbNzMj6P6byN0UOsNXC7Sql/dRs5p9LDyMM8V
z4PUVslxfHk7oMMGsRxaH+dUYAtnid3m2t5Wf+ozauc22TAdKQC1m1BCSM7pE/W0xsc3IR7JOPfl
Vu10PlJ6Q4h56H0qltUepchNVSFOh0+Fi/RwPpO+CKgXaeQgqbITgd5giaxsRglAPfQhOWSmjrSR
mGEfVr0RQl7WVwJl4yUkg2mP+G0jYsYez4opJQlUIj7VQYpX3QfwNLGll/m6Z0MnZDtOde/e6kbF
2h34+50REQAbEwVeoRbdRK2kdlYzTFdG/49xyAc5KIxJtGy2ORz4DLUml7ljUKLK57Z64ErPcJUF
N+pdNTA1SojSsEjosGQy5kh8tiZvk5BwrsXilzFtdmWWhxKhI0h38sWqgsNjyASBrRBNKnXx7ag8
D/YxgWV7HMh4D3PvG+kV3+n54MegWYbnLeQebVlPSiZTUgQBIE7aOugnwcsAu6oI0dRaaRXzFIjb
Ws/Gnh/y+Nt9p0aotuH1m8Y3Sbs50QbNzV/27MEO1Njm05JqWC3pZ0jlWCh/frZhEuxePHP7Pjpc
7Ynv2mxOEksycMARDj13wCGatRKdwZdz8EyrAucAGDaszMERAooJd7shGC+0ZLnecGaQKro0W+MB
st7QcIu13qByh4AT6VfPw9OCFgSx9+OCYLcFKIv2qiy3rY2cdhnQExgrdWXt6vetk8zO25TL4caz
1ashlI5aFUgEtRqScfXfwVPSxyc7sj+SVmvONrp9/+nWMHY6PfJEpWzFFTlWMAcoqgYwFlJBni3z
wb5bmMynwrJ+hlC2/x6KddYZY2vELbVNcs08/rRFcQ+aR5s38zCRg8BajWlXJtgX7/nSSkKVn/EG
WM9GTaEuIH/ySl97S6g2gAF/yKnF5SNVOjn3o6glpK9BXXa2isWJzGMLHPyt64/SHPA6bBXBj3CS
ZQ7TlAcoMx9rDSG0Ql4fMXkDISx+9CaTglcdBwhmU3YCqCMeHjdvXpmryh/cgsJQSy1DCpk2NNDX
wpFvZ4G3DBZwoHvUGTAAyY8RIherxO1yY6TfJpAJMxrGM+1szlpX7gt2exXnaV2yrltq6SNzO5nR
2dHAECvdiQEafYp7kvPgwO9vLrT7OG80DochsgvJWYJ83cto7tEFeJPhePhSFdBixH3F+rgMkofm
JXYWyRpf3GobAXZsQf7qtxr3OlvX0EJ8kv83WjBs/jbpPWq+4pHoMRAoMSF8NkBr/bxTfZf7b/rX
xa2rcPZYS+FGLZE4tUu4DTeP/UxjihUk/T8lTqy65LXFKYj+4w4Ka2cUf7QO+zPamSOY6xpjHwbM
bni5aL35CNVddO5qbdutKvo1tP04P3siKsbJZ53fd9/XPZDFOkk9qLb0a32f4AlO7if/Cirjfwh+
o/fkn9I9mqXAbOQ0dzrsjT3GR3bcVvBHpCK8UxqUZOcSszO8U/rjFmkmQ/CGNeAHmcqJd0TihZUC
pmdYmun45A+MJFS5jA54LKZnzWscy2FMsCr4ENZMTKZCfF9MY/j1vXzHrfG++Oz6ByD3jCSMJSgp
sUdKY6IJXSfVz7eWhVFSoxfQQPlr12W9MYiJgtPF/9JJk557tu0B2b3WqyUTV6kkFQDibwKK/QDt
cnCcfpl0g0dT+2sBtefpowUviA+e7eFRYerkM0H+2KuBQFew+mk+2MQ3SK3bl/9zmFROG9lwX5Wi
WtGUX9qgXWIidh/V2J/vUVc2lUxmoIzA69TNzNL841cHg4iz1B383b/6Agyyl0gOptM8fOqBfvNI
9MxI6qPDadf5wPMhKegrztLJsjlSJvtyo4hkruH3cOgxo0vd7PiAzqf4PVRBjs78TfVnu+yYGbZQ
Hn/EGk5c2qbwh1l7CdZhOu9T7xe5jMCoKmRvQ8VjC2TIeZqpgWtCo0g9zr/YUWkTgO/JeC+YREDg
yivrSEA7WPSDaifXZq9fzXAbaQeT9gkRvwplIgEho1/Ik6XFNWpcdgu9IzJdUyPqa92YLfYD6b3T
alGhpew+uf52i5J13bxV7j7h2S5nnsVKNK7MLuwTnhIDGeCly+d9ayaJjhdAqANqSML+5Xfu6tHc
u3h52l5kTkUOy4yxT6KvSMeINsAq+foQ15/d+ufAzQhBdDrThs7Rx2rI3VVa7gR6OBXsahNW9jU5
sknZkDrmxq40zgzDItXK02B+W5MAnVfk2o942dvLzxnQcY3m/EgyqTXdy97xs2gN7PzXNpXP3u9L
feyvgxzCzsBmVogG3Cq0QLe7O5Z+xKDk+/oEmJtHc4oxIAJwqKB3Tj3au6p0D7lTsaY/GkrCvIPT
nFGfJnUQ2lcLXoGYcNn8b40KHpd2pClm39yt6mSCr6Jce8DSlaPqyaazsJ6D86ISA0witPY+pnub
EZ8uamAUazs+yCXVN8eEccvhy8fe21PvYn7HrAKX7QQ6LxQsNdDehuFJ1haCQXafEf/+ZU4HYMgf
1MAU2gmF4FSqXSWIUzWCIznclI1Y8yzeUXtcWWuHSGSYIAN4KDsr5mIJCQfd8ydlW2znXDBf+sSz
daSJ04dSABwKOc0v3mLNL6kCBJSBbzgVjxZY42K7PyB2N++iOmOe+SsYorhA+nVWnKmlfpxQB2Am
5qeRLMSLcwjFDHqfuRmwPIlZTXL0QBxi+601BU7C4FaY1Y3otCz9v0rlmebhQM1HmbKYyBHJVNZb
H0L+nedw4XRw9B8LOu/IukWwwBZDjgb6aMA8HPs+LcDaeHKKTXSFioJHBdIpVLtems91fFnpSeC6
6XVox2l9qYlJyqE/Qn+qtXII9iOsqMRkSSwtFZCAi7Bb1Fgj62yvzvCgPWIBSYZxEjY40IWezJR5
squa3FrpPsW9nGxtV8aQUgQ2acQvhtIma087C8fM9+020sF28XxDA/Jbmv2h9HyxdwDg3Bh0V2oE
5g7SLmen4Li1rX0GWOj+vIo6ltAAuQ8gygw5IK7c7QPuUjzvvTkcsrc0H36SBaxvoN7pB9wzc1CV
YrD1sx6Ti4crEG90bqkYR5/hmRFallD6QDUamkasuG+0VKl8Ha31cgYVbK6SZWMIsRkyf1b2Apk6
HSbjFL7NBBzxZAdafrSgOaxi3FEO4wXanLbKAWfehawC32PHE8phCP5obcezZSHATRAdgHVRHdA9
PYnBMf1FZvMQMhccnQwGslSbEAuoAXL5T/y+l7N9CPEttWbaAEbFloOGJsEOh7nZ7HaXi7Z8cnBr
ENe6M2k3cqBtUSl1n7THzTclNaW3mY+6Rx+QPfnyT7YS6/XG1Eh+yZ5ozmXHhexhUOzJdB8xZtyV
3kmLGaMw7loIP6LdDUsSnMFrlmJ4ZJ5sRwdOxB/Zvo866HNzS1+5dw3eDWPmVotCdmn7pU8aICVS
TSuSx6Nn1vS89zAZY2jEQfF37tnAvEPuzIDyrvxUGJoWaKnxPwRuFOenmhx9uU2fCBymbjnZ/D/e
ydHI9wuWAsOvJrt9OTjpuX1lAMviPDcNw02lpi7USxKIEdGyHpIXXTaI2IABZD0zze9G/WHNwhm+
QcFAQKonmAN8A59Jhv2RDOk9yjtMRCef/QxZb1AuoDNp27N/kloWnXr3Lk+h41/+I12gq0Ux8ffc
r22uucBt1w2XpSI1vvHzsUDMszXgwhtOM4K727w25nsBM9Epfb6lKwYQpb5NgGgxAGfbwhTYFSrL
dHRGLqMk13b3HYUzj/FUXagmCIllAqbTaHMvqe/cGShrx8QzfpVNmOnzecuJwWMtk5XwP8vbRxXz
OL7E8YPrb7b8cAn+XMxw2v0V8+GWSXiMWAXtKAS/dK5w2FTI8YEfKOknuH5aySL5iC6gCl98JA5s
GL2EKKk6RAheoyWZGReA76eshRUYfMBMVTquYgg0Tz0Hu84uttBs+ej2vCHJfMAr+kydNd3KV3xw
5DxeCAKOsq6S0ww/QS3rG6fCR5rMbrAhpVXuK1pO3EEJFnwxTiqaRZoSfmMMXzsNt9A/0W02GiUw
tkDvyFlCCZNqh28gmwrgSTAzaInOSpDqHezY3aKIK7OfBYWPJj46BouXfjQm8vtsF0MWJZXdorve
5RzpH4Gfqe7aw945zQjIKVoFJncqMAre01eM7Vp/i4/J6LEGsHKd9MzQ6KJRtPkwfK4vLJRhqcTK
qVwOATu82SHBCpLMYs0Xx7ePegQuN1UaLd3IawzqwmzJMyF0vW3qaL2felObFzFc2AlghD+ebZle
1091k0grEnLkYDcCNqFcUUu1mY/qGXhTYLikLgjJuPvKzoHLJ5zcJYc9R+DfposAu6i6KWiU036j
2c8n+sGdEI9PoU3ox99U7BIIsrg9K0I/H5Wi1pQO9Kwpm1npELcFmdi9JfXZc4aOabaD9DjFXufQ
huxf9fuLpij4nZaWcPK77m42ZqYc9gvIHUad0XGFb/RC8hDsz0dg/75no7JHS9sJrJ3tfGkd7/pY
tqCw+GWOCEYW0Hv3fRH2VFaEwR1t20umfEUalbAWXZ4eLxQ0xuG6EehGD8twAA10/Yw2HuulqzbF
4q+c6TGNHRU6gjVLekrKWOM3WbG/cFrdHqXdeNOgUZYjtS82oUGSEwsbtl2oNxbKOAeArhnT8uAS
eiIKR83KnRjoAiexAA36hJtYGJurQCUeKVacdYpDuMJysDYXD1XCkMCird3v0xuy7F074nrOvcd9
QP19Y5l/Tf7Ttzr7pVBPChMWCNyRlfp3lQnPklByQCn7f+QpDY9xurg3TRxKOXtC2oaRrOzkrGGk
t1jfFqDbDVI86NBM0+LXpauKs55vS18aRHxT7Fie2srEKBQhfdykgPrMhg4LF1fjj5TPS3Jq/coY
yD9YAnOCTEbh+BIXF3XBnmHNQMdTuDRWsEXpw8QpWonVay0/tIc3unhfiYC3C9Yt7I9Kn4qyyNGl
Sx3Jaqk0Wkcg12GfjwSOWqmmRhvxd5wvTDBCycdCiGj0dvoy4mXFUDIj8Oz9wotIm49hN7wpwkzo
G3zwuk40FYCrPUAJXul/nVX5X7/JZGaEOYo5L/flP3bue0U5fbrP8VNUUI70CzXtNragLxVjaTZN
46M7McJbiSm8YqkzEm0W6oA8+0PGK6jx0EI7GSWAj1xCaRdgNNugtDTc5JWyvCqCXp71EX0RH6rO
/0slLQVwSunIdjtfqFWYp/wKL5w6pI8I6w13DRXUU4b8J88agh73icOXx0k39c2kWx9Qbd20aXXW
4gYSNSQGPmxdJa7s3bI8XIrhYvhxV7jhgk7d1XKklzTkRlOs1FahLpEObJxaDDV+Iy+93HxMn3zq
x5xd19smvMQ+F2a9a8/LxEirxUN8p1NDmZstYBO+o5RvfmniLQYW6ECB13dUGTUnEm0FLoqE9Drm
E//m62bgyg6W1e92dkeUJPmrLgfw1C+HBqYvLIEtt0NFeIrsuReXFi6k+q8ce3GnZo8ZoJPEP/zM
F0qIFqGDug5TCyJdcOrfruC4eHtZQOAaEdsoGtznn3kKsfp+pxEagTuyP0ymseCn2SDHB6Cmr8kG
LhA/iDQkcNxwm6qxbMcOjpkV6I9VlLAmtpjnpE5fnDL7cCKdPudXv155EVsW9LU/tKLqlrr9vlUA
ZIkbbR3jjnQkX74QjweSfe5MC4qGotzKfyGCLAbVPabIdEO0Y3a8JLSozEBlJ0Nc6LC5K39AKx/G
3Pz12Admrm+HBDKint0jdNrujffbZLt0wN8M8BCRXgcemqyetva5R+rn4sHRq8a0akrpfH1vLE/d
TPmub9ndIzH8O5OX5i/Mi7oDJZEKJlYpS6ohy/MfwdBuYp7fofQXh2xzdx3JUaM+/DtOD/vrw2/5
G8nJRiPTQZ64Ai9IJ4JZnJ97gJNl/HIYMuJyWGaI43w6gDZIL4sxfXJLOv2PZFf2TGt2aHbVQbkz
4MzOg33eOpILzCLyPYc+Po4f9jKjc0Td5h6a1eAomLEEVEFGLfT4KIcbiVxue1N8zIN/fAV/h4U7
hsOfApXsYBCBSb1XEiuCyB3o7svBiAEYrJNuLO5onh9chjbOWFy6jPohVoqj55UtCi9NtBQWzEZK
4lqAxY5v/S4i7KaTOQUvx2Dh3Il/3Qf8tRdX9jrf+CCgeLfQpHucwtu4NsK9eibbBxzp0+oqhR57
AjA9Ksj6JKcq4eg810SX9T4qQ6NTqp30cBLayZYPla/FdWcMLp77a7ZGwHbtTZJHKdF5gZY8k3RA
Xw5//5cr5jqPU6LQgsd9dqedJq1KsCaVkU0EmbueASb0aF6AAZHfpk/TWqGwI/n6wCgElZRX9768
gj6nwjKQOnj23rj3uoac6pPSKI4vVkyyqZCsufSLKhRDoLuLBz/MXzMV7qmC/tYxXoVYT1MUK9Tv
ztNczBApivclFJCe/rfy8BA7I37lGadxLtLTGDPJ8qj36wdwgtjzEDd1DAL2nkcOdtA8mM8Bb2mI
PdtyU2Cw24laJm0JwkUBW44V1X2pH+4j3P3DbwNrQFowDTIjaelWG09hsvcDZBIAeR3ShEfLLd1t
S7FeDrwIuNP7AwCaAXo954GN+QHa7eWW2siZZKPfbeQSqzIUZINfC+3V/y4StzsH5f32G6yvv5Pd
o1J5IBFWewhT8eV7HMxHYTcjU3+7vcyAJ2tVVhXgxSp7WyjFKHWLnP0Hbm+LAp6TodRaac6Yv5GI
MwDD+WiVYuAzrb0/HzUDrlLUOSl5AF/L+N0mlsQaoS1IdpACrh362chG5SdSbAPyh0TE7jZPmkYf
xEOYRD/BQaQuKYHnlTuHSsbrJbB4Sddwou4hJwxFfYpiUHZ9gAaY50BTAT5mcylSR/2ocaiC5neq
na6LG+F4Fw5xH+2BVrdGinD8YvSkyXjj2qYeeUMLAIyy94UaN14AfLCnOSMcffSkHcx3MBUjmceg
XYxwOQJHYh7oaADCH+Re/rmCSUpyqHFldHCAHs2n+3sfnTlu+tPn2gw+waHPcXi8Q5xlFihB0fy9
HaXGK0insxUwHoQ5vrsRvouwzW1KmVDABAAX2ZxzZ6LkS8SP+e2fSF077thRSkbnuk6+b6EFTg6f
eMGrMumh5iI25tEJ8v5jgAZs3zmTK6Oz+f2NZ1yGQHcqBdjA8OfE9ZuJYKZIxqagRUv0seqb6c7i
YOPO94fu3bbMrVLl4u4rT+4jPulFFsNCXyPrjIC+Q1e/KIKoGYB0c1AOElewdBRuTiy7odteZrZ5
CY6neKRASmcZgbxgXgrMnPkw17/jq6U3xs6tpzsFCIhS7RRVBzNMy1Lyn9xLEqZUaRiiFYmP1n2b
QBxd3ZHqdhvPk+OaGeqaEjxEjxOc6hylk9H4JnthnaRcpoC4EjU20QPR8Rfl/T7uPAXQlKs8VFoD
leJQNyYoN4g7hWO75692YnJqti/U88gTUUg5OGrrkr844ksP7cIskY8TAlEjnnK+bh8S7ZMe47i2
FBihC9BopE6GF1+vNbgWzbnNx3Z0SQ8T+Sn38s8NwF9ZtQHVkWt+0JAXa1ShEya3DpSCdREeQ6ls
V01lCIDZQ2QS+YBiAfjqp2NjmZqR2nVNEOHSWzNuFecUxNpCPQY0kvZkT1OhOseBNm11uCZE3WS0
6Gs0OYeoG85p++/7PdxC2gEbsIla3t7ahXPLgfZeuN/iRc4e9F69feX2O8ygYIG2aOFTrsS1w/yb
ZdkFKTWeCkLwN0ncpMvv6z43U5ilcBgaKK5cp5YTOS3vxQ+FTt/hITZfYptOTeDCMA7LVXRheoMm
bBYnK0E6lwyUMDRNFj7/2kCVQ1V4RzbZVNUtHsMPQ2izM8TY2rL8/k+iJN9ri7ZCu7nqp/DlpAh9
cnGayrk9WWsskt64sclwLheOqsuPv0XbEdLShBjhU5K1w8By7nT7Apeb/9xZAz46hOzCuycfUWvl
tBdA5iC0CWaR+QNusnPqoZqqg+EDfivUQYD8ai0DWTdSGXp5G+/436fBRJLpImuCFCxdRN4C8xxq
FZFvgXlIPaPwEC065Mp1SZ9kC71YhrcIroNCpPFPBfa2qQ3jjRls+S2K2QpoMvo0m+900v49+AsG
QGm9uFErZBKNDllDWc2iF7aORfgKsEWuKtmzofmhyTn2hrmNSFtcMcjmryDzNB5fj18O74mooT4x
XwNAqFpS5FIG0H2VHy6TNiixruPZmKBesR5LdX8hdVSVIs8su1CIsIij4K9UiRksCkePU9rYAPps
rqY30PqltIXSPB36ycKFROTQMXLeWJtiT9Mj9pSMF4+ArvsV5uAN/9aYFaNy065+i6NItFSP9iJL
TNbqLKJLzEreyLgaivTtkLuOwCGBE4ElBboZQG8FKQQ21IFkJw74SgCh0/1ai9oDDvDE24UtF6fk
xe59rWeYad7ox0JJ5SKjQQ9pjYTTu83rnyaT1xw6Jo6eHhqq+fu7AXNLWfLyI1pRwjjvJwTocDB5
0e8oHyFnEHy2JQYZjiDTkqwR1cr2jowHwQwgw74YofBOxxqpaItyQF5i4/SlSDTjRPuxQb6M3VRi
0nOZViXc+z+CDOkxx2jqkKZpH+I0agFGNtylmjO5C+l4AGFsfj/eqFRs2gML6ZHXXQ6bvLSMRxp8
XbDsr7G6Y8sXRC3lzgJmEAayU4chfOtuvFAmNdkuHOpL0mhkaeOuILzQuLA+H/leGpfGI5Osq6Nd
XAePdf6uzLq8y2RapNdBue1CWIofoJhWanEcthco2q2xywpujBA1naURCTnJtx+Z6/gTRFkoEqzP
Xe5gypNegalVMW1l6Xfdr3VShq7/D/pDn/jlmAdsq6ySB/oOhZB7Kgjo8z1k04iiTG8sbqrCBLUp
fzz7+AgrCxX/aOID787Aw5kAXl/oX4k9CvQTsh+DCVZOmDgv8yv5QxTlJHuJdLKy6wqgIQL0WB2L
kSND0rlAiGcC2Sx4i2qH/xhb7+GdRgKSdcPHZxt0a2KMz9sC+zKEVcKEfLVwrMQyTXz1b9n/kUu6
r5euKrsKVR6V8Hx06LTFc76jTOO+D1KgiYhkJiWm+utCyfspCDKKJWN3ZGjZgglPv6n46vinQVom
CMsMrW9tWJui5gfQudjzjBKXEigX2qOdKxI071xguwM7DqGMNk+TZRCjbnCiAmppqBeC+QVa1Pe9
95wEowSxzLAoqrn6xS1OZgu0CD68zTkS0aIj9Mp1nz+yHf756jkXyHtcy5z06BcRLufDvnmya7II
j19kqs/eV4qZRSUYFxdqCD5z67qqO/SGAj+03JSrFQipNUTF3bMrKfKQjA7VdQd97ffVvJtcIZLV
U9UJM9lxOPgOLTmuRTFHCLnX7EKrJoKDmELaD17da2uWKvfMMlITU0LVEj5qcGkuSh4dXARxSJmq
54PIYjV+SYq4Cyes4d93b8fSODI9SRr+tjLdMs7EQ6SwW1bs0F5pyrXsC0xHuy8B8RuYU3qBGzVC
tZQRgCVFPRmGz2X9tG5UTombCk0ZC0p4IJtk9ZObbN9vuW5a5XUDXdvpTktbWXRiLbf0zYiA3apj
F4mlqHGMTH5wRkT1aiUamd7+hMXw7TpTYF2nEuqQid0td1SvjuY+ak5AkaKsKkKGrW/yRKjePimy
cw93NUNzZmUh4Gn0PHyAIRUbpTGlU8YrvD/9vIR1rKxa9UVL8KhMKwI6pEhxQWbghLq1y3s9nGN+
5a/0p9pa7xAFpu74qQAHuovG3CeZjvnv/29wYmvHPhDgfN+Yz8hH+eCcgkkpvdomaXaOKUyqkk9l
rmUgfphGfnpMrhK29xhpeOTTGGb1Mq917jAO81BI6wIGIe1AUSlzcG/09NyERbWB335vCHrTy/ck
OosDt0tPw+a30PXG/JS12aylqyeb9Gd9J6EV/RideSBn0qBk9if7Ts2IREgfKJcQw08j69qZNEk9
NFyyEdLNh77XP5tckwax+pptoH3TqS6PM9CYhM1Ly0+cD2NoMD1XhL63nB98jA4FxsoiAL6ElhHB
JOx+0/ZYCEZvxXU17M2Xf7eZUqhmSAZfXBOTE7WORC9Z5wQcMeGUf2DwclCFy98LvjoXLBooQX2+
8SGEo9aIipKbtykj7sNQdk0avWrxtN1prFpKFex8Q5AlyAclPrylE4tvyKo13PIO7WuQ+UeM80+r
3ECFUyALpA8M+jAm1Jwzu9bsYCe1Nn85p69gHOWgm1XMIn4gi0H//0aTRq68P0uR6Ssd2j/JpX0q
3S/RXEXbHJ5HSqrtN43yLehNiZmfVbltmpGc6gQGQAVXGg6R0vyI6srjzg5JYn1bYTcbibXTMdCY
VbcXvBX3NS0vpVDUMq07/v1CJ+wAWJd+F2w7REm2eVZBSwIbqhHiMF5jqq9r5EIDe+F2b7OUD2op
KPj8jmhsftG5xA+N0O3RtrYndRaL53CoKhE+vdxkkDStANlHk5xPz7tfdCXr5P2/EcoK+YjKBfMn
4wZyl5hlkwgLRzf0xh0nLT30I74WabQSUMSCY78jPU2ODJ3/fZJHO5et/tCu0nA7pLHotv2ngdOU
YaKjoZHerNaWCCKTQu3yUTw3R7GVFFCxuWw7+Mh/MGRiwVhwFFtzPPhAelTTnTQJvu+QAZxu24QT
SKgRWuarCcAibOcx7rdsORa7qnl366Mcf4vjhqMSJH7OBDF9J8tfBNW0mFNVWSQOYOoiwl2D9OQm
lCKLZX5J1C77JLhu+bJ9pb5JemtWsL0ouzOoruoifwaG0LbI5XYHai3baBbJTP91CdLZRpPd52h7
3pdsO33cGxKYW+clyqCICyVh8uiW9YsTNrC3LkGlQAQfyUc4gm3puuIy09onF+ShQjbLo+x7JM10
s8khpN3QCxt2GxRu194XHbaoR7cgU6l8jl27lFZC6oCtRaEeU7HTLgK3JyyIcwIH7S518GLIjzln
v4u2w3mg/8P0IOAJD7N/5mJkBjLQ5Yo0zvBhR/Jq++QaYdemusX6Olv6Xvfb8JimqoOwmd7Prllr
H2W9kSyRLhUsvE03rVyLpKEnrr3EzcPV5B46DBqd6tfYaqntB2ZtADN/zITBdR/3G7gup+BJ5mzR
lRjMm2rKSo0Zt1Qrw8N6tfIJSSE+fhPwPHTX2h39krK8XowctqEoL6s8MAOqwJCkA03K8u/77ZMU
feqOgEF9kya1vSZrx2V1odIwNn+Bbiw4qCRQ1uPzl9z4QpTpqgix77/UhogAH5NtdhFBF9PxczTN
MJkzf8EpSUtxIW0Y5gTPZPIUaFPkwebEfmOCfV20r7OUNHckq3vT9/B17pHFIcm/yFNOz7/JKIvx
dHNIFc/ufScWhEIaleytDrucyxGqCsxsBh714BFx2vLw1ctvPzNv22aMecUA4a9JSkJtDrJaEdeW
Yp+eifx9dqSbR8YXfuqWaxGSEJ9XK1r8R9TOAcb57OJnpK5hYI+GIKf8j8mT5cFYGWuR9/AjgtWk
+/T2zqX+4lUMjezH/msD3ipGQt1W+TkNsjjPsh0whCAyTdv2x01NSUPFYRgcpjWcchpAhnqjoHRR
zVRFZnAmbI7h14x38QoxJhOPg6hbzZ016WSxXT9ywrToGNX+dugTb+CJOrYXU3A3HSyH3tls9Bcq
wCl0ATWP3TRDO/TfrEfKMos6vmh0mI8XR+5fsdG9gVEBliTae5IqRKhfTaU1tpQkI1Taj2UlqZRj
UhTVlXpwsqOzi+ArjrkVd7kluAVE+rbTyrLl2GRq2lIgdH94SOwhRROoJkivjoRGtXB7CbQar1AS
OKAC2neKogU0Y/7Qh8+1qzVcaEAf+GJITY6yoqUJOF2nLGihRW7y40chpO0MYUG1NXBq8tgpTSF+
2pgh14++Ouk7tcS2i4OOUdO9U4kOd64BbeqHe/pSKSO7A6GCTio8bUwPW/AKiZwgw+qI4WISNfcm
pEb7ZCtjvgTLUpj+U/WIXorB+bHi+lOZf1GPrDeL0xan5l7KvY/ciMtaH+1/mt6BJGsiXL5x2plC
Oha0k+p8kI2AQMYVAt2DUPpxUjWTPQYXzMo7Z98Jj28xu/zF+8xaHPzmcNX9UKip1q0rGyd+dw9R
SqzOL4ylO6M1YzoAXjqPiBHYHilB4FUZHIwBQCFUIbRMfhfFe90jiuYZeC1z3NIiH84qZOaXzuHL
PSZw9lxN/kn1GnoQ8yGeraBk8FLFe0ZPP2JkQQ95BG0kDgUq0yKdHPrNoMLFWKSv93BC7xiy+buQ
vakDWpbjAeOB8uZUj8QM1u+vjv5mjojrnzW5r30XIst168Ij/cXejRnvin7B+X7hJ7rUTMvQku4K
ipDFQwIbby+wOLktbKhs9cbiKMIRtyjLn5CnqLWGCj4qTv3jvgZJTRNdsE/sRvW9SU4FmSIDq0BT
YmkufvP+mWVT3gr/j9dVMBHgF/xO29x6H6/oj6ccd7ixU2OwBF+u7fzqVKcypTypfAp/KFakYOit
5Z/VEVHpIAHQ/HR9uTBuNkOaeYDjlXwkHQvzbS6cuuoBIYDP0xpD1w37Xu9KVNYWTV+Gjp4DWH68
mSFgifbfjgWLd2sCIH9gp2WlL8Uh8qeoiKb4bR0bUKUuo/U0N8NpIf/gHNPOABxNtPEXWPvT3hX5
5kGuWFfNlPUnqEgNBzv08PUAzYHqqD3M/i8xHvrZfTEdzkewpKICQEjkVsWk0NKpxqGB/ErKzRKy
g4E+m80s041vwKN2cmx/4/LsT48lN5Lp8gbVFM+s8aa3u/g4EOWkp7w5bPISHLtS2tvCCgsJaCUS
ke4Kt8IeCK24a7bxk2mY9qhZuM+UajgM365Cbtz6/qJz1a+2PPrLfMXBepZKY46LZ3+LCfcJX6wb
xHZpFfimD0Myfthk7uc4iJ9JAcOVkT8Wpze69prEWujRhWHhLfgBqELDNEyLVOT+SXMdWvCCIK7s
PsP/Tn64IXt7nf849hkRwIriMtgLYONuXCEgMzKzhzmzndbq7VUxOV6TqDsD/vrDj5jpdpI+VYbi
t3MqCEdnzhLMlUgIfWIc65baCVNaotwUllWUS/ih/JFT7QCMLwQUigmp0lkxzWxTzq6aza8P5i7S
ztPy3k7G9TFss03b0p8G/U2Mngft/hgGAmH6BIpaH66kWEnMz6y5/Fou+y4ewxvOX4M/1jJsX5Ag
zu/nhkpL5rEmw/cERMPGeuf1ZV6gRdRcYKmxQcK3ByixKn0hLmpN2XR0ofe09eRntCVUuNzcK8hC
ajQKhhOio0h0emC/P6MIqNCRENbDHvOfwAvK4XPHG2CvnM3mLU/NNKkwg65R/3mqT0lHvI6RONoZ
qQB0KFfkjcjUuy7f1QeWnsg4h16pK1zRhH6Y0J0fxuL0B25ZKyVJPnr6d7vvN5GgGnzkxqFl7JX4
px8yRveMx+cbFAkHa6QXJknMDJjdqlZNMLuiT47ofCMn8P4kQxkW7lbbjq+52WN+NOxMeg0bprt3
vDSekxSDmpG4yNhZD2V2o9hJd5KWvx+ky8JoiLpYzvoAfFIK1lC3BrNIkKwfpYizyKlGXolI0L7V
AUSoY42ed7QWaNX908yg7AnA7RUKGbKDuLr2C/Yy8LPwA+h9XpDn8oRdxtOPiaJo6FbClboet3OE
4R6y0XKTXoXLu5+LadSl6cmyMjvpNywn7RE2pXSZadA4LNcg86ELK9USIyvXkQn8zq/u7HUUL/kK
brIhGoZtFaoinQf2lUUP+to2z1eH1FK+vhXrqjqo7/M7s/EiiV3nYBk0SrrBDz+662cz67NUni5u
aZDBnrN8R/ekZ6XfY+Gh8AKvWGKGGwgvV8AmEMOliJFDnG6gPIpO2UPuAwHd9XUvzdg26eQQRMHZ
z6/41pLdLvJPEhGVd8lEwSg1OvEesbyRBGmg1JocHBwOECfipduWYYr+WZNsQqHv62eH1e1Juaut
EfV24/i3FamJOpLzet5hCbAWv9qWtqBO9Xg3qcNiWGf19rX3/TSJsSqnhmbF6WC0A296LDcGqofe
dyn8MxTb374Ii9PuiR42HUMQ/uMauSHJ/+VGr8j2eEeAr0ZQ3QOKuh0cLuEQrVGAXSfpYlguu96Y
UTZvZGSxGSH72KzSEHbAj6HKHZ7cTuWXvxpyoO6Wu4wVwqa4KdcoxVNozTkhkwoUs1o0zux1gdkn
O/5isx4pvmH75kV5SsJcEJ1WhuUTbX7njbfD02+OzNdo7Abpb0/tXJvcPh0GU253V7DGJtKlmOpp
XjKrTJr9FUnpqQ3Bnq07RXSr580edfqRCC3Bq1DjAWLFSMPMAxo4w+h3QJia4zIJAr4KUpr8FaJr
b5tRQkKgpPREELI9PzLP1nZCKU4+u8LPsK9XPnW31geY0UqGHGrtTKMYfv8GIQayD6cacZIy/HI5
uMXrRjT4bpPPxYVd0zS7CjhMp5laDCZAKMeFswzqp1b5bh6hOromRQwmXe/VjtBY2oFOCKkaJmdZ
vyi3evRu7LtRZNJIyupobNRQZWc2xtxO56N0DJwgSRJ18qGg1yqJoIRnkWu9oUVmDuMXF617RCLL
yVMgQGjHVBYNS8Usu0cWTgksKZ2/n5RPwiyDCR5v1/qlkUZhsJVx0AlRZP0BIFCWWZyoPJ3/hJOO
AlG7MXjkEISu3rw75vGNQwQ2CQTgSm33mXZbLiikIwHV75sX+hrT+eG2T2SJnOaV1QPyvedaMrzp
XV85wn9YP3HFjGmTx6Fxa6cpWxnjIg9z6LHP2dsSzQDGc6Zwdeht3Z2sdRtMLqeZvSWolSidpoSC
XSgjeeQb1jvojU7wYoYmt3/bjMjqozIHOHLkKnSRI3vyd9sH+GQW9KCTwzIfzf4NUkT8+1QpkHFF
2ajhkfeSQbR+eixGdYaK6Q9SmsxHVi9WGHYRYtAg+7R0X8pMMZzVVKp9GiijK0nAleuz03MopUFX
0WmPUB7pA8lD3CJlCQWp/1oCouu0tzem4mhXPDgWKVN3dkrccVkXfAX9Ayv7A15wHRqPEqGt/kqd
yAZLF2K9tKMxkBFQxiXJnocbFY7auywhOMXr/tB7CLOjbSG1xoXM5vZCnDddLkymrkP/dQg0Kh6k
TV+Xu7EDJ572ni3puJMDe6lfP3pW2wy5fmE0SZxYjAWcfjW/qkvYhNRCD1pExiN7Ay0pxzdGWK+B
6O7bu+UIKgnUpwMOAacBPX8v8RNJEmI7Ks0iA4ijm+/wsvpXZGEgo1FnrjW3IYMkVBTK16KCtb/O
r7dliZD+PdZgruxb7GlGk3b7ACKkEI2kLqwH84E56cj3R1eZKA6KrD4JudFX7Z+EtxFQpX4k+UIP
KO4/rOsk76p+oPke1mXr5MlOPa0UrHgvz7BQSIj8daHP8BhomLi8Q7TlYITRYxbGLlb/ytm1pVw6
NV7lYo/QfhHlq5KWr0Zl0xR7t6nfCFJyQSPha/W5I+CrYXMbSaLhH449nzpwQNz7PuxhkNS9TFBq
yiqBSixe1htC9C/10j9lrO5AEgs3UwkDDoAJ5bI3DFgJ6teEnaKY6PA1h6X+pAASPH0o8wRklDcl
+FNA8LShQACEHFSyYwXl+hssqzQr6/yLKi5y5Vm4IsiJioTy9qAFoAe0CvL3o2LDsoxhv3J1DjQt
cDEkRn6MEzm9PawlsqT9++BfvHO3vhaPRjWj491T224MsR26ojzOgHNuE5vcueF670DFsN86PfPL
DqOrz2S6VBYqJXZxsIRptHBgohobPSOkdjMrvA0d1fb66oXW1Xxc/dpREKdYbj2bbpPhHq4mA7Zf
hdABF+wpbS0AQ3ynax7iyDZyKDLlAdfGh2rNMd/fn9NNWyLHDjrNcBlb3mVoY+CSg2F84muNDNs5
d9jH4m1fXaBS/T3aLqEQZDf4AbYZOSnamYgXGjnoUqk9ybf92XeKV0M/TYnRODDiMCCsMhZRLWAE
cACm6rxcwKnK/ybSgKrmt9EbFMFQs+MYWSwTbXHP7xn8amJUzMJPdbF1xVbP8uOrBFBjZE8vtbco
6s6PVeXf51WtauykALYc4Lnwj1jOQ4LSbiHYZaDH2QX48o+LvHsUnE/Jd8gKtmTGzw6vsdRJf/k/
YONJMeNgxAB6F95BaYe9W+1ci5f44rRlftGf3cdc+U9sKx6Y2ccpGC36piVfwHmvvMJ4ag/crAzb
YdTnCEaYfS3/W4WaBIvqLlACL8nmJ9NzIStIlkiqxpQjkIZaCmWHyBLLbkDYmtdU6ZBgKoobdxXY
G6llFPRZkPa6yV972RUyI80DkpRPwWkFMSfm20enudUp5nNP3+UDFV38jgRjfArIBjh1zcF3bjOX
Ox6O1FgrPqERNZ0zvLS+p5iZ/0MrHEvnFvKpVgIaTaxOVBaM0XnXt5t/5M29VmFauiaQvxdX21iJ
Ew8U3lPOMxWYB9I8H/n8zGXdDDmD6I6exWgyKvbNoOYt2eQpUJHPaJu5ZanEN7Ch/nBvqOiXUW3K
iQnKXi5eg4HxsDCzQ4wVv9wVULQTKUQMjSSU2tkFTXmBy+NqoiA0CxCLsHgoPwqZPCaOAk9t+GQk
gpXYajoTrcMOyrKxK1WigjINNSYKdvsHU+J8UTiAUvEPvAfizPNBFvrLaJFH7h8za/ujZHb7nQJK
AS7hx4ghz9Cf6msn2mWpGdvriwf/G7gX8M5AvSK7NPRjuy7d+PLNmOr978eCKcoqtsJ/0rOl5JkP
mWjqR1S7XOudP9jp60krWEywRtSaQhYJ0AjgcSk5H1gXvyBrCOjC/oMFn7u+cvvaz1qWXSqZEaot
K5M/jNwRiTcQuBI6R70fKymZW0/5fmX6WR/GmDY4tOHQs4PhcsEsW8vEOQMURcY8/fhh+Ud2FeW0
hg1OvGh+07djLIuJk4vZAayY5O+HrSKMFTUddGC37lTOP21k63DowZeBUcPtjpfGbk1/aqbzZ828
yDOakeZEMyk2IYiQFd8DNrgIJGP7+f23kzD0rSAdaKouOjmnYlDhODp83KX+2xpdqu3BC8UdrkeB
bSdJUOIxwE67u1BoCBOnG45+x4OBGaFjBgX6566F/yeKNTYQ5F5muaWg2VpjtxaYq/4VFoDeuIo8
bAKb9EP12nlcRKTx7Vl6itAhhCuCjNUZZW4A1uhfkcTxh5RXNLtPV6/oknlCZzjCwZHWqZZh8ZBj
CgX0F9fcfqWpI+uTBSHW7MgwbpKz+6rND8KpolZxZrs9M6JKUSnRYa/HqKGFXM6/V36APecCochv
IK8qzVd4APoMIdwLDIdqs4RDLLJ6YKSMljv8R47fAH1aQLuddkIXWzGvVvW4OijvuqL+8+ru22L4
8gDmDil0nUescWV5vp03U3Vsnl3E5ZzSrmIvJMv5fPznP759ytd4Z5084hprL4posd1HZGcPBub+
KTzRMzSa0A0mQLR1vmhsyR/MbaJ85DEcpZeWcO+6UMXnRmiFQ4N+0xB+8yVgIo8liWeRoxjgpMVj
vGgOpI+ckL+ld62ENLeLaSKW7SBRae+ZnAPfSrO+8vhXq3GfAg21ZqhL9/H3nqabEH0EyNa2aYJj
pcUlUjzMQhmmd+5229cXcdAb/cPPMY7uWok5sD2ROOh3qKOUF7X5/s3ZqxBlo/QNjMoGEcwbTyuG
752SfBVCtAS9Kaxxz5nT+AnjdlUWxLSYQ+GOqFS6noVsrL1o8u2h+asiL5nMZnbtOe6j6D9bPmpE
Br8ZTyA1VIDwqg14rwGkQtS5vJL+0bAV20SStsixi9JBNv+9FuwsiqZvpUL6wWMgQdGPMKiwDgC4
pWbTKH2nQ7gTY9T5yWBeAv+FXG/vgHP/wqb5uVQjEpw0yVi7bWetPQf4f0g2yTJmtj0TqdMM8oaf
myt7VZ7JpAg1kuQdQU8lMr1F+A8TZI5cIF670cvNpsfTAMtad3Iq2Cd2OH/4P+L6iNaaWOf1tTFR
T+5iWcQoP3+VwxvgthhxPIdyzQa1y47FK3PXqe6Myayaag1fFy2bAY/1fjRcOZhAGwg399l0IGG3
b7nr832KkLBE4/Q58KiefpPQMC+9DOVQFvNr8iM4bnP1XedYzrSVX4YTMmdSo4bHfgbNp+Dsh9Hf
QEFpF4AjCWJM+iDdsAhbmlrewgZ84Zso0p0PgCj7c3ufEe2rp5MUFS4dK51S9TDWpIZS9Pk3Tcta
v7ZQBXeBIe7KcJXaOY9QKJjS3s6ANDoMhDwbMN5tN2hJ4lAPdygTfRPqmhlKKES3oYhuQ6pSgk2g
g/nNWjJPQ+oG4w32brCyICjow9TD5uktspS8xVpOu6Ru5yRS33UpRDtm8ZttezSX0AAY9baPsYMF
urx00mg4zGozvK+88jEg2HoAxO8OHK+8luagOr0Co+BNU/wFXc0qOXrx7RBdXd1P+eto8s5dsTYd
L71L4vyLVnWJC/aOfQ981ZDydKLYYQdiugHj4/D2BB9kquUQZgEDzj83uJoYN4P03TQFPp1HVcR0
V3H292N+u6TpXZRFt2vg4ySeYoDK+1LEeU0DyXGVx7IqFbRbIgZzYCRL4Xj/S/iWIUegsZ3vdWBu
l+LjVtQJwjiyx1FDwUUCmhV9MFCCTJ1BafOUtNpUiKbxq4E2sQFdw/ehyqtMvVM5BViszK5nEVKR
nINaZ4pGWHI9+lvNdruPsqXA+8CTVZzGdnBOM02tyQsTe6EqPRTpvI9U7eF9Y5a1TgF3GHOvNRwj
hycLyJtUpxFxr/EjNoeIbhML4o18wsV9jcF43RaBuWDJUOHadIwG7ge0Q3IxRiKu6C1lbaFkdKj/
7dckYoMDzWQP0JTH7q07C7A79B4eOGBkM+/0GBgiwVUPtWd+oGNGhB618t2eE2mG8dyx8Ovv7ak4
fOcWNUFbKqSCWsn4Aj9B5AhRP+ODj/4MHdw2k9ltFz77CTtZSw63wSxrtsQIPmpume/vuQQC0oQ+
DiFKN2P8HIIjIkXdilgdCqh6b9ClihVO+U3ZfxqJ+NzO4nCe5bOSuWXinOA5OhCD3Uw+tau59nDG
4Q17l71u9r51iZ6qPvjosU4v1zyvCsV5MspPjklQJc5nOPK6Q1RVa6xqp7E1F657ZQfDUohk8Y/a
IwGeagHla1OcGz3dIZ9j1AmvobEb0wZJ3vk86UxYxYKqqPVL6Z7nGfcH7QfTFZDwbDUCmAf16xK/
u/Xv4yJMdAu0kumZ196vXFRHVjZfhp8YY3x30VVCP73W32Cd4kuKPLzPuWhmDDSa3/6c1BH0vIjK
34WFnzRf7oKhXYNlnEn84/c2iNWsGwPqT2f/QYFIB78f2uYG52689pb2c9sBmUz0ew5oRvfev2cX
JLKPAt2OxELnRsE//eMfFwNzojDYTEntFsUlEJTlxcWk1qcI0QyDMITshr0zPLCWj9UOUO0lN9lK
J26sMXKxFIuLwrTGY2B7i5G6yo721ROBBSKz+d243k72kXePair1ZnRLHqdOc3uhV9UEGYUMhguN
+5fOKJ/citoNk8Rt3GEbHJBMU7MCNtxYVsM9Gk8Xl3FwoI+G08KxwrrHu56EWpnwHnSSTJNiog8Q
6z/P9mYF2+I35xBq5KpET/eoIPheu22AX5m8WSRTpLBJEsGLFdbA42hzCfnol3SarpppCy7GuL11
aFr8nMFeS71w8Uv3F4ibPperW0m3bMVjV+zaWBX9w7bUteuwmOzi4MNPsosctTErO5hvbi2VcZEN
keJ0tPytH2xEKQwljqmOgnTSfop+T74UenWKmh/i5A+me2VhbN39J7wwDmfIqgrHNiVqZoYJWRKD
LbvuCESy44htj/UARqO84zahybTaU87M2pqFhaAu8XKK3z/M1pM9ewI539bSWI5O1/FVhml0FPLf
hYob4rdS2V1g4h+fYYdlZH7Oepb68kWxiIuQd6o856NzFpn8HJYaZkue4lYpvi7cdA3yshh1qrY1
ac3uXndoZC/IUdPaWALCwPINHdeqWF6Tyb1mcVWbKwifjE5fFj7qLMq8rJPN9ZHXdg3sb5EdO6tq
fDA0b4exc7PiHhq4BveTZXjonGF1qIyHv92fRttaFdUACEfF8j64L0K4tGtO+LzgIjCRmCofy8yq
Vp72m/g7Ks6irc7/NZFZoiicVPSyjNFEV4LHka/8uyCl+2HHJjsSeTqitDavqM1w4VKiZQBXWXrH
sTB8F4i9bAjGFMtKPSc5pDdyAVCx35rE73Cy+q/b2ijYTD2NTLt8lS0AZjgBHT6a5O5FCbi4HKLB
WSECHXUEcySemiohoF2IVll0rMwNAqdz6mKzW0RYOyCg/AX/W7gfHJwY5YwdM8mFRXQT96pJADDh
tYA76Bcu0hsF6tyINGwwYiEQWkin7kVMNBeUHDdv04WLnw7CGs9yeskjhlUPKLDPjIYK8WdNznya
twjixfZqMCH9YXcbsTuHB5g2vF7yIJGf7vQcg53LKEk4ULJ655ns6AzsYAu6uwfN/jn2u0wwZCEa
1EC6qzQUokXBzxFh+SMlauy1tpakPbn2u5y7siI1VLElmO2UYowlCI0JmC1wafC4VuRG5whPS5KS
hIVhysVjdB68lvNAoKpNXdEEmeg6TAfEqGZ7c+F7KoMKdiL+3EGB93rTCDGWL19ogFIscwT6NdHi
VXrJL7C8f1jGIwvb3B474J+6qINN+0A+li3wFzV0Kj6oCH5JBnPYtCkWBjb/zhXyxgxCHdzGIidI
yU5eh4ijgrphO4uMFuLdcak5dtBmoe2m3Q0XTX8QBzOYf6lp4LsYt5LC9uGlWXriSQtMcqmSPD9K
Au6rbRpGqousSSFgFKn8hPRkA0DSBuT2PhkDMchKsDsOgGjyzVd+lMA6lPOt58XjxBL0nrQkBepq
jVJCjl5WhE355sTQRCON7ZUVqK5+IIUcmVsTDdiTTcfoYjQAroz9IPYKu9IwwTIwh1AqRqg1OLfD
9BF8ziphD4me7OW+M9yxYUjwBF07xXw03w+hzS+yJFwI/dsf937KeMRhlUOv3MRhPK6RTTOAG879
CBGJpxEiGM0yXGS3/FUHxxxXcSInUAm3mwc3W5CKFaN1y3NTs7ojp17gGJSVFaTktUVuNQLFitxl
HA8SCaVNHtd3cNlmoFL5Ghz3UD51rsLcqMCcoxE83lTxc4BwjSXowB1FX1NcRHQ5XTuhLvUDueS3
4swyirtMF8N3wQlOBQKf2x2fedc00oogYGrxAG7v2lYIBGLBiMAi0Q2uBZ0Bnf7DvDU6hATme+dE
rNCTx0XP+Bs+MPlliTdf9dsCBc36c0VvEokmDqhz
`protect end_protected
