`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
H+/W8lU1c3gF5YSUsGejG07/Zey8qovlTGgeQVnfjJVTpada6ywn425MC+Re3UpCUNxsUmiNbLou
8/X8M9GQ8w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mg9LoQnG9QqvkHfwioahLm8RAjQykinVqYqXixaVwcLE7XJjpV0iqTApecAxlmmIYSeJfFMVhkyV
j7d2rm5l0UQ6dsbhP9rDnEsgY6XlVZlGtZMkd3/Cvv/UslNjJoNmU0RqAvr5neFHC0C8tPDgw+T/
4RkuK7mUzoqQpXzDL4k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jl5v+2WGqsNEu4wjmOwIDZui4wl5yJZmI0hiE7hWVU9e+yakpqa2fNSn345h0G8Pb6syohAYCIOo
x7+74i9t/v3eAkjPR6GO1sCsQbcrQbVpcusiN7L7eqNuwB2sXoCOz9eDWNiGbNUv2an0ciVwGvGu
xlLkn6c/UrIQVaFtX+wU+cWNvnjHjLosQ2WEBf38bw48zmTdp9YhbrM3t5nZlN4c+yUK5cijl8zJ
4ptWYVDzPEfvUbDLGFg4Xq2A6LKiK8TNIs0bFG/r+i0n0xQNfFvJFq1ePsnCm9d6TpAhYFPs1lZG
vsVM6RowS6m0cu07SOVkh2aekwta/X31EFTwiA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oITI3vRvRXu6OJDbgOMeffqRV7wVJd88fj5kcwY4sjj5xRMX3G1txYMlv9PlbAVSz5OuEWgmM0hP
BKdyZR55rBQjKtrx2A2QdSYaAIJv1eyWgen8RgUhCDZ2p9Ut0r4vWq/I9sjAZo3eB+HBSNHriiDi
Bj5dD4/P5WTrDq4xTSE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZUMQHRqVyznaffBVXnjoYjN8QtkR2JFBnUSYvSE1AuNK6X2WF0CYP/e/nOkH7b0o5w2EqvuoxtY4
vkpf4QKnKqb2lSN8dCpGYR3Kq6KQJ2QCBqrcKyYwZOF3iWDv2pTUweuUXZnkfkjs56RCSBxA8kpP
A6MsHzKGPYkBIkFX2Xvvhj3MXVaGQn1n3ufoHwMb3G7muNYZnR50W7ztLwAqCRMtrzRvB0HTaudF
UEZdRZgGTSwpUd7PSpgPaLBeLiiwY1mBJuNpbBtMGywMUuEhj61rtunn3e+8g37dPw9hLeX5lKTP
bJVycgN4acRTFOCgIaOOygfErfWFAh2RaRQLew==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52864)
`protect data_block
4TeHLUc9awWZJe/iTM2TFo8BWdbAVu09E7SOZjNsDO34doZJ4ZYwYuQtmjN/hGZcFBTKzGpqAh2C
2wpW6+FMGPyDD/FqOVWYC5YJMW8A7n0TmFLZDZVUw0V0qUbtp2mP9x1uNKQq+zK4TTypoROfubiA
qTON06wAtsueOUh//GKaln9YS6hj5gKUIkm/u/Bw/KCU+Lo1l34kY/GPS5rhZy4cYVHcFSAaeykY
laB/XMU9cbvQDS7msNMvysUs5PDO77E6jiuGxK2GFSQzctX+sTCDslhUoR9IGOGnRy/V1imjtD+k
r1EiVCQ89OhXM8iipUajHgoaMRhZjpAPsub9rFoYhWfSfsPQZPysLLjeqxY2ZcvOJVfskR4PGVxR
erdQYSCVCRbgvIGTOi0GaKBYFQG4GrZflKd1sy8APH2Vzl88I6D2aYgnf9bPmB9LgJvkgBxaVN03
2sKqVbRuC8rlTikiRP1HxGDDdQB19MRvc4PdoT7TuL8OHPXCAX08xL3cuvOv7wyDduTG+V9JMZ/F
43x5y4dMvayStgPuiQmlzqFSUVR16+Q/nUjnPmnjTsmhum10YfzMPBVhNTyNuJzsl+Z92dlC27WD
SXBWUX2TytDZwB02IJyt3x/I9q05qMFNtw4EdFCszmJ7nxjtv0znUjMEWQ+M2mUcccuEJMrY2Asd
Ezgga+nNkbKP0X+RL/Td4xGlXP/IMMY3FDfRWl05KYkYEGCY4gy1B1b3d1Lao7dNgKCdU7ekotTB
MM/p2zebNL1MzBIKAo3+h39oF6Vo+3iT/4BeUOLkTYBpXan2kkypSf1CbbVa2nMfN9Xrdv5PELwN
YJDVuRHWNSaKylBdKUX5a7s+O421wFDC6erIiywDO8sTMsBYiZXZPQYq7g2noFBbsGWLpSwX+FYV
0A+HUBSAwfp8mHy2MylBm+CYYRn+1QYAjZ4giTL+47ozJRTPuQGesq/b+6qwPM493YmrxrwoTII3
xD01ePiUEg1zFGao28zEwD/4ky0ALSdIMjqYMnmV1g1vSgrQbrYsnIVRdVXAhlbmyk7Pv/sHe0EG
OOQY6ua+s5AjvNbkgE84ubR8KA3KUeQlbRF36bhy4oP4hBynUS4bIBGbqKzhdOGdyE4D+Tt6jbVi
ZSCUMnXyVodsQh52ydeZ7j9MTbsErhqihjThu8bUpTf4UfYv53G+zQw8O5HVEA7W4EqkrrusH2o4
gyw2lolq+y9jVSGD2xvZ/4mmmUkacuweFOCHvIWUyz4I9boRXFyIwSi2hao5GWaRm5D8n6rNFOLa
G1qlMtpOd/ORO7wsXmHxVrW+X9H837jmFuAMsTX6P2s7u8AkgbyLeMbVvmoGlM0WlQUxwzh66ymP
peoAo1l6cU1wD/TJKoK2ynmIU/Y+d2S6PwA1MqJDi/wSwC6+fO1kXU222pKY58iIKLl+UMUuLjnr
VGTIAjPit4ygiKt+A3xf/9H8DCq700RmbxK5nclRQV3F/+Q8f2b6b/mA+9n4YBBC5+9YCAwIMNZ5
vaVpApRRA8ig+pJchWx3AkaoMA4PiS0CSPxt1XBHSPfYCwOAskFAA3gXBaxoaCo/WRYKNdIltwzJ
qgmQiYoOh5dIZW6S0tB6GG2MfdG8hOlOPYR0LzAoT3VKIO47twk5DMWTO/qrd2oqclygG0tMOKIQ
LGIVcUn0K1prjk5BRMx8W+QjYCF62GbqEAZtiiw2PgvFYXpJnEv9Q4KlYDwBuvnt1J7nMnizuR7t
sxWrsayjaN1XHeTUrqzFjWGWaqTRnic9lseMRPJNEEvw3lDOeIF4IdlInaEY2L50O0gdR+CLUDVJ
XVacxptlAVFYUZQOULeLzwUe7RVx7gINqon/Op99rB/KuC0MtAVUcKqkqqtSa8uv9CIj1WYH0Etg
epvwu0g2lrqT/NjiyOmODweE9oErdtsofnEshrqKddahwvxyEyNG07oMGHGKY6+bBCYgkZnb1tEN
80+zL2CZLygeOvYF02mggnUO+s2NkR9x5eXxb9EKOWUkValZd47AB/XTbcoJaZ3nUWdKGUUKHR/X
JTgYvLY60rtT8tM8USRuZiPc5qcyflLjTFMneIuB81JOjxI9OHDZKuVqecB97WougnGdXyiaUlaZ
uU4PHegFC6MkIyWOiZmS917bUfcLQjeZ1jL8xf6TgWrpAtLZl5S3fVaimV0yDux1HehpbzhJWa/5
Ze8MUcgfs82tFXRUclAws8ELfI3ExiQiI1reD06uWQWE8f58/8qII42/+5ufHtQ1FBpghFWDLg/2
zlXH0YcowwnWT2IbBOcvVl5s4iMxt0Y/Vali/50zae4WtKhSgVH1y8hXzSnjwo3O6JiG87SpbWBv
yStYgAlk4NeuU7OJ/CQquEQJi7BcgbC/WabuX0R/QegTrVcKEamwQk0cN8dk0397E46MyfUU4ydJ
eBWybLGUlhJIz/hWyWkZEC6nR9MyCEjIno0uTldpGc8QqVA67zXcp1tw45QZXRtosLI6/KYHBNlm
AZPN26uEGQjU1EhihXVGYBid5H5ChmjoEgHQmkT1Dupc18k/v6IgK2x6y33YnZASWOeJ8Lv28wQJ
fYvN9NE1H6csnhwZj3OmWdCuvvqDEOGl+eLjHDutvzdne+XBgh0wLXwTUpFi9PdzRWbnFNSAfrdx
ZftrfmLqMoqLQ6Q3hcjAGy7DGJXiiVcNfvEvD7p9WE7jwizbHzSBW78IxAwGBO7CEbUXkdUxuwvY
ul07Jf42KHzw7avvtC+dQJ05rcpI1nzjQvpWXR1G45d1wXsW4ywY4thf49r7hHPkUGSrMt6fjuHh
w8B7X/0sDFWFnXpf9qIQB9j0tjho+cdxLfu1CGNQNLKIQmp49gJkx4UL1m7UlFDZJgrIaXceN1kY
hL31XMdy1U+mf77vBdJByk7leg+VvCWddGX0l0epkfmp3vwOfV9AxFYvOoDJBXbGmWdU3umzgOtD
GlzDGIrhXadnaVQV/9erlfusecP9ND6ScrsWb6J+QV5fgnOGT3xaIhl0OR9MHinQptvS4flg4lmD
TAz0d1NoHhNlRv19AArx08pawDbrUDFUkb69OpfVNvISsXqfBriPlXs1bELvmUsa6tFgnumSW8Fn
u1CabVM7z9Zd+fFicIfYTTZLNHA/i9oeb2y87QAs8ANem92ykDP/46l1wLQiq2l+JGN6PeTCwBG+
MoHnwh+7d3P4w4rYgy8GJRXm5KDMlhIa3ShuYHp/dNJWZKlzKGiYe1nQwQMQpVZGAv85/o8JCmso
2BlWHC8wy5UnbUGsKh+IeIoDPyMLMG+Ik8a/dtWRETSA2AcFYkTjPzU9vPC5+Yn/WAVmSjCXBvcn
Xn1tFCq62hHge8hsMikf3b7iGvM/9XitZZTGqOl9dxtX6goRac8ptm38VXLLRMOIg1bULNiT1JoZ
2ieKtMU4Aio4Dkv5Zrc+Wf0xz0LR56gcdhr3RjUkMXnYfAJx4VXh2AgixdObiHoA9k9TTHNcQdWU
MUYoxOkjV702LBc9+7x2K3bJeqVQ706U7c4KEqV06bS/oAWBHmv+xN8/+fAKIqt9WJoHchuS6bki
JrI4kRuUlDoL8aBIVP+peG/traIOeo1+/fZQnXFixkWd9KNhzYHDm18zmIkAo8cdxCnZIVdNJWWP
fxHBBi4Q8CKYinHbSL7E2//vWlseZZ1UKQPqSNaRzXKtXqy3j/pAhPPqHrUgHQuXzxBZrNLDOsYv
bjMp4aIxTuoPy1i2IR9KLNj03yKwYFllLQP23/kGHP4LYbQuux1Uetzn8ZR0Kc3cnznSEJCNPO8D
ZUb7LlDkoyLnoqY4dL06Dbh1+lKOejsuayfSeMlAs9suMWhQX6wDV+gZJXe0uKApSicbXCR0JZmG
QzPHDe+J9uGQMYwplFSFOTm22OIQrs9h1dGKM5HT9ajyuNyyiiqVAwAPv4ADIDRtDEaRKhYswOK4
NWxnAChWpdwXfMfLYCQrGQSeg42Qa62I7N4tC5iqRnk7jfFpXKVMdLZiwg2trmP3YFahwFR2WDht
wnR9JzE8+R78EmKv7LXdeiYmNQl62UTQDyWNq9kOw2HtIf7/FdBH0fhL4yvsp7nqP/nZnyowXdfo
ImzfpUlKQIIw3rY+d2Cl58/DM6zvM7pfQRE/RnGF9rwMvo1eenRfH3MAhauYRIwJ3Z4D5O/IJ/Ho
RdNw7OQ8WIzw1X6vZM9EPZUSjMZL4aVF5jAXYnnqfyYN9/MmPzQ0Aa5JS6pDKyd3rEJX2d/jd140
jlvM6rO2TRXLeHqW7Pc1ztfFusQDaayBJmL4rZU8Mb8rgd2GR0N+A+wgYIVVjWBPpzjLqKCXdH6A
EvsDaJ2+T5iNEsAWy5cLo9D8CHdFzPl+zeYyRsGrSC46fHOKX+wNeKJb1ELnDjZezHcljEpqEHZq
BKmmQVaagfEla0lwCSYuexzaIn6OESIv3qh0L55II1kpk5m1DRu/h7bx2MqBQxYP4Ilkykxohg7+
8df7jpObSahZ06h2z2x7m7jXy49q7KPrbFS/ZYzRzbhHcZZfH9Mqw3rTxtObT5Eo0kgua3SVlC6h
eaN75WNG6icQYOW6n/3/PaIEqoGqb9urVkooHp7JdwDp/Y53cZ8vptoOWF5Frj6AMeFuU4GdwDCm
qp/Mm63tgFmNYMRQLV7s9tbqNEs+fvo4nLzIUW2ZVPso3yrMVKTf/vVILZoZpiHKy8lkuf4QGmsy
7dHNTGY0D5/92xfgN4aFEvGgQfR4QyShGjz4G5+6KjkE0fx3tTlhSvyHU/98sCnUW71WPcAmPJbZ
7QKKLa+zLxgQbXqMZ8NksvSUtNbJLHP7vfElrGbv/bS6ZcZBVpznO7e6zl7j4ox+QioF6njdBniF
QSwTUJFyswgpARl0vr1ATCo/fLXqiwu4W5kIlSqENoBwH6F8eO75qYRC4uayPofAEY8Yv06ewZBa
she8FM7SkgiCzsnkqpPo3AO0SV1ggODq+Jnv5ipGGt3XbGvErPCrDBpNm/N9uj1azYve1u3DMzna
3+i8KQmmpqL6yrOWZMJNWR5shOFFscfVXyR3HTBSPz1gjL5CJJulJFjMAC9ghf35xr/boLgMtE1y
i+FnBO7DwJIl9DPrOeKmImjexfc06UQ+nFC29IRqJsI+5zzV4EslNheS4VpszG6bpRka8TUe01zr
Rufof04aAJT3pGpqWF5Fec9qppD4syY79pIzGY87axQbqwlVfi9OsstuUiCvO+RkJoJBv2+yrvXm
TzAo3pddGV+ED9MgktU0S3ulM2/MlCxMqvzR2SATwZJqpiFd4WX0kdMMNv/ed/4nNrm3BcnkawvU
s5kd8oqLLXK5gVutSpHps6mS/EthJoL3sF9cuSgBzJqjBEDBKIkI2+1sxMKqmgzo6f64CAgOWk9W
bMUWCDgMrgZqvqEDgdxX/jKJ75AbPyKGqekhJFj1OGECuYVjI5IhD9HXsQ4stkv4DHHBDLZgdsbr
Wo+nAyQkVlLobOWMifF9A5pL9XgUKnZ/yAaTagCSrkUQBL2OwyUUrMmyDoI79rMUxFt+NRA3/VsN
BUaCCMIJfTTBROa83cikraOry+GyqGIWkEI4U1xY6BBRIye/tgzBYgyvW2kgeJic2hbs6/V56Asm
GkSld7zlEN91xA90xmifFOZPaerxgH+lo4DQ1R2FmQ8foliQiTMtH1sZIItSHRx5IBHdDBiO1LcK
TCWS851nZ8KHPBU+wMUgzCJ3gWn4fZRUwHjwFjy+yeGyGrXn9Bx2UXKDo8zeXv6IOMaNZXRuu/TM
aq3eo7bLUN2mLdYKIHh+HR83U5xUoK0X7qsA2bGfB5AnOqONW8qLpgTj/a1nzy9uSRLbVZsm8hoQ
ZqemyKV8ZEE+eKdVBdo7TXSWobuu+fwQMqd6igCW2pwdKPskIy5CDE2FjLShSmbyErrFPr4WYrfP
hux0gXtam8jZEYMRnIxqrsdmYLMGaztPcQfKjnOA7Ot067SmR1B0sCOWm85EfN8AZqYHuAHGNdmQ
/LWNjAhgiaZ6Nnh45VYFUH8qmm66IGBNtveOpHLYH26rvvDK82AbUby7oNknNedqiIR7YzXq8KdK
Xtz2T7G0UGDs8GZLl2lr8PveMFaT3Wc0C+6PsbnRb/FlpJ6k8HbVNRmDy9Zd2Wn04DY6Bd3JUPaR
VXbI888iGhUWU6YVoaSTTDHnToNc0uenz0N+t15E4YGU1D8t/mABThYkA28pFs0EMogiqw69ZyNT
+TBlCxMf/x/0l7qAZWs0taHBV1w/8VAQwaWxu8piNi4YTgRnnC0wBirj+dYfCs+KkUaKBgCXMgRJ
VGsEwfDiN8lKbYQLlVQCLPsFlQc2lPBUIWbHq7MDjlUERCC2PjAiPATVQhhtWJVdDRrhnqHPLP4W
6/c9mW1TWDZVpu/41MWrV0wWOD6emU6rRRgIW4I4l13Z8unpqHVaHN4B4x1vFmyMkmsBKSwSLS0h
ZPfpfTQy5rTfdte7ZKD/ndDt+bhsxhG92gjH4fDr6X6gNIOQlyDGMMGXUkKFuUBoQCAXMy4q+oef
1XVKcelNPKv3hx8MNW6bGnrb25WeVs7t8DNr9hrm1T+BDWoKhg+5C58K/uleOT1teTnYWGHGtyk9
oKqUdYhNBp5ReZMzfLKd+FRxi2VCzkbNsXnoECGMnKz0sClH7nUQZtOqr022t/dxSC1+k2iyw3jd
FIpHKx2nKML9KFoNTtigXLGr1FTfhxdL5wnMg32AlhWGuMZy93c/FbW41Ll3LrLh79x3cbM84Kdi
tyScUJUhjcq9GkSYOXfHBJ4OqR9TUM6GON9TkK7zaF50kfqdJhuf2s7nuXXm2oCybhURDu7uE02e
f118S00bU6M6XEBfa/BOQWTDKqvTQzs81pnpxhq/MY/XIMteSV4SR4wkwPjF+lgrwTKUbMp0ZFsq
DCoi5zUciTQTfYMVm6Cvwp0ghx/eZ48zVS35MVt6p9Y0jMM8FidQ9TSMAPU4Pkpcc3xx56gnqeRD
hG1DbEhT3JTgDLyEnlvAOrFpZsHshoiowOyRimJzdeyB3I+aX/6K6wYAXMwuXKdGcZgGcj6KHO+x
kAUL8yuXDQisCVefZFe+NGrsxD7wyqDPJ1WYZHfYIG2rUSiVNU4uhAl1t6BdouSlF2KRe3c8/25u
XZxMJ8T54YXegksxqf+wuAifB056rBtSKUQ0nDIT8yY14DE9RXVTAQzXgUkqtqwgSztLv/Vf9KrL
q87sEcQ8Z+E1ZUXuIKfFG2uV+kGvYc72ehGKooYXltOHk40U6/d9ldc4KbKtLtC1ExyYJs2mrPGZ
RpKcPaKqlondnDkHfcdyCjfQGXcncYnAOiTU/P1y1pWqPeuXDU6egeMOwhCSnJBAlecFUncnMwiD
9fh3w+bOqG5FfXAfcyv3nATN8RC6NNPggqo5Z50rLPjRh8qHgF7C7XH4eevuzkQOFfi7fY2yfQZE
xGsSF3rArqC/B0+t29UHPvq1rXSds7IlqCpQ2WAExWGzKSPFqBCtr7+nHpq/pdNphXx2l3bUUVWv
gRbxB8E0y9ELyToRRgSWz9Pp9JAKJbDh941lhc+cb6txaTFF/OiDFkGf/blu75y2n/vcc0Rq/bIq
UaX5pQN+497202hDneLO17GmGtYJ1rZUrz7+Nc2TYHofA2gorke4jJ/JaewJc7alUp+cxySqJOGw
RL5AL6EhK3aMgl2Vnd6l+rL3PkN2or52LvvvFLjNACQAFEUNL1/2g5kdlRPvp8WJ+JB1PwkmwFjw
45SH2g7CyPPQQcFjSM1utPGV3ZMuiE4Y58T3zVK1egmTnH4VFwdSYI1hqMIC9MgvlvHicphZ4j1M
EqIfbBsjL1Of7+5E34DOA0KIgSUjMANTeU769EWNGhXi5HS+yF1itFV+iiPaPavuVADXhT3hOOIk
/Gvub/aiGAMc4PdozTJYUSYqM3dNZaoTVyc0e/QEi02uR5IsRl4LTaeyTT8kWr/UgzhCJLEdnAY8
uMTO7YRjmFkyAIZBzJi6Zpj90Py5aXX9gbvo+OnNkMyjZQlWMHBbqEicpDkr8kBDXeeMDrHrAxa5
8NpqskNz1jPYw0Umlnxz/XZD4PXXqqjV9v+PbFA0vlSS7VJFGHXyLY0wlBm6L0SqXhHvbxWJHlGL
CIjJZWBRA/tk0eh9bYPxoD6xhYeqU6c52rDAUwAc4M5cNJA6sI5nJlGSQfk5h9/pV3NWATFgHOvi
W6STHb4ouN6R2qvaQwCwIpweSy57UNBQeYa5JuqGVkeLfx/deYLG/5yY5RRHT3ixwjQ091KA/wJD
7B+KDfbmRk4c0iujkuf4rfNhsOauFBxLr7mg0q/ZlrO6Yh6/q+6H1NahnW708gMXlE2WK7kb3zCC
2jGIa0QS0QSZQEjJ5RQC5zLNYCAZgV+oXTXe9S+QwNwtyDuXqQfFOfW2fthzZAM6kz3j0MvcrMc2
5VFThhqgQ5GBaorla8CxkqIrUGFsLXKXgacUmmXqA/on8SfTKoSwFMSy4DzXToT1NNe1FGFDU8Sa
MTumRpd7+3+xFt0dGq+XVkrdI2WsrjswpaQ/9gUG8uUpIyt+kpfukhlo3SP20W9OEAgQiI4ByOO6
Kpqa8F7vD0igpjsCtxb6wrqINtJtSISU4GgEtS/rOdhEZTqJn4cO4isFcodJE1GLuWBnY0hv768X
hKk9anjBi8Uga+eiqaxFQ/aUWPnaSG0C3OvDb/24spGXFRkXzmt5llGHlI97TRmYbLk9+8SVqeWc
eWkEEZ7tW430lqqEmVeb+owPJkocl9qLOWykVsCsfPYo5xa/WBYeIJrB77hhNLGAYFugg3OT2xw6
pC5rq9pfEakd7LOXv6NLXe/7iQlQPnN7SVZUPLJ8lHq3Tt8ymrtRHEmqHEmsBmsU6ej8hFSRd5Gc
qwXtSH9qjq0zQh+Qukm5VWXu3YLohksIGEL2vvWbtkQUn97uAsUsbT2eJ4Wv52OpX2q9NBKeMlrB
/EOOv4TvPDIQ2FfuSuI+JPPpSxxRD19sigvl/uJ//MwgZNUl4Nzj0Hj8w2eOv9zcTMuUpBkG7h3D
qupQ76Tes904SNLYcuES+mbyM7lkVunQBMKWyK/n8Jq3P+BdYjgETAqEpdr3Fut+Rw5hijGgYIQM
oAiXntxmQ1wqV9p6Dfhb/6+Z31PZ2PPf3AJUyEhF0aFuJ/dEmuOw8Y9binETKAxRNP7MRazFIyq7
rgEQMAEXx0gOUGf+SiTSWvINDu7ioxNe49DBYYqTxu8R/cj60GzJGHxJIzN1tYB7HBXp2uYuipvW
reqOcsKzAVFjxr2v50d3CdKYOaDv6p7folf2mABsZuZMYuy3ABnupoEV1ynY/sJXGMXe6pp5BDN8
rBLkRbi9DVg0is96ZneJQIj31NPCaRE2tDNTRYcdR/hi7Hwne6WtU2l6exVORCCobF2nWrIG7tAj
e5cqFWu0Jf04kkwMmgzyzHXyk97CdZNG/8NLAtJFcCnJeeIwXfXtcYa7QCy7r95L/CuymZSqhOaE
PvGH+49dLQTxNsD9FdHd+vmJ9MEOgZBtssUPr240xbQTd2U0jvqczcb8y69vnNpnRN95uEAJbpkC
y540xS9A4Ez5TlPkXrTFCMGCm0MgSnBBMx1SXjEjj2weDe+E6bGL0ZG7POlISDcKJl8G1UNJqVFW
w4jcTD2C+WwwZN1fBUSHQoUJMJ94TyRoZabEPLFEh+fwvL1doBfGlP/LOXtyJMGPACW/fBRTqpgU
PRfqoydQn0J/ln4cICbyxUcmD107tsyaaDGSqdumRCTY94Ei5n6yHrJOY/Gj2RtI/MC3ewyVwChz
sja1FuL2inW64i6J72E2wq7XQgEphE3/ScKlRZKM24a2t5spL3VkGhUQEXMVTwx4kqqT55dxc0/I
dhaFt8Ev+tyM/dG+8DYmcnu+JG7Kh7f1L8r9dwJC8YNJ9azcDVSt7GAIsPkNm94qHMH+EOWsVaSH
2jXsjiV+ougH3C258iAHEbKH+3jQRL1WAuvtFOp+k7h0H6K0bdgkn/SyNzeP25Z3TzkpdATdkhjw
C/cl3EDsrj9rwRyitD2lsKupVPwrxHZcAjmRqepMT2wF8sT7nYpQ4qbrgqRt8fKJmJR+YGCXv8qg
HdcFr+WvT8hUH3VyXPSi4nVyy4L/XKPseXIvS0WHRLj0oJ5z3LeX34WvB4xvrRqklHVlOYEIS5WM
qO8yRDiuUb8i4LZZ4DKfCcLlXjUQ4qxIZ5Rvmtvjz9HULjxiDYWoOh1Wcf0O1nIFmLttdaeQ3S7l
AvbQfcqEI3lfPths3XcqhGwZth0dvMsvhRyzK9z8sTj7iurWXrSg9UXOC/Ejr0NMlT2P42mN5ma/
8bywC90Lb480h8GcuQxo+sz4N5IpQWodIXlb5m0U1lFOLfOpWq9vYNZRGYNma/sVZYgDI7IaJ2d9
4kwCGVaIqikFZTTst7urbd5OdKHAwscyIQ5jiQUS9e4lHKQZRaPRrzBvNe2JKHTgM8QLi8mJDsqk
nMw0pVnr7BDdxlyR/ONIald7nD6dd0UDbdOvOGiuNXnYQ0u3H9tGfOdsRC4T74ZgzaEw7ot6Io+J
ENYFPyWvg0abXyv/o0/8qU2FgFQJ0hZ2AoY905H8155DamgHyXg28w3STbNESMXou/LPA/fct4n0
mCiFWs9VbIirqzsJeu7FpAekihYH2H8CnVcF9UktVxtYuv98LQYIv5sYI8dnEfzBBP9G6uhShvtl
zkkg9GHIydA0cOR7ic+Y52ixsDZ6Thi/T10djd5aSsTAD/lOdsEfyAQ5OrN2r9aCkvMx9whO0vno
105n1CwKS0hJm2tGr08Gjiiavn7EbpTuhxfm6JW+dTHlM15s7r5AI6ZE/5PMBNbRL3U5kVIitq3k
sLzrqnnl9JfstE7xE1FxRg2SMP699FXvY1lx30TTtToQGfxrAF8MV54qSBH4USj8I9VnsD25hmiC
Yzhj99o5CIqM5P5nsu7rl/hIH2i9cPXMFQU0YNTz+wFu9QOSgwhv67bDRv4pgsMaK6xpATE6fATB
TGRGjKg2Kjt4Vhp1WhvEmnaOFz7SwjvkwR0L17GscswsKSwsQSSaP6Gc+MOU9SKvRwvYoRfnfslj
nejdWfwQq9F5s6f169ErieNENuN+SB1UGJMxFivIqzbldQW46ahxVw4MUW4RK4j3eSRA7MpQ0POp
LrJwdol+B7ECJGyRHJ1ftxC/u3elopIC629gsuvEYAF4P1vd7krNtOu/p4gl9ruhuLuSlIMoXhcb
OZWfbZLQxy6UrW/jQflkz8Cn9LnecBQUz0VacZgPOwJ/yr71lTrzlXVLBkv9LRvYTwKZSwkTE1vh
UlnwZNT1UWUMF2BYHLq/8rdhUyZbF1hlWzVP75OZM2VMAEKEjwegqjGtWIQI00HhuwJ6YnAdhbq4
nkgLvJ7asSk5EbLDf3AjJdk5jONxZos/rVhHNgV+3nXbTLpsn2RHAsQguM/V8VmmZSyu6nV5qsz7
0WSJs5WgwX0pVPl7wBKlbO08fyRLmGI/tW7yapCRQp+W8yHs78EA9h5PyHGWaX0uDLl+EBDry/tu
e+l4ra5gryUrcYxYnTe7Wr0BkCAq0krARYSGxQGOIl6VLP2f9aregBOTdL1v4aSVGhE8/nHZ6ZPu
+ZzMNbhCk3ze6J20XQoyofY4TuXrEaoDiDlSRbhbnIAEMwpvw6goBgM6v03ekBp91BfCAn8cUNry
rk65yBioMA1qsBfvHhNs29wkFLiSqyERGOVGAyu+sD0Tj3q8WO3kK20nYv5y6T1fXs9CbvPy686p
S0AXPbb0fYe6QfVHpEBnBFMLFhbg2yzVw7dYKALAIUCnnbirlOyQq76o8xiBqryDpiBS2qTSvBK/
dWlZhSyNGsjmb89xbXictjau1b7dWnxgXZyzBLy+ruXO0MCCpu1LLbY9XCyqtkG1L2ITB0fLoGpo
+BdjfpCVGQ6BACCAbtetpHWJ4B+o3NH/Bkg5wZnTsCsKQF8p1JSbxEXQkQ371R1NqDUQT5NdTPRF
D/Ir/hXobfXfipKh4iS6z4I+HDfp2nQHZszmQ3+NxFyzfEbmCOw2oQAVonmg/m+8O56f1uoe/kzY
iC9TDxKW+Fq4wVbjriKCJMmTZKtRM9lOrAgjl4T0QhwMwitZg4jZCMx5fEHPmZSieEgdLUZIGGIT
oOX8X1sseT2zsL0VVKIGdQuqA6nV/I5QdlHNGpkX06mAA0lAHrc5JumAm5ACaVr3fbnte4JRTCRo
zWRNgkdJwMcKZH/3QD7SAdkydoGB/tHTNfCvLt4u8AORu9sN5uHZ3vLTgufOr4MmWIWndXkwk4t6
hEsokLPvQFn9YHXDwlAWMULs7m8vchLjd9tIwy7+Qiog3SfYdmaDv3g2Li+SgVpPToVC1OeK2gH1
mg8KNyJvP32g3ExX1i2bcOn6g7/oEMT7ffv3KEzItk0l7hftW8R7UXvm17HTto47mjZp8dkwESmg
oK+7+dQzybZ5gTP5frywNxEgMRlRYJ6aWE7kliKmj6UsaBYvYyfSFy3Q7GREpG85DAL8gKDckxc9
g1DiVaws45TPjqMCJRsES4Sk0a7M+wWsUVtLcsbNWV1VWuTLH/0HlWwMYP90uc0t+/iO9lUPisPt
cAwOiYdbdc4BouTrMbaXerjyd8u3y74IY5cLLPfi38Ijep+KiuLw/iya9xJpqWU5kSlFsPujF1Yr
FnkkisfVf+UM1Z4NGjRiEdLPGdRyFGAHUsKQcBP6aobmDASHc3hB9gkrsv4m5bAM//nr3exJEVIC
qnSab+cNy9WaVAbwBhGJHU/GkpO5SSSy5d/St3I3ngALO00H+Z2sCM2az07UfibG1CYGMCccq4aL
le16TqOtFvSpJE913g0poCbsHtlK+Mozr9NIuobL/t9XTKDVRJ2SymxKYodufYzSyOGSwZe5cz8h
rfM0dPQ0AVg7ju5oKbCM5hF8bsZo+z5xgH+wmrJbkN750R2HsXBjOVhGcn50AAWG9YfUbHgJHIAO
d+Ozw3gt2dE2X1jlH1i5mKBGpcJik1yroZg+hkmZEEqZE98Mo+LENix4sk19ZqFly1Q7400kXQdR
cUSuTwSwLU3IaNcwAsH+eK18L2Gm2VoOhcBbiZpgDfxjOHT/b4fLJItYS1KIZ86a+Mul0LDeETn6
x35afgvRBDG0tZJgq3dgEnUs6CM5vuevTUsHjT1SYG0X6+Z97DpGWbqzwIL5SNLu2i7IzTa6fUHq
oqAOg6ZKbLJ/xIX/MPkqndC8LtHDC0K2/abhF28BkHdm2L0JF6t3t2Z7BnOoP1I+1GddGlO/6fJ3
V4tKZumRhOCyQPJvgU/A1Y9EYRrMLlTMz/6pmCmUOufc2I2NB68orlkBNZtqGDkorh7cOBLKpe01
f+PdLWGyQT+oY381fhgOMTCuLpdBy3p1kc6fxBG5KT/VVzSrMQ4uxd41wBKUuLvj+E+yQfBJXMHD
M+mPGQ7fgth9GtH3Yqj/FHO6AtLE265QwJ/5A8iQPt3uRCdOm5RHR+WM/eVPFdR6MRQyeKD26sBl
T9WXtv+zUYvLGEnw+3pMMCkdroV7FQGbArfPNbpChd8Oi+OECRt5hMycAa+BkUpoWqH/Zx/2lZjP
UdNEHTpU+Vz4CAyNQvrPFf0iIJ00Se/SoUpR6ixk1RhMRRYDPyNZt/PFyJCG3RJzHj4aDaqUD9FN
QR6QQ7XX/+enGrs9tjA1ZpTnpc9INOASGgaF6EKw4oIG/SAmNXrP6kKy8tBXROeI051bB/FTfsgF
tCZHCrfae0r1UOk5SxCeQkt1CfnrKuj52qiCqPcjQ7qYxOI3TRT71YzKaHm+aLvnpgepAZLPcI68
sPmOYnlREhMlm/hUW5bh6npk75ZB9Uit2qHm+2pRJDsrpLGiJSkFewqNknNqIv7+H08SlgNuiPxy
nFc+r2ke3zKM3bboe2aPhOLi4aEh9x1upJMXXY6toTrDsNBtJVRw8J+SLYzoMkkT6Pdhy4nVf45g
OF9NweZl8ZvcEqWbHyeb4xQJebAxB+xrGqKOab5fpZrcXxR/ArR1ZIQHsGOro6dmK2C+zIIv0vfa
UjbpdBEuwie5HQarxAcIsT6R3ELJgs84AzNYAWdojoJJL2TBUaCJ1Z02bt8PTqtBIXdQXmUS9IpO
b5PGFrxd5EQ7INpu0H4H8886aQmQl+P1YayAzLGoSlAwZY5unbixM9UWwcb6q785EhKDb/nSaHpq
+mk9Ce4D8CLEOoVXx7SAoqMJX+WkkMeQhfAu97UPWGoBBvxiJxvoqjZqiCDUUR4Ty6muvdEUkukI
oVwUeY8wOCaWDMSyPxLD90bb4e8petil5G8uDNGXva6N7fem0B+8q4khVF3RvbRUXYkWvF4qSinm
YTwbrvBCoroEmqVhd8YluDNUJHw1VjujJKQLYwZcd5sMOTKRES0ATSmUS47Zhh/a+vKdBBpKT+4u
fLeZLE0jQqZVD0hmL5oQ8qf4TY6pkiHiYjTo1fiq8AlYPT13Th5zkVHiQiadfM95PCPL32CzWN2/
oN/QcA/oVMR16tvpKvnWo9OFM6jh/qwqEVlDxqmlUkVM+pe9nW6XOpMPS4xSnYpHz49i42hQdbCB
neA28qTNDFbGOMdCWAzxp5kFRnwtXvpI3AuIK1DAm4wWwXikxOIvikKw85/zW0H/XBTDSP3f5KLb
vk8Gpi265LLlYN67Cd7NnNxFGszkX2Hvlmmby3pRL5REOn8sFs1XniDHMIqGD0BV8aPKWjJT/53P
p0OGmmrHB933N/1/bbxqBHhQ5AObk4ki13iSOu8vzcYz/KyDb2TmeL2MjB0cNIk+SwIzEgNQVxKD
ioqokgJ9aulonLm5MDPKwyaWhlVXm8HLegAMVzDDCCfMrLL3BFCwgRTTJc9de5Pj7bgOLx3OrPkj
weFq8rHEdwVpTsnA9FYc6bbdgF594T/+k9H2OpteysGPF+l4BKwMTmxX910guIQNT/gwlQ80ujA8
I2ruIKfaqvvIYotJx84g0xzE6O1iJyBK19ql4AgC8aVSKaMVj5EQFCok2km4LkJmX6jvV6Kg78A1
NBaW/BzFgMffSoTQMxzHbNhXKYzWrbmPaRS/3+KPUaQOJZrifqnfq1CA1lECg4cIUrbiN9WpI1oe
22PkEyQc3DJ+3/sYUzJ1fTNlLLoFXeFj5bdXDDdQHQnAAqkZWqsrxkXWmDpTB6+Fe00PRuUd7xRP
hyHjapmpeV1EseNc7nLxE6SD6w5UuU0sTQieM7Jcp0YK/mPeIAmA3hH6D+I7WK8yaG4+N8dgFR9t
mAlfqdCGomhkzuVfjmf0WsbJ5SlhjUoBRwBbdPjfxn391LJHKclq9dkBZM9A+0fk+nT3vq4eNvU3
2r6gZfXpRWDtxDG7w0lbf3uKVubQK8pu/y2NzBuUsSAUE1KPKvRqjNzc1ehpfepzOhW9RcLBu9JC
PqMBGdo+sJQucI2tsWiElmgm1XPqbDVT38mXzarWHY3GWQUm0VYWmwzf7yDDFdL6kcWjHo+hbhBv
t9s2Dd3XDUxw5lAO5zovJSjz4pZ7xQstsVOV1xvi4Hs3bAA3fmgaeXXauFlhe0uM5z4qWo3muq4E
Uy7ykPLfWzMJv9UD8Io5NeLG17hieWmdQFX0JNIp6whKIbS+gIB5i4ZDfFIAnBRObtPaCuoYDCfb
nKFGhmfInpSAo14ByUcxXLUTAYkQuQc62RJ9StT4ZRl+EdL9WWLzNTjj5DKv3krKIpEGjs1bXNG0
B8+LIihuSlBhoCzHJDu3QltQfwimhHIIad2/5JkB4mwoEzwiR/gq68MvPqvpxaqFLbOp1mWQFEhO
HIcFNihVq8fulIc+GVqtC14mI05CXST+g3nVsSvDRZuz3XMILSQGb8LDIHmSc4CJ5jBnNQlJY6sl
AwzCDzIAK5Ls+s46Z1CYtHaakWjRsqZJ4iInG9+50ip0UlEFkmyuXxpqy5PzB+NH1bwzIvSfB/d6
U0yLXNCjKZAhXJeU0kjDo2IAFZAxzpuEWsDIgDbrCJidTrKDVm9P0ZXTu5yH5KC6a9EupKPsmPNf
v1HTXXKvwCbehVcDyaJx7PRIczXLMKABL0ZwQ/rHHpnoXZNGQeZ48KP9LcQZxw4q/AyxMdwQZXQ6
HwovUYKZX5r6wg79yLvQS4LfrplnRivTJ7cQ5h7NFV4TLvYn5B24XvNFAdCMdFqIGRpXkkp1Od4F
QvNcII7TPOYssTM1RkZECfR6A7fqatkmZGJcmTSoEtdCOG6FFeoWpAwRqYAPWt9dF/wE0uVlS7rN
4jfrxG2/dUn7Ef8wSNl2POA2tvtXyyUtfMp4tGibvS7gwgYpDHRiVRakWGiXsUficNKm+XG7Ed1C
fOctRryAPxgwRihCjZrZiFqJ0OXth03rpcTm3341Wktk0S8YcIo5AZhaeNPdeQEsmDC6vvqOLvcT
vGcloEawdfLw+dW6EE5MdQDaFksFwcTBYvA1yNitEexYT70WnwUjvEL8GzLLL309BR2CrKNc2pG+
oBeV+pV4noDOcheDQdIRTbebkbg1q72yK1GTNVoRc69/dWcKlrHX9oE5Cc3Ix3KK7nWrmhdVXe6L
stONECZ3r0tLCPylBEmXgj2XqJrTBiclsakyjcHg17U2ysN47dQOrYsnpqe+way0hYmkcgucsGRR
FXMpFQmdE4YTqXWFmKnnmtrtv04fyOATdfngFgtue6edHeAtPRqPfZRMZK+Tb7NnfdpBoZeTRr0k
7KBbRm8Qd3w+LU2jnyqTuW4Mafgp1F0Go58dtbPM0ay2HkYJ36Z8yqX23tl12YVz/qLm9otNzyTH
Uy1VoccK43OygaXs1kx6jLgSFmejCxIBPmCPnuGZ+mlNhPD2BUzUICeL/iXTZl9XLNFVc8B2FzZh
ik4+R0zHMluX+Z82cdkA79emkev39XlCU/wz6wXGK9xZVDzi8eDNAv+AXpBh8I9i6Omi2rhDo8iz
2OT3cQiqaCV10Ns9N/uJgFBPZg4+4jLvRdf8o8WOC5Kb45msQPYs+7DlBwtvHiOtM+dMiiR8Lm+W
hwJhAmaBcrkQTNl2BW1JHSyAg5dH/amMVqN0H0D7qgkB/QWZpohlHWAU+F0KqbM2okZm5ydc6Mif
uaQduoaP7rhhaIwFSFsktKnzZRlwMt82luTs6SwNepMPjKsqbyV9ZKnvPdqa6m7aWOYTWlWcblOf
UAPZwLsGe4Fiw8qcSbzWVy26SLXCXEuQG4Qb0SSpmm4jfbZfivAtG4XApSYzWDhxTVUtb0D3Ytdy
ULrBmoIh88km3IsN7pDrsoxKTZbAW3xcvkjJDe2wmKzKcYFr8rLX4R4rdtvkcu6G7lIgf/1Mmik9
7uTxtKzSG/LLx6Ldx0Xrctv9gNNbxmjXz4vCBOGX8ys3/6n7UtcYZZfNVkZ8XMpSfQ2f70Pff907
uIZ7JGxD+KkQhDIrDXcl4JsS8NUR9yeKDTIMHrsaXt3P0OzWYSB4yeZfJeNs/OvkfzoEhiog5eI2
tQYFSQA0wcXdsCNyhwjHtO0bQ0LIl+Sul3W93kMP2zqQ9tSDGVlsyHXw2CEsWIxu3UkvChu45eCf
vmdxpqtixP6kGuogrylJ/4o4FIkKKBff7J+mhKRQ9oAa7Y6RMP/o6tn2LhBqfAQ1n/lIV1cAJBUG
xpQMmyz/Cj4sYqm2J/32HdmJrCEPwjE4+uYDrnsEa/yKjxsSr9j4L5sF4fUcb6s5mJ414P++GqbP
yXgWa5L7fAoQQmFFfZPrrTNZpNAT6v/G1UlZ1JatCZ4QOK9yxex45TApwwvm1jaoySy2c7BzU4D3
WKAL0iYbIerom3/3Z7KlLhz32zo6y6FRhFKCbvvqBM7q6UD/fSB39kjTNEifkL3wX0x2hI+qMDty
7eR+OUlEwxlpWZNPWgxi3XEgp5jYxYacNx16KMIn1S0aQcihKFbc3rSpbr25uOkcM9FcSuUweV0T
j0CY71ejmtKrd59+XX8WftRPrZsV5ogDVA/+gTM5ShzCnfwmZy4ZQDDmfQONvtJeXzsyuy5S0w1l
0KBUywWg0dIvS5/Lrrri8LVwZ00BNZFE9liyAHLz55gTnOGIpBrnP9u6+c5jVRlbdtVoLBTKNBhm
MSbo37HBZaMOWaLx3LV/6APrALFLaAjIR14FCPVLbKri2OASP2Tdj6AHeBY9C+q4GukfSbmIG/bX
L0LMOnSDXL6HacbysiuDRgfY4G06LtUMhPfkbrcy3pHO/MW+rTcI8RtQNqEDYbUi19oSkJMhZKjk
4xDzJ9pe2ZAxoKr8N5J2DXDoTDgPkFygOp1IWr6+OnEPM+f+00hWaM0zjdbJccFAERRt4BojiBZK
7ASy8ar1WIoNQPWJKCuR1ZTw/BOLnSRK1fbukfRqW63NRclxNBvd7N4v7uZ70rG3H6Z2nn+08TtG
Vb1YahWWLUAZXDL/v1u6FTazsKqzjFTrFuMbwH4TE57qhGxMqMJ/dlk6qhYiahiMnQvAhgcO13Lh
F0yJfGGvtrNbZNsK7G3STqNvLxzCkomWd3RP2mHTWYwAS+bFFaomr386JJrWE09ul3XuH9PSkR/e
0YJzEh3tgIfCbZNFhpx0a1E77U+snlhUaGCSPyILzx2GN9J8UgwcjdYLgwEsUIj5HeDD/XkhB5kk
JNQ2cQRHPcrurAT85iKACMGFEUSJAKNb5SMp7j7YGydTXGxI8Z67WjiYUaKgwKhS2ssQLyp8WoqQ
CGqLNfb8cmXh+QjwI9YxHAVtV8//RfjjoiWm+HU/0LLbDWowRknUiDG2zuBh/8omJT2Aghd6YXn7
w82/gXYKDGDMaicL4NI/3+zcpAuCfsqsl1NdsxmoUAZJMhXkiCZCVWoZYDhCmBaTMTn/QNQ3IC0m
qtIbnPN/05aPPsmJCU2DRngEjjC55zKTCBh6fc6E9x296AjwgYTihfmwwgu9zC2c6RbzC1a4HqwF
YvCN8GHT8VtGQb6jfw3Ito7nq3KFKtjR9KRo0jvlam3eMS+0n/sVlxXL9NOIiJ2+eStMIgKvPA4o
EJ1+iwThn1+gb5GxZVQw5tmzHL3fgmm5f/SL6+/cN+neeUq1zvHTHZ7pElcOHEIJF1chq3YeNEd2
WZeJRfJXwb/+4fF/cb+Swg7LcDhCBonCaXDp9JSsorXzhiaemZ6d9m6dK4oR4H4QpYrQ8id/oriA
UnJXZugcO7C0pJh2cuGTPfBWfLN/LnZ7zuzKJ2WgOm5Zv7UuZoAJjRATbeURmliUnk1g2hZaOq3h
yGulDnXVe9XoOre1TP41Jq+j10ZWOxz8c4kxz3eouPXfVjwPi83cWSrXQ0a+L5g808Jn2hLv2w7r
YPOc5R6Ar1/t+Qn+OkY9cJGIA4TsAQdQvWPD+Tr7Dk7FaEV1UWEad2kLtp+l3QVUfYKdo9OJlH7U
OxBc2C0BphWKoAGszUFgqQgPiE4wy9MvUEcTuLBI8jb2PQb11i+lvCAbf8tse06r1pq2FEBD5hp4
TYWm0ZNu8d/CumK1csP2RQ3nhRoC7lXpqO//z8om4WNEnoQcCjVXTg3ZxNFAdj7YsSh9jXlzUhhR
mJMpHB1+FvxgXYP8FS7xV4TPnv0exl5WAND5pAZNVNTNgnMkDiZsoQARVm7PfbK1VxcE798bInMk
u/7l0mIUDFw8G8UOx6s8WPiPS8/QUfKzlAajTRa3IX8Zcx8aeWbA0Fau+onJDCjXUQduuFUEj4lu
Lq5QokGptuGzBOepwlHT5ABafJgl4t15nyabvXQ4L96kE+8dAtVvvmMc3bOlYkAg3mzKi5QAIGYl
V+j3/6FOp9y/DTGv9SJubVjn+0cszUy0sruv0uBqAqjLnyUSmjdTFKR6dSt8g9B7jbG6cqEByHBm
NqfGZJDNdTUq7kTJeg2BYAlQ3ZcxtHJxdJyqr1YEIVP7IfXJ8KNQYd8nb6tYpUSskmENf5/5jhbv
GihR59Mv0+t31j9/liypxIWP/gaD1C7KZhnlY7+8WX405IwcPztXPoYQSzTmBSF+ni3cnxNflaYd
OXaNRYVUCEBkyIhnNLK4OLLePcHmQrBaL2VGKbR8sjkZycvFDWZl8Pnjem85cGNu/NTcPzw0Ui4e
I6Vi1oFEiqBCJZn4y7ybyKbYmQR3htj+jhqOxyYfGCQBzzmSGshm2VvP7Y72dpN+dQ6wdRT95j51
12cU9ayE5TFp3YtL7T2hmm1fHTqPSv4Fg7HMzgRBix7VL1KdMciEOYMpDgHTfBYFbI7AYg+J8YSG
764m/Dm5JcMLsM3Ra8h94LhSk3+kCfA7gYsqW1FJM2NLXkxZfZQfy8HOAh7z91MPl6IOXRjU+td8
T3CYNwOJ80uK+Tnm2P1gJB7V0L1NrEDelhfv5cjptlrP4q6TA4D0rzbKJFprV1XEgw+yUNJc4QR3
WNNyZcIL7YBJTvnx4gD7v5obZw4swbS5+5OBgrXQOnmO2He6NNgZLYCWIBgT9HRyIkchj3ojBoBR
Do+AaI3skwGb4U50KJQwBvHP/qI0RWp1IkWoWSgD1BJH30qyJ2dmhraJdSRFrONFlrGZWwlmdgfm
Tv8u13KgKoQUJB0Q3XfdaPiBTwsUGHiU5BG9MJn5HJkfFv78QJs6XYrxRJ0maFTH9/8muFCqD+Rj
9+pgIXvSWg8phUHOE0yVSTFWJWPxwBkcs4MYRs/8kjRzJCWZ18sKNXScasjvqxcoLi+5+GlorQId
vo1MBoHE1MQfcebAu06E8ijITXPXK+qP0bnapAeFjwznPvQUxm/UF5aWqQucHD3sm2f67v7LsS5y
zCmEEG9qPzvqWl+ZPXaV5B3xuV6WnVNpO0qzgaDHxOyPCp4qge6zs5qj/70eqRzYOFEs/4/GHt5e
XY+/AGxV+DaV0MtQcNEobDFjW7scKIDl9PTrb9x2hLIAr7zT91fhdMhG7zHEuhxvAnWNP6NKz5rl
q+Td+3bLYYsAz/f+l8Pbp2M8F/USslwFPH2sPgZeK0ikd+iOd80v1rS1XUPA7fmIczXr9ZVpG87L
sAikIv6QQHaQjCbAMAhlWWrlxyoKHBEfoWWSljzyiufrzTGiOejHQHO2dDy4bV1RWg9n+qsbEpIE
fn1oGLflXcBL7CCs5LoFS+Wi+Ed/KjWDV+sIOkpnOD/5LvAHvWGVyqW9imBVPMdL77uR9CXI1B/2
RRcOGRDyPRigWNBUj3e+8QUSXascCpVLTFv8owfLoRWLA8yA/Fl+9LEcpAIybMxJB1w4YwomxtVO
gxXmHfUr44U+uPpQAwyXYmhRM7hV/s6j3nZG8lQ1jL7st+EfdHVMvkrJ80U6hxdlb9l6l8XUOW7K
WBF21GK5/47RI/uF+U7Ru6jQgIXy11n6T7/Dw1nGCETRvmdPQRrH1jms3Asv7kmf6NWdIJnf//LD
nRb9RiPLUQF9r0gTx7blS7PnCO/v07L//sDvMfy6sH96gjjG2AjFOvEWhBOFbY1SMSqYXG9Ok+vv
o79aQef9sahqR4EXj7GZTRn9vu33XS0Z4C9Yookfo2FbhyY924SNpBG9bnzPHJCewhrEm1Twnek9
PFsdA3PrLTckiB14KbV3C1w2MmYxfCVjBq3oDPzAVJ0JNdxUXwW6W5VxxO0ryeIBCPp2F7ASVFkd
ZzJ6qg6Sc8OBfh87iUrlGJK3WBYjvwIGnJlWQzxRovub110K6CGYiAhbf2E7dwy0NDrhxpOt2F70
X9QCaXmbPeKvRzXCx+MtNoX/75Ocp06OTqnqDH+ai8Ss8gRQLIVYN1CW4+swsE6WFvN3AvWU7jrw
ROZ+eZm9QRlDVsJFRI66ybjAWpS+U17rrPTXcQIPn7Se85ONq4dc5v7D9rDgWv5opIozz90L/UiO
xpUOa5tyZGMGCDC78rTEtepAFXMC0oKZNu09LU7RMMzevp1YUDBIoTguDMhuXyFNtgjnsov/+eS4
tk8v1z8QRncUnWFusNxpdlR2GIdxBirwTC3KD030xF1/oBX4ZWhX8AThHDBbFd1vCUgh8qkkTX4v
YL7UJSNOwSP7AUcgjXoBBH6f2VuCwqUN0G4A+zUQf4tyv6iECI8WhVRuSKv+hJHiypf/a0VtVjGV
FxnqT5p8laDkU9vvqH7mn+b5C4t2IKJp5amTaP3bpBuo9m6M91jy2LbmGZrMLaFNdR4ldMVYdqUZ
XrN+0jzqwufa6tW2M5XAv8XkhbqY08dfIPgVpq0aUJZUUr1nEN0pDtFM8aFQtb0MbjluaOgH3yKd
ZBG4UvtWMeWk403qIrw8MEcP8KOXmyozsAIuwk5IncgUDtUMZmWeKmT8Rd/Pq2iV7XMvndDuNxqD
eCVdbdVRjA9VQQFDA9MTPqX4EWSJsXBU8oKpd5cfBhlZLGcNxA+JdAHJOSuGrDcJbyQSGxA2WSkq
atPChOZHbwSYLtrrFqNaaqYX0I+//TOWKPutVgFmUA9RneJEmeHnlYbjEbTF94rTVSGNFCQLktnd
fNFhFTtnMV8uhZdCfAL2FwbvSpzIIZ4ndx+B64cJm0oMt+XtAhLmQ9TKzZdGkRhqbP6AItm004kC
QEm3YgNvceAy2Yzx32XkoPR6RGsjSN43BO9mipJfq4/dHsnVsTVs6XOtGM77OWWqzi8EHd5IOfc+
npSOJ0RGpT/Dx+HC7ogG1SzsqRUWXDN+ue9a4B9KiLD3C6ggvRfMLA62HDM8iZdkKu8/z5zhspfL
sj2LXz86IpgpMk43RIkblwSomOdCMmA6rcZUuyiPN68faPRRWWl2JU6P35S7awgyTyW3oj+Pgzpv
G2UwYlCpavwH32YIuRwnbnxn5Ul9NWUm5nFfhT7Lr9dSmahlAE2GAgYpZ8S3g7HZTPQpTWoLzAMH
bOrTj43lsRBMfNewI5e4kymr7HPqiyJlsmSBYz7Ccu7PLA0dQqzth3XPKbDar8DLrFIgwLYotHfR
tzHsdBW2B7pEIxBp0xwfV5Gf6soKTI9Lmf8xdWJzhGO1jvWEjVGJdUEX0fliataX/L0E67plYi95
EM95/IUQHcC3kGzyI76jT36tSOkGK+la0K8OENDj0sgR7h3hLrTmqhf5V5i9wcH0nH0naISOA8Qa
Pw52Q+cp5oYxf0bb4394/6ylTit+JjIzwrwZ5Qwo1L8Q3TUbaGX3AiwD5PNlnLKjmkJNTqFMGT/m
UYb4IGLEx2reOZKBdiuf/Q+F/XIbKM2ZpqwpR9+g46D0EJ3s4FDK1CoPmkhoH5K0drm9HpBnWBPJ
1yOynIUPX8SFRyptA7Mau1U1W3a/iZxKSEuVGRmY0m/QNCd7WJ2dzaIf7LWOa/QQmpL9Re4IUg4F
LrM/hWn8bGbrk8rZpoRgfByoQw6qWCv8vDFuRVs7uhXXpfZpiYkPKNEfcN0HlmeEEIPAFSS+Svu7
d85tpG/hol6yKRBfk9sxHbSOjgTaXLZr06ufuG6Gllm8G1VLm60twr/uoDaEsPBIYkhLbRkX6Z6N
mwNppKN+rsMNKw/DmhUBKUqqfQumat5HWjadvZ+JTGDi1w25JfgFJrXAl8hFU2dQMlkO/lXoiWCZ
utiMOd0Alm+zBB6ZWB0IXeigYIB2atxWwLxHgGmNnW+FgcDP5rMIIL30hBFwbFjnTpLPZndE8l0q
J9XVCaOxn2EJzEBd9edfNfQuVfaMgJQ9HrInVYXmu4p1zCuOnwPZyvqbmSsyI6Rm5oVYmFBTwfGU
4YwsKJ2Ptp4Uhy8pJJ4UHwkQiLD51+ovaQUgZnuXLFtXMOQ93LCtckKjnlvVrEeIIJo5vFRAH2BJ
f+z8oYrd63flibxRd4IWuXjSGs96jRQ2o97nyHa9mOloxbqNj0gBY9PsjT1fNB2rGUcU3nRRoDCf
O0YAQGaZUPxpWbkLeCU2mV93A98TXoMXWS/U9KOK7ZwfSkntZgasuTlY53hPcHiIRPRImNQ3xbU8
GSF/YdMxOOKGq9LI03yAH/VP8Xkibj2klWlznNTomeU0xma84cL4mycQylotcEUEV3hcobgpcm61
lE22+7qw00TNeWL0EhOI7FfYGr8/7uR66iCzh8dZzLAQ1qqMSESvZlBbZj0tcNOPCHP0d2qnt6hx
E/vRHaCHzbIEFHBjveVD6eGyfpl2gF83OhwzD5l41ohl0vW6+GVWNWDMnCGpBIeihuUKWzpF1SIt
yoQuiv/NK3/3box6c2U4ZCkw6M/AhXe/B6+Blcqgpv1ES6gXdYfJTH+HA+4PcLxS8IgmB6ro+vvN
sMJsvh+vfHYrI4i+9xZSJGbbtLwnpGDIusf+0Alk3DcnSZWciaTlDA4TcjPE6GkuuE369paBfRCe
oG/7JuBrpaQ3BppoMvSyBlS+NfSUu5CZi4GMgEhW31gLKsnxIpOppjgWxb/TLlEsKT7UI8v8eSvB
5WC32N79OSAcCXWTZfrM1mH39NGgzzVBsSa0xXODZIWk4BWQvaXCxhtluE63uuWuUZwUxC576/Tb
jinSgRhshn5k5RS4EBgFTjM09/4aP6nT8/SzB79DKpSDZezgw+zpWANLsrFRAKT40maH88kJF7XG
qODOCv0yZD/RsTZb2R0d+yxHzYN+aVSeS0ZsrAjAYHKqSJf8LwL4FidWOrqjP9ONFVY2h4lhziae
PRsBOSQBDdS4Hk72OfgcyRs+7HkFfYv9WwD6o4j8ulaliLlALehoEIcsq8GheFg5KV7gZNO1TIrB
Rp4TnOtcKCcifZac5HAhE5UUOD6md6W3E0roBydE7/Fb393oBzNl4X0dm78KXHOwjcJ2z+RP1fIs
V7nZXtale0dzxfGAwLsFIOrXdHzeiD044ZtVHpK0NtGmVKPQSlVcYAhp3RQwnaLvGhON0IPO1ASx
03kVYvq4AM5QtfepOTuXHOasZCOx9IB3BDKFvadWHcov2KsBwn9tGIinYFyIjzoPo9W8rMO+1c6k
0JvQvdI7DDK1yeLf3SA79x7kVSlW6OOQkwjMrH86PsyTsvKzpgG/gN5oIstApedwD2VGVMFZogr9
rt6uyfSHMSxjfbOcgH9zUw6ar1N9N7mgSguZvYZjc1XQa5bXKDAXPfh3V17SqvK1BoIsNi7YzjBP
kQnmPczDg5ESpagr9jRjsiGQ5+CzZTqVn2Hb/iQRhtdliJPjML42qjhmkGmZzb34qTpTrhS9lqtN
SvoqVAvYqlijrtLnVLk/RR6IqgGzqRgQ2c4Sr131aIc20sbVHQMrXAGxhD9ZsVu10ajgoDsJiUc4
YonMn7x0CZcGPVScmZA9ZUxNx1faXBtQxR4kS8kLdJab2b8OuXVF6uRyXs6q5DKDjocb8Bo8f3JX
ujpPTiIdyqflBLL8+UsGmwBZ8m4ArafL82z5MX6zg1rlgoc4xFAkcQkKIIS/dTm4y+OVclqetDa0
9nnZAyZ4zC1MM9FlYn8UFHOsHvo4QgToSz/mb8UwWXV83FsarwYOrhBjehHwO32a6DOPGy9ncCxM
WQCJeaJdq4P5EfoVMzbbkw0QuCmRXe3Zs3fAnaQoc7znqTRLtpvAK9DxaxfFjk/aZVHmbea/Zgzy
3EoN306SsQuyY1et3sJQbl2gdHKalyObK3CpzYTPatJsicjNh3UC0u+el9thmT5skmQDyiiQ2NwK
1iUFIrTeJj3aSlLxGXMSsM7U41tJlUEPRy8VCcu+zJTwDTiXhLvsc4u6Utu5kZ5rJF2CUbbvtuqK
5jUx4Y62qL9VMB0Ym3czO2W0cgfsQz4T+WdvlB8tnUeVhV+cS27OkfGv2J2PRc73ySGSeMOGR0O3
7snZXyAUFP6ivCmpPoSf6kSM6MyP73D5J7Kzl97CkrN2G8uY/fJ03z5YI9bCSGD15D2f/THXKcgo
l7MYInXuKyNRJ38DFIUlkW6WdA7ZQy/iVVU49UU5JF4fDmObkqU00CSCjj1O26s4+5TlIXrC60Jx
m2JUmIUDho2q5nDu5riTKKgmfDijyWdUdgDFoyoxCXbNdanUL/rPynNYZM2wE5kX1i6B6eZddO+9
SX3OagtbIjslnNUTQklJIA+ze+DtxnRoTpTADP0RhNqnybYPG3PmfIlQLG2tqxt4wwSnBL/ZD9em
JnSWGReR5cR92ajYo9GN8oCEUG+Utqny8CTmK3pq3WKi/3j9Dk14ow/w6nX67Q5Tzk8DwZvdGJDk
UX+LJaSqWGzANqDhXZTNEcOnpGzorj+3lPxUNc/wfYoWf9TbGZKJtbtttLF7UYHOQFXY3jxqXtr4
je/TM15DnDRnYcbFSvQvAAxLIEK8tISKKwoM8Mg84P0LL3pJYYZbIIu/QE0yKzu2HG9vA38Ilql1
+GVHAVkomlU7khREM8yJXRHktVilmBssHRubj++wze44Q39k5yjNZbUucbjsDv5ww9REIMVeXbA3
1T77yfTOpmXFytrMU9LZGWBPM89awQ1rz7CfWGy4x/ja06CR55jQnAtCD1hy2O9cZaqjtphm+mYv
NevRBsFzJHrN10YWX9aZ05F7PnK7b3kpkwihbuGCO+wpy7XEwQmsMBzmy7MnYw/tVqie8qWNXvCd
87G9L11/HlGF1fvWuCTvviAjm3WjfSapWCLNgQtg9O1zPf2WKTwPDbzxYDPWLd9dihRom+zVlylC
0firB6ooh1I9eNykoXX6tfbFufkSJaXQdh8W6BQBH0njUxqMDLGEhmfnN6G3zL3s3U5V7wJhRLa6
jLpZDckq9OpDViGVj8CE8AyHJUAk0E21QYFXq9x3LH2F9ZHX6J0CnzijwrmlipKLm2etljB7xHH/
/PcK5YqkGfIVf04BWNYgXdjC3MKbNJpenmZkE1Y73wby4zP3R88Os2GTo9JrU2Iky+CSqxBQW3Gx
VWVMqIhDfiwb7WergWaevvFwWYUs4U+6E84Nl1BxIvT09i5ehCyvrdXu6nRXTuMne84AZ38ZLHDp
s4uvMGQ8qSo1KTWmk9+Tqb3qokFIN7v0Xwc+IBEMfGa74mvMqg9UZRo2lwdIvGNKzroEV5Myl96+
9qHRg+jZERSSxcGJvQrpsxxm0gBCx2wp16VuJlZLa9sINzrgBIPWFP0x3+GJHdDGKQk2ORQXARp4
1eE2JBw5dj5T7z2tOfpw15g/zqZCPU6GV4XHOC0Gz0ZFYayBHA9SoC1NgzOUsNSdAZMmRx0IB5I+
K9EfHTVwqauFrwmgXiexyI/eKbUYeO8UwONHAubmCJmGnUpaRMnud27+A3upUd/7HcOr7TrzcxWW
2UBMEPaqjSlUe22nGdLt9Q6T3IyuGZveRgw8KuVt5cLdj/Kx2HgQ+J0pHvo3fvclgjw1WhVHcTCr
+Q6zk3taTE6cSmx+dhIVQWikCx4ZcmMqcD+hTu9qD+eAiU6f9S0EsDnwzhgBIUs4cd0SBiPijo0w
VSdBqGt8nFBi+t4hrXOfIcMonbIuIiw/51e17EwsNIpr1qca66s1nMuUYkwpuOqcVahcsDnOJgYK
+hkUrOJvq/Nac7z+HsV6OVKQuT2Cmk4rYYcy3WhocOUGmXXiRNh1UnI/ldJp3KZ6YV5Xk8d+WnYx
k67ihPJyqVKZV9aTAPgk4JCqfCUS0HLa4nTBE9RcgFJRN6vJNnF1tNR7GYc9na5cfL2XPms5I19l
gyIc9gKflP9H0g7fzEQYN7XRCIcRkOy8wtMOMhshxrtfS7Je0th04TYm0ArQIixLjXbKs4GCZ+mX
WFXsVEd+L/05B9zB9NUoKcpy57PIhYktAqWgxydV+n97rrLWERMIIfIKBv7fjjgL7EN7sMkxOkZJ
eVP/B/50qIj3+i69DezqGZFurBqoXXc7+b52Wjo+vuUBh/vxpzCRT3D5up7Aaaf9XXSLCCk8i4xW
3QgJDLoTsM98jXvxw3ODGwzUiqaiPt4b5tzj2NuvIxIRwdoOoKt5oXH3gvcSy6zRCSuasl2/mtER
yZz/765T/yIkDermCuqrJV8CrO/GCYYjhfC+G73PD+nBf/rDR4HtRzDaW5MHmgWqdU50MHcvjU5n
HFkSAwbKb/+4FKvKvppCNfkcptnKOaImiUcn2+NQdteljqxXgBTFWrHuhMMHtKzy/Z7UAkHiIjLD
VNGlIvm+ZAgXkw4u6ydoxgWxwxOnBxiOBDiHjWRzrRaUVySppBIM555motjyRA/eZBBHnB3UgZ1h
uUBwDIqHMG+MiOdwWm+zPczT7u3aYemuQM3MjP7uFMwWdYB0ELOG3CF8FHYwagTne9b9FEvGgbBn
rM7hvb5DJjue8i6162xgNi6nckvCC0TPYW4VGTzj8gel7bv8T+ZkNVG94FWW3hJ3oHCaUav2RLu6
wxSuPPy8NhhdXjBCGkk6c8bRXJPu9A/aO84bAYZ3JiQEK7QcRnkcycnPPx1YwpGMGt135uMZ3/C8
Zm+ZL3RoVATwMhcOHYBkf7gW4b5vEQsSSBNbgBd18TLMe3cBNCCLzb3XEOpyALQm5YUEsUciXMwz
sGAyPRQRMc5ZLY0DL3F+NrB9XAttO9zjnXtqfDQGhK0f9ZoUFgPVTqlMVl6uN6vJWuvQ9Z/JaWjC
iY7cg38Ec9Ro+cLnstMIMUvyUyBvUMEwtCkH3YTvdgPwnMS5dG3IjKBnU11czrJnVrdE5ga+Yy1K
guhhObnJMeGBOVmmTlplPg2GgFJMHuC/2aY3f5mVgkWT6ZAvTeo+78gJwUAeHDWLN7FnoXsLEV58
prVTZ9s48V25mzGcNs3NoeZoorr9Xyw02pLzIGXG6NH0ol22nQy+9vJmI3PX+JL743ZlND/uoJIQ
QQqYHRxSjImevYMeEcbn67aVwnvMlVIv4rfe2Cy4xy9hQM+d312t94JewzVY8h5pf66hAdugl8hG
qu9fb14+/nKvPm/l3vk1QZjcBu2IC5Lp6xxd4JaPioO6U79YJ7fAZ7xe0kjEHTR1LaVX1cZJ8xBk
ixLHu4AOutW6E3vhZEEnSfYoK2L38kaR9IQBMnXFrg5h5AdfUIYU5lL5mk7EpEFrBoupbRz3+6Pd
R3H0z5inCO0dftsd+u2VRtzwi7Xr0DEkbPXUyYw66yLCI23fyqNkswYgF3wCQ6k2a47TS9TihWDG
JASWc9c6/exwF1HPcYg/ugBawNuFDapVMLp46W0Lr5x7/D2ImHCaxXxoJJav0oNyrc+OTdeuTtlF
PivG/H+FvH/BmkACFAVhJ56qdqe4RzWo1XmW6atWPsaes9rgyQIlJjwHOa/V3n9s4Xe7mOznl/e+
Wq9OUJwCerxnieYRTAgshiUIiilGwY+9fXuDeCIT1GeDeEzkRrZukppW69CxA575wIAcnYCUAHpQ
fsFu5keR24vofcjY5UZ7yZqhh+ED9K+6RH+08xlOvt62791Gf5RAG+XCx48QS0A9bpN2JoXi8YlJ
ROshh2Qdwmq/UV4yQE9RQZPE+04tB2ViO4uamarropR4Dg8aScHMKdtk2LyxGUl7GOKXC1esD/st
Z+WJHdHpAn1GVRhfSwIWHVvpXRHUjEZRSduVkttj+MGPa4YcniougsZ3zNFO9Obrf+lTM6Ad7Nn0
udMvGDNSlPha85GYp9drrrgibSMqm5SBlue6YSk7IxZnPKjbz86vscn6fl/ClW6gpwqJi0zrzWgw
ctnBip0kaCrrX3z+KrlcAnBwKURo77R+kzixP2KYZPzY9FLEw2erCd+ZRkVsjWskfJWFFftsu9Q7
CdZ3dPCTGwPppcRlTm32yz1UuADofp3ctdz1z52vb9EKZIS9jYdM6Rfh9MV4/uBCDEKOE3BglMes
KC8JuBtrNKd3Cpzqk9j2/f7dV2g8y9HONBjF7cETgcF5MyuqPGns1e3QXyMT4yXaCNodJugxuXYD
DqTvatcEbcxzHJDYtO4uo/gT1FkwFprfpuHkVzIfB3+K8+frzvtqUzTjfdAUxZ0uKfldiMl7n3Mh
GBiHH0iXUySeuNtbnO5/jvvQ27FhW/RUhKe4wU/rKtVeFdYqfZ0lbT9CeEvF/WMYj/FIzwNExy4b
QVctVduSqDcjSwRbC2MsTXX1cuRvIZWlGWbHZD/j4cTuexk46TK+Z2A6PFZJcDJ3ks/IP0Si5JhB
DOSqX6X6ttpf7ydnLK08FU4nLfpYK05WYDO3Vam1EzdUV26yTWdaFKk8I0uTjKKPz0sgjtfyEIzk
+X91vtxRQYFzbu/+CKWUFmi1BWNQfFMF7Jgin1cSHI74pSn9NRBavyug696ufJ4NwyDCg1CJ90R/
imocIZ6EjcddLOXFKktvCwcPt5QaH+IxG65Z7vkJLV1qQ6qRhbgZmluaaqn1nET1t07Mjdf69XX/
ndLds6IsaZrdlcQ7lS7LT6VnVPCucOhlgqHRcrXj4GHi7NiCUw69zCI1oaIn8UEqc0f15FNqzs8o
5+UL1+dzg2vfrXDh6YoOw0cm1IH87+wi4TX8iPoQweHwBipGCEZ/PsSLQExR5njgfBg7/n+kEpJY
UOiUFSc3wXhgBFaNGD39KYD5TxmCyyU3KGO+y6+jbHT33cg76nLUDz53mLyFTPOB7a/q7T3tmy+v
GYsDH7g/T1+NVrDqnJfexZOT7xoz3l36Va+TD7rxNGjDwgSiSuDegIgGz2l+USfL9W8eKu0B6duU
p8vGCDNNv/AqggsEjkAS7uwXIoro+d2WsPzV8sbc/qWpK5s9TNo3oryTH3j7r32u5dw8Q0joCkP3
/xvv9O45O4+RfaOv4aMcuN3mzMIQ17yNDktyh/qLfzOBgFrmtvJFrGxqmQRTnlGv8RM6TYj47kp8
iRozT1guwIC6iHTsyFMAheivmwNPcC7CdECOW3zJ9p4SLSHVq8x/MnhUu5r9RFM62vjKZasob2i8
B0KlZl6gJMKhCoaPhG55XkYQwHtsm9JEEqWYy3S80uD0lNiQSixLCBKNEeECVDS/DZUhi6AbqTZL
guMsCpJv/+6kKd64/noV32aylJRGXHflEl9MY75Mya/wxIb5kKAr7ftkuK3NuoVoIYWy18eWWjfZ
k66bJzrmv4zibiBe0H+g2dPszZZ5dGenFOpH8GsVZtQ46wfdsRytVd7BUmEERpOy/sQVXdzyaSu+
7ufbhDr/ZW0ENSWU/zvpgIGov4Rf0d+b+7D31qE6IzkgR5DG4nlUILI3qMm9iQCmf40jF9Wtyxln
jcAXkcvasT1xjqvKyE57x/A8ff1GpPchAQTx4fQ7l6h3VC29rBIACn+qXTgYrLcy/3Y2JTc4bJ98
BP/pV/kynIcqc0i08x+8lOh2QQJo1HLL7jIEk36kbKw39oHGe7GPF1aqHIVJMJnsNjYvmUnem3pj
eBw6hjxO92rr+tQuXlHb4f0rzJRBlLFnwDk4o7tBwuLMbF2g/XUrtspNEMoFqSviasDPRuwDtFxI
pzjmRI2Jj2C+Mi9G1SKlJp7PsmBp3PN+ZeLHmeaaFjKoSEp8GNpNNEvs7nSpLfZKrODQ+Kpzv9fa
4G18WGHy1dgsgM5BeImlf++2AVB0xQazRHl3ZkaF6JmOd31k55iD+4DgUk3LKLyURgmZQjQCbaC1
6SzBe+00/bAsjskLEMp4NgcEPfoJ1zRJh+OKMST0Ijd1/wFBaJSqNw1DBgPpAAH5KgctzSsW47iG
iMJtn0OYGZtt1HdnKuGjkWwABillTbrwfg+tueQDDS0/TXcM6Gy4L3UpLpV4h+Q1860350xHxbI8
9vgdNq8oEDs/5gF17sz4Aa/h1pRPeeMMCJTtXNHpG9p2wI/F18M+i/dzAn4no1DBwjsOjH+H7SiO
K/M5muh40IdvL6sOtmdAr4jKRQN0ijzJX2vRtFE6vlW7LGgo/ivmO1rxNvsmA67wzRSdydF8uFnp
7z66yOO702DQjU29Gzcj/MzNAtFuE27M0u0Z5kIJt6UbWVUI3/ARKmI41tt7qhClFqGL4Euz9AYY
hZl7zKp0x68j5IOkk7d29h1UF+/e+DmJ/GLHTJWo+JW2IA3tvDjlstKB0topqtuB9nPCbCLsFO5L
Qj7X4auMwv+UoGnau0ELnEsKYiEHNP8OUlXw53Jv4Z2N5cy1vhJQ7Ot58ACPkCZy+i92ixIk2YFE
TqwFG3M2HgHr9j2hbAglbFrvWzwTkJ6DF5+BkUSo5H+avrb5wN3WLeHQE46Nlj/zjRglKVBCyalh
dFu/W+1mjbRHUQMt+J3eD6gNBdN5roknScGuJgMsOLpilYO6AzvXp/HXm54/axrGT2ejExOTRroD
u3j9UPnt3ou44XXcwuU7n1q8hjLcK/US+kCoxjt46hIKbuHFdPcKKrOMmaNvfaufEwldoXpg/8du
sikSxz5y1E6x+nEnnvtOZWxr33UQVuqPXjJ6ZH5SzAzj6bvVXe1pRvVhBezkpWlRzomrE0KVDwkc
TsRQSF0nVKxy3GPihV3/jtQMVPuM0kHiebyUTcFErtPn5CbAFqdbrAEbqgDF1egDy3RjZEN1S4jA
GCcpF4mqNoIpxUqiD9RuiOrF5QdlNOp40qCjK7r0NAX0bopAmRamAcmDP6AMXl5+YDJQe3JRjTzw
+NmfnOXa7z3haBrptgXFirUBpKLJ6baRQDaBE9uoyHHNq1o0Ocg+i211LZ+ghOooWcTKOIcbcnRY
pwfwc+qBkWj+P+xtmBAX8AJaCUSzip7tPDt7BsEyaiUn2hkS2mzZElycdEhY18DE4qwuzrRYwpU7
saljUMxfMRfy1NpCRJm6Tv1sbBK6PrvsbL+W3znijziJECm8OMEXlnktYa7Iv40acbgSVxbPNXc8
3EfGYfjn6ObTPEYMiqZdTMnJ0vDyPojg05Up43fWh9DU1hgL84K7TpxCqZsL9PpHUh6NXcqe1aD3
k72hw+zpkWtaGIPIg3VY8AX8wSIug11nCDqQ+1gFfI2PX6e8m+uzNPdWo05d2pyXwm9ffIU5tQFT
JWOgLXQ6QB2k9FJNibkrLWkgkhBQMjC26ascfhpAwGd3af+2DRYQhg7XOy2F2eaSZsPQArzGPmKe
LO9f5dduiwcL4fdWP9NsnpriaINNbT1txuYM49hysC0CNpd8aXK5obGHk2x2xfhWr6vrUJBCKH6r
VU+yQks3BbNFnAi0zehpOxJw9BDqmxZsLaepRYq3rWpCYYazlQTL6u9PR+OI8RQpYEm8Rv495K6p
qWl/i2W5dW8szkq+nuFCPjAyqBuQLWcE4cNS4h/l4J+6pp5Y9bUpM85cSjU4LVAdxhxntQ0NxqUN
LxdfozQq/+HJqG4zsPVgVltvDmmSw+8wguxkjnnBLSmkKdP0VcZaX13zHmOo106t7xb3aSiOAwzN
aFJotmBlqxTGaQymeLO+evgE5GWLJ5ScMIXWBqLVS3/E+VmyxFAEuN5Aum4HmJJd3rumf2mZVLcN
7FeYRiQduGNDQ1uJSUL0AMzXFnrmUSZ6kXgIWmFat8xIDx1ofLPTsbvCEMYlfc/sRFIHn+mgThS3
9rTfzP1W8KrIUFf83375/0mIGJRLU62BQRnGVMmFPRHpXPXgTEhbzrps2XLF/tALrxKp6EisFeUt
lpD2zH6n/hhOKYHKN0X+TrRgRMz+FF92FHpU9pPLNTpOTkeDmvpffZD8ryByDY/XjklWonKZXRA5
q6+8UlkU19WBqq2NT0KuEKdwZZDlb8+RYnlE3gZYMBjGErZ/3wDjtuQn8jCBer29bvs9GyLRgBse
cePkfemrzJmdL5CLcpLfP1EU7H08ymIJoZ3fbItbMrwSW95e9ukdB+ta1Xx813H1b+znNVk+4Rzj
o5sHCJkblH6yvrFgqV2luZTcmdYftXMyQwIRoBmm/vDtZ2kDg8VK2imysk8SMEZSKMGAF2nVult2
5kEFNtRcu8IGb1NEiUQBVHO6ouNnzs/Y6meGrCnq6pwAsLFVDXqL9z+NTbbZzhwFa5b+haFEQDKk
C+MLZnzEwnEs3U5fQJ5QHRQ6VaEX6+3DzRrjVduorpYCQG6wRcoSOzb4zcQsFaxCOtNUELzC8uGm
e7fIwdr1rNEV38j7WVS6RAGGOptaZIdH25miIbFBLMpgwOO7CNl+1TdtAFApcrdBjIpbF8Ht61v8
2b3SBtjLY6HMXG6xEURZmHLznbVm6DA/inWkt8zIaxZhf8X9CU8cJArt9ilpWghfw/QQzLyTvhfN
PZint1BuMQOMlHf/7OHxKIUbh3O0rEgFcnEeqn2a0nEIdPNSf91nbxZ6sTv1yj1F4iqFQom+IAPU
cwfYOpl9dLj9BOiEwCBL1U0cstn0CxyRN0uhrCA49gTyYby1t7akYIL2uD3uy/zV1vWEkCppWr9C
j3S6oo9M+TKEvc2GjfCjceeesrPEh73WQyXsZgExcEUppBwDQJcoZ1iumzmWRrAuPaf5PtUOajXb
StmBZ1w1ch1zjKSJT/SgmzmbiqPCUtlmdoKZnijGH3Q5g86OObV6W4V/NRBHgObWbVcdjCofRmBc
S+kHlwGT3HzCuYfdgwfX52CMh6pD0/0G+q8zzfCw345+GmIOgif1Ip77zD3uuts4PW6rhu+z9PEc
bdZgnG5a2gx7aUR5oqfRnCEfEVwcczcaVh0Vju+/+SCXZAd/uW4aBl1LaF8EFGwTGno+ahGvMFHk
121icRmgqno9BA5LrYKVI8Bp4kyZfXuRPIcOOx0kGoQwxrynIGMBe1DpAyYcZ7t1AeR9UYufIyca
JXgS5+0FdFqElPuDK/e5+hlXt45vj9S2EAb7KBJZQbQX3HNTizJXoWjphmSs2ttjo/V/ru00Kyg/
UfmIv1l3QYuB54mfWQc9VtZnXpMpgqYewBBOgC6acZWHeF4fgSWB/NCwT+Sy5mpd3iBP6i9fUJDH
C6ekK1C3GWn0RqN/wpnoRpOuds1inB+eL98ynG9u04NDhZtWnMfdKWJ2wfYyW2m1bXUK4/y0wXlY
fExHeg6Q+e6/Z9cSlEXcUWFesPG/yiwU7ykWN6TKuAIiisYl2CUl/QkXqozHnkv4hY+EXhEAHMlP
Kfn+bySLVDg4ZCYRc7YHOVU4GVsdgw/yeKznb1Ony6t1M9s/LA8qo1DN0z2m8oZHbBEbMm9fgwCc
/aYT/oiZi9Y86S6CCvL89TTE8jvsMXNoK1qMSzZ/j0elpX4qJ45EoCYOjFSIwYSUMGy6TrXZUBPL
g7neDCa/3YoDh/8yFem+mo+Xr49AdoSdqyhMqvhDykevZaTcvR4hCZifT05d4/JzfRL2qLb9jfVI
ol/mNdI8v/vZB6Brw/ryiN4ZK1RRKsyGqX16QNu1azkDrPHxeIj4xXXDX7xNKWuHKto4ltmqzP5X
awxbcveNvkwyZdGPCDlgpjnm8UcUsUGgKoTtDVS+h1PRWCNvFOeSKYhI2AJe9jncQSCXWVW5dKb1
btD79SWU2ZzlHzsye1XjZvSrEm152PhEVmcVefz2DFBbjZN1jVanTADiqmPiLZQRnS7mm22Iqw/I
Ov7MnGSb2B1pOD+OFtnO6cZ+j1WyarRuj1uboSNF0mYBTLk/W+tNQC6dwSVDhjnAGoachHf+gVWQ
OWgrlJbrVEZ0HzHNbXlFcs9OKoFZcsoZA3Zm1QrFN4gD6CTeKsVgymF+USefbZOKFsBQyyW+xv+o
XI1ZrVD90yh7Ej6YiDfoU+LpGezo3FHBh6IiOgvLKfuwyv+QZzZG1o3rFl7QP9M02tziMUK5pLuv
2DI+pWTlw2FhlD4jXhJ7JqjxkO0AlqBMxc6MZG5ot6K1u1kQYzmFAEbM30BNbh+CDDdUewrWicwG
WCQy5qIPg/3Y1WX1jAOA4/lqznye3G9GAu7KdspxViPxzVL0dGxJIwngC/WPX81SmH1kKRCJ5o+l
/vBOHLOuwkXs/4Bg1AsCp78GXLv+06WyOLlHQmWJEVXrNz28Ro4xUPiz3sA4PU0SV49f/eztPicR
TV/k7hN6A/GSxb9I5vjiQ/xMDeWj5LB/V0Mj7S/ms/7NZU6k90fh13zToe2g8z8ez6meQzG5CXLZ
G1WVIZ9I9pMV72qhzw9pcaD4bvQL21s33sVvUaRtTPUrkO/6wCQaGOR0B3Hmdc6M1GbiAEb8HP7V
Py/ftazU+mX6Rhgf1iMjW7T9lLGPu93PVxjd+L/u1947dv3JEXhkOms6/M9ZauL3Vq4TY8Q2/VdP
rL23UGdsCrV/4/b382g4qeCwFTaa3X6YKA9esV/XZ2kQiMDveTXZ7AGeDUFe/ur7a5/Y1wqqFbC0
OWU4y/ecDw43VTbrPnB3IUcEw02gLqeVVzgX2G5kRWzrzI6mRivS4a8tiTtaQcJgjOm5xZl2GDY+
4cgqgh0D99rffYTnobemRFWoFzDIRG1CoesBBw4DS4b+SSTRuTWCto/Cna87p3BHU8DE91pAU0Rl
mTAGza7z9+U7KQQoenKtpy1SXuTnXQjAt8q2urqwRhLDNVXO6j7JOExKAWe7jxgxIurmmh6HP36T
iSNTrhVgVMY4fInCLqsJj5Uuli31xMSn7yjweQEvBCLQtxenMAL2nKVvuwB4jrJ4qffz/3ui2RE9
KX6jS2t8GeMbo9flovniFXHh5Mqq06tb//OjCMonqQkZ1mCUKjQ4JE47wHPzsClSbRH36VgpqMQm
FXhDuWUtm6OUV5am6ynQxLEx69ds2IHnGku1fuycaJI4KPPsCZ5n0BepDmtBXwCdIDi/G8KkoLwc
B4apk/mZPvjRe1IjRRkIEWt9R9LWhP5K0J8Su/pSO+0BsG5ctH7K4KlT8gMEnsvzdfAIwk3ZH4Q7
g7am/ZOV4J330AxJZgF8WFAFGACVI3LDt86aPAMzO6sc3bsZxoy223/ipegwB7GM0y7D1IyYf1Sr
HulEVaPM8ZgfVkDKscUmfQyMit27sX+NEWX5uLoXPy1eMAQUWzsMHIjMdXZHkxrFXKOtIpTWHGRY
3qnFEg6opwNdeDU0WA24EwUsCKuaePJztgSbk9LAZk6JNA8opZVu7XVKT6cL0DCoJa/BwDCt1yBW
3volXKapewUr3g8QM2OqGf+CpUZQUkS00IidtwQI8NOkAvVKq1N6lBwFG5XXTE+hQwKO9t8VzPNO
ZBMYS4j2Uk0A3WVd5Ns/1sb3Lcb5a+lMRQyTzJOy9vRCHrJbXiDgZ5DQknh/W7uDnEOjawSW/nrk
kR+ErISqe6bqKbLuxFXswjfqSUiNJwxmsGAvHBeYNRtsgnV6aafEi+h9Wl0HFXftzgw2hG/kr1qT
Bdozc+kho89DBst69uczlOJG90k+ZeOzu2mpmubY95O2m3kCqrsAjiFpKDjzjtc2IsuzKYEG1Zhc
4RpY8Xan84NUQ9AsyTVqhwfm5vHguJ8ZF3oRYoQmbdOSO4dT5yUm997npfq5oeZkun22YPBtrk1D
c4oRAh7fV9sNQ11v5GhX8Kif9widFGQDSvOSGtTgkU5kDh0+HidNjLEo4LbVm2S/NuTwCo1mO+PO
jEJSdcw2YXKUaDCs75Ub2sURGHihtjypVQ0allHSoQVdKn0tRPNSS4+iI0NR19p/iAJZFx2MjM5U
6vFeUtj2RyR0usabAOpAyWyI8u2Pkf1IXGdR16JrWzYf+EmagwPcvHSRShEQ9KAhekjTH/cttDdu
/UETh1BLFVlxB6xf/BYAZGR8UWjneCZTh48TBLTQlMpr9cMVLY80glGzFQvD4NOyYSF7j0rPaO4x
AxcHZtHOkB+VQfS2FTvBddaLpGOI0jq/UQBTOBvBgUSIbSHE6vqAivaxaOvORP3nwWQEUuvaQ1iC
+nZB4EtBs8QSzGPv9KWwhPlEUvpcbpHw48XIMwoj3ztXd2OtTQ0KItvqyLXoVEobaYtyt10DU/fX
f3ypoQq6qyGLusFUfqznOd5AoS4/1P6lkRhwizDo7iCT6DeNgmxpy91/sy1fI3HSkjU3WasMiSIz
eJdVTo3CfukfBHy1Eh7Bc1gabXCZJTV1og3jiiEi1RUjtonp5SP3tiKT8FGM8Urgr38TvbySTq31
J8ykUN3wo2RGbx8cJDggKwKVgnjqsmXlFDFyGAyLU2+wFGbHYuSb4Tdo9eScBtF4YRJrnqKY6Y4G
NRQ4BZfSqFIY2ODB8mOr65PTBGeyfqw9EZp6zBNVBKihxFz4Di2OC15KuNUQiLRqHRvQUZRVYCR9
N85m4Qb9zYGu37uZwpqYbIFKkgIAIQFzS0wUnhM86gtsSPIk0IZYH4Mwseq18bU6m+i8/p+ImGXy
Og30p36fwtoDqEmhbQBKVKSzsrvxJmnfBhpWvQFmaxzYo8q3JzMtPSWDVe8MkRz7puJ84SJy/l3i
bFOKxUS/WKHN+2fucAD/I1kA6OMF5O7ClvPnitTzVjSajID+v13/2WaFVQEHn+hULVJwCFCOMb0S
Yg+ftZxT3ViZuHyBjAA0XutSs4B/ZwvMMqvXUkOYVg+sFg24iiQYfgTNjLiQepgnsbWdWLiVBopi
Ii40UI0jPaLLY9K16WLnniItKV7cFe2yQejqOsa6I3JHO3idUIbKFA6MxGd5zRWqnAbyT3rTk8ct
rC1LC7JUGQpIi3PnNqrClX+CR0KVkblWg1D9Y0yCw8/0IVNcirSJdOSWxJnFa9PKGQKnkJdCI0bt
nNq75MjSam9Pl/iQSgjtMaPKOWrRQ7t4H/xzq0EaOpud0O12tvPc/gP+ltSZR/LxlAPMUj/cBeZv
16L/tlZTPSqI0bOXRa8yKKISb0DQNSGlYZUmrZVe+PG/644a+AgMxVseuWsxhsuuwb8OlE5MGDcu
eYPdsNFI8wdyUTJeJvfFPRrX7x4ZcGPb/Qplim4+ZEl18kzknaXIv/xsLsX2DMmkzTaVZoItAMgr
kTGEpkHjzEnQe9JYUmy4kJuaUVZ6u1jrTtUhhJTTI1fHPlj/OwvIOoM+UvvC3xgRBKF49XcxpW6n
BR5qgR88dmy+MFwHesVU4Cbrh8bSp1T5XZuSLjd/t19dIWRg3KpMKLFNzpe1kbsoyI9Rgf+X3Hrx
r7nitAWWzVNKAw/TVAgfjGfZZrdEj6l0QQhp5o9bDEymvxMazzECAxxLZkkN2BmFwl2s4A8etYKn
55Se6/cLSWZJCvVQGFMtdax185fdZHDrQEp1Dy2Ov2PMelp4tDQf8f6SkuEHFWKfE8VceWdzFe1t
LeKgmRd4PDhwgTyZpMm06PmtEdm1X6k4GkFHTVMHh4sUNHjoon0/ggiFcE48HcEkZMOIb2Kl9NMI
HEaadNVjRgBvMaq1eawbSkdZbmGfSQzXVyRShWCPhLEe0BBP+03X/2JD9Df9U/r5Zt0tyrvCPi7Z
CClXzU5oESil7Z64WBlb9RlD7oRz4I916owg4+s6MJi2Zrv0zJXiZsgD2PD6X84dz3VvGH7o06YV
+92lRdrt28urFBViVxE7c6gc07SWSQfUnBJBBrlKqZipyaTqUeN06F+00nQdRTAANyl+g0WCXy4J
E+ryB+jcqstVLFYHr2cBJdINwU23YfhBQayjv3axh7GZLcWuelCGxqkMPauvyFUEWlHXx1Iefq2v
P7g39qpGTj+v5h3lit6MG2d45oHU10V1IVkBrHv53JGTz3/7IbPXafBwTnd+uOlMdhlwGlHtLGRp
sEFXEnIl2Z6ZkBTKpFdyVvE+nC8V/L22lfMRQzl3+GWADiFAvPLDw8yCQSK3LBUthhK4gZA3/xAd
ZAa3bivPGkOhe0GF1gsvVchDXDT5dsiPpjXUgXkPYYaIi4TC8VBD3R9XF+Cj3lxP6/zthfacz/7m
3EVH/WbqbVut//Wqy6pXITLEzG1VJz3Ar2RCU6UrSWAgZ5bKUpgqPF0zyRO9MnkClI0N4XFOPaFd
BCL+VYbOYx8p2WnQhqYifuBggIN75T9U/D1RRnS2Y+rhBlzE9dk+hSpKfGXexSqrb7VJcf4m8ulp
//u3n/iWzlMlTCq+H4rHm0qGeGCa1M4sb4S7dyK/DrpyFx+necXmMkIhbjXYE6rlDz0bne6Yh+Od
Xm+9Sg8kHeUBpBAv6ieYXt+vTGH59ek2IY0u0FOoPALb9wuKdDLDtdaCsB1mymCzzEBHTaqw6f4x
/ddskccqrJ+K5NU3FiUuTkMYbtIxX5YAuiYfqB0XrHx0vaYEptEoWuztfeZ0jP8PovhXednYcKw1
ii3ZJrzKCjaxietBqPbPGSwNSeNDojFXYBXoXkYPD7TbhyVk7TE2s+fY4ke6Ghy1FPoAyow1Ig+1
FGZvM5LO5SNDnbXuNzYaOJNRq3qkR4p98ZxROaI5EdNvJZJKjZBYKNddoQSIN0RCuvotFotpxY2k
dsxX0Y19Lkneh7kLKVicPB+i/v2MdDy+hHX2G4hPmd1aKP7MkiUApRHJSt/KLNE0OXijM2FW3MnR
0uIIRErk+Kug0T0oz20uQyGq2ELyxcNVvaeqqMLpJTiO6DT0h1JDrIhYzmXzJJsXGJ9nbUfZPmyJ
JGwF91PfeM2mzXfpqH3sdkkZZ45L66KFL8zF9WWRkj5S84JRhMKwj9xcBOxu9zk2uwH8PuZyIRxk
fCxkf/1fXlKgYQidLB0r+/Az3X9Pj0rJHfYTr9Ydz3JrDWT7MCMawn4Qtj2HRQC6L01EZnUWLQUg
uhc32C4n9rg1df7fn9pOaxeN+Z9Oz77EIw6Qw15S+plBfpIGVfY3YO+6RJWbhXqXmobNqR1khwxy
knSmMGsg/rHCCoeFJ3zJouXtI5IQ56/cHzn0hwtca5OcongKwufUR22CYu4qSQljt7a6YRfzZ5Qm
HUZhcZWN69W7qymseIe0wQx97I2DIAU5wYcgF7hmhUIGoFjFEkpVc29bDU+x8hq8A/p/7iEgvJx8
o7pN1CB4gCm4+CYFYaYEMbUfY82Ei27MhsWtEuxCOxpD145GHAjnZSnhr7eqDDnQtm0fZrJEN0V+
CkxuNQxGTlodzyTGBr17Oqv+Z903vDtNUTtmZqcv55kfchzDDE0jibkGApzPN1PBaDWB2znzgZHJ
Uvr/WBaWXDCWfD3wIi3dEDWnLtHBtRZLu8ht26LrijrXhVw4R3iMN6pgyIj60eWQEpJJjIpovQsG
o23ACm2EbOAp4dM0DiRY0K2fkeqZ7n4cksC+OOxwcYqppmS9B9JfjUXsjm5NqBnHu4fqJ5veo+SG
W+Sg2BtVYV+Vfc9k++JgNRVqU4EylgWhRgolqq/1NHMO2PjvhGKe4QsZ/wx+7q9dlexVV6zv0cet
6jyNREJrriRMEpeHGWMFxA7n2bL/Ds6iNtpEI2Wnyz/ZHe94ttGfn0wAAdUfRZHkHOpD92VV8Dme
yGhGwVbpQM83bXBqFTIhLFn7KzpW+gQTfqJfEWaWLZh5DGqh06UrKbQqlEU5iHqvZEIoOmguIvVu
cpnjoNOk51AKfVFnviu7uyxKRcsLVus/jL8mtY7ArrFykT0lEbbEGgeM52g7uqiUeGauCC8Jkskz
xKRV5sFuSR/M0nl38fgTQwMLmbc/S3/ZIUUB2o3lhiWqIHCAT/nCw6XdeP8D83G4a7Xa50DxS1uU
XY/uVFlw1WNTHSOYD+iiB4mdfabFGWV2bJg78tLk54tdKR1wpfvlGjbhMu5Sj8CI7YGOI0KrAaGv
53I1Ng+n3w7TraEBIH02+nTHl+OQUrCU/N3QrELEj9wmiWJbfcQUBIR0c3fhsft8BNiqOgZsZXXv
FZKQV18isOCx4pHhrH7k8n74wBRnZlNnQUoH1youlxoKjd6vBn6Uum/fBPERs2Psff400YDgPLiv
f3fsXXVwfIsBQgrc29aoE4atFAQf2n/EWm4ejlKCm+1GfS3iMF8fPB8lv/T0WdPDMBd4uM/F508G
NqrOBa8SQcnaH5+cbWcIWy0vrjeMV7/0utOrslEZ649/nMAkP7rLBpCX+74jXlypIuupICNhVwyn
up+vCwGR6f8Oknsw5geXC2wNw54aN3X9qo99ZtHEy3/sMYEEp1s+/DUzMsFxDQLz1oC4BFcts8Rs
nXTYThAwkeqwL8AtGl5dOiqvt3g9LuD55qmtJMomuN7+XYim3gmOZEuBNjKBZs6z/c6SiN5SPHy5
hE2BD5YhkazNq7xaqDphYOqK70NtHGA3RyyMU44bxu2juQrVbiLpm5IDDbx1nhRQwZEcwMC/6n0j
xerVpgUEkud0fozIpmhdY4CjBvnxub/MY7nVTqgS1v2cyQWVaM7+a+ccQ3xgfzEp9xbse9YkgDhd
iVlhboSf4DrIDpWz1V8qvbKRuaxJWrHiI65Ley12N53k4NGEkBCpMrLxyKhtR8nuJYdXUquHm8bz
N2LyfjOdRqnq1jXZ/J5GlzpWbwaVkf/HBgpG8ZMI0UjcX1+4Qaczlpts7uoQAkIAEkFbr4zLC8r1
hw/hp01jOiJFWxIQKF0sYYhoFDKlzfFNPbU/p0Glnn30zJWMMDEoRdieu2XkOpS+3bl/HLIgXeX6
AiNlEI3a4x2XrFAy/Hi5n0gT+9+8rL4IAadrmm+U7u28U/mT1nT9n4YEddJVGKK0ANltY/HXBmJZ
Ky6JabteBk94RsqHn9gvWIcOzHk0fZziZyxDkFeFAuJIOJfVJ8cpEqeoL3VrcOQFKtZ56a2/pxE0
4vgL6LWG/CJECyRcwBt4ySVQ6qnAar9AsbFVqtw+gQvqPQAgc0AEMSpJFRA161qs8d2x7fv4zsGO
OnIIy/IY8UvHaOT2Te5nBf+bwZWOSgslpPDlGHVjw2xH6rSBUbgrEkdP4avW2gZAtSSF98YdEZCi
VDEEmeWj4VQ6qukhMw5RIKai6bJqfHzB0Qy5z7UWFwaZAAFg0+A+vT7pe2DCkF08Dytn/9l5qNtq
6LJG5wml/QMzeGOXgj/KmjoLbyHHZdwdAAEQ+a/kwozIBcBecwMxn0o3QLoSquayxwPrh0eZF4hg
dYhb1O51VOeBQ+04P/8ccThz8hsiOKStlYMgFDw4LXnhnC7kOOkwXcWYwKRmJFf5EPOC16Rlu91x
C1IRuEkdvdsVZ8j6l5MAAWrC7AVj6FdZzT89DblQtUhrs8F+WVB5ksrtGrgtL1gFYx6RO7KByUvJ
tf4hOORm48AX0sVSfMQ7u+N4J2vBf3SM2Kt/WkTdtx3GRnOs5xYf02Nj0PYGeKXyWvQHHI+h//7L
ECOQi01yMKiCQgbCLtWNYUxoExPHlw6jCUE9DOyrk4u4+/nA+fbD4+o8MkHs04VC2gp2o3QKIC7+
Qoi7qptftlGhrA+UtmSvX5FzdhGjeNyTodjFpNyxDzH7Co2On98j3PjyEb60RqYUsET9tMZld/xj
l1veH6DsyZZgS718jSwGtFQikbRvuqRMJpApdRFiftU7yE0s1goS7jboYiAN3yOk4y8v4SbQWzf+
FbmH2j9FWlTWtVwUH4+jbfRuvtltZueVcPoriI9R2zqxUZCgfSuvro7kdOCAHmvIqTS9tzjqJvHy
n4B0fX84/uInN9gyBJ66i3BO8xxkeIfQI6pQrGuJ5fs2LGka1Ca0z2z1caWPPu0tGnrr7aU0AMxG
UcCogBgkR7hQISS1lZEkK/fwrOuvFQROAv4suJlvwhQCIKSI1JEIiOL1sH+oZVkek9R/TrnrW7+T
86tf/IXPcnbyt0+/hHRloIJjmB+HFy2HskfhT6nyMHqszSANBpVtlAgs0dNXrL8sdmleyyJTF6Xt
sZpcW5T3O3C/+ELrhq8PbNQixD6qXQPjvJiuAaVUUz3kljGYtknfyp+iyNzuR272Ziw58N4ACyk7
RyroYhKD7tAcOPFOP4WzGnqusT8XlxEcZsVydmcJilwNdQfggYObqYOOB7Df23Yhz6zc4o3d1pp9
va498V/NXszbsAIbJcCXSj1voUTFmwFM/fE6Zlau79RQ+otlfZHD3bPnnfbIKNheEDy54ya++BZN
t4YQH2ayTGsaKPii1cwW19ZDk1eyAjT1CWOM2R2C4xi37lcGZD5JHhwXjz7SFBVjix+bUm3PYi3F
wLcveWPoEysn0YjA6YX2BxwD6/zEbBZZSzTAy91sRAaoSo8WBBiy3Z5M5m2l3X6L/AxgEewgkYiV
ZRDyid5yRkf/6SMss2Af6pFsswoGVNl+qE0ip3MKppgZ9KjBXaIl9GRV3H3nAD9/CG2UkLQBLT3r
uhlepWHGba7nMMJnl++QRnQhaCbEJ+Z1AbzeFzzDJ/JgrQEt0Hu0zV5ITM/RXJ6wCboz03ijuxuN
Rc5bMOOzzA79GdgQ8djRhuQVnPDT4vwXW/JiVLrRcSl/mARDtQ1I2vQRjjxoaOe4CimjE62EgBcJ
3OD+sLEkbK6ZciSkV9OkP4fC8tfebgbH1+e+Iytteamb5wC7DsfNzFEV+GXpOBcB4AYRlL93TGUg
HQ4amL1vmB9+bN68BRV9m7vDPXnRt4lcMoWjd99r9HJL93SSoo8HzVUUfkUKUp9HyyobaRND503Z
fqg0fE0SpzD+tyul2oMXfyrl1HXFW+bJpBjPd5XD8VMeCf+BvabD3vroe97TP/1KKqaPlDH8O/S5
BOU2+6lXmFosCoBm2yoGRAy0Xst5rIV514cYRovKPdySo2IKS4JwIjUcJhMTKLFpv38HbKTiQpPc
luszCOpx/rHEyba0nJUtOyFCyAjrsWis/u4lhmwgfZPH++pIylTElUVLur5fyk3RRF3VybvaxW77
/yRLn7s4ifffkBfbBK/lYU2kAVOS/RFDiFtc8Q3xKR1cHd4R6lpEWzCZ7hPvXUBiHX8AANnRvJXS
ZydFqOu2DkmqvTKP3ipmjf1/NKTB7WoWHKWpWVjdaZGNS7VORXyKzA8DzPwre/WK1Rv30s0lH2VJ
QYHkI9ontKaz+oo7PS8rz1v7rAIB/1lf6SToiN3fPyixWW76S6VnO0a9aqvu/Ohg+ru0M0UfyfTq
R/6ZvJ3aToZYAZj02EJjHuhGx8WXp8aX3wdyydsyUptTuFa4uu1MMdEj/4TrNRcQfTvwBzt1qEwF
jGVQrQu+NEXzgINlgW0S3hyNS1PPL3i1MC1zrps+2o2E9Ga/9T+ghzTYAzZT9iJWbvWeV6c2n9JT
RncMNxaLbZZwOaVFIreqgypBT9qlGh4h1vUMHRg/BU61Bo3culn12fYvCsFkkWNXHCQseDawi/BU
k2p92Uz7cnSJi7m0WPtzoyJsEo/Hz0FIWsRZ41Mw8DZhXMNB3czv6lX3INEGzUrQITbRHAzHT+f1
/moYoS/uTNXEyWwjdT8Bcn1Y/wc9xLA80GbWGxeBGUvl7Sczl56DNWM2kT4PromvoCOqLm6pzOdZ
B1UP0xXjFPAypmoIVY7KVSP62JcxUtGIENpQ9kXhCKfYOw2IYzQLDbPcsSvG3EBKpismwzh6yxEs
7U8VwkwH88XmGgLdIdt6wu4GMUWg8crLvPTFVD9Fb0edxrtxVriohwr7XL8cv8tjx0TcSbe3Ir/d
mZPJm8X6+GfO5Oj/STyf/8l0y1huKQgxw1YtLkqYOYxCcQXYbX2aQV5p3qk4hLB/SBJArODXL/99
1PyDSSSzld0v2KBSueAfa8YzDP2lKMiQSYlUoIqhSks0Iipn7Azz1JFN273cQLNkm2gGcNDF87qe
lgcBoNrRpkTRezbAGZxThsjzOsfvv3N0ojuNqZKQ5g8bAzVAIUWuZPsFqkcDS23zbOeasJNi1Igd
dS/Bs5+fkAkWdjgJrkWEdRIQ9pHECu06kX7nwv5BEcCGNgRsNgsflj0GFVZRH+I+vHVfrNlDeXrL
70P/XhGkVNAMNigh5UsL6sLuRsvU9bU+Nog46XGDgxN4OqEH1mXuvYU+0M4YeKk7NTT5fvvlFK0c
AZEDB7Y6B+/DQz5ejazDobMC2gDUfQNcShWqiZx2ZPYkh3rrvZt5shXU2vmiUpG/jYFVttk90L0F
qTeF6ErYE/Etn3xx6izUW5M2zgVfa/KXLsg3YXnKqIv5QmbmKpSbn6rCLd7l0QWt4V2orBB8Z4Dx
8T5YFREQ5psZJT8JjGz/r17CFqh9pK1vuL23jrtfLaEzvddGm1DrP8I1sx2lGWCM9ku8cDwa7yaB
Tfz76e6WPfA88TiYLZvi5YsYzCOJmNln7vQpAAMTKn68n1AfQ1Kd9ORg7+JrlSNKItlUw0OGzN49
jnSkEnon5hV/6jN6TeVzlpD7m0Z3MhcGbqVBQZyrMdBgkFxzMJpYISIOWVBIc5sOculkxPYV2OMq
697CY5AWl4qYDO8tMKgcq2vV0pEw+sAjAFCXKxrHS2oMZM8zv9o+WmdRQjwvZwi8WumaulvcYjzb
A/+LUgr7/pMKbCBEIrEqHfEOYiucP+Cyt8SJh/jjeByI8vveth8DhOjvyz4+eWy8f5jU9TqpIHm9
lNuruagfkHjKoQK00WSkd5N4zwWtWKux8vGrKddURp65BHx6RF5QO9PazkkaouvcV4G1p7/l9ogM
YyHMLfqFQQNZV71E/XmAUZq+EcnJ8Jtyv6dv7lk6ZOlhuWp4FZlnldZsdQ7qm/oDhEmikEN3n/D6
z7fd5geiEY2LueKSegx5QKD4e6HcTaZI2qyMaw7S1BkDGE8DaiDHoUx8iZtY1g+QaztD2TKmh5cB
LzAAa1QTdeMsKbvR9Nx7vizNys4fDGjUuttejKegM20hfOLkSveR2iP/58sjkCSrJPGH+3wEP31r
5HAD5msMHaQh8pyA/eFbpm9JrxykMnTnnpN1hy3Ud368+VsVDBmRQwD+JQvSJYJflbev2CJ1O/Fd
lPA9bIP9mn2XLBj2YCX70aq3+YoAzgjnzYRo6D3TguK263Kx2K3BaOyzkbY4u0WBzfyPdX/CdDoK
+MDyl5b93youRh+5IDhTrVyhFTriJbeiSFloVuwRQWlMFQbibXoSB7e89k3/dxOflRg63T6Uv4Z3
gP40WRYL9wPvTKKpQKVv7V4fMWzi8faytV66kVY8X1TwI6Vb6D2HypU/ux7C7bGkX+mwOJD0iSXw
w//aJJHYOV8gDjQ3hUJ5cNB/a3mURWf/QpHVOOTyGQdVlnYbH/DoOC27AC/zNsQFJ9n0Eh2ONe/+
YTaru/nnGDaeSEmlO3/8CSue354aSXBH4tjSS0grgpcI4iS1raRuhdYUnDTEne4gP5I6Qa/qp4P3
E2zWSBSmIsAerxNXWxh6RmDxkd35W7SyyKc/sbPOObHHYrMP5Ms392UeBbTGHUKIfFLMW+Nv/Io0
m5de8kWxj3rPqWN6fp4vXTJET0zrJh34MA2ThhdPkXK9efPB1JZgEGMP+zkHZ7TJHvrUutaQGA1N
UufvdZiigFHPybD3aqQlNGSYbNODDw1DLJDn60MGs8Oq73d/WSDU2uafjcnL1A7OoVU3X6HA0iRZ
UULNaez5Iu9VfmfcT9VnHpeeS4Tfnz7p2+fMuw56OEaPmFF39fa89VTRVaf7JsUosAiWgBDSp1lL
exSPKwuaHhD8nKnZOXRgRF5AhdDN+XmL3ckqwgMqURfl0VoHd7SWW0zKaYiu0z20dVKbTHQLUgzE
Z0tAnydtCDhld2xLBfaQZ6FvszVycqqr84C4VoLJyQE2P6NAGISUh3B5nppX1S0Ppmyr0Hdedoax
ibAU/gJFsH5wBOm/2uNUskB5x24RjkTVzqVQGOgRXPjzh81d0mFelL+smkjJplvU61aMl806gjOf
XUZb+xC3q1vs4/6AbsTcouk2DXXx7t4ddenPU89DnZDrTxm4rMpCytsFlWpkqxVuSkuvEAAOcDrS
yQ1HkfJYj3bJYspz1imxjL+CeTL5xzzxKCgCTfAxybqZ7Aquz34irImLCm7RZwsTjwchj9qfMeOV
DFwwkjZRMQEQkyl23mymig0XXx9r7w8CHO/lAtWz9BtsBs+w0t/eqiKbvEDH6f4Qi4HrPwRkoWCl
10pAPSJYnvP2un8wLY11nrFkNMPiWzo2gGOcf0KRzwLTmnLrBWBOoHr6pbOg8BY8VrKxVIZ/ygeA
IAKNN75prcbjsifm+wOLzqN7Iy6W/1ArS0X45yXEyl7mPYz38Aj/mh5ESAbZ/zK5rWygKghCxe/3
zwhKOyimkC3SqWAJZfU48NUgj5Fh49ZGp03c7OIsT/3OrMl7jNhwUL+qEe8ZpI5oBgR5eUodJmMh
AommaWhtNwvyVtB3oLm4BEvQdGRUHt1N4NSeWw4/mVWavuR6F7EdOHqTfVd31xv3iN/EwQe6u7E0
Bp1ZQwSRhNZuQTxz7BRVUOAgrEX2TYv3eUh306OBhdi91HhohXsYyGhP1/mQmOhsUSI+pWepDMt4
j8NbbUJ3HSKVaFaG8Gv+VV1sauMPWyBA8+FG9zNZrDJau5l47cdrffLcEB5pMF4PUj7lM4eWP6sd
umV7zEgdvUTdsUKAOmXx2dN3lqrN8laE+KOfQp2NHFVRj/JWFpq6wW5zAE8smI+9BgR7a+mClEwp
P15jqHIPP32d+zUw2u5Mq2y+Qh+RITSvZxfJE4l6h5RXgx8RC2jdIt+2l9VjIDemYtze7Os285Ys
MxqC24aNpjho3ZSvznDhsLDYbORo64Xet8oS7NJnugPgXtM6xPYcti0Ugw6WGfPJnA8q+g0ewum3
XlFbCgdLPrPg+1CDP51AD56/RGNcvoXESzdeJF9D7Z6M04e7mcZhI76536WZUHRLZ/YYZkq6Z01G
JvkmtrGDskc5LeHSTJsSxt5fWubP0omSp1LWIJodcb6z+vBG4RDXfJzxeO6K+DkzOsXAf0HGkLoj
rVN+BimIS6WNv5CHAc4l5v4OytsfDoGCt9+BhjBBv3b2KveWRm5abl8W5JWzVYQKrGm1FIHU3TKi
4j+hnbzCFE5pwsyaJyFpL5KCZuvwnuHKn89Y+fcGEGhk89yGXVu2j1qKHxz0cdN3CJa+iicYf+j2
p9xPct+3AnehSmWD/LitzIGwOcNoe4LQEuhisnpShIi/mfIkoVtCj0scAJp0ud1BJARTAEngUTC9
BAyhJkInbqiT03Wfv8JbFJQn3TB3H2X889yp7rjh6LuTgQBhaYfFn22DCF5mKITtMF+be8UNsEo4
2jJK6+8Q5RQy+HL09kR0R6tOdH7lwSm8r1rPKyu/ZD9BMBjucYZhdpv7pMblW6cnyv7vBAwzWVMI
nc5WeDUr/LLnz/WGdvOcmgtw4Nkz0g6PSUtFIdOEoddg0ZxVL1WgiQWOAnLulKS45sDY2qJONGM2
Qx7k83oDyV4aXzmpEtgbNCsBAUFPxjQ8JZ4rkqQFtq6hPRwTUZEdUycZdqqBPsFWfKdGZo76psFo
bbL6Iou4/7gfPK3qL2yUvmGMpJ9Q/mgdCN89wpVRXl57OqsixtyMZGD8XFyzWY2AH97KGn0vIH4K
JMYBPMFe3M9e9C+uiCmEg/tWatcmsXTPb23+mftkQvh+Z3MXL6r4w2D1UUq8xI223jkl6WC2mZH3
5Y4FncW7lC/9/WcOM1hEfrslNTdvPV7N5QcxoGWymmYH0el0l4FoEfPsX5bxfCpWYUEYKOxeSaNU
W3oaVnM5c2SvM4bMsefAIb3nG+B37KX2HVbuE3Zw2Q/xhnBywuPLvpfjm/oM33lfH2tblpQDzZUF
1cOW4aNoctDAgSGHpReGYnYrTFzWiKgt6jqsa5duzjT8eCcb3mcC9pBmEyKfwlFh8GewmkdWwI4R
uiSwY9kvozU/Rwig1thvGFUqPXrP+svpPwY4M29dTxPDpQeSuIo536RID3tbQVix21InPVM2H4f3
qZYuUraliEl7WS27uTi+1Kk2mXlPlfr3yxibpmZCwli5MWs8ykyekTE6UzfJ5ehU/zuTgDCB8njV
ltgQovq1Db8PsN7KzY61LnDLe0q1ohmDl9cXrCi3E9ajupb8SFc708DsvoNCZ/5sXWFlcBEJqPIM
EaICT/v9jAKcX9/kQYVqohSuLNdRYtsJUhPRLGl5f+DVYOgpbzKaP4XWI/nezSCXB/kVWzX+WQml
ZP+i22Lfik5OYHqA7DGAiNN6GKiQ8TJ+ig5ThUcHC2LXtGE+sFKZH4SMvToyyhALrULHRqu8aa7Z
/IkwuCP8oVQuZaVSlUuC9eE0y5iTv6JgZr/jMwAG+2BJIeh6VZmmNLHx/wPOjIs7+rY05ERat6gB
KvKP2rshPr9S3+CN+tWaIf5JmxNgpXQGT3YnxlvdBZOMzQqdbfvJOb7aTONMqCicpbuoWMDK5wAE
TWbM4ShQTT5EFu5KOWrDyC5Klgvv7YJ9Qt7zezvQ9SnPIsrO+vtLm8ir5UGPQ3xlA0U27BaV/zcK
9Z8+F9zL3jyiNu0H7EQ6zCm1ZM2PZPQODFn1AUhLqSb1DRhMig1uNJj8G5V9YmSF1A0nbloGs2am
744TRB2WZWY5XTkdbr2KkxYGveZz7IOFAwaXADUFbtfLX++7dcbTXqdVUnPQBQLpGwQZhBPrG8eY
JhJDta/scgKwjFvQRHAEgJRg9W8rg1brU2J62EbJXN3J2vRSFsoupmC+f2cUr02KdLi5E/Wkgowt
29cxniG3psPjGokdv6LZLlUj4cjey3MYvIPJjZJa89Ar7qwclhee7OPq7XD945VeW41PU7l4G47X
ntqigibsx2PJqvQZd7YdOHQc2JQoXmamNWoWDG84Cj9Hnb7FVzxSXqkcOByVWr+0Moq3ptretFIT
YZbKMpEpHKAk9FJcMy5r9nlwBmCieLwI2Z3YIxANIJbVj4WhRe8cYZfUkvZy7crQXZjxM04T0BDX
GjoIC2vO3cDZUzZ5litwfL5+A62l9TeEgUZkqDW8kyxWrFdR1r6EG3I/uRK2wls2EH4AV3dBtA3x
yQcXPgvTht9bJHt2jzGgZAp/YvDl1czujT6sKf+sWEnGNGOzslloCYXO1Rpoy8a0kAGG18hZGWZL
QFiTsvzLk1w6yoyTZuUNkccfYwQAdVsi8mra1PjGbeRAF2v9cyoBqVT4QpYy101ak4RdYVDdd/vD
1N7R4AQb88YYWFg+JTAD27y8oTCkOBy69HyzHkw5LCkPVemPPTOW7vXCGokfrOq4nYQHK/l11MbL
zhWDKehZCAs6MjTniTN9zHT+37S4h8G3ZlDzatDZv1y9uCWxE1ZeouLv07bc9T98xDc03AwsB7aL
r8HGXKchGkZ4h1r2Xk3ZorgkjZPUaW+usUBXXB5pw3IlbV6KAKyvpOGW9uZz62c88peDXTaVjl09
fNHiRykQ0WNPaYu7uBTMp9uwBBFdB61BCcxtK58w/nih7pM5M6rPuJFwlrpdg2dNIYGEm8XtzdSt
QoPqiQdqKxUgpDXomvbMXR6zRlCL3tm6Jv9oL1YIE9iZ35KpmmzpktgEpeIUDm4RyNliwJmRWaON
4GmyXrgLIKL/mWdp56QtG/QxSeT387spW+y4s9PaRzjU14qoJXeG9ftPGcMVmayeB3Pk+PNHLaKy
D/7RkM7LscQnM66nyqvg9XL2/qBBidUqV0PpH6NiF7TGV/aoMnTaOlsGQYPTCbbdUOoc7kPyILJa
hGhtOjSomXDsXqRvTCc12cZM9FBQVrfI2yqDK/gMuu7AhmPutgXkR0oxFk6Sspl7LeHkgDoHKHb9
OfVsAkgCWLih7aNN0dEKfnY5XX4MWaXw2OElJ0LBfbJj6f2jc3imOxcwepGttAAxMz6iiqfRtekS
DhKVDi71batfTLciyflwwh7sWb1On4UCQbQ34JQWU7dUfH7rcN3mjbktk6c5HT/A14En340t7+n+
4XtnGs1QaRKEl9LalAs+nTGGpoBtPvKb0vUTRcvByJwfJCU9WhnHrWrhF2PLGVeYA1+ys1MCYKC7
9MrLTqP7bF+xZKABHuWPx8CjKyqm5+uYZnD3Gj2H+uIIl+E1FB8752eO/dMMZHOrrv/kChbzhRhz
PTDJkvrEEMNVgzsaoFYfkEE6apobT9aU6yntCVmvU/Ka8a6Febmg2/OEQRwjtgdIdMHyxP95gfNa
0mKQoJ7R5fL+4AD+LjgpHDk/RnB9pnTCqcd5nXZzyiB07jOqjtPxrf92NIu7XZU6UDndYUhSgu5C
1wObcy4Jwfwlmk/FFpI1xd+ZEDDg5tj3gnEOu1lQSMzW4crgGEn6i81NaRUG9oJfYJuhpzRJQeTL
Ys1ybIGmoCeazEVJgGdbjbDdn+DP5/QWzyDNvAXZ5mjf9Hi6u3mWNHuxY1a2t0iZ0eOjB223cYAo
/Jny31XbZJCXfcpggYmzeDYYjUa7MPG+hLe+QYab7Jdd0wkDupzAB9w5tOnK+RSaRon6dblpUBMn
W6juEq+lq7ub+yFCtB7gPNyJrQrlNCE6kXaWkcO2+rQZsm8SwoQSZJrT5xCUvuTmcq4AH8SmzQo9
rNwrIZAmrb3dpGFCK0yh/YrdTs18iaBxwsmy/8fxypCllmEBHGOjebbRvaIHgDxVrltnvhxZ5bOa
Zcw8bxxzmX9gB3j+U6byJaGO93Q5Nl6wlD/q6kI3k+tZ2PiLhToevF5dvlj013ZAHzdU5NgJ9eGc
WxpEbhqMDIknQdv4hiQvnbj8XqgTkOm/m1FpgYouHmvOartYSLBbvktSkhWscLkfPzdbWAw2wSoN
RPVrPfpEFQrEzAONJCh/ivYU+Aaq2mbUC1ZpTtLixhf7QdSf3WZ4KWRHon/dk1Ycw45shJwH3NWv
EhCUgWKVMb5NLl4MX9KK+xNS8yztRwiItvrQDRmJMEU98gzpmTv6giYLc+Xak2IZy1UqNK55FESL
rUMOQ5OkXZE8dDtmdi2NOYx4gK/9EncuiEd64TVDihcqTVHjLtjkdllcDMlTEKHZ/Kdvx91JeU8o
zx9GE5AS265pG8LFq+0ixtaN3Zci5ssmd4TXkbgRp7qYE7ZBGA2UbGPn46aZKht2/+na1F1GgO/G
VvxG/uhqKl4FYwxXsQHYtv8o6WRMDHIaqnUeys+fEsr5ZASghsG5r8IPQu0Q+8Psf5QfuIXpNGgW
K8zpUpiYqg1w9qGFNRGTL7YCd8ElvMBVgpnGMk4s/y4avGaK2TEi00/Wcp5HRGvUtcDCLmRHOxWW
o07R7PkWXq6t1ccZ4QwYSuMKV0wM/rFh/tEtJNuJBdN1Qw6k88YtL25bN2FY+oBafI1KVC8igAZa
SVpz74xbfDdchXMBRjWHEeEP5vvRdTgGEB/QoxV+ZGEV4y/eZCwOM4VWyymwuHGRvf5lhLv7hIMb
ZOd5OC2jL9xvAKmYCYMSEeHv8evLPznkylG6cMJ5dli38MY9NnBCn9gt5HU/kFBJwjoP5wFF1V8Y
91b/WFuaAYG0SMpZsm4XvIwjCm24ErJ8bBGwh07MPDzzwG4bVlP9OdGt06IEAwwebcxIy9G6KhVD
+Ih1sZKDap5pxbSGSfGOm6Bfka1d3x8GMa1fh6yBw4tQLKKYgIp14f0qy756Ay9o7VQESteOUFtw
z+FIcjMbdaMjW/3vIK5Ji4x7lDnWK/6n7XhBlOeQmq5YWNWpguSQNmZZLEpnIzSix9ZBoubgMrpN
xjRZGRRGgVawIBZ5BXVk36UD85jEnVmSAGfqbh4U5cXL7RQOoMR0vGo4rHvdyuANKnCaoWysGRWg
96QeelZh7Y2V8lfHaax8AmoRPG0QTWTGkaWLKGDAPlkCY48xfjaLq1K5m3M7mTAkacc4nZ1SjWfk
W0NhV4vmeu8XBVlxVEEMtIq0KMVa6PaVjE7/hrPJqVPUYD8I6xKFT6Izv9BqfF+Wojzzs9kC2+Lp
11H2x/YiM0Y+UT5GHWvRYWi7OYLTZ9tywM2O6USa4YHJ3y6Z8+TnOzKer8A3rH6CF1RHsyaC2hvR
v5PrhTlXTyNuT7ZMo6ISzicCEvTlEdcPnDFv34QI6aCD5tCfEpU77WukAx+MDnSrBZQpTbt4+w4A
42onROeybhqzBLohT7IGJf3rJyT5Md/3EHKmYCesjMtS+V5RveZbFArQbyumH7PWAMuz6aScvtO8
EhE7I5wCXaz8dJfP1bjjZkidFoLRxkNgum7YCZaleVsCD4Anc4hw8ATs4OVj711nIyksbxXB6dfb
9FGnqBpJ5UxRG4PVSTpmdPO+0dTng4O1QnX0LlptIs9fUmMsOhYvKwx1qSwph6P50NaD6hvJvuFa
pryWNcEJ43e93r0zOMjrxK6rDf0xNlis0aC3fOpXeJzQHoOkz/EAjJvjE6AwNeRMJUc+rFklGPej
+PUZ4hGcydHdgFaTAs1vjDgHPyJGN/3PpAUtwZWEwGjD8g1ubSsoyeL1ahPOa+rN5QBYdTTjF8et
TeWbMQ7/6SMMWH2QASZMRZPHHGBu4Z2KOW5ddznjJbI6OmXGgWxjaMO0cwWonM7J+Kao4blltBD1
R/3gN+DTmgRr+Qtn9QkcIx2t7HP7CINeHl+tewGwbiJdpuJVrB5i6QXEEN5Fkz568NB8eZcZZcy5
XN+d9MNVcTVcVOPLVkrdJl4ybzbMTym9urmiqbscSJhIFgPZFLoSUdCnnUZbdAJGG/5MqBZFDqEd
A4gZbCTjcXfk92tilQvJfLi3/OYNmOc1O9BocDdNJ5b873ZA2Ggc4Sf5wzEUEu2lmjWIlkt8zRph
REJr2Pyccx9jtvdNJTSBTCS1HxNJcu4SeVshOLEZEFJZKm9jvL4FljiVmWAZUqZywEUzTvv5Sonf
jkG9SPwppdEyeH4vd1hrculXk87PEZaPiEQrXGbLQPdDX2S0kbAfPlGWUu+dTM4WZdAx4wQ52M9S
M4WEQEbV3H8QvfKZqKjmwiyJeB4VqZIQ1cQeU8cslAZdbe48XmkJVYavEu9OlNgb0VCYPu240Q1G
VFNTfS9wcaPpohs0R16Cg1WDVr2dEffsyxA0zoR3NR+OcRdkjgseM5q9oKjN+kr1SECHARk/NFHg
/MgX60XpBMFsmNRPKlDomnmT6IEYB1WvbdZ/sgH+L+IEDVmfythrY7/z1Z0MfKe9l1znYwg0Jxoo
9jKCGNZOu04ZjOvVXz1KChy2H/vHRK+Dkybhl3yp1DNGphHW/a1/nOAGxrSyDOi6upQnSQuwM3JT
zx/M3wiGZTj8NqdhP9q+opSgud//nDOlDtVBriWgLBsT2e5qRChL3WfNyRRZpWpJEbpDXURjlr5n
sxBlnWdXGaiRTW4FhQo556MjQd8Cxdn/l2K0ZSHnR3uGmA7nH29JXPFO4XuLnPTi3PX8fvty0mJQ
lTBH2rMjX2vJQJvG2kLrveb2FvLn7ANVY2s/a8UyGFaKME/huVcOJNJ6DkSN0s2IKeJQcxxwVUrx
k1ZghogLKyMD700uAe8JJ7J48SZSTWHQyPwhm0WwkNs13+Ag3z4VlrfNzVy5EoSm3eLpJzVVDNRV
XdogcY1PeEMZv6F49qlWe1bfnBT88gFbTrNHX9qD/hN4/r1KgSqhwMUoEm4gtWYxSppvZUCWj3kr
ZqpjGa8VqrIrX2sYD+QaiOMXHrhu5IEhAWx3CP1r3RNgRuZFB+mbs7otiyGB92OjT31+bX2kEJyp
AF95esZ3+hsxwmLwVSJWk4XfwU+/7bDsrN4AA0qM5Pi8SVDiTFJzHxQoyhYIu3m57pb4WFLfUraf
6MxWaB39+jgmLuk3UUAQb1OjAqyTC8It5rhLDNyX+9t7Ex+XKUD0qc/fOTr7By+pzlXpdiimwHXX
2qJ3Z8ZZ0aVgDKblEgDOeW/tagjt4enzuYAIres+eYuzGmEuGjqq+W1CAelqqXiQKpzQy3i9nUte
T62sMlIfFufiqGgKlTg7hDoh0GvmFUzrmDrwHsYdtRq0iZJ3IV/hhHnig3JKDGaUtJ2ln4Oex6p4
txFM6Gi1eE0elardmECHdUymjdNvhHaOpFg0n64gEk1WjFqHLratJbxuFa0+H8iO9br6QZLjxvdO
su5WrYKfWzzyFmU0OFnMeT++/J49AwTQnwo2P9pJu+aWsnLN7Kuuw3bBFyvWIWWHyiupoMKAyHmz
HuGBRyreRT0qi7wh/qV4wBhgYNC8rtU5kfjrroCanCMkLEB1SKCJzBzzgcO23lS/NiDcoxagkHz2
Q9kcgU0WDJCn0/mv+dWpjxJYufxlmy1bnU9a/c+t98xlmXkbQD7KCbXOpf1y0WJeuPfTAG1MIHPm
9bTMZuXjxVNmTTGm+gIUDfAL3FDDh6VmcPt7uTdgoajgJ1x16OXS/KqdwMoWO/Do0IRNH+xFC/8O
sXKJmzNBtzPYHJRIQtzrAY3mc826fo7mEGqOykuLWS9aIJaTSl2mXmwh/dqG2xE20dnaz0mUZbbr
TXKawrbwV7nbH3f96Q+1Djfk6ntaqekmSMwLoP/aPLYFfbXmo2k8IfYoWn5ZWC4wQqdBRiG1TIyD
jV6ce+w5vWLJCd4rKKveAvD6k7M/h7uom2U8J5Qh8ynTtJyqjBAHYuyufOKeZCTpu2KLP5bQeLBz
dW8Q36Lbdi6+063jFoFaztZ/EyXFUt2JnObc1tGdxH8fQiTgvr/v3feiV6586AfEE29UiIbRaLp1
YYA9NhdhNPfgawH2qHV4VV7BgyiWzFOSZhnATunWJZtlgMVQn6bxT6/UZ4TL0gs5McuZLeRdsd8o
xa+fL5VaczVJSROh2dO3RifP989Vbv6nczy14ERh32T/WX90WtX8UzHaurB3dWHxeFQTOzYJlBkA
60dsWdwfXHDz6eWMDc0LPgUfRJqnq3GzNqzRu978tl95tCzZhwPBbJpYp33/ZULIekZZsCI4Ieh0
jlf7h5a5k38r5i9XBXHNZ3x7dFW0fh3DqW7s91Z1oYrOOcpYsLSl8Vy+LqTF+u5FiSZo8ONcnVY1
OC+LWABem4OVW0J2PwWo9N0q0ioLHoT+oyQPr1OSEYFkVUYXE2WDyBipqLaqZUdARsy+yx8AuVj3
rO49vxx672fUYUAwmvTwl3gXfn+7ob5mNMMPfxXQ5YD/Y2vlyBbrjdXLwyVKlnTaI6j8Coxue4K1
nwLRWA3Y7oHosyeupM256iFRPKjYus6jOwMLLMGkiOoWlJprdxwQGPDrBjwzj1dbEahFreQGTBiz
feC6JD2475QnveCEh9pmVyPt8KFQDn9TrzR/UcrMmBEa3X/NG1cpcOowWP8SnvX8X9z9Yo6HcrEF
kzUhTqRzLzqUHcmooCGl3ch0+G143ciSvsU+dtSgagsACk5a2HwsnqEFCQIJNOfEpKYJVF46C1iY
Y4V3sAzaiYgUT8w8YQ99whBjeykIGjF2mtQrVvlGCSEhnBnng0eNIbxUAS+1xphX9Q++AQ1+j1Gi
0pBKZCJtwCJsh7j1S6UzdamVz/vPHVJ3NJGS8zhB0evJ0G5CUyCtoA3MW2kONTqH0sUp7kvTSBIK
/B0biw6I5Z9shEQETAAgrUgXi8D7RB5cUakP81wSG1rz6tvBKr+2JGgoZPS8vF/CqK4htQAOVZam
MLkPdWHt+QXmG1K+m+HlDPIA+wDPa+qB3fyYgTdtl2y+iBnxtyI4R7C9+kvoyQXG0CHcZrTmZ1DY
uGtHhGwvwf6zbIKZf+UVDgqiX4Xf2U6E7ryF3y1RNPNI6NquFFJKsDKF3kHd7eGPqo06+veMxA4O
vR/4zoPQSdZ4melCgzqNHjWTTHjmkdP24pqGqQx3xHVdeReb72ibnOqp9PALsqKoFy9tdsVCfYLs
jMKdtp4mE3XYrshrpwR5jq0eMzdTj4Tklsw512s3Ux70R4QFit0tGKtzJ8UqXIQhTWeS0SROG8nv
0zbEVHR6ka94NhFAdXDPf6HZ4ULAUM6P3QysjHk+N2Wew0+uzePkfdkHKkX5etBIMU0zCWehac0B
1HJJy9iAilWoC53dUvwGyfZV6ALf84A4eOk/yUZU52aeRzcWSIK/KG0wOfW6cS9AtAMVoSXTaAB5
nTMZ4eC1xR/5wp8xPqj1mvK3h0pCj0CHGcQ1EVCwskwwUDOsKD7Q/r1t9YU2UtvcwsUAo5gTVsi7
ydJHmRDBHEiW+VfxAwF5Yb/UQHmF/QnmIMeCwc9gSIUvxungmPfb1bdnqEJ5PwzPgCrK+ad2KbEu
G1aS9cyanuBblW/OX9XKbBH9fKD44cmOM26qhG9rfb+4GzpCdV+k4XjjdKF4CXpq7lep0aNkXpwa
5TwV+/FAYW/aiH0yxu8qyMiii6puRzuj0rHI6YnCkH+0ewyp403VUThL0AXdw3B7Ey+wT1VvWdEC
6PBuLkOzvgwSLELVtOegSzHyh2qGCR0E7WX3R5ZVjQmyq6RF2AfExzhWulX619RJ6B5NswAjHVsX
1Ws9xtSdr9Ptq5QNLUmRGtUgdgOULeCX9a8QAl+uHde8NPEpuGfG1KBLC9HKefTrV6x3HKfUfxRd
y+zboJced+0iJHuv1YY859PF6lf/z+Y3WLbF2Hf12TdyAtBYOE1MT1icSU9xdQD1aqmTnBAyF1tp
8gVbDOAs1GoaW6+5/aZyiQTauGTy8yaY4tUp8R5dmNxRx3VAoKgYYYPTi8nRcGfNXnHDt4AKe81h
pulbfhVKforS8sLrq2qDfRqOPh+KfcOaWcvcijBtyjbG4+rwjwh2tGQ4lZp6L3TOBruJ81REbJ0S
0zBYBKI5iOzYTRg8yUUtE1iOVRY7vxEGuEsvKILXgMFgheW1OSsCiVkDXUdpxGRVLIe+h9DlRcmV
XtuxnGZfkkvHpAPL3PIxQ0Vng7Hu/OqTNsSHCC8TD8I/mJbvLZySewj8f2+7d3Jfc4WhlHQRqmqw
4e9+EEqf+ZMKMsm8QLRiya2JA1XspxeLjQjAw/ThgD+SmOEtVI0vCBlXHb9GdRFY1BTLjU9yxgaU
sRdKgb7jkX4tuSV6qGlUSG3wo9h7i/72cn+Km+w8UkKHQa9kO/Psb2CWlSbTvhuvddd5Pqdcx5FV
iBtOvGjM36Wrz4dAKl2u6mdEt+DAUNZZiJvZQb56sIM2lmDSQT4NhTRi209PU+bJmOw63rEw4Qzm
85boypXKQFNx/hq+V3iwk7zbsv8y8N+QA0JdQHaA9LryrUyB1eBUFvpdZHvkP4K21S8EcJ9Rd6u2
IKmsQrK4PKZsgENetQXqreMM4aLx6eLNsKKXtw0PMNrQjiexeTt5MyHidXmlslZk7R/JVg4SMlkS
Z1UWDAl9Ifpg3mj93WI3Cs5jwFE5tQEzEt8O9tKA5kzFbC+e3lr7YQwBkFakf0RkJ3nCykYrDTsA
ceHfoktrdK1H9NnPzGlNzQMa1dWhIigHNoi2bMhN/g4zFskU49DopGXWNx6OPUcztGBk4sqeS9IR
gzw0IMh/u+8UHthxioTZZ56kkOaW17ogkkcJ+JgjVzmUvyGhxXSfpbOzmPt8byFIfvQd3gira9+K
Mu5nASN1lVKhUa6urk0xIUQJYUddGxGA3mdsmG7hM6MsH1jekdaG2n6HWDIQdGWPMBKebz59OtAs
Ux1wgPV4YYsa5I/5k6T799X983R8Sf5AJCoaela6qqVG+k1djm6qYfbV0zPBDDmgKBMAtcbE8CAa
GTLswB5sOWUcKYzo+Zmx3vZZ6edWPsBbW/krJb7B6yPlt5osrWubMF/XAidvPdMauhS3W5Qp519T
I+G4uKcJqCT8eWe0uDTEOhd08oOR4a/TYslunSJssR5K8+l0pIzGcT+LGqnRPFaQ9prELI31RZiy
NWV9vXcqF8j5kD5riaQvXYHl7cgCmv1HYP57oxbosDjqiTpftKiLwXn2CrrFf7zhOJElBa01PLDS
we6ef3SLbndiphDdeKWnyzKntL1CLZyWhTFDjTe4y89qXVYGnZhRzti07Nw1xkc4Jp7tsOjMqip6
kX2qKovb4fKgR3Gd985ejQ2Zg7++CVKtTXgQ8nlgt0/1ScdXg86Bagq2wxUC06UREjz9Setc87p6
/4358RcKj/ZYz+s4IQJfi712xGQrC2PC51ltcunMpSf4/Y+YAM9EAwcv11crp0WfC5X99ql70VcJ
b/dA0qzxE4wm9MwFVpqDRlnesTC2MkNZ8lm/reKuiLClG2/YzCYRH8t+HvMB/CpcR2xC40EcbyoR
XDpD4IA0BfzeQ3PRhFhPmAoUe9q/ocMwhDsW4L8UpEHCqjWAJk10ouWsqIbD0RGRoownc8nwh5nF
5HecSCld1VwTD4lynRC5vHUKAbHJwgk+Q8GyN7uYtE3XnvhAicOPJkvTDJzQ24VwajnVDCkbGrLR
oEsfMJKwMDFiaik+B1Vrc6qFVi7U0jGqmOuaTZMvKaMvRu9AA8w/jfo/2DbWCyYmTwH9DwD4oYnM
8P73djn8uFwM3VKCA+oOaDFYCctivYYpbMEi5ZDcLMDDPig2zmkUF0rOImK0ahIwZ5lwZYAv3X3F
/7YdAMhw2egG+yUMSNMVfhGCG7HtRsSv3uW5M6lUmrtm9Q3qgs/looPhAhEuWfJC6/s49F+FTo1f
KMrBNOg3TGo1rXdzgvAAg0gIUFbYUDXaCxs4QtZbsuW8D29NHFeVnhHQq9q5273e2geSI3JM2aR1
8hPCp+WhVAn0eIeFz/5RtMdt5MaFM7+C4SQFHv3uW6RTtrjJKB1tILXTjHy0uJ0OPcnCwWA5NBTY
RNQPzdtsytfx7Sm4HRRlxz+8gJsofLUBXl04Qkzty4jrLlXXpNxR4o2giJW+NN9huw9A2witnCG+
A9pp3qo/DVhrnsHboWcHIRSjjrOn8At4sSG7GznWctpP0vZUFI9Mr1nI4HWdupvqv3qAV/ql+dMw
OM1UAtCmvNkgI92p9NxaQCd7o5lLJPXz5dBzAzA6PTok2GOXYNXETylj22z4V7JAIE1QwLXRsiHX
CRJSUg9ygtEGyWQV6NnGORm5uzJyaHa3DY5fehhDUsZV6d5cC0t4g/42252D3ezt9LmSi9Gx/V3H
6hjp4LdapY594Te1Z5Hd60ClIiQKyUPwpwD7/UyjsGZzH3j57W+kgRKXAZC/TbFDKhqJ4XDjcPx8
Z+9Na/A4I3l9MSlK/JFaMQI7J7rJoSN6BLeiubaicxsWBsvZib42YKi+qDpbl3U9trEKB6LkAZ1A
yehr7lBPM75vz9u1GEk2unDqN+vFf1vQb4FlSWBGWEPmKvA2g+fUqMb6TOFu8yDPs3mZ0sYH/Lvy
rHgZRTRLIJz9tyNgLzfX6v9M8sy/5BVCuHhALdgqw9ZXoIcIT+iZgAG+9depcssPQ3J0Ij/d0hCW
nrARIZyuSa2meMI4n9lbk81/qc1vYWcj/qBakBu+SbKlgp/Yft7rsDsJgVakZuPDcpUn8Y0IM23k
y/n1yPeK5+W5UEunfKw8OauhK6vsx+ihZl4Ii1KPwBSuVWhLpOC9OIbo0DZPCPYxxDkLdi6HTI9s
OCpmEw4X4g1K3jPOcwIJHHcp6arpXSwZb/Pvvj2dgUZ1Ujnx/4tKqQrrXZxTgwWx6slSbJfF4OzI
bwrQspitb/WOVkKBQvZsMrDy1pPY7Hefa0frizk7pGpDLc1M75jZxgGqq8WKLdArv9YBP4knTMhn
OHIk1EMzLtQyvop636FgbDl8Y9RPE5qv6LaRb+7+lXxT2/Y0BEeAHLNtBqLz34tD6QHFvGP/Zfum
d7N0ZnRRKcFzPA3TQ9Js/IpoLesqrn4kVt/UuSTBj3iYzBjn/ZXdg8o+MaxMCXUj4OBC6KxH7xCI
zWe/whZTvXpCjEDNxi+/nfBnk5+vrcx2oozdkA/Aia+AXAbGooHHYd3emurlDUv2BPml4eh/Pnpn
YkTuiJRP6zQMG2hcXH2MFVAc8Vo7c2K1A5ZmpOq10zhO2wxHvY/Sa+GHm7w+YRVyO0VqFKf11OhP
pJ5f3zhdVrB95KBuXx3EoUNkvrygfznIkbFhQNKIG1hn1KHtwetMEOttWDWYargu9ODE1gsrBFb4
NddL+h1OL1Wo4nWf63jZWF1SdGar6TwvW8rTbJAr6nQo4MY83ZVj/x/WL3ciUusM56BPidH1G1DD
nX6wBJ+p99AXoEOCS+IcSX9o3raoZ7nJ1Ex/plzf4KYlbwMBPb3yPl2uG+xn+rEFWH1Y4knWTof+
7yCHLV3fTGC+9UUm68WCOpICd2R7mZMIZVAH99ZlZgM2AFCJMwBE+cZAYoea7wMWAyBRzGBsXmwN
xplYJzNKkzbLR6mZ+6S4VEMyBanGt23MHi+7GfbH06hhsa85Pq0VLjJv9CM+xaHuUj2h4YW88iZo
lhn38tM0MPO7cZw8+qqgY1GmQHSnVlR6CaRXUKRFVLtNjpvIVstyEZfpAWtkH1YmhaiuS55kNxAI
IGHX2kUiUW8rpBWFIqM4FPSj+E47Zw1yrz9KwNXmdSweKYlciy+pRJIDVYxjUMUlr2+HvETlM2XF
VPWihqsnGd2iFMSIngUr4rQ10QEmLlF46zZ/fxzdwT3uaqs8g8S7ADaI2SKB1TF1L4/PTB/cgqxL
8tjUAR/cVF0myNMD8/0GSwfQ7sQd6iVKwIncb2OUNXy87JzNhShAXg/ecpbukbsJH0FNe5fqUKAp
Uz2tJfNWpE4Ojhd85we4nQsuZ/2jbM9XevUScYq4hTCH7QVID4WHvAePfqmijR/xKVJYGD1WfyrH
TN/doAYt5jiow/ebwdHBmkOarz0kWYpFeB8gqdKu6YaDeSXyEiVTS/Rb8NMcyBbLJ43hxMQds1jN
cYJUGTZMNhhgYrAI1pLhTVPDjFoMiAW7vRPcxUynCQClnXH31bfuuM6uhvKAu+El9kTyNImDCWnH
l7r8e6D+Vpvg3QQhdDAHsGEiV19+3d0U8Q5SAuHr53T0OnrATwPKzYNTalP9nzrQ0PQTWKdmirO6
V5/9ofVThA7bDJK64+m6DQv3WOfTu8YyW/T82wxLtiU3p1lHPNvBMlgMg2nmkJ0ct+Efrlsf3oCc
9Aes7Cx3ngQIKMrt/4voCu9Y2x3CcCAae3wTbc05o5+Y/cq+4RTN4GguCisoQ7e5GIoxZtPn1qo8
uNWeT53eF0/hLgMJZ5uWjcUgCuC9iafg7QmBEff8drwzI7d8bs8sLhW9a1mVaE5EnofU+vJ9ccLS
eWmVXWwW7n0nuRPNqrglAZX3RJ9HLkhcgQAa6L0/ewEQ8b12J5NvrWyV1jMMKbRdCw0NWAEVEaU5
funcWwGnwlifrzfp9qRnN28aRsgs31VzR/xcE7Vrgw6rxnHZen+Lp/NkgSmTorBUoBei+tsdyGSe
eJ2RYJm02vlFGgjg1mX1GVjxW6sGVQ9OkXJue+76fbTcDjm+UmwYpnOUspPlvRvqKuET8aKTlwm/
KNvye04C4l+KGlwgCEIfKRHh7OGGEqj9pBrcdZ4tJJ5xIo4bHeo/1CJ9sTfjjPDBZFph3pL4aRtD
O9huiy9EWS3l9eZRZxGs13OVllLq/RegyJ32sb4oi+FGSqu5bGtSC5oOrchmyY9w8SHYyn23zoGE
h3VXHYlqVPgq0klYvMzJeu3UyvZUq+Bf/kWKVo1OSdpZ2+6PJrDP2W6gLilvRS4ieT4TYRyyMs2v
+iAj3EgiI9b6EWnsA3ayk4KgmmurynBieDDpXqKgC3LnNbat3tC0Z0qqBSwmQYvf11pelITKAUHl
FpAdRMdJMUvb+CgISRpYWP7qsCNEwradwMN87Lvox6Ju3HHjRofqxp7+paAdR1sywPBNBWN5jvq3
8PADKYTddOqjQMw2AMz0NHnWpIWA9mKLEZIXCzaI7Hq9WCYvOTqGFPR/1nzgpz2jOaJDlsDM3kjz
bvpMCwJonc2jhs0Wlc/UTWY76e9symU8+waTrfyqXUBuLXIa4B2HWZR+akasd7HU/WwLFaJnqhaa
2hU4gYxHNxmJF1FQep/df9adufbn5PE4tjDzael+qeA9EZYxv9Pk47DLUNcbx5GK5JzTn3zUUWM0
wmQPwKP7pyKOm0tzw4kBMy7tOtvd0Il84HsB7gMP3mNHwfsfN1fIa08BGL6vUR6gBjgP4YtOBV3o
LWFt/xXV1oRzKQv4yi6WdIwmjXlDlx9zZSeH/tmdoyS/FV/7k4kgbrizle9Kks0RPKdL+1leCAet
oWsJB2zgY4vvos2kEoOqKwYGO8NV8IAstUdTir/hPHsrz7xNiZCjKfuV651QFqmMCJ/wDNh2rVBL
BKCqk/MTOeVc/01PsCXslpR8e9RyQRYMWm0e5FbjSbXtaS6p4hYQkmV3CQqg+D1xdnkOMNxzruOq
2K9WkKi3P8p0fjT3lGIbrbdK5TqKtjOO00xmvnFy5hnsn9JoHx8xAHt7ti5sM4FbmRx7oy38R1Gv
iHxcK5ygdwzziPgGTt/89s8GVCjvpNbuYWI4jOIlhOenhFd89QBB8Q2sqUoHNJ9ybw7AGSp9cMVY
Ih6fhkTxtkZM6Q2qXGWqgoJVognsWKYPgEE2pZVtKgEWjkJL4z0ri5dBg5R3kp6oLI89JqWWOwPW
8YA9PEibaOFycv62n/iRQ3yBgNtAKHbY99diMVyRf8j69qAK6Sdh7nE9cCjthz3/CmvtLKzAU9TS
Qp4p7WoqcrUE50X+aLCeCgESsggwYTWK6OoUGkXm2QPpLjbC+SKZxx3ezicBVTimzYn7L9Skwuwy
3zLlUteWgwwVV+jybu//yaWJs0cPyw7xPfOUS2xaqbukACV1xTRRshcHL3LdRHGh2T3CtqDuNYdW
qv2DXlbI5CyWcypfpxpcSL36AqvlA/o54rMtXTurFEbxu2uy33XZAfNRmYOZq0nW5OGr8Z1aGSV8
Htx6JrOEWQ/vPZjNS8tN3XJHF+BmHvV9aU2YF53jXh9IkHjpFnBESHE2ZTJ5/wQQbGttrbptOnZo
9pSLR/1B8ratcCSJusx5DorbhoKtA0w6eQB9vagq63fLvzyRpcCl79/rDhg/MQBKfG8+w8KueYBa
IWPKffjL6eCJmvrLUY1Y/9T6JTDCg+6JlG8ZnzkDo2jyewgKu961drxTQwXpD/mqPyaVTmfCyrym
nsJl4v18OGepymNbwY3yrI5AlRrQUabZT0dgCvGXLrC5iFPzOeZP+bhTayOZfxi26K2MlRRMI+ki
/bTlmM4pFLP4b+23/CIKv2LWbZ5FZz6jhLPk1ASGUphxyTudyYSXLoan+W5tz/NWM/mEmgeSjSOQ
lxGT/dTAmjj9g+MykPrC4b4CyGubsxZYWnYFFQKnxqluQv9IbzWtILW/F24OMTytmY0oKrlEscqo
uGowqKUfIDaY4Z0kyFrnx13933QIBpz2J9yO5ZzmoaiWnaS31JvaQG2ilXiO78EVJwzwx8qo0Ax5
yas6Ta/oNunjqHNpQSSWHQcilYzdpDl3WouBZIFYk8RlIeZTaLhgr4UK8LLIb5Imwdo9TdMJh55i
dfvK4ZXmV5ICjqx0ocd7IqW5tntuaVQYEeze2/yV2klg/bhUXckIufcdBp9TigugkUkU9SIK2yQS
JNparezHllOZ9cUGdSJZ0WJnAKw8VLs/odKIaYLiGX45z7AFJ3M2GxQ79tCh0SD5J9iZxfbQ0nuy
Yy0rep901tH45hwUiOBJxcl6fysq32aycion85oEi8hlbnKstI/XO6miGDqOJyA0bBiqcXVV3ldH
bT4v99Nt/KUleUmLuUndHVJ70+F6JslvY091d1gGeNUzshvmzKcq5qJPFmYWwbxOWrc+4mFW1FwT
KDqDVL+IIXxG65FF61KIXibgn79qKMQfaGm/3jafsXTXRxFuxpQu64wWvQorB7/nfLj8sw9KUYbS
vkDZFCVs0wNud2QdROPID52itd9KGajt+7DeJYY1INQFVn5wI2Ff6TnlhIuZmKtTOY65Cx3UFeFa
8Ccx9ueGuopPsG1Uoe9sbTtKgmJ22BnkDS1H10Ykk0UG6JatB4BhMhcjxrw11kuTv/zL7CsL1aUG
eoH6u/QQJO+nFrZe53RwHrtyAp/9cTG5J2XALWRrAqg5Rst2WhspXzG/M2ioXVRxM/Kxo5rB1nLD
k8xRxY2a7kdyZo1BVR84EqzSnSXpz77sxK2AP2y9zludOiLM+2GNjWlcAyAfbPr17tDoGDSdxcSF
6orjnih26neYs+vBBylHg1W6Dds7VhacvDSNca41deiLNRY3gN3jNyy6XvDsF3RVMs0Lw131ByIs
gu7PKypFRRvUhsS2Eq5/VWEG5WkafANrpPXohpWQrvvybFNrmVxZzSDDAgCnPPEY/62U4lnnm5BX
N1XEk3cpxaR4Y6DjeCNomXRQY0WjQ/jlYkBj+xLvEMlUE4hrNmruXxQUeJzRokWzhA+fTSkhhhYL
+OfQ6I9IWGwsZoNrodyctE2n1jTbxuoi14H/WlCJJE+jwUcTJhq9M7IO+2Nd4NrYH3JCuDfW9ESG
dTUBlKcstMdMxiZYeiKuTk+fmQAlFNETXUPj2oLRmxx37jvsCVI+/iDfclSL84LXL0YpZThejsy7
dAJqW8ge1LTzWRJXDxIqbwzPDDV7BN36jikNxgMjUFSQqkVhX1qzsvYtuVQU+mF41g2sszGP8EwV
RfbzWlcSg70UQJCXijRym3UEu8ZXsI0yXu5c2xnD6YxF9TVheVX0rrP2PHJOLx+t9z5EeB7Eu9LD
Y71XP0oTnPBwgRQIWmFfseEmhNSbXIEEPxJuTcJTk0AX8mAHTCo7PtIfpfLWrsi6hF5WVMNziSJo
srqC0BLHJDYq9I1ZqMfmMYDqo/e9fUtrdPHlEGtQ+oD7Jxy0ZNWp6awC1s/anOYDD/pMBLgg6iY3
Zo3oJIh+vzzev9p+FOVF9CTKKdoXVNdrr9uVXQYCM8vZu2lV0R6hOtY7DhS28k5b2UDfbvG4mXOr
LhL0N2auVwxv2yQEGdpLckv7E8hnIkPmFuLGF8ufbmibjs4lJ2GMadkwqsReprEW8zhTBnIh3QsH
O9pNgscO0fUcEht7DH4J5ErsWAYDHD+4tF1tkaG45fIAmxuqlAarFkgbGVFrDXKxNvhx8MqqBu5J
wTrRxouDOk1o81e6eVh8+WrC/psPth2RJ67yvTze/X5R8mg2PpgBNKj7C5BmjmYpL4Sb8XlYBZbR
iq1I+huptxz+NHnbreofTRyLz7my8W2rNWUxsTS4PQZYryFG5DVwXynHoSS92VHSIhHPw5POtgH0
GLdEK2mskaVBhz/acO0zLFhdslV6lVsRwd9TktgzC0FvqZuUAZoUM816asrukt78o9iuxNkAjCPg
ioXQI4CB1sAeZSJAEa5cLVY9+M40aUoD9jMywQE+lKC/BP29l/jOj6ZIuOQyMwuFFtB/FhSLH0hJ
sT0BeZDetjhR+8DRFFw6KP+2KggN41TotKwaavPPkbD3JrF+DJFTVtzIyW6/XWO/xYKaDhaa6h2K
C4isd2wOiaG8VRHwJ0TAgWL1QtXaQ4AmSULSO3ErWGe8/zxO3OEkGN9o6Jia7Q7L3gv7/RciYJ9O
wsf6uHkNfx2yiQ8Siaam/YVSJqYOMtHuVjWpL/Qsj5DjNGUJF4rYvD5+H3HNkLR02HwalBHIQ4IB
c+uqxDwq9AfD/yloVe93osM0czgvLJA1oE2Q/3G4ri5JMkbdvk99LqIGUtjB2gI+mu8z/joZhi+H
EBVySZrd1Oec8/wj+UAuqcwAPgddy9VEO9ypGY88jTRXCiirNECduLN6SnSEO4LUmCceSma7nYDJ
/LYnCatTjJEXAxrPZBL9gwnM0W9gohZMWT/+Ub7cBDSi1k6ZO6gMZ9hgTKP8qU90Xl3o1XmlrzIQ
U0Cd/anQttE1ppe74WRy5/nj2g37jtzFvkve4AZJ7VTWlv5VDj0GXfDGzRU61cpZL3CBJP0BjPe0
RkY25KPXoawkzprqB4nxuz0Gf631B3BcNRBpOji+GdI10aTfVXsHHKbh8juXKvNMkQVBYL79eQQU
zVw6GPXPYq3NF0PlQ03ucRnwFbRJBxf9ACJKcbkTl7Cx4BIVq5rcj8kkY5nEesNZ+XIRbCCmiD3t
l++BVC/exds/fH6PU0ckqkfIG47nO0kHKoqjWNxx+W2s6fqZzMtBG3G9AtK9HMBdRe7l2WRd7/rm
gkmjMmzOWdAgSB+Ubu0sWFUZj79kCIOvd9u2GtdcqTdthCxfjPi6vXzd5qnnNnhq4K6NXaeAzbhe
l7c2XL7hKuRr/OsoVSNbakXHXjb1GE2gyVovRLt5gJSkL8LWRecR9xX0qehddIHBJj/IntBB7woE
GVcbazAdI1ML78drcvfYV3cYBiVsrLxtBhaVEtMZLGiARq487YTq8+Yb3g3Y+lWEsqFfgIeY8qHF
2Du61dgCuqC4yfUjY3JloD+Um6Z7AEuM97kKz5l//6AF2IJWh28mCf4X7u8LWPL+lxO0U+FkO46R
sv4iLBqhueJFv+VVS2E+AWYMlpesHuyKC4r4b1gh6aTY+sf2CnbUQCyloGu+WsXl5AZ6qJOnVzFD
hQYiXqURSAxzM114G2OpFmBgEy1rehAt37xZlk01MDIU9H9h6sS5s3UHoO+BjpyS6SN19U+IcLca
HNeVB1SyEpX6QzGgRTM1DYddAniESRHe6tQlq4Uo0y47sptTHFBUHFoyaMPGFfZs2LslvfD4vpid
HLhAkdcZRCh2D7YxFZlUXicdujNHH2R5GPqzKlj+1nCDVkcsnhW8J5WLpzJgmkgx7ahcGH+sPInd
5LEw+eDIUs+dtImxU5E0RI8fzbe71F1HkHgpOjbBHvPD2ma6z3Er4wxXvl1c8biogysr/8hjArxJ
Qa305ITt/2V/DAX8NDsKMlNuxzlfG/HuYrAeuXjVntpctCtNgtgWN7zJi4VBTpCWE1ep7VIShPeQ
+CNb730q+yf44j1VjqxEROlD8ln6pxMHNitTduSkGkG8P7mmXFVET3L7IMbT0er16NOUqr2bzpBR
nO53d6Pu0FmHsx7Pjf2miNAXHT/ZbnsugySK618cAChozV7JW6esQKY+kNU3YKYlEryFp//YvL+z
UaEG+WaD/6CCSrYQ2nt8TvU2ICcmea24OLhcQpXWnQsnbKkfQjQtC28oRzALy0+weUtjyDETitMJ
xMVATmjZ8zxRhpUeSMq03bAMqx/wmWAVxGoic/H3H/WL+WwNKxbiOQ9dCZj4t8hln2qCNxXc4D17
okYC0ZyacX2m351yemXYVdrp2v7MlxG8zOWFVGKU0VAIDVks60PlpM+sYFs5lYXjjYFjTiEsLj23
my8Z4xEqnJBipb//NNww99KnnYyBDvJe5g9FteJKLrmYixNXKj0cj5zsGfBeSxyffahb13pKX+VG
sN+Fp+GVtA1pT14qCAmlVixEPpGRQrDgbenrmjpgno6kz84p6qgk2On1rYZ1UIp86vNZaiRte5Hq
z4BChRyQFkpm1eRgiNwygN0W/17UanxmIVJXvnJokN/7CkA+LISFdKZjPG7Ujp47Jznvaa6klrm2
GUA1CWq3YRNLN37BPuQiZ0dgitOihSuBopjVXqKyzxzCfuL76pkO0AuI1AwZQom172gOwz+t/veL
oZxeNnFGYwwDyMhY+pLMJZyq2nIEhHRk/OF09KswW/j8++5ykYLf240wD9RwH7Q3Afcip2OjgDve
eg5nGdV4+uA9eNl3pIgmRta+cIASGcVuYGxlcjRz8XKbwZzMbq7Ha/BlreoVzH7r0/J/HzYXd62K
sY1r2DFzuaQ5Nd1+EKg+TE1vHddbZ8LTC6RZ3Ypu8S+vnqd38kAxRmEDbxObHU+ehFTKCT2dVUcW
4b1Z5UdXHv5AMnZNSIEcsF9z2fAhJ4tHeKd3vBI97I6KpFJLNcbHNtxprPjYu8WMEBjyoHAQ/GWu
9COi76x7jIqg6xHtVP5zALY6Uk2DdXU1bPTMRlq3/VauyjrhhYEzfErTEokQc72FdQkvGAgQ7cR1
uG85KBTVFFYXy1YeM6fU/6OTbztFaydydfVMu2t1ykwYq87fTZ/xNo3/vnQl2u6v38nr/Jc8GTHA
V2XGIm/alqjBo+ndPIFgJdTbnCaZqrm5CTwYqvRG3LtBKL4a0hWfToagAhW03/tdoY/bpOKeqqhH
37dG+6/7tzJeINcUGmiAz0l6ilTS7ZlcJV+aBZEGkIAjZamc4ZOCM4QXlLjaSPnD5IeMhOGNQcen
FVh0OUE0Kj3C2puq/vNfBZPRJFYfQYL/FcDxUsH5+GcfR9063Bd4hY1/JAUMZDNXgwPSTei90528
9tpDnNHj190bmy7KJ8iy6CGbYXYGfIhTD+R/4VKAw+sOruXM25q5+/R0oyNjh022nY5NIM/6dyWK
/sq95BWHuqJC3a0+In8wSEAlmuS1Twwqh2U6HAlTmOWYSa3talCYEiEbVISTuj1IvjryVXhqz2Ew
y2N1g1I/WnqTnbsKhTjPUoggRjECmd4JFRlDUSDZtfgSBtcmR15u4jj8pg5gl7paaVR/lHdiMBEt
whejJe3MUbGcShuxOqYe9iFBNP2noOgfAVB3J9j4HKPZdnAXhRreL08PJ+oDJIyv/spsAwFxUjSz
b081NOaybPuCayepkGISZHYZ4vtm5Lw0OA0PA1ZgCZbhKXOfSkQtKexNohaCSNUnjE4hytOcA9eH
UP6JZRStCJfSsLIdG19mgg1vZF0nL9V0LMd2v8W8ly6BlrSNK86rdlEMz9T5Hz2HfbsKO56jEqoo
TWRDRjNrf0c14hz8CtEjcDgFGRqaW7hvpq5B9RvSY2dG0tNqqmpnBO+mchgNIFcvjw/E3zfKYUio
MYjBp47eOG9Jp0SlSmGYRbVXEL7c43iuTz8jhIrZxUIkaUIWPtQQ5ezvSNogeQyeqptfo8Ufs9do
c2D84aK6xMzK0N0jQbkn1cUjNtEEhBtwwTEDK7iPYXWDBHVKoebtWqXDaRw8xjidaBwHxn22IGvR
OrnnUn/qomAfkXkj5MAbNYduG1sRpLt/C64YZSgZ9MinDWG/k1eewoygpiisUVp3N5P+r6IpJF1/
8xIeI+a4UNMKUET81tfeoeAM1+0X1XstZ9pqFcZE58edzzj5B/FxZtweZJ+HkrGnkpBj12FVLWjT
rr+mKkZFAFkwIMCcqg0fJ34f3qZDRvKN3A==
`protect end_protected
