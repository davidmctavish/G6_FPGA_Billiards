`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oPKtzbrQOC07sGQ/iTGWF7Oky4sqVzhMNRdZ8uHNcK6vhYwVWtlPlAcyT7aCNgtijuoTjX4kL2Wz
aXXFLzGBUQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bKOLvlVmB9/NRzucKbQlgVqx+iVYlI+7l+zgJJ29pdUZaDUYLUmFoB4jAroiJdaV9WfgS+V/YukK
56kBzr4YbvaixfIG9HNLYSzi3czAt6rCIOzCCqYFLpOA8nUeVXUFmRing2DDDhVl1CMAHSbQq3hc
9iBIhz7Ml7VtV+zUCiM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
op3Wb0Nqzvc2I9dzCJ/SJxs2kQGosXJSaMfd1QcF6jVI/9i0fOW5gh+gJ3dsENDZS+X9FDWkllB1
ieP8OlvCUE+mkqMr56Md05VH6pd1uwX0lY7CeOj5HtBRX6rqTxW1l8XpVZlW6CbywoAYv3UZYhz0
SUiePBP9/BsGcjSTFl0RXmAwVn/pTt4SkhfKq4U/DCu5kXT+KNfbyhwsl8weev3pgm/oV/8oX55I
TTpGpTh9yq2hb2GkJBAwULvT9KcLA7PhdfUkFAi99jgh1XXIPBwiGMAkwqOBQF7zTn8a9b2tKCMC
WiNth6JawKF6usmPkpAk3iG2teAUsSGICLdYIA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k99fUYUJWNQ26iTesoaEAGjGVV7mbQ0N0PputyIo5T0wQA9qvndBGPmv9mZHaIEgrMe8hE9IP9AF
VXNKYGRQkGmOZ56PE9LXUkRD9Z1leKjAuK6QAP/9phYilO08gzRcPXEMzy6IUKHt14oxouBWqfxz
EVPObWByuz1xWcjva8E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jQw4aHNhLPJM1lDfzyOlfK4BtgPqJSu5/LkLDAknKFhQlr+Ie51R/fgdBNV407U40dxcXBZv8Wuo
d9EXy25MmLjJ+u7DzPLbpDjcuFUKsyg5xcBCNvV+HQyroQb7Ige3DIYCE6rEnyiWNAgQpIQUgTIh
xl9iHOs869nu/amtzzFEy0YmO+mJ6kLaDeY8smBgBw4NivSVLpzVG0XDBcoGHdrclqcvyzHJWjvI
ke8rU5ubWqe+JoFksVcNrPrQjceXHvC5SNENzACwmmu7WrT+NwiJs/OArifD5blbuUGbZDgrnikP
yxaTT55KEg0wPy6eXDaMiWxd4EGqhcOshHut4Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19952)
`protect data_block
mqJtE+0o2tUf8mKbs0CmeD5EGpUI6xE5LYvpeV6PY2rT5g5n/vXl8KNPMKHRDmrY9Kl8cy5kMcg4
kN9ywNsMT4rrR1RhSUhtCBbKWcNp27I2s4prF5CNgT9o8tGZANhR7engYwmTdcKd5tTKky6bf0K9
UF3EtsZQl/jiDFpykW3YVExRXhVw+6b8FtsM0acgz44naRJ6oWom+nomnJZF2QrcsTajvERfm+mz
Q3dMaCRAjZOzoABULsMC/+od/4u1sCuXDrB4L1i2J9qow7UgWrqAJ6P1KEbiKcNiELZG2dpv2JOS
8yok99xsmQ7JoNCS/M2bo4KrtrksccHAaGtG48kROWGckc0YkG3WWNU3jm3RX4CNELTyAy+UYPWW
3MXgFq/wf3oAeCB//FRvdbWGZCsG6UlFOjC5T0yG+5U3IZ9e9Zo7C9/ntEzMSfv40NN26U7qJe6w
XeW7wa88Lu1TaG99k4pPZfFJX5oLC6jor6mn1e6eX69uyelCBy7JXU/OABcNAVJ78a2sJsNJvr0n
ch/QnbAr7HB6m0N8Og7x27lsCDE0yghI3kiseqZS//d1yIuE/oo/azGqgAqVxYEaG0p+2S6ESGtL
SvL0iYpLAK05F5dWRjK5qflMcUXBkL6TLYLU9dIXz/+bvGtcYkUb1fPfKNMgXkd1hKzqwbvuaMdQ
V26tl4C/BfCTvJNBvOnp8btWyFehH44voU9SSzQUCCpY3bVluY8AmokiNI1uBcQ1KYxFf5nPV5E2
y2AxYcYhcXUjQ7Sob7Ie6VeZpqU/HPf7YhHg/pIZVLYUdVLQjsVTnua3AQTJw61n3+Q5Q5WG9oG3
p0jubRIZFmWFW4sP7h8NvTrBLMGCHfcWSixgt6+Drtts6C4pX30I7TtNC+qBZs8uqFMrhxs3fhW8
+r29goxoLamPfHFJTsmKQ/emx7VYNrAjwvMRjrw6Q502XTD66Cp8TibuZ9ZTjabJwElDFFnAVxAR
sZmpFZnjDmXTEtJi5VvB5C+4v1WZKTUGmzC+bs+Z6WLeofrN/Dc4yOmhlUbIj4EyYBfHzq29FeF6
WXyjFL6UoqqmbOlUR7SKj3D23XjmoxCULvKUyiHxAsG6ygNERbK5hY07r/7KMfttAFbcfLX9bG8E
Ejh2cc/63bBLMfUKHVEdKZA36NgY8r3Kxk3mjYxSjcdBJhkeRNxfVS4O5B95D840Mk1gSjYQ4ZSN
61M8hZKkhN/x4TG/ficL1S34so3v6emubTyDFA2BVTCU7uVubW+urzWxckZZcjRA0hFnvTxK8k+g
fkBqc3E40l35ML0fxYrf7Z5sDE3ACLKfyZsD7caQknawI9CF0OKarjoCsbxrOlaJ3T1d4UCBSwMB
gWBRFjZimk7O7BnFNfUcWCrVOde02UjZezmdHszLy1QtRMO2MvC/FEdTEl5U2v1gLae+aPj3A5yq
pWQ6BpehS5mqk+2EjLYRLAU0SEN8JESxQV3yKtoh+IoioBSYs1l2K4rx/boOyxiMo4ETZZeB4mNf
b1ZrdcWYL6/7aK6GeSAJ6k2ftq1CmZakioz7gfE9do9xVR82VO20gx8kgyDRnmJgtQg9opzezYS0
PATiNCZwyh6dI2HQ9FHBuNykEG+91AXS7y3MuOni5FclF1FxZGa4SVP5qx1+J9jmOLhyqP6bGHhX
6ToQKg7wxjw92D28qVD5UUlAalr03bloYy7lDaEnt66JWGo7gSXo5PLl73WsuAm9otA/HJ7xrBa1
eq76nxhcjua+4rbmHAEEi/gq7K7CuHKcGTeCS+DJDtmRbKWUJINPMtuNAopdfuFb6TAJ1pR/FhJy
bYcqsmhqtO7rxf/CeFP/YZhDZEsAmtUpYDFrim2hpDyMiQ10xKqLh7rouI/BfU4g6BXhlJP4eMo9
KXVTM46E4ssS7Swr0DuoqmrLEhQLvP3fKJ6uGHIyhYroKSv73IY/FvXnW+QqPbqdb8kpfydcwc5U
ciM+1YZwkCTFYiPDkTWCD/2/pXFVjJzSKJA5eucr//4J4GNSA1+TCZoMgebXV0QgrxI2ziIWBHUz
bbTUz1/7VmuJEnOQT4qHdtJJ2AZrTx5wi73QynnzC4l7l9pNSd9W8M536PS5p1UyOeOrkGwPyNgC
viKuqDxOFHU4o2oN88JQ5taQ38CrHEFLOrjau96O9WpxRI8xRglJE+UTzl+JVqKPVkxGG3EZnIcp
UuRs4AMaeRhA2X8fqaSDdvKh4sgtrCJMvYSK9tuX0Vvrspa0JcScN3hX2JNZoM+gvAKFqo4/dDWH
rzDUl3iUf9yh4qgcgi3CwtxDa8xgYvBGB+/jf6UJEtnFwm+OZQimxLdbW8ePKcKIE9Ihk8sDMq/E
GM3bzzpvy74iNszQavH+tgAnyj35fC3TDdtaxFQVTnqIOKYYckZB8P90qy8fXkD+7QX7jP4Si9YS
4Wz5T90fll9B5k9EjsMm8drtyBgTehr24EdL4iwd9ZIq7I+M7O0NXxjgS294aIkI3QiOQ5Kk1V4o
Q13pGf0/di0iHVfm6L1Yp9jva9WkZvkXWKYDEruETSIVtyYnAteMTBtTmAm3ZOdAMk83/YRRY8hk
x54NkxhdHWnINdl3PSiLC+z6RJA+DBRqcpBNCWcq83lmvP4A1+lin3k+IM5ER9QmmQMtMFqo3qsy
7ifWuSsayuCdE84a3q2VlUAkz5DYM3b08KtfZ63w3FPWh0Qb46Jemyx1sGqF9Bn1S8jFpsXximMP
54cgD6sDcXmGDR0hFtmfYXHOofyJ75R6xYENCoZmLmFPfl8zwrVjUuM//vZY7+GfPkNwtICiOwKG
to+Ha5lME0IUWy4YtEEeivrO7ApW9fPCOq4P2/iueVuyLuFA18EdJ2Fr7K09KrX0P0+x1fpVmJSk
fvhEAG4yEiKyY6ngS62UuRATpnXgY9VZr7cJgtH/foCSPNhOEO6IbA7NkVH/iBKF3JHBXBNglYRY
Wr5ptQiUFu87jtwSZWDV08LWSz542Yh4/kgAYskne1jmsIZsGfscjnoGn4qhsbnTpynxeeX30jxE
eeH+/iGgyA2S263gI+zyQWnKzAOOGYo+uGXwwiQF6ZTA81rL28yI2eDFcGgxSxJZJqEl0TGk0UG6
5NaaRcMaPyEmHSkfHjj2W0DrhJXpE2imNUXzfVy3YvzuYhptk5HL9qKmJuaCDuLxUAH5wwwGIFRM
EkzHI5QX7+BtfzxU02m9NWo1Fb9aSa6Du++jjoWk+4MdvlwWl9zKoDN/QvQx7DR40/iiO7a3FsY9
NV/ASuuoAF2Jxj1hViUIIqO6hwm8sW0KPK9HmchYny+KTO9/eR0fDD85+oits2OOOPZMPX1ITRXx
CcskMWy0atQ5PcztE4Y0faFhoi5hRxUpLMX4vg0kK0GgdM8nCOoXzTdHdjxyWfsbqGGhzNAYJNiG
juCX5a3ClZbb+achDULPelOERItzu38RFJUxWZf4MAEaW1ffk0mkNR+K4/MZPou0YrmA80D53Do1
JRqK54hq7hjKW0MOhoWHHNcnwyZvumUscdkECMwqOpvYECFw2gAWFuPbn+5KyhzafXoOSHBsibIk
/4o+N09HyjG1svJWwiZuXoGqMQlE8VVDXmcmJgVDIhjwoFWkQMVvmpO1jjpR2shhfTlpXOxkUqtB
wVBAeENaPYehaPFa9G59ByPTsvM5MXVpVmudzNxaz/qSqwvFJThubmeB5S3YbRh0fp/4ooIMW70X
A+nL3sfBFWHl0s5TW5gZEKW8QN7wjeK7ESbnmNkD0c97hNFci+bxYYuuB9opyBI97duOTPqksKVl
Jc/Q18dJgc8u+jvqibeD47n36jAtlJ9FnRhgu6ghKoHzNiwvJj9xcFM/hyP1ul41yi2uS8kp1+dc
TSW2228aqmyKzkZCxkG7uNrxvJJYs27nvaRu0LCXZtZeLZh8+nYwjfV+UJHH5VQbqrClSpeltakn
rHYIfPWryDjAIv7Vialo7yn0n2peSTcxhhxqbw8euDbk6gEtrz3Cvskw8NCFjQuMSijB3pHmTW+A
s4jngl7GVAxiR/wNIMjpHTfoDqsE+t+7/tcYtSGI7j2uK546tqVdl0S0qn8978C3Fdv9jHYAK2hI
xKk4P5bqLIP+wl2xefcigW9ZVUIjIM5W5NepYBgYC1fyBS4NbluvtEDctqti6nevhwW1UNii90bS
P3yOICN2dBW2+ez1szGmCR01mL5Q4Psti+XXVF7FU4G5zkxSxd0qUHlpNKE39uZasrHsAZwpB7Zt
31Mz7eQfefHp5pfW+KJOXZ0RVrV3I1UXryqOmDKgDSd7qhxO1zGgN+2gbrzUnSqAAzj/A65TTKkx
yy6KUtdfUdPtizrukv2Ri+5gdBFB2e0L+VvHeipDW47X72hWtP3VKNzZMceq72TaNOHSgvQ0XnSv
2COPNXTtJcWWaOVD5XWKHDTAs6wgqkelNCJ8D1z7NrVEcfkDFNCMNiRlSkgDw+SCTd2Pax0UvwPp
Cg1jClcCVB/G8BwKr8Q+6zZOF08LuIxutCCZ1bnuWTCI3LpDUoodjb/kyRiqHDTC2BvIEJv0civx
CCa498cfdrFkzoJGcXc61eC+5Vi320GsW+oRWk6QvQawnW3TygatXZ241iYbAesJGRengDxeRRIk
7aGQkit6rCfxNGRRzx07uAGiWtJBIi0yzQjkMXFCDiz69DhVrbTN4FtfxmM0VYLEzax00aJBDnBc
tAKtIx7BePTqJ8vRGHXcUgfJqqPyGgnHkSrONXfd5sCe5Y9SmEEBUMJWZRLtGr5DtizXI2EW0ias
TsIX1DKIVS4kUOSnABKtblujDUj+yKucTmWDJm4wUj7JlQYvOBPurKqExY+YDiwsXX7M7K+eekIo
Q7bFknPk31mTPs7Mn941QYMcDCFybCS4LY1VJd+8vHBVifMeOHHJcjCrjj8JMqoDJhU4zMIrYcix
zddLoH+bP59PkGLs2Nb6rUGCoWo88rNC/spu0SS8Ekn0RuB6aIINWPb5GCcqqqsfq2h8QdMBNxB9
qmVoYKR1e/rfjlCpYzEdIsxceG7KCVWxFBFafUFeUPCQmydlaCDgi9J3r1Tu/T3rxSj3BDu8j35M
ErF8c9kOiyTHa5uJ3Cckd+oGszBIsMZiWnI9GaoJ3J2OseNpR1/4EvgHo36yJo5ou+jXXZ7DpCCb
qIvklEvZ+oGXYmsE2RldDCmLwyLyTxMHshTVwqo5B5btVzrevPliY3rCBZsxTm/SG7sTMbBbeVfX
efv0EoS1gJnbR1Xw0wZ780NX3mk7sok+4JByfGwbPKSuA5GclEJmTB2qyAGXYsH1X5Svjl2L5sEI
miNjlOwhVzn+UxDPT+J0KP+HuoiL7Whp2mbFz0boEGM11UZ7GnyaPN9zE81tO3F9HD6R3gVvnpZK
JuCX70Q35JRW22JzVWb7ZJ3BMrD3n2nj0x3gXYE/PBWkCH6H7yNU3bbxNN3/9RjqH+1PaozONwe9
cr2b82WOH492FPH69eg0YY+1ICz7RrU9zWS6Yf58zqgtJUmk/VM7yaHbpGKaX2N9JtO/OsdPTZu0
CuAqkuwLl2h6laNXr0MI8rapPnFWViCLySsjCdG+g1bUbpTGemF4XdoVLjTFBsTJxOoVUtl6CGI9
npNsPbJF6R0QMgvNkxVSQvWtsgmcPJXr5Lwp3G3YZs2jw/uexidiZ1X/TtJQy5TaxzwtXSzKyzfM
tdQGw/cxUmU4aGg0DpN2ME/OHA29tk/P8jfyMcGT73Rv5cEDnkHxRt1Nlu5gAGfElkrOH3j/F6+3
Q2FQkDv20hqmyGxXcxq04F/304ZVVKW6e2sZRyYz+fIUXDFaib4igIpyZ+Ma/4SOgdjuKJcZ/E7d
XbJDjqROHelemgu6QpBwFgfg4d/LBYi1jbmTy3mQoJOvLDLezSwG2n99x4ZWwvcosAcHHGkjSne5
6A6yteUwGhxWGY/p1znf8QZXOtddQkV4mHYYsy/vkO5xkXtqJn/1Nnt8BnfrRaQ3fmuZmQ52hLXP
gNB2/brxaJ5m5AijF34sRHnj5iz9JaLc79/PJDvXwvBE0d2pH3twCp7fynpGlyudRfBKmfeiqig8
Yd0aIrbQy9/T24V3cqPzbcUY/rcqemhU7abHtF0Kd3+Ly2Vl+a+4SeIwUGguQRvkoax8BzvakQKe
zT44Y5yo1DaT1W8Lc1LwoMirpn42f6AY6CKEi+7g8vmpZzpRw2rljopFmpoMckdqHZBVM9Mlz//V
a45NHC3dUQ1mzlkmauCm21SGZQw2BLnd9oRxMKBkIFEoFmyx3CyF6gL95HuoK/C7K2st74rNaSqJ
AJ5sY5Ep/Fq1+lFC2u63IFyCPxF6IjBBqC/xpahrhr0QlzUJZltgFgHhqvLm9NgssCnHrMsifFbW
ohw31JDsKO8f+utKfF0fw3jRSzvTz40jSw2oVinfXuLVMniYamTdHu/JkxMLtc3kynHSVbhgXNYr
zKGFOyxkhnAlPiqq+RyVX7WhL7Ch+HurrPHqeuisjt6j139r3a1l8dCSpeoUb0IPsy5Ts23TE0u0
8xW0X1zf2kAiZ76wHc7o8Nm2PccecfHZevNd6sv4b9tgAADV32WFj9ENUHo5bRpT4dDLjyO8ciId
p0+5AOBMoxFpgvehFwpj1wb+m18Yty8ULvd9cVox3qkKYpmQo/PXJXThg5McCdgkMNHLsHIU1Bgl
bEJ+PQETaxbUmn9qWTH14b61TRMjXXWFXkbTxY1OtUysamqgmjnWIxroh6arwqresYEj71DoNxje
zrk38nV3HnPjGvIswD5foHe/BNMCJGdn2bIaUflIBa6zVMYniBpLlgHQSoLs/4tILojf5ttIFP/i
98DfPdWCmPrEtuc7C6Ea24Kg/h/dQfiMZGhAWIV66YrzQDUBZzCqmJ49S3utXyyptcDKL04zCCen
pOL6spEetJjCf7F9PxtLSyb2rw0fBjCI8iHozhoGWOeJ1MFzZf7KA2gqI+s0Z6Vin6R0dMgqZ2Sn
O2ph9ZN4FiDQTG47yMrDfKsRBkmitZXSPBScsCNeg8WFVh0Knt8B5tnktRXiep+PtgolYd4O0gPf
u1GWaI8zWJVVh6usIv1HTn9RTkvrNvs9sq4y8D2cTZi6d5wECDdbWESglUtGFb9YACyzzuWpxuFy
vtgF0bGsRH2oP6x3SKcXQFJsCdr4djQfgfYWEHB9jBSWCu4tDu9WmXtKuLj1bnyxAJ36xGvHI40D
+x3JFnquugDEylyJfjc6EKCCRwYXnPEZD9GREWDx20DUaezhleE+acoVy9uhMWAm9guseuLlk0Ks
nZwrU5mP+RskrEhZa0aApNvmPmYNU2z4hb2py+nSiXcByCP7C1u8pOqoq5izvVivaX61ETBANoxe
N+4T/tHQOFc29+B+Tgd8BQBIeDupZBSTDS+KbEps91uguOdKIeltTgIzyovypUK7fj76eFCXtShH
fcUjJyjsVApEGiZACPeAfG9rUYdn6pRXaQrpO7xZDnwSfZ98TGlp2qr6VWunuHPuhM/FJg8g6it9
qfX/RbJipEFus0uv5qaEwGYxlRyPe/s4bKFlVmT55AEJRhVtg7Av7y00lFp3ZJBasMUSpOm+e3SZ
LEAo/lpmxTAxM6OlDAShiHYBNTkgBKlI007cniUANQHm1cnhQAgRhtakmAA/CVvjhOJDs/OnA2in
5gsjvEIVeresPnZDMx/Eiy4mKjINK2YiyMgT5WVevJmNCwih71mkzx5AMo9JHj1+21+MhAk0SqUb
hQqa2zl+xhJg6PJ0rmQcPfRXjuocmdu8431tBQUS8YHdHVK+k1+V8nwIEES0H5ffIFHewaWVhuIU
8xVpYLNEaN5ywe/dpDb4YmttjVOILMRiMB/geg0nYlUBzoK4Kc2psP1jdO0fq4a+xRK+A0tgdern
GBN3Q1XX8Pk8NoCypA7ChPjBLsY8Kih5xpu3y2wFEFU512UH+nprDHf4NINCiOBJKH48OOH64hY5
Cc/yvp54zVdpEX2mTBLm/mEv/vxMRubkixb1RiCBNdmbh24Zynrs1MsYaHYA/KQOnTp6bXMJlYEe
YhOkUHBX3b1yM/BybbmfRY1nkI6YK6DQ1axYKMxnoZnYxF8JHL8vI5i4lD7HmwA4kJJdCPpEOQHm
iwqMef1VxU5zEY9G7hO4TZL+ESXwOryKSQ5xWjQp3/0K/UqKDqjQACdpRZlOmen2nqo8BABja0/r
9l+kYNS41tw6oWx+C7VnTuXv+JwY+sOm6As8ZProKuCwsYEGqWoe+5YVrpjGG1Jjt0kdD4D0tY04
DHFY7szDpJrybdpX4ufWbKnnohclHHni39JdsOzt9Wn9jNFjla30/3MnThIgOmTwum7SKnFo7dbH
FiBfuIR0WYiMn+/78bOLdOZ0RWpuaFmr8/MMxnCdSuRW3aDyYqrtdgdLNMPtacD9wNqhiSrz7KeU
nZ4bwmnGZ6qA7/Rhsr56ova/VrTu3OcpDtpymGwX0p2PXOLMkCF4ayQX2ty2HUsqAsaJWs93uTyl
QtwprnIaVXVaUyRwIVUmy7q9WMoly4hUcWsnRzHo5P+4fOw7PV63Zi+QCUiuVl/qbT+3WwcPTah7
lxOI3EH5H9aAE/ZVxqvL9q2jJ5k9AQs1WMa8hH6y9e4K4C/BebXbBwa7V/s9KJrmpIKiM1N+wfvi
iMnBgQc6kMRU9dy6xfRw1QM8LGmvzQV0Gb0asOX3UeyK68agEfgryv62N29UU2tW0HMvcKHxBlXJ
kw6jj3j3SVNYfakS17/5eZ37oYOaikxBmCx3PRjhi9cU1boeae9up3l58SDKd3csjo2y8Sr7tZDS
yZymi/G7FbMV/woaZnFH2Je9NkV8hrHaU7002H2hHNO9d3rpRpYMDwld+Eu5tjkUtvpwfnsuOH5a
F2E3OkCPKIIl3e177ta8PeeZRxzedIET9lN7h9OpEEFj0f9J3qpUF2Ff5Fa3ZIzpurZsEaQER7h4
pekBedOXvCGY3wJ+ZnYfzDhSan6iOwgs8RfpwVVUoILj5c9CIkDXE2FNrKBPbg58ErOWqPlbU1e3
zxGVV4ZuOs4ajPx1SxQcHD11efjNQk4GjxSkiASCDHe4q/EPjjfJ9hIJGw+HG2MZKT0KbdRgiboJ
d2EObnnq+DIKwWQASm4XA1NS3NYoWYgP99itSRFlYq8cP4qv+6bbkRHH5qZLv/EZn2/5QPZ10L2c
6z1e3PF9UrqDjOUEdvgXFvCOoA1ZJHBzjjXJRiZM+J7T0OWCf6MaFVbSgLjaIw3s/3bra3eHC+dD
56ZKgUIfnQQ1YFRYk+3vtKsQugR2wOblI/ZygRGXio8zUO9I/+fi/S4mHzA0nrt3MNg7o1Dkmb6T
N5DdowaC82fpifKO3gueG/Ch8l8A4R+MFDIBMsPw7z2UgGG2JUj9nWWfxJTt64241M5xL2f6gVH7
iZ1AGlJI6YSys04392YWtaL+AbJfeTBOYb03Qf8efOPdtCt5n1v86DN9hOm+FvMu7BQwUwPPW/JL
00d2CPTWxEsUOMlA4Zg0/gXYYSLKAFLrh4NIxIzWCnBllVFCXOKmKH1XaNbmfd0IrOWYoxlhoWyZ
vw+VqUENaimuewptvy4dWZfqnQn9TsuA4uGizmqYraUR48faDxwzSRpZ7qgMQ4SJGNzY4GHD3JX2
pLcX0rSaE4dz1fgsMN/gXeW65YJ1qyupubYHe35hFla4rz3BHqKASEG2HlwjLKeha6FTqXADBrMV
5UxX80PjdR130uvdt8koFXW0ageljKWOnhzYG6Z758RLb6LzqjpkD8686i8pXHfn+AahFCHrg3jj
SUfituN8pJIoRAyez3+MBqsy1lTo9LPB7kdb/fhE1EpeRC+yXw58LCpQNsEEgY4PTtoIcArO0ZxO
CFiL4dBrMcmnefojMQA98JjYWEWVKjFDK9vDXJj/qlL0VlTU2wJFXEFTvrTV6sZq2VHGD0nNlLn6
QoVA1vDC1fUwA+LhULEiMcLEKGzhcAhugNMzOxQfN+u5e/vrMAnJo0KAkj0DnjkYUdM6CFwdWB/P
3ESeMegzeUH8kUJTM2vW+vzrYTzMvVjPTRVQsnpim504TqZswSEjwuAQN7v1IOB41dwpZyHN5/Jz
IVVMombpW9jYIdI7F6Q9MmIjxB00UkMRCw0C8pmJSv0eDH0/1GF0JD3TFrip/IgwnqTofbAOeKrN
MktOdhHUu9ngrAWJS299C5Aumfa9sg5QfCV1j/1ast9+9Bjm1y0QUzkJVV2+c4gDlWm6rVF9uc4l
r0Rzc9wnGebIXhdr5hgifFdpI9g4kzAaHnybWP6vfoa1fWd32evmy6K9tfTrGKfp0QhZn2rGevwU
5f/JGJQ+aBse1hFgydvWajD+rpEf3dcB6A2DsAoJzYDWjbfcALs7C7yTvXKSLmVvLdAL36OvDvcy
MRf3HnrERepuPz79aQqU/H00vSW9chJgEi6E0V2ps56E7wcHXEH55NlS/TOnEP0a6T2qjgFm4gZV
MsXgBxWi6gddU7CL8PZPc+OuaYs609zzpugJQN6riFn5yGgtafLfDziJ+EXuURLaLgqEz5R1cbrq
aa3f1J/+1+GI1M4NToWMrJdO2hdMW97S7xeEr7hFqiTrBrPGwWMlxvnd4VpBQRdARxSo8Qu5OASa
Thhf+tgOUAt7mapbTh5uE+a6DKHrPCCJa+knoDE428nGHmckJvDnQzsDMHOJEiQ/fydZqMUcO+g7
8N4ZbaNQdVY9ZSv2cRHvWzmKxBtjxwM0o17qVZOfVoiaA4YlnxqHMeC4VYtEw0ChjBnt5RbEEUm5
HeJyt3EhzAP0cLixNMl1YgODc4Ee3yID5ex9wweDbRlotnP1BgXSeizmDF3xjYZIvY4juILebVM/
Eyr2HrSwxNarW2gpl8QkfJHIe/whRe1dNqeYtLLPhhqun+KzBCFKX/AFVC+OTiwiv8YzSfOEpv0w
nnk/rllmpeD4EsiRAm0DiqtRympapfHWEUxHKOshz9jCcVrE5f0TauZNy+hLkyyvCHVBuryt0Y2N
Fkw+CXM/7xGCdZLzdiR0slYAAAcI8c/96PkEYV5L8AfHvavWJYx7YYxAPdmLXWD7Fes9Iu4DIXZ6
iph+fB0g7YjkPMf4tDmRxCpaYvFLFeNDcNS6yK+Vk/+CbdcYsZ+AMGAH8gcWgOoNj0kXFq5yWdZB
VRQpPHTVWEHLFTjMC6c5lKp8cKcAMa4Q54zONyP1ux1ON32khKEvcu6meWm2sWM6sAgo3ymE5JIy
XwyeQnWfjQgrbTgbYreg0Sh3pIpg2Gu7LZjRCiOeNfsEJ+3IYEsvhVfhxCfeEvknn5LfYsmeJ9aI
gsytyBUa8d/AzT6Ut7q42tLB5oXkpBg1HyY6vWYEndnnUxsxlhB16ZleomShVZ9U/cEuqRZsSaAw
8PK2uCmNqkhVnZMzP82coQTERDFaIkbQIhTyxy2YShis0LxXwdxEt3etWlBVtjknXnSUWAbfLMhS
nDAR4x8p/bYPRoBq3EYNQoRCDw4wP4OWFm2/BeTLI+kMRhIVNI39hDIf+gMekuQZz9KAptoL92Eg
AlhWZRC9O0T0XC05EnxxESI/82zaU0pXyNf0dzYV8TpzsVIF7R522Jt//FUxWpEnOFieoH4dU23Y
0+zdLcaXLqBYfzlIzbRung0khgZfys78IE0b/6zm5TA7M6vjTEjlnp1Mzod33Hrm3SU7T1iAZTLH
pQbU7DRvaCuSvPOWznZnsV2AoCe+Q2sUmQ474zolXNTlJng4dVgzGSzlxxYuiKaR+Cof8Mm84wV2
DDa6fjGFFtGoAiamjwX1B7+1hqq+HrCyfEOa80JVglkgrZiUZgz6bYKuKFzxggkoeKG4jR4u9kyr
WSCs84XnRuL5Qrmujsg8jBBv8OFOpba/q03DYyivF/EF90w6UnRq9pLQchKc3POYcyKYiDGSAR+E
H86+VmLaSSdzJd8tPKvkYQpvNPeZPe8AIbPF5VL3jkgqNeNHxTTXjgacIYY9uA8QmxTiwNZ3nE6l
mvV73i/mPJp7Ok77gZyZTYZEIsXPt9HTMzoXkLzK/TXAo+AMmECI1G0bSDTccDHeAko4y5OA806v
yJBz0lEFWWGoe8EZqRIHvdQIR32Z5axQpbZTu3gMh0t73+O7rz8KHVr8iufYemBDoF7bGTMKPl63
B7teZ3rKBpIjK3m2YLq35xRepjjAxQiF/tU2+2ZCABpqGWHZ1TM2lVxtafEYHUVPTfXq8KACO158
URWZmlmwYlfbd3ciGdsoNxRcj6CjDoDbXnwKMkKhMqimu4nkoUzU2cM2wSQvITN4N805IXGdBx1c
3TA4UELyv9Ln0hlw7LFmtK8s/754G6osViqdLE3j0Oj467MHIrK8W5mYB8TukcsK2kfOKYK48ZbK
K+9P6/Na/CnvQcH46I5UzCWxVOMX1ZNFZ0FQAClse76bWmx5y75SrCdQ4v2hEUjdNanIPZZqBYHz
Vw1ckc8pJygATezWcK7VmcRJYRdq/MKlATRqHIzi+i2gNDTjnZNBNULh4s7tDoG2IuRVciCgfoSH
BnoJyNT9Gr1PalojdeqouHXBxRSNN1ckeZbsTmqmnLohzvDLiJltD3b8yJaNrayJe4IrI3iGiS+F
OTRfJ1EhfWJu4d6CP+8gwgH/IhmaZerLpdriqRxFI61/V7SZ6eDsTAN2itwKeXuKUIRvwHsK/KnD
rjSuSrMDN1VTFpjptNAjc+/3vl96nmTtLlojjjwkmsDxrzZ8H7OrVo+oZcInsK7TXeTb518mbCJP
v/3vyIiwKCg+0O4Tp4tB9xoK+8WgTipX8GHvSODcK+snghZJLUFbGC87Mw05N1dPpTaKV9nMY/0K
3NNaybsKqikCC4BcGajXA3YnonEkp705BLSSiqaRvE8gRLme94ww57NGLGRE422o7igRFhg/MnhK
8rIqeq8SNST8nYA0XLbU5TtQOZlDdf1HwFLpbgYjeGuutceIqD5HEyExLsJlcSxZ7jl2ddwO+3ZU
1/yqrwR7RILF1E1hlwCZG3qooQx+PnWL7RghgrXIGhwpBugWMnWEQaVzVKSV3guD8XKJ+A1cH8KL
Ss461vQyobPBYrbMLHg/9Y96EP4M68xzt8xluoK3waoHkNeBNI96cn39HXbx7MEXcq3IlUaKqsze
iRZvkIOs/5mS5J/kdoXpSb6ujr80B14PPsK9Tbabx51B5qNstXG0z0ywhDyxoOlomehHckqoCsQU
lI0JcrKQ/Gde1YU8+6RpnpjirQT4RVOvE9J82JtsjljaWZPDrn71R0qx3gonj7+KFcu5oxaHcCWQ
lYBpsHCMHOe0RqH5KKP+OAb1p8GgTvVuEbov5E7IEg4f5wVsRd1UPHubShGa27nUal61x+bcXlFF
3OM8xXG/D8Y5e2SSGdfeHrn/giiwyJufBIuQp67Kr4CrZlpcDJVt1Lk8UhXaCM2z9jwsb8uzD6rC
ApodOdnmcvMq8JFMK+kUFXZn/aBxpKq2Rayd/YvfkDoaxtmwnxVKabCFqnCQ2NYNhgizCqT1ZlSX
fjB7x1oZ+NBYqT3kXLQ+5l9oJvGEZ48QNyDobMq9foCbuXNnzWVeJe68oxz4k+CX98WMIoCmVbUp
7DUer0mfjzjGUUsbpX31c8ywnngqSp4d8fl12OOQCl6f0xk/01YLG52lLwnPxKewR8FQhTT9mjLo
pWxSNk2kLa3d3lJ/bgQOx7Fu78DE0DLaXJei5v/Dunbaf7oFwRia1Erskzhb+SiroBk+0IktEFIN
uNohVwZIZLFvuFO1EGY6B9dk5yI7/smfYXd2jJE0PJ7b20veTUuGjrkWB0fL0UrqsmFJRzdWleZM
ySTZjOTUmcm5RqE4728uT695KsYIgXELqo6Cl74GUagp7ltg9JGMOIJMrWaFQ9hpBIINHK+QNmRT
jOmB8CYRTUACswBKQK9PipIY8JRTahQfMCMg77MWCrmxddeGoUOSJ631Aerf70gjw7qMje5jDCp3
tZRQRFKqf7POdrf8wsI2Q5kQVQ/mFFgMrsL3ueJn0l91+3mlOOZLV0HHdyaZSfzCi9RVbdEzwDiV
CnW4bk7avxlZrYlrs8fxzPj1y+J0zBIDz0YyOeLRXhGsL2Rzh7FCIYZw0M0Ar9X6Yejm6QZR03eN
29qmxav9kJAJOwd0LJuTyXPOcTnIvIrakSkkGV3mnDB12hl7dekisn/3dO4koaPrMKdbFeJXldmj
LpBpEphPuu+KqjDOXu6f4rKWvIuPDskYNa92UJrakC/ZwFgVrzezT0LjCLqvpF7eVJfyX+03fd9U
J6TzrALcU3wN+g5MXnpdFVC5N3Ze4Etw8e3pF5Z2U+zdGCENzaGV6F8DMLPQuT/mhfyqe7xXDL3z
jRsxJogjeJTVsHbFRpPtvROyBR0dhe0UkGf7rk/KazYJ9sPgD1xr5rqFa8kj5GdIbz6XtNvJE8X4
/8qLgVkFE/QbgUCRKUQ7z7bTGsA7Qs4BpK5vpOWRWvAU3zz6DdisBhF7J97rBdQMn5bb9HxP8iIO
rQkFJe3UsXnj50sjDIP7f/8w9R95hG9Mk/GFbGi1meuPBFscvKj3yqmaJLH/WSxpPLZSsMZBZrq8
Xh1F+cSx4gtpayynYpO8BvaptUo4YKFyhxSZFoy5NCxNFwliS8npIdTNsmUFhnsfjpRuiD2SdlnQ
2CrfpW7QGGy42myJjBOWjNHW0Qo48rpz7DVnMhJ1elIPu+vhlnRM1V/sHj83J7srImOMTAmLNELF
gIMhup8MnnuyrJaxpS+lK6bWscxcEzdYswuGIIlKpVJMcy+zrqw8XDnlHBh3zJzlPU/9+lZjT2X3
E7Y/zgTybjTEmJ3TO+/I7/cLelOV689stEKeyP5jLRe5ap4QFcORtizcggMFywvufsM7ogXQ9PY3
3htpJEsoUGERoESJH7QFOlLftrLeda1UKrEA3QuWCqb38WN9y0CuKZLtU8UFArNf46fZBGGIN2T3
+Rxlw3mliaNFjhsyPetlhcgZ9DYv+eYGbYv3MMOjuDorXrVjCzt7qq6PCM5yYzow0I1bwKqzAnV4
CSlhVzRkhbPopBrRB/Kjrd0tt8u3op+rC5iUMf5tMIiEZHgfrEgb/M6k2Po+hjCrTcnR5ZVYHtUA
48SgjflVCGWcAALMtWtEW0Me5zwCYDefxMlxJyXCWMCahkucyAN8iaaBzQSr+xJSIPvSPXO+4CVU
TYG3C0PGn3tOEI9PXfsGcriObbjgc7yZTPPFL3LA6WNfqCBpDB3DY7ZFgH4tlHiVU+fffQ/c0NbG
CXPfPHlL0Jlek3nrlJt+b4OoId9gDyxgKVcqgFey/76hbLzPk5WS0ZEXUdt6XRRXZmpyCQnRR6qL
AIxgURKX6JyN2W53lAalccJ6XQv7yz5ZI2IhbVCwibP6Yy+g/C1i9g3oQ68+M4hfCGbxhJnHPiwv
BWkFJzZbVn6LmtZ2PDahj2qQDb9VxTEe7LhGK7OdUd6rPW5u83PKhV7cCLLZkRcbEg2M3RoXZ5Ry
cyF5t8yV4FLVgZIODNrrGTd1QKgLAHeGI6jiosQqIp1M6vsgvTOtnWnd3Qp1P+woK1SNBGG39e9e
3TcLhdhi3/BV5c3NeBy8UkdgKxwsxu4+EXFq1QsjT7XR3/n5gduXf0Tt23XCt3XwiDnYUzktcjfF
glSNm2RjtT22tod1+DmJv7sN2TPUuJaAD/68RbTG6m2SOrIvx7iZLE4GVhEAFO1f055KWwRWqaTp
PnSTnHrjoX75nGKCFP8BgpeNxe3a6829lTrKBLRL81sRS75EZ0lAr5iODq8ay+3XwwQOK0ZdZ2Up
l8v350b+pB4HoE7PIlScglchcVtsk3FtNpSAuWCZZXNcpYWsIBlNiz+atzN9Z7phwoq1+x1SDpqk
x6Gq1FxBHhm5ymjL8dYoHADK8hsmgiATMrvNt+NqxHrGprjpUKavW5sMHCUi43QBmqN4TIdLoAh1
5hYhZRshRnqgjLD89PJIKUHTLdAoNGBeB3w6q6JPiAs4XHNSXLECAx9iz+GlCBAPP9P03OwqKifs
iICug6TLCNr8OYqEpHekMRHSKqK4w6cwbexltH4KCRk3iP3ys2VCszqOvEh3OkgG6TNpiK96Mxyt
OISE4Cq6e5XkKlPaNMRfiAjbpXRgoW1qCwt6hIQPpIqHsx2WTZzqssDA4Hlm29/JtuSlc7NyoQ+c
LBbTEZ9ynJU7+8TKEJyB5C0MjggaJbNeyO7xdooxt+inLT1QG8B2XpZjd7NnKKq3k98Ec2E6yurL
fNwNVXiwquo+b63VLAcwoclpQRsqfHa5b9QnEB6O65eVTeAyyhl4gJB3dXvWYWw33+piyp/y81PB
w/5EheOayCE5bOaQ1reOayFW9/dq20ejzb3iZyyZY6uAvws8n/DwKy6ThwUPCzFTakLDWGdy1FgE
+LmDpHZNo4AHwUAREQclXcueoTXre+yn/1YHUr0acbF34OVKjrikY+1iqqGjoXs6LYYXvFNo2GxQ
/geJi2sOai4CF9w21tmlPwUnDHqiclkXMjdttNmQ6xRwAAudp8S4OnRPS8aw7V+dksafKu6j+pDa
Z1pLpHBOXysi2sZBh6bBszwfyMRZ3mEbARmNoaussmE8MlqBT7uzuD2PE17TxzC88kMZnR00+7nV
JnhmLaJACE7DdYuAx+Exsx2ZtWFYuZ8eRv4svTml++CLoaX76bIWkgWtz9jhbEu3vZTV8bAsRRMU
aZL8WSV5cW0ZSdBYffZB2QK3cgXi7FQBpzGPY1tQeN1Ze4ZVaX9E0f1lK192s2sAAlLXwIbAa+45
KdXs6U9OFNAA9NYO/Ay2hCE55rkN9Kpi0ptWBYJnGvbkBVIOIqxijL9k/P9qW5f9hhdhZ4f69jE5
rcTBN07gUtuPOmyCd/YRpzJe+Ls1NyersRd8OY5G/CYUgFgYgYNB1j02XAe76GdBqknx1PTumBJE
12AfUTWmXmXek4Ug/p/pDRtuiFXvc2ZjMJ0ykkk+BoGc5P6CCqP+5hV9PgAEr+p9Y7Ojioqtrxdn
ahOn+qjZrVRdrDw0OqTfQARm+bq4yTfDEUAJvzGNoZaKOzBCNKCZ0fxkm7GNbOxWrRRjqF/j4118
je4kZEOFazMi6cp8z7K9jlPb1m7aRMufoq/xYnayx7naQ5wBEuzbDK1jUQY43lXA0/8dP9LoxnwV
GQm8AvP/MSRyTKy5kHCd2ln4Cr+60FiM7eIz/IYhWGF4GX5dgKlvH1FMs6G4Eevnn00cB8kePcBJ
GQ1HSn9ayz575MyZJb/gi5q5YP0MiQLLisxArJtRcIOt0cmulAGlBcI7xsNThIEzuAZ+nt5TaOAG
barnWSxO2Mg11PdU3vbPxkq842qk6lnaIK9t8WiN0BrksssVy6f6ED0iF+wDAJNe4pSZDRG0Du+K
IsmMyLweR9m2X2/oQSCzpfQ01ekUo8v86cOHQu/EZ+H1K2Jrcsw5mFCrjQwf3lBzCjK926AEXDLP
F+Lf0soMmpN3A1k7366W4wpnwoLEvrSQ1ao4LMCBiEMbfx8oiYjhY870xuWlvKdGt3er8ZJ3SOXM
ktrYcWw85+SfkeeVaV+SkxxKEUbVRhQ/U2aq/7ZchFx+VXXfPmibnqF8QDLVxAz4BOgTYqkY5pKL
QnWHuVbzPnYPUhCGnkyDt9XYU5gTkyEXlbMWt3NigwROkzSePB3lIdYuvLt0QWdBVunLO9j1JPgo
hXKQ3/T2/DrD6wsT11JWhJhOkWyk0gxLNgRkCTMKpGl30I/TNjmKbyPQw/FM2otdz2plU0Cir8sc
o77jpZ35yGyXxwI8PyFSbx4j5klRXMx6gtIkFGUCs2vw+s4nl0RyHrldkmdI4oFqw+pkuHOwa36j
yYUS00vXFcMXOeNecEmr6KvwPSMDPo9dJdnRwygOXTHXTWF96TE5lZZlT/w+BkkXXBn62HJ/xQqy
nCteJlp046KrQdM6l4J/ZEcfnClZqe5xQhROOEQ5tgQvl3uTn7PiLf0hzRQwJe4gvuJbqaptWbgx
9z8h9JwbSepkMh0dltaKeMqE0nt54wp8BsA2BZWoEhUf0d17YEjk75G3fDvEAYz4AT//b0+Z2iKO
JNAXIXNfAGnB6divnLWZT87vWj7tk+vUXpGVsltYa/3l4IEGmJUewzYpCdTp+ATdN7TyPzZkux4S
j7hccfdOooHCh9+eyLEB4cKZS+qD7pIxOvIXqhzPy9FlYv8/SHn53KexfQy65Kx8hPJXSFCDrLEU
KrLVnW9AjyGMegWI2B0nb5S01evEAEXlVKIodaicl5bZgGbVgb/qd7+Wn9rLRRG61mNMXcPqpB4A
VYB/fbu8mh/4aurAydlGVXvxKwmwUo0Wo/xZQwSl7f4Lb+o7Aa7GgHwMBlgPYXL/2BQ0yCetroHX
QqcXOrMrj3xIc+Cl6SdUGcKdZwpWpdq5IaBSDhO7IRqZdqLkj0oNcnmn11b3csygk45qJC4ZAK4T
xHPmaMe6zOD5jlcvlFpo6dag6A1IK0n8Ojc5d+/TRSMJ4itoBj8C/gUiExVaL7JuLENJzTgIvI5k
MA27PwgRsZpPdn/7cqswDjJQLCNlXAcL7PaMtoS2qODHe1rvXgt4vzzNU3+9HVXMUK/D77fex1JH
OW+rEMvUznAH+ICF6BROTO0lAXDIbq7S1GpUU2aIhk77Incw7FzqiAdNLTzAF5glBNI/q6cakPLr
H/foxWST3eWx092UXgDtw5GbgFmARquRcb2JDtpZ5lYci6Hf+TnunAZdl8nEKmaAx4baA1z7GLoM
38IyBbZtHzt3kJMAaU1+5gqag8rqxf+AkkN98d5Fc+FZbQROdRTeSC/rcU4gDzNCYMspIA/1ooNP
Jf8ybP46S/vB85gWnVIBw/X0bmBwfD6PFP3Z8Ius03gjBMEHbcBEMs2UjYoNavXnq11WY4/guc5o
A2Fl71vV7Ya8FasFqh6Bm93j/fzkbaVjlNu8k1I2ysCCdFTofdHtso8y0U5ie/8QYMbK4w0QbnQf
W1anqGbZw4z5zyaS5rrDXIoxLrv9Su77M/OOpziQrRok0PtY4AqODCheBlNRrWfRuiTLkAKqcZP3
vg14tpGXqdzVo4lE+dheChlakUVpLroDsTpdgu27wB2t0zpjP5LJt6cYxy267PFT48D3XGVbulSG
9AfcznSe+KP+fwm6JJdVRmyeadCOMdCaJNkaxzzJKbB2q2obdzpcTV/3UthY89twF0WXFt1LyNRY
xk6bWEpHduRZbPHA8k2K27bjabWa52/j12OID6KPxV6wwdRSQ3OEhyGUNw1ZmooezP8sviDsOKo4
2DqaR1EJ4Wk0skNSx+hoO/OD9wxDljXPx5r1u1AbW3tI15UAgnGxTOJNcX6AKTKsvNgmwe6BSCoJ
xxdNaffEuI1/hONTTAjDUvtPkKwb6lQkeu1IiWGYnMFgFZrkD4NC9Z2qsr6jLQ6yvukq8e/CU6hc
6k4XOhfLmhtEFLn92N79a5hQ+tGVHjC9HXO4EBxbjwbaWB4yt/vZ6C1aCEQ/ug6Qzu6ljDvsTbAh
E1LwZUK2v0Xqu9EVxZnKvkf7Z7I12p6ACotomblQB1gE0jS+GH4CEV5n2AAgvQsr5ESYV/8v3TXu
6VKoYv2zqBNXaPFUpcK2opbUQ8SZ6W+ojUknbSq2sUPnJ7TeIL+PVyGXJyvxsOw+CmeV9BoZisbl
Q8gIfYHvHgBunseBU1tCSNfUW3K2GcjaL4+RtlvjMMtk0fg5OGYDbz9wTivBSC6aBsJIYrwFCDMi
+dDkSCHh6xI5Ogavd0OaShQFIyEezioXSr7oaYhpxuB4ToEv5kPwiKg/tG0pMvFG1HDYut3wphqL
nsujdobNPKJJ3L0yU/78GixNiI0dA3of7nMTOqwy+/JekSfx331OV+dA1SvlQxcuhTRLKG4JCGxv
aWVllMNVm126ZZx/CFMxtK+UX8azs8Ep5VVFv2mL94v8wf6iZYAEA4pkdM4eoNUwECc8VU3Uirdz
Rur6bMILZGMM2Vc1xm/Eh39ABiDYCBPkp48RfCdKT37CjeHkN7DarXYluukGR0ICsIz9oWKIXwW7
FdWAeApoN0DBBGZ9yOC3tcxATt5fWp5bKqxEi1pkFMxDie+CK9yfIqmI3DqWm7c3DhNUPLfVbJv6
dr0OAPHDgXa2V+EPd76bMtDRVW+GXIDaFJGQuC2lhgIoBjBehRhuBXcnAEVVWD3FPhe2ZFFYGnbs
XpW+hQcmmk/k7p1fucUs+wAChqvhBYhbdLQAp/WJDXzCQo5kcaW/4tFWd5l9MRgnihc3vFLD82yY
TAoJYHa7yO1rTWc2e7RPrd97ljHxVLDDDuknsoGFzRpD9RsqEEIlWx9RTmbKiNflZijxCr3VkJQq
DhEHSlZhiQUkPZHBEmXi7hy4KvsDBAvVDeRLWbmDAQJLsRy5QijbsVBgab751GTsmc/nxnOPQRnX
YyR/7SoemTgxNFr+hMVbF8KWsZ5k+15bQohht7eObapr7TJ4v2XU9N+/0WfLZ/9J+lpQinulpgDU
PtQOZw2xftQjxa1xl+lT+/kyEmbjwtpCHiVQc/XHugV6CftwrPlrtntBM14uFYduj7UXQA4VkHtk
urQHj3jFqVLOxfU6mQsts5YshAln3gv8QK4JhIDH8U3vVa7ql9svXQ5Rx6dRFfiLK1f0hS2oktlK
rJfG6WvS+OHeAAOl+BfzSj87wUPL3CoATC+YfnBwGhyitzaiSseg4D77zZE6qfOLSj3sMgpv1U7c
VFogSeLb8SqzSrlXlMYol97kh1Pj6vq2Wd1K6PEtaqw9LHxxaTfotSuafB1QQpzUfn8Cz1U71eZJ
vtgRR0HzEjPHXy1yi/Sv8C6OAyu/3B0v9hlibcIr2ikUKHMaUuOlm0jxGadKYSBOHsU1eA4vrIeC
994BMLH0JeFH2BbW3xPg53DqVeiKMJtJNm4MX4ZDzLJZtHsKHvbIBaZ4u256EkH7w5oKRaOfulNY
ivFKFxoGtHLsRt6YpgpcZtsMHtnc5h8KHm/ktGru9kNj8+DGYujNMkylI8YD9s9tfP+bB4sYmvqw
bKraA0Dqparj/0mtexHW4qnk8XuaIjC7ZGPcOim/HtUsw04hToD9REcl1qhYLpLm5LgdB4wpP1DP
VzWjjNQQm5TAuI0P9d6pfDzoE3ethCokJdBqzmqaeV8tYKEnare3FqJqRhlWymk4enH5IMXLrJTY
ACUHw/u7bi/FTHZH2ygvKQ7RRK2iaa2PK3uOIDdNmhxI75Cu8CYCM4DZ0OM33cQ6QcgzHEamH9EY
MEIgzv96ualhu/2nx3jd5xoV9iR0jsV65JtAcwZkcC43P5YHCyDD7L1VJtiZ2hyF1oXmA92oRwVt
wZWURZmLjA9ah6T4vjqLcLXJCPipcrSUh5yrrXT4NkPU/LqnzL3VisVfHVRUyW9PK7omkCAIjV+s
YLRN4V5JzuaFEMt7c/rSjR9oqlfA8mUBQN4W7PFTKCJQYbWbVrt2cml1pzrAO7vuvFx4bU22giqc
1lCEU9afL5VpS8oxt6IpDtIZfW3hw4bQD9QECvGpoiFkCu1fhkX54NNCba8VZ5HQsJlZ4B8xlp3k
GA4q2ppUQ9eiKwvWYzTlJgye8BEvMJwu/kjiWZuKzvD69mKZzGVU6K0iWgEIou7/pCYeQ6xMbpNx
FkNiI7NkGwj430mAoE9o3pBHQ03OHmP1IILYH7R9V0bLYphU+EFjn1+jFTCCqrrHfTSmsmVbKPeJ
H2lm46cOSJ1Ajq4oU+I/jjBInmTcNXwPzXbnGuFXvkW6nMI0Ron/lgRIRMsq61q6rYehtImvL9ry
W8xezRyOZmOLr5JyGaBebfYLul1/h08pNz57Kp34JKc4LqS1gKZnLQiA/jNyOEY993Bm8DcGSnW0
iGrjaZpL5ev9pGt80rfc8q5MIxWZhayiefL1BcpVTusMBHe4noIg0h2UeczjtsJnnq+f4/Atu7xJ
1PjvVoe6aIXO6kZjv4xpvWL9tDhVRCt6zMttz4iG7ydaJopMXvAFYQYFR+a8iyv9FdwfUPT7BVxM
+C6N4VCqN6mXYIvANEwr8GAgX7dfqd3tRHaILWWzkkpKtMu1+N9vOxrqbHK48BB3qwjdbcXfkJmt
SVtjhTynWHX8OYfk1H+X3RXi3KWufhFP1IBJw5bVrczsJGhl39h7ogZFoS0JLC+JXqSH/u4fSEoc
Z+DIJ9f2oNy6TwSeRDA+8P0IYmNzXgL+HLTshDkidxRpUn+CQeWKwXl3H5Taj9N2LDENlAgw3DBj
F1z/9vPPBFDPD0KOx05YE96RfcwyZmGjPyQRAuK13hdQON+iPkf867m4O2Lu+i8OOfj0EHVmt47O
Ih1PNxQopEb9Vrzr+5UUZIjRpHEMwAdEAvBYzwOTZUlbS5lGF1aZ6cleyv5B8CEx5xjw5ZvZxMa6
IcXNdKuxjm6GdtVtcyaYpV3XHYpFDDjMB3H1+XTuGoisIAM8F7WGBblkVtqBvGyDhXR3XLkVBLMS
boH+bYOKeOutHgHO2Pl0CYbIaoj/GUZ1yWDd8R9rbWQEXprV5BBABE1iDsuV89xFzIBcrZg+/m4M
SGVsC/QUTlTaM7T/hjjCbz4kEVBDq6kj975FtMoleb7KacyiL8e0lgihWpB9NDlb4GmaC9KAUGoK
NAGzvTyrAvTg6K6vIgnp/9faRVRYnNMQIsQTXpS86ZFs1Slq7ZYB3Hqnepsvo7fuC1MDLLDXdEV1
YKhePHNmboljpnu5BRCq+Q2gsIAW7KZXardqVDBdAGWK3ykASpK3KHNdgI1iATVq0f9rmAkOql6i
gZUA0E4o9FXiMVfjp4tKA1hjpa3/VZWx1zJP+lWRqK7tg49Z8leTdji1YXP01mIE1jIH6hfTrSCQ
skn/a9LqXpsEFcMlpW5jxYvwB/pW+p53e8JsuBnmp/hv5w8lNKQrBtyKjIeJSW7XCXzzLNdLWTnl
4puGgobT2FF+zNPGdv6aG8lV+NMeRTQB2Pv6FbBe5wE/VetwEvJqTbZM9qglps5ZV8E+37aEQ125
bzgx1zNgXWI2gVmwOGV5EF8MXGb7CqaLdij8A9vpueKq35MxTtCNGivq9u8z+HM/NsrpXKw6FkWc
FW9ikCX0FL7ALH9hMi+LWAWTyuYhRV5JfL7KEp6/+EKlXk0VdXRbD8FQLaGcyVUns/i9lW7Lq6Bh
nm5UKRzQx52uTQTKcz/CxFJ+8Lr1tz4BSxwxIo/rA4YDexrsNX0bKs8Nm1Z8lmmzB7wjC0ulfM9y
4VYeJoAI4fk5kS/ZRNbdoGNvoZU8Pmr9kN7YNyKRljpPQzGjwfwkD8/XIMHVh1zHEXHB1kTIrItM
C8j81MbFvNEBxBBetD5SkNfp1a6Mku0fQRo7JhZf2j970ZAHTJ6FoUt7xLS0uV2Sf+jSsu7k6Ydl
Su0qPm7aj5oHMZJ5YUoDjAurclKJ/tscyDGa6oGhV84ium7adZZz4YOcUO+O2Zj3X1pJLgwuzBkI
t7LPHljRSLy/dOZ00b1HPrrPuplz8bY3tAfRW8+MRZbKM0o8vOz5bwOau54plTEM2+qghZywtunb
A1EDILpWeqM5nTO8ecMV+q0iL1I+T/DMc5jXCWrhx9cQT0Baq9Q1jycyPjE88nWXR7GJcuzxCfRL
1v/0lSIDiROx4Op1bf+pBtxHGJ4B+aLIT33BcifecxDHSa+hDCBOjM2pCKUymJEoFTl/uTJ8TWoc
aLgdU6sKhywJ6z3tO/fHIbqtOgcCXCsoWBFV3PBBUWEO33ZGsk96Dp0soYKk57sKs95Zw3lL6j/+
nWZ5xux8Bizj4iJUT/I2wjUs5rpVZnYNa01ImEuCxjN4P0o2qBAA3CUXXST2WMdK6+gQbRuibKh9
1pxJb3T6BZY8z1fcwb2YCCUS60OYAhhv0zYOxm1YNTKHRhq5fMcdVT1gtVs37hviKJodiHQtIc6i
h9mSumXnKMZwekQN4p86EIJA+cTXtJZWAZyJQuo295XMrxEDAD2K6MAXxrYwal9lvtVtrmd9s+M+
WBAdIx1sKrg58xIf/Vw2zhtgdgNK4IKA/rPytrN8DJXfBUJcUtWCT1vHWhmsovAXC1Uuv9WRWh2a
6U0taxoRrKDL+TQqZz+Y0InLRZvzkqeqxRGZbJ7lC0ig4z8W72X1Hxyb2PtgcSayhx+kdN5jygyJ
OQR4vGlSHdYUDSXlspCeFiuizAElOXSHMQB6211HhGMPFHePPrjlxKHh8twPR02FAczVE4pusOz+
fAOHGoeI+pC26bqJ3FcZTaR8Jic9yn/78x04q2m+65GmI4Bz9jBQ+TEI0kFcbHBJDwsrq/rwVsCf
5z+Q6mbihKaY1BZ0MhSAKYO8OiIRsYstz1UIy+Z5LlWGXr+ZZOqu6nhYIMkX7yImkhK2MojOvKmG
IJKIUb131+zpaGEDdJ6D0d7yrsFhQyg72dB0AFNLflSHYsknvC4d6WO/9is72vf2cJAsqBNjxges
Aet73yCfKZn5PG9a1xOdZcIy5CmJ8/DKag3qqa6CYT8MMLM7sE535RSi/7zDV4rOtwgEzZn3nVd5
dxNyIhg0oyGeIfsw39Lcg/WUWK8vTi9faCPt9N+DztxkhEIpampviW81/v4Nw6C1QSg3NV55jV1+
Hd43aUDtfkQnyFrSz+cznTWmPLZR/FN4viyPoOJY49A4t7fklu+LNH1njGnq8XQ+wOUZqAq6FU7q
vonzqNc8e16FuPlqiNepRSXWNmqJ0C1IXZtNx3CPyb7oXvl+x/kWbQ1jXHDTXeEuJKFo1eSMtoS9
u/HCBq6WRCaYmibpN0l54b3dTLXzESkF26Nak1UYF8Mvt0+EbsymhriVBiBP+REoEYczs++tbP7j
l/PndS+ya5m7QBrJJhscsDEBGpQ4tvvOMqxp8EqD5eEoG+fRIMAZaG91yDJL/Yo3zRPHp3+AYJTF
sFMK5HzDNo9LAv5+Pax1D+NgNRYUnCtJfdLorCp9QOjoSU2fDqM+4Qgn13dVV0z9BBm+aLo3C+VT
L1C7mY303rMWqNapsZBojoWZpLIeBKjeo+hi4/pIS/oYhg5O4es31e+k9eCCp6nH/jgsmFJ6pVNu
LAVoV/L46jZMF3qilIUgIgyRxuBCdasRMF3y5GvZ1X8oOpNduB6KkBCAl3x5FNI5kTRdclsnFadO
yIcWhoMiZpZX6922cJxZ4buaMRmdaPgp5bO3xAsEAZtayKLPMaQpuLzhEz2myL7r+Epi6Nou745S
YdcVRuQXDzC15UxVljKBB3wLWgF6xkUJnqNsQ/a2Af7Zhz1wQXreLYpxQ15LM0r1ihpcfjW/S0zd
VGCxq+iYZSQMpbbTl4BgqO7fQTQ1xqx9cft33E73ZrwTHHznsKHJsT9zcJAX92PToiNUwrboRMVC
aFdLlp08xus2QVYTpeal+tsLmCWKgRZ7Eqwh33TKbKf9OXwm2YO/ra9k5QUoI13AeEc7d2ETfaQp
lJXvmP4Q8pmdgk1N4ISF5kGFnMquHAdtofvGnnb+VGshPFbaMCDYPF6RrNSstYJFkQCDPQIu53A+
pfa/wCkLg8w5J8LuMOjLW38DO8VzUbvQzthGrXnbmQMaoPjaJUDgZty9bjC5MbtH8W4Jf3J8eVfS
9ya7w4EIV50j/Ujf0vAhNiooRk36Sk45TKt8LoPaPnUAogYaZdootcgT8jXboGuR1jV/pwNnvcdf
AgQBFlh7NqrAhOX1jKl46xjyupUNpwp2JX6kxIjRc/hQxjwbBPIBWz3C0YKnEjfmo3TQo7VaBiMn
HgXqSNfV9xAHW4BhC77DsiQ414iTwQikfCDRxS0avOugR/HtSnvto9Gf1EUCM/sS54BKcV5On4sh
9z3dCY1yLm4GGlOqpGeOnOkbZ1QRtdMoan3ZpbNBPvVB5FSSvGX+yPQxtmu+LO5w/qgAYyH4xDXd
c/Aa5pgALg3xQl2AYMBSxZj8KXKxoMu0EHtVMfm8jORB8mLl//5fqQESNoekPVXjcaW5NZgRdWCW
tp0bXtTXUTiBTu3ntXM0+kloBwK15R4nnFK9H2rYNJjMAcSNRSsCvlKrsy0XkepoudIh6efNE6VK
ZiKx/bEZH8nNurgVXUDZhvU4OM2OXnpQRca4GZVsSRk972mE332e1aH9brq8Mbm2pUyWIX0Xadko
Q4NVFy0Kavpoxs2DV+JmyiHDILM+f1nut57tHdBiE+zl86qXF//Jo3OHW6z7FMJh9eJTLvFJQ00J
j5Jmp2zn2DzK6Eu5xn0Wic3Gm56lejmCT5/NNGWbZgBdgAYpFeZ0KRH725sgk90y7m9flvw7eV0P
rGV3azumcPuYVxt+Qi87rKy93iFbKELYoxwuuKARfsmW0tZ6oJ/Tk7QPuuYeIspyBwGSRSvQYSqt
5pmQWApqAZau8Bnkf6rm+WUgItiAZG48ri9etqqhYR6ezIIm97TWbGef/PPS73uh5aVTM8hGuTD1
hUcFrXW2+0J/OtXn50NelpI+utyEouon/zJxMJTNzz2dnEIyifx7+ZPsfhAqH/M4U72nt8XXrhst
MIOp/cudZ+9bxFJWfZvf7RIbBaEoHimImdLqdL0o4qv7xoDDSqFNKLMhM8OXT0OAYj5JRMfNEdL5
Cb8=
`protect end_protected
