`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n8JgK6wVPP3+wlBIB5hRneg3g6SRaPEUvFpt93tzulO0sqyUGvXnjnZHIJqDO5RfMCoBHfsSTgV9
wrYI/9czew==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Eq1GKe3ONCTv5oJ5hldVCtK/ziP0a6jWmLWz7ggIS3AdUF/EFuERHlnoSrdxtYtTdWZ3TRBTSjEv
kx5kClN8WCCa/dW9IFePhlEW/1lL1Hk15NUtrJLoeq0KnIm6fLOVcB8zur2alC43cqi9Ws3hv9Wl
Wji07zh2gBw6qnLinSo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aq8QdomEwQROVgt77ZmTnxZwILY1qmjZDwwcyj7inv8agvWcv8ndJJll8suCRC9hZ7bi+7XSi4Rg
c+20ZEIgIu9SdxzJhubfNI0k8tcR0y4f3sd0HL5s9ghYRYMTdQ8JfYcEUbLN6PEPi242fAYgje2K
guZ/Fnng1RKZfsFqW5kH1bNVpJasfNV3CHHZVacfbWWLVs0fNZ3j2iKX5LeZ3UmB7H3GkgOc2czJ
yxvSrtSCSYdw0XsFIPotnaO4TySAQedLQhiNbsxJljJFnY76hBkwIjQCf/SqVvbyMCeQa4KfAKW3
uj8nI8vEXdJSpIQ/kxe4xzVcsIljYQ31Jg5c9A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jAjh0mbyo33av0MEk4hSI42t++/FMn2dKZOX2AyEPZUKCHUJp2E03uozYquz1wpMC80jIFnp69rk
DgxSzxZcJW0Ru6MiwHSpCaUGk5JZTEOMQldGFZ3OL9Iq+Otabk5uG5mXKofieN+0KR/sf0ycwhSv
om2kHxeH1rpWUuV3Hag=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X9HljJxE70++GAxOKjp8kwNTa/AO2w83nYISk170tV5IHWB2hYA2cRtsn21F7jDAoSxkkANqEBWu
NTsNQyI+JPinw7d3/GY6rLwdVNOgZdwiCwI4mKKpz6AnlJsA1WdOXsJLxnTOpOvcU5Xd4UHC1mBx
UuelivztKH1VgLss0HL8CA/nf+G5k3LezabKnVNoGupWDfqNlCpt/mllRbvf/qWCKwZS1iI4lTVK
L23tknaMVgfM6LrYKfkmJRIBV9BScz9XRepqtxZkZzMAZzDdcHYN8g+J/HzHL0Cm9O8wOEq60w7Y
HfR0FQN9ua77x+lprTK4rBsMl4F8nn6wy1JzmQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9104)
`protect data_block
y/FmcqAMiQbEdx9RVr0SH3AT5u2SD1swq1pEPQJIGBu5PnG+/dHjug5kSYU2PJCzDECU8zWdkiFc
F2vkFv+oswg4RAT53ebd7ZF48uDOqGOagOCvJ1XgrpCooQMRb/LXC3HgyPPt7IuD+/qKjvxRt3i9
AovmSeyfObByGfMQjqi5JMHB+vMl4iwPZZBJqCbYYUNAcMOkERV9CtPww2LZAiy44UHgUTDSGV0G
8UB9bra+QPXdS1xi88tp1Kyh/NDuChaYCnNT+59pFmoxyQ1k3D8OwAsyIElHgLxxBpmqrtCdmh13
YjrsWebqX8ddkPmEP4aV4y367fnaxynfNtR8hB/4XHF5j6v0v1huabph5/A9gOyt9Bh/FmtOJrcM
oSib6Bs32/CV2x8I6fcfMuFp1+e/ipVQK/VNqXb5baE+piKD9OQzfNjQOptrw99PZl9wbLrrurdz
DyNWgefP0f43ksv6yKFP0cUgpkSylzfjA031SNiHJ8P7O5Pz1mIbDKxJv3qdETBEIbDX1Zc1RNVN
5kJhavOi0Spa70yeQsJbMEFKvFhKotsPJT2oxF5h+qMYHWuQtvi75wAxhgCGl7ZbJ/PGM06ZRMN/
nGI1rnlcD0TU/fdCgpkTwcvs2IA7dPfJ4V/uFvQ4lr2lcRT+DFKDUOI+MUlOCeHPbr7qWvkUA00T
6bqCWeiYs8sAzcImkHLE9qJYWRGy8PtH2U4FxwvOYgpMHT/1xZ8VSCOGH2z4GY6hft3H80q/dk4W
ZR2wtcZf+pVxKm+qapBHovVXwBO83nphFHlTrwgDQfdcgPhPLWg8tK+/ShABRbopPS599uPzrDrh
83YjGLi4b5o3IHlgqBWlxN+ZmW6B/cnPfaJ3JoZTF67cJRFOYWS7XtJMP/zXEONqpfKqUTCDyGrk
EESKEvauHBbZEYG7t7NmPnWC4Zwb3tIxUke4kTmBPnLavWUpOKomCYnwQtcBA0uCjViK3+6iBS+n
HygKb1egSg06kZDm9cwcM6UiMVWCYhgpf0h+DurDOW/zkozDcDHpDshZreGVv3J0QPcDnptf76zt
k3a4tlnSicmZzFqmsUy5uoLhRle/q9OB9b0lAETPyAoiX5MTOqJokzvpzzVLdBt01ltJ3BcmSPtc
wB5LbvtClog1IzknG3NXSsWHrAoMXQTIqM2HufVEjMmi1zey1KFM667UOHP0RmwUscBCWvZy/Tn8
epsz0XuniY335PObPyBp5YC4ecIsauATumLLOqPTbkT+nW3idS65jV6bLpfh7gkZ3ON+iaxakwy9
uU1Ydn6JN2Fi9JA43qHKxEdv3q6zUTGfWrmcIl8I6Y6gUXT14Ac+RtYdQFwW9F4OBwyPTYO4sv2s
5KPgkbx0wq0V/1LbhhPpnQP6lniI+OXWRGOB3YFX7H4N+30sj8E9goEfHTH2TjeU6laZPP4eWjlj
vJIfrGN7H8nDKiXIx8S2wwVEPhGEGpuLa441cqiRQZpGvlac46alYitKd98td1Nh+GJ16EWPER/W
VUaVKbcbubAbqd82eFsjBn7Kft5POQVhS9kEfKYLi7cb6x384iSJQafl8fsaZyxh8T65D0gGwgdS
uaA1UotYpeYMb9+8EYDMTn65G0Du4HMdJKixbOB/QeAgsbLRLujMvX1CBJU6i5yn1QYAiErubfCJ
1cpzQ3OE4nhw73ZiUvDQjVQvvSp/sGKUM4QgSZnnqgQtNMYlUOKNkU8WqakFBRCyDUf74AkoM04/
g8E3r6mCJR38XhQ0BnDbDb+ZFa7t7Nsd07nTseDty2LK/BUzCmHm3FIxQ+zEYOLQzzTEnPR/n7N1
gLPsflTFSGlvI+HHfnwkoqhJVQQNOA7HW80IdO24MKphqi63Q54b8S7BcRq6eQEjdNFBci7ZgQLd
q5DI7/nrlAXVOnIZFHlOHghvVBQat79Yn+qbMiUD/m0zipK7Wd9vmWhPnDXOWuR7EEYDuu0GLFCI
2F4HqpNxyjkRIA/FKjshi6AYNnjhC7FdoZQSi/Bu9uGvT6eI3oyXyJCHvaWP5k+UpVs2cb4/FAdM
dqJmsCqHQ7yocES0fVPAxLeDkQbR+bcnRCrzf7yqQyNBM9kU8OKhcKPttt3cFQacZ4GC4E0Ql32/
nPYkeOBF9z+Rib/UlVNniNYlpN35Pth2FdPy/wrPx+lteqGVozhjy3q+g+NELVpdg9BwOrDH06Xv
FfqTXASz1KewkQI5KCKJkK3qxCoaSBB4oA9v6EENEapcCMwfKyWeZAGI+JwgsDockjjfiC8AViAS
yDmS0SJQMjarV2EIcZK3y8u2ATqnbl0qxPJ+V8qt+JYmpWKzof6TpmpavUImxhrNJJQhT12//CoN
ztikX3FRUmBv+zdkRsWaw+GpSAbBon+SsMs3TEcYXDHXgmbglGx4YWOwUsaMYEWmeKvo4snwPEcm
dCWe6Rw9OzNNuw7TwTbWPr9iBMrzhOSIempFhnH7QSHr5DEQun5LOJZjW/tx3IsY3O0q0jRC9kE6
gqmFKJdSK/KdP2C8KEk3blLf2aiwZWQNakvXqlPkORXHkQwBdDS3iJ0fN4XWx36lKrYLImBWlvHD
7NjabtutWkDa9+3jYDMLKzVRaQbABrtiv4Yor8bwwKad8eTMxjBKWpn5hcjS2RQOpi5MQ8oAmqT3
rxdHlo95KJ9VzrnIaSn5yCYgjVzXl0CYNs+GueD27RhTbB12UIPP2RiCpwGdzfcSOe7+OspC2j9Y
q1sdtADOqJAZGLB0XLm6MtzMXo8GymFR+glh304dOuFyYVJEQG2+IeXNXJOnquN0VYKPyL+YGySn
RSeQY0Kv89gpNj7/RQ0EcWZ1Ib7C+SyNrCf9WlahtWLatScIiNgv2H2Aygwjvr6xKHGZULPFzj1t
Y+s+qTuTpUacnfO9KrjBHiEr2W+imbXy+Y1j50vQv/3Da4owqJNAAiIiP19T9qlvQVrRXjqojOjS
iquwi7IHtZD8vkKSkTZCcdBCcxCz+DZIF9IpAMNarrPFsdxOlQEF5F/SDB458DnP63JIocUR6EGB
w3fsiQPCW+veruALT2/REwv35vRp9kjtpChM7p28Xpe9JX75DyWGCpOQkc6SYYlp6hvrNFGLnw4h
PQ0R126E/jywh2CmTiUEoVTyeJfkIHU1dmQDm5gwZ7PlCRrqSanVLR9qEWQsD59+/ThPUrBKwWeq
0vdPB1xdJly+I+bfvEx/JwCPKhPisRH5v7gTLHyYpSQmCA8/XJlepEHmOqF7tEq3gSnxI7/3S2/G
ZzHe2upCZ/vFMPjwxW3srZTGYTbYNUGPw9TsEkJmgbshDKPJ6Z2dKN4vum+BfsHmP4PpF4Ig/8kE
gzrma+GYlHH5yFqBOfLtKDlqoyZCkUnKTSVRVvxYqcZJVRONUBsPgzpq/XH0jjJT3c6axCp3G8h/
N0Dz9tPZnfBrBiL3x85903AA+4OubiB9FSuiEgTYWF+xQGmN+T3T23ZVz62DxHbU+CSu7jHdkTgU
TS4Tap+HeBXYa30WIShJHU54DVQjIOxSIw9coHEFJ6DEYa68H9oKg5GmMtdZyGivZbgKGJFV2hAH
nrdJ0TTWDlEnZxH4wZ6uQH6cgCF24bwGOVWRS9/aBbZ4vnQgDbTBswVwNAipbIB4wnRLbBKYN5Nl
Zv2kSKaa/UbkzmOmJIXFuC9H2tATufFvvkPhfZ89lplefB0L8dPnbOnbqiJ6PWITGak4+hTcMvYW
IhWVL6lzCvwTG0o3WgN5bu8ftA1up9uZZfS9OmMpkM3Z/TJomt3K+l0O7AUjU352vNJayLzicudn
1fdYm+5FcadtvJQtBSJYcyIt2PbIEmPCbOJIHM1gyilB/DWklshBKp9jcgS0WBdkRZVx0+nJHP9L
xAOgQlXfhKWmYOrphPFxAPCA2moqiqeX+ywYRcweOCkC7GdJPznMOfGhbovctn0wL45yDtwFetZ4
xR9ma/bDK976zK2XfEHp1VppZjnxM9gh7uyR0R+0UaI2Zx4D3LCyPnWxDjEkcJcPDol11/df9lSL
9Pd+9PDwf477Pvn9AYe6TIwGYtFEfXsxXUq/w8gurzvRiUem8h0U+nxkRv0t9RB+ngH68WKPfd3S
5iI3lgGOkD24iJp1CuxXPdLsQgK0M3Aaqz4sifLmLxJ5k+a2a/f4nPQEJVZZWMH4tpovQwSou5T4
gUT0Og0teMCdve3xM4RSHX5W7PkXaV+jZcZQJKiPlDfWe5XDXPtMpKencpGSXcWPumP2/2AVJhaf
z7B2NMDEcVxeWO7GP036jSdcC0G57nI4wE85l0nrSButVqzttsyi6eTVF+WfjhMvbE7khnB3o3+t
uTbEqriSqPwPN8rFrHl6LG+1ZMEulr7ic7vRSJHff1s/oK3/T2BEn+C//Znc3yFst3vuUtudbf2t
VqOMAVxELZTVounHKefsyaJYLbmb+Xn2sN/ubjehMMGVHQ4TJafPKUnbU2e57EFPS9TARfAoEC8V
qLAzF3NB8yUGfVwjR8iBpXyAXNOlb2fc7FcXawjHclU9uLiN9R/fSM9Mza3g1WNd6ICGkMKuPSIr
1QmG5qv082f+GnqY6Kr6k+kCKiuyXv1lY4LZGa2FN7HYpiz60eKSnyVhiWeSqONZqc3ogkVFhd9W
ZF0Y5EPeBmHWcUPJSXAW+ONuJj6zbHIk9djmR0c1pm9wlPxNIjTcgzLbjt/wteqBzIn7v8gHTtAo
6QA06ZOE4zLTXXhrTeNOjR/oqcrA1zlx3JdmnFMC8J86mKt8ITh6WocMW+GbkErkb1ek2HgfXqNe
1I0XsESRsSG2cJcvO73f9/1MrF1xnhsRNY7ooFnPYrWObu/JvdZJETF6Nhq7ibZCzfCOD0ehgZOD
YuBxUVThmxB9CZpebneNd5WuAQnj5okyHvs77IAkvQRuI2YOi0HMgpzyvBNh1APZlmYR5q71J+AU
FlYDov6QlAOMdbrl/ozMsF8codbLXF3U80noRwgxDzguIVFcfGcn050UE645OhQRCTS3aLwJ8le2
kgS4k6ci2lnMh55UM4f4atWCan5p/6e3HmUpbdHudRrB9Pa/Gkpom2hki7Hk1nYpTziwXT3EYoqg
6YMQWfT9DtrTOkTPiuE8WGPAOWvmPxomxl8ufypezVS/SiWxeeXjch4Pf2NidH1uCBIGHw9ppaYd
zBhk56bBUF9vXOI+hfVOc6hzWc/JPpccWQh2ftpUSeqH1rx1EoLo9t34U9JkxDtb5c1w2YDEazkm
9gQN4pCLbllPw+KkUNPHpSMB9Mo4lNrYqqmEavIzd0DI7hTuv/lT0ooye3GGuNFfIclnleahb7ua
DvfhSgQoc7vW3GO40Q6U6Sa+3+YuE8q9PIfT1tgeDeq+7gKRolS/qlkmybcLSq88nWoT17ueF9s+
iSJypsSM1Kp4700oh0bvp0J6US3Ke/ZBJPgHVdDOUlnGWsZcy6Ih9ziJSMtX8IZJg5GPrRkt0bQ3
iOIr0aDbvU2enyH4k7T+WoOFJWKzCN3+R7hS2T+CkV2H8L8+8JVnKeLuzcH/R7uAUgTmI+lzsPhx
SH7yYHwtjCmC7OlVjmxMAmTAGV+AcBuYq+6tacYTtNNOw6E0tSLBHpAWAJCoVeJY6L1GWx6F2krt
EFugeMD1ebSFkqTxDtsqDcHISZiTPnDOOOmk9OEWdSp8Q94MtXDhM1+9pZs2uNUPkTA9uhxgT18S
ELuLZOMDJMFcB4AVRZFAUwWwx/KMr/PZgyxHy31D9GPhICuHbAFiQ/jNk+Vac4AuafVzk7CcHJPr
cTkeMB33yPJm12rtVZMNicjjZaIN7U4bY24wtlapED53dYX3EbokamFPy/iYjUU/MzK8zgeJnwXV
8QNaxieNBbJ3rNkNj5gKZ4yZPpbc73IMAw/SR06+hGMgcelcreDZ5vJU0v1qyuA/UJQvl5VuxXO6
w9200chbQQ5d72Lzt6jqkX7wqtTRoIBBrmo2UmIPYzsydkp7C3ZMGF6Liyww0t/ip2Gsj/r2Ap5/
04HdZLkUxPPqnzLWi6H3KNGcL6EZPGGgBnItx03bjWtT9rm2fZTrwICC7huwfrbbdaBy27EQopal
dvHwdKBBYtZpmm5n3VRA3kiRn0J9gpwywoRKBWlDIiLTqvk5yoMJOlORduVfGusGBn8TuTv1jDea
Gc55l3+49h9hbSVw9DpdaoPEafbncNv43C0A6Z98YY9ltICNNjPdfG+RIYYRfzqFWnYEjL0/ZyW6
EeaR9172WJcFNf+bx3OS9OdAiOf1Y9yROy8kSoCJOPmPDIKejRLcSy9ctyHb0d4nJulwm7CuoTHO
XhfiixPJJ6AMb81xhJuqDh2WKRLu8Lstxfw4yUVklYD9EHIjWcR73+2apiYCknbbW3/rEryfwPzV
U848vjq22vM3hU/trcJ9SQXsQCLxdU2YAxneI9LfjbnicOx07Lbqf9nnhm0CTn2e3EglF7tlvu7m
RQCzZlSd0+waCA4bYt9wLwvgdhCDxazmxElirGMOZJZVeLIBPWsyo2hOE7qNH8E1kccUHd0E3/rz
2feGrdIdpAO9fvqjWodMcjoHScxGwj1gGhIlDHgrzpm8AsEWQ1qb8XNuZHwuLZKbkjTGCL56314W
jT24GlA3OMwZg5Se9sUclstOZpMNYHo5vyPSkXHXImPWxWEWz74IAOnfVlLX97HLXpGQE10Yi1MJ
HcPWn/eRMT5O+9ggJfaMY8mQ3bDahrdzg2OFQaJAFvLUsdgJHmSYTlZElgyeHGxnrSerCoLMTlCy
CiNHXBisHH8SqnE6jYwUittaWTpjTZKDvGxgLWvFsR2LHcyF1bcSyD4EankTZU6XACF3tTWrwM6D
y2xqzTFpwbQeD+OM/S/ahtG/JAlqcAhVsSEM/YzeM88BdXoE8Fs06VgfQ0v9AB8qxHyDlo+GsGq1
8RAX19Wm0hyAbbVvjPrQ03dctR4KnoFEHHac/xJL9ngMKNTJPUJOfmn7lx2yFBK1Xl24k1QkLJgB
f7IPsIjO1KqY0K6DAcl0B6wRNSnU3hGDufFXjBuxyEErT+d/kMLQDyn5ZOaGmGUkmHFOySGVBa7P
4grwtWIkYGbJS2JPm+tiDRj0O+nVYv2pfVITCUbf8Zwq5hmIhP6gFUQ2agUg/h5I52gWBrvtAH50
o25GMB6BsjNRAEAteA8SlSoQY1gyRT+DyjduOOJgsSL7nW9ksV66K/wqR9JWZeg5ViiC6bwI7EeZ
dKEuxkaKKFvkNGWCg6feRpBghmS3Jm2RRnI4//VE9tLVpMc4jy6JG2sO35NNtoTCD8d8zR2b04/o
RAvML+oMlXcwTEEgtyK7QN2tYZuelDLAVOc/GAau97C71vnHI5lccTdt/CxajC5gvi7hnFXs0BE6
DcRJRjWEI5ATLIT8XBoh3+2d5jDpqBKxaVaA6SNb/T8b7/qboAVX1DxbNs0eTqfJE3JvlL5cvT0Q
LsPhyzX1nYhYhUbFcDG/lLwwRL2G8ayy+nCQO9DsvMbyzJhpXhMFsMWiycGfEppmKIqF4Tnv0oaS
VGGY9RbEaLPG/YnMEFGtBXnxztd5CdkC/qD561TB2QnrY+9NARoLByEM9FIN+O3zAka5CAw3/gjZ
MKFv3VF/an8idmGjFRrkpocRWLAyOLq7RAs4WBMc8yElDsPXP1DqunQWZBO9sQebufAO7DBjWKNe
bflcuBEZ2FfqVfvb0wCPHcP0O1D3jLNkQWmhwg6kqRd0T7hKByzxA2YGrgMNoJ1NCPQXGY50LRBn
VWK5VEkD3PgOatgo1AKVZwZ+uC7aHS73dxg1tS6yYZGmBmsy2tkne1RktwmyA2L4vjHyENuOsPdN
dA+7pDRJGarAvaQMDFMGUuoUzrQLxitv5aJxExZxT57KjyONvf7vylYqEZ8QKHqe7tggPITSRNi1
NRVPEN8MCj8admTacsLqO2ajs7T8vaVbq7ssCf5PIJgWq7KGpKu8Qcaifx+Fv96n8GWYCiYmgGyW
ApBzV3/sZztX+2CK2mi03Ylr6YLP7P4stzfTmsZxM3MnJoY0BH2ZeihPmxbwB9bhOkzR6cP+qo+b
pURIglxHUcR44zGQYFhBxd2zR+rYEZanS7KGk7dr2ME0DSyJR+2DFOFL43iHda1VsUwQM3FJ6DrW
Q7F6PhHIcXHNscG4vsAT4s4hcLn1R+J6VTOdo2Uz1VV1xzxHrObL1o6UitOtBqi0Pc7AhjZIIgI4
RhmvxfPvGeRVgUsZLBHW1PZ6N3/Ycv5MW+/osnP8P92dOTkvH1gC5YapHTz6rLy3bpbA/1pRem0f
4xP2OxhDCAVIIOBlW07agLLOTeeYFFwYMzmohUG2AuM3P3JHdjlooym4OvNOcdo+8Cf4EaTNjpeW
L3d2hE6sxYFTKTvbt80CPjT+qBtVppCEdbaWkc7ItFzwGPiiJBhnrnD9ffeF0F6D4km3PpSk8Khr
DLk3Tzu/EKKVrDJ96maBE/oBCT6lxBAsLuBY0GQ4v/E/llSChZYU3JE6p0n/lUOcGaGH/JOu/sqF
alrQk4ciHIIgm0ydURkiuDuLVpYUtZTFkT4w7bAFF4SRFx6sEKIWCYxwJUKp1wDD7X1PLf0j7Vyw
XG8QAyV3lP9d4IQBtaJXhQIf2XbwEuQU/5kG/Hzo1MtjM3C1zbi8an55pM1vJpdsv4sEY4o5aVnc
33Lr9Z6yNqUp+mQjj2madaY1E87qSi/Hy3IH547hl9SFvDmz/dGhVOcJcWS02iyYs6oHIRte481/
ne8UWrllbewzg9NisAc9QN0oYwit3j91gZuyABrv3siXG/IVBWWRFIXK0bNnzh/08AZK31QyuEjx
aikNFj1XXzrzOTLMrJMUITnvs3RrPRR5MuNbyldNzREPKebI5VLs5+cDpM2HYh4oCL0zU2pT15hd
p3Uh9pTNGENL5wJcZkKgX/HybPwXkSFP35iKny/GmfXnUhonOzjOSgb4e3E+rc5NbEdguvNy8xMb
TPvEsBZqCpz+zLwu3XkYYy9Jim5TMr/BegZeeNNFGD38esVMAJQuFBUe465C78EDhZ65tBmc+lvC
ThWRfvlmSYQ3KUYhNg7fSXjYbQwyxmCaz1vm0uthFiOo1q+C9BjXDMLvSq4ZjPEF200ovznzvh6i
VexmK70PqtZJgYWkpbsgn0ON6yYd4yaLHFG2C08kGk/Cu+BiK02kePC9LRlgnsfM4QpYQd+l3Awo
VjQdWHIbhNbtoi4uX4/OQW07ruJ7cWmRjgA4OVErL612YlWgFDPHIy8pxc9EFjiw98MyHkVAnNGR
0WwXxidi98dJ/wAt00HIJ1NbSsx9Jpa8B7j9UfA4LVIEZQyc+2cL86iwilF+v+0F6zJDEhigthX+
ejV7GZlKVEUZs1CC7GnVp+Bi5e6qUybGBqPCj4obM0wHjD6eAbcppF1d36/3O6+hW7bJyahGp+YS
iV0acOpAGF35Zt/7RCoWhesdy9p2EcUUFuilOKFag8ZEenRUkabC+0TL1RLlC42XtP2+9IgTD6M3
j0NOJYvnvNxnmwmrusl6IsU6vXODFuKRd3NE1eSY3EiRYR4U5ncXwDywiVQwuDLR/nl5rZGWDevP
tqMbAitLVgc759VwCyP37KzGh5A5SKw2i1gmeY/vqwi/eYRsM6yc4vTvF5TjvI5ifn3oo4ydOGcB
gU1RbNImVK21dpXaxmYUW3uurCNkcbcZ/rx17V07bPs/4MAWvgGUu855khsnGztZTuFBA4JJZMwc
9Xpd7T4dPaHmI52XEdo499yLhCHodrjUWn2lmqEjesCRI8HkuKz+Cmo8mV2XobFb12C8xpDMB3hE
jMLsxyAN0PmkM5pEMHWUvXARBGM1EHkTmM65gaqObRwLBGfeCHrNjOBiB9snMhs4KfUeafoqERjp
U+q/omT87LFlJWEnywJ0wwhHx+aTqW9Pt1qheQiTemR+hUPYokFXg7jGJMVweENSzBUF4Q/C0BZT
PWFu/wJzEs+VcWZTyJv8HaTq781Lk9iDZf1eKZClLYu++MqDTjc56aqhkPKsH4kFjWs+kujfMCxC
WWVkeQ/fnKx1499IfHMhS9kMaDkfnpWPtXGV51J5nKi8wfGRNHqlZr5G8Yx3m/Mr23Yt4wQhGou1
Qk7dH9sMn7YbGARulmYAOzZEEiBSsxbpGTkNeoYtVK/osrd8BbBUiGugi+G3SxmZmzdddC5pNyun
2mrMojqIHy5Z5T49p1x+fhaR1s9AYb8Sk+ewc4903vL9iwH+5//bKEiEZu/B21qZ2eSe2nthZe53
JgEMWy5LTKahY+jQTy8dhzia/ELfpFm4UyQxpxGCxnYQchtopufeDnxeaoP1mk7Zm7+k+16VDRBB
j5wnl0BySuBHT/Axb3Xom6Wh45vIdeL9SMsY5S2f7Cp9WF0TrpX312cP75SuT+kNOn4PdgddNktQ
etrtHuVZXNX8VHQYFXfOL1pqd7WYUxd918jFK7NeMynUcY6q4hqWYRzED0NHGueZncKMJO5omvgm
e2kDbh64l2gh63lrKhmU+quLIfQ8FFf/7GUzO1NJcUSfLDf4/+e/j5eS2KcKFzaL7kJYnIkF46xh
JNa6jJN61PKsXUflJuya5zCoJsYnCS9q/3x1RFTIQ37zxQ9HIGOxJemBihY53kui59zh4k1AKH9Q
oj0dGrPwFGO6r0/oAxZ+aLJr47cPigy302SX5/XVMfLcIEIyzYDXKRPATOR0oh1nFZp+xDluk2An
JKsjjihvBRuOFPthlTgGa9mIDT3DIray3HpLhFLM5IuCgtQVGMwwzx7GjEZWyWiUds5kodA2i3lh
7skhPBN5b48QwLdfD0TAx+5EKJkHpFxYnq/UQupdZ2kVKrxSE47EpTx60o8ix0UGJOXQNlGWP75n
B/vU7QYRG4JXoGqqVb78BRZCz4VK/Z9n1fZRj4rdYlBjzYaTFnq/B+8OeMzetKz/k/Pu8DFbWirJ
3K/4iWuCYbAh+p3fa69ulxmpJGbDyCIqKExqmLOnqdf81GxmtmumpflMjuOTLvNnNCGGExpcNxry
jhJTpGvdiBxGvIlUi67EBK10l7QL1ERXQ/eweHHmy7vp+Dj0uL/ZgF1Nk8XxzA7lmPTdwGzkrd4a
q9ew2igFWGw//qMRrrEmNE5pT32IZ3DzpjENTgzzy0X8CK7/YjO4eTYT0EqE5RgKjXGQZESXZozZ
bx1t2GU5VQW6JVWBDHR3P4gLDzuBMLv55CuH5XPlilBLm/KXCTLr/V/xJO87keAkHkm33k2Je2bx
BL+tnCFYLls1ZJH5+eDOeCpMeM1ifwNEt7OkzwoUUXxRfmxEccO3Iq7vn1x6xG0ehMr980z0AX2r
BgbvzjYmWT3WGXa/m7WJ5HJnStY7jZnDeel19ivLuiHVvAKyEztswuDHjCYWbARW8LHd3aAlaXZg
hgJQuceYm+boqP5CaBaHVQw8aKrk/Zly1t9sxTiAIvFTjDMrdJgYfq0Q6g+6jbE8+womm4mtCjO3
Ui8WOTesUjQawRXydoEH4mNPk+UMaV2H/r66ukXnh/gsNAAJnnHvySaYwPd+qpyzu9sg4vKc3wau
thnsljPN8xVD4qVN7zXBM/5lBJI0afmuEApBcB4md01TUYfszUvuBV5EO3lIkpmaQ7XRXSwjplKS
11eqsK32DIJDTCxzL8q5NoAEnP+AlhMLnpZYZ2yffvBajT1IYNzGXa2kk2XX4zlJb1NYChSBcO/D
pM5QFF+3n4lib7vtoGLcQbr8wVx2es9N9EgIu8vyBvYmGkfw+LfjGDaYifEiFsCrCQRnH6DIX3LQ
O+972dU42/r4DjPti/UGz97qqIXYs4y8RLCnHW4m2P6pLae7sIAzGEyqyP2nuM2OFtIDcsb+gD2Y
PWOPXGLZF1n/Tnnztm1F8RbP6fCIhva55hRvGuqQ4sqygBBqdj3ZBLQ/1OgMECSPg0u+3bH07ySE
FK85NIUT8Cclg81OEvGa/zcJ2rO30hoEGMGNPPATwpOT2v5tNirQfjeguwlVTkZSWeSQZrpf920/
FQ61ScxkvXyQ3YHdGO5B3xPCfipLeSI8O2unTSH5GT3RkUc+61R38pFLL5y9O2UiwghRzblT33MH
34dkBIC8PSBYVF+wfVcvbFomS0va9rZNSz6Xlh6bMqsWoTW27bS0MgA=
`protect end_protected
