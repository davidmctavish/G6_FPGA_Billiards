`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Q/0JcanrYN/RnPh65FxF8+TrVPIxo0wjE+s0dO0IGxk70BELAsbas6mJHK7YoN1Ee0RI4siU1JRM
RGhPpQfcqw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IdJm485tL8D4yYCTCtKm9rkIWSqtzE6XzNH9XpCBKosqSjr7GXW+2mt2JYdNgQ4ZrxW0sVMEk/KM
JaL5bOu8v7LpxrOnmqNttglLolmnK9yRUMZJnkF/MbLpbn/d+50AE55Dm6I18tiVFOdN0gGfb0ZK
b70GazgThdBn3jx49Ug=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Q2T+jBxEUK2J7OhfZmaY6UMx7F6nByTOZ68/ubVU554p0PCkKsj+56t0z5IiqqQXWwdKfmisUtLD
3jOga/ERXfNsvE2hyMVbQcsO/VpKPtu8SmSHIcMhADNrviStkE8FkWixqGw86BgGt/GvxwLVV29P
evrCpVL76Rxb78JyPcHMXnLbOV94HMVK4l1xRg+CgNrN1qUW8VTXbFqwF92bjCvXAcY6sn23HubP
5QqAWNpgpEiW0iaJMCAjUR0o18WTfwvONEXktoUXLQINZRkEKqjLda42qJ1/rkaeAiKvZ+5juZsL
wBM7lXJ9ANU5brX2tohdcD1glfPk/Eo833qxdA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VVr74oDMypvCtlKdhyv438dQZ5FQ5kLOw1yj0yaa7THG0kyDDXp0XhANnSSlDrgBcjRm7L9hfQrG
ZtipkSl48oKR5pLPXtphhqzkOm3r3sVyPqYdY/vJlAI1dYSunyjXlcWdSkK/6BAJ9d1xLczHLKtC
6zMKCjQkLvWKNdfmgfo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DyX6jl5NH5eMcsmvmuLm7uvkvql4Ob3lpcGjUbtqe7l+mFUpbJPlUzBIJrwTrBqtigCEWdFt9ByD
Uqel8trtgfufY9+18ySenlPUOsgkQBfvJmi/F1GVvc0er1C8w5A9d42XrLavyV7TbsDtZbxJsOeJ
2NHVo8okOEp03LZ7dV3ur/5tCNDiD6dbf0Mh1GSNoKEJbhacycFxoyS+eUS4lMFrf4I4cYGK6ykE
cP2UxJhc+US4rQ3NbP+iaUbDOFiD0BHd4jOD7sahTFzuZ5zdh4UBgRNJg7ouBC/T7lokROt1G4jA
p0bi6sh7tx7D00NbRaNH13p8mIJQhfClKbnfKQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6624)
`protect data_block
Iyd4kJpr7HkHtznltUv8inrnFQN3NufgcsEJxtY3jW94ZcNa39t0RwOzZ650vTtlylf+HcPvpPTA
/Lsbdf1g3Xn3em1JyCCiqenxQrtnZ523CZTvo+tO5dSiNSdl+/AmdHyE9Y1Z1drlQX14bpmAhVC+
PLTKYKmAU9ig5E8wss0APZdr8Qwx6eLwJAjNflQqhUK/U2MVNNzTBVG4QJvwK7Qgp8j4wt8GrTuD
06lX338xonvJzUitubAIOZFeBHWbIk8fwHBrgn8ik0YCsYhk+8Rm//48WWNHgY45WjvRbJbreu0j
sNDW/R2TDhs7lboIKYRtaO4AdIZ7fJ+JDagJ4MFKyDST5gFCIFI5ha9MrNuBFsHk/ex9vDwb4D/Q
U+wXCL6Pnrs6oqNPeyV1no4haoyz4DrfCmHDfp0pa56YAfvMOMJOeCl3rfLPEX86M65/HHNAttEU
o1fDw2TT0/fZl/rnoszMZK/1peQJlJbIlI64tGw02JioCHgNlQxp5zqT0OyCxryZzTgPPSJrzePE
WWqUnvr4rYk6UHW/C9ixMF3d9Q2XP2UX2mSWdUQsjAZJaTXFKiJnaf+93PZujkbocqfqoM34872N
E+fkJ7oglqXaO1Y8lWQjXlG6+G6WbasvSCj0tuA9XFaeV0US0xu9sVtrXEo7LNcx9WfTI/1WCM0D
M1jvBsSy6WGcr2lf2Ehh6iQ5EDgEjPp6QSARnRVJr4JHwTfrX2AS7x6y3SNscenfXOOCxB5FP6rJ
N0xTTC9jQciYYRXU1/bxSxHDJtEJz5JHUE8+874I/NHZ8Je8KKYO/Q5eIWWrIY7nm1lmQXGIguJV
vwNFtRfwEBnpAC+nQfg/ZXb7H6FhtNu113hBU7hMirhCy+0odtbEKVEEdH2ADDHY2Q74sEE6hbZ+
PErDeHWIVSQ5NJ+MXZPXrGPwRGmXowm89+bdhhm5K5xWRb+kPytXXLTFWBL2t4aIdUMza20kxYFJ
hGXjsnrIUOXLHpEhTA2Bh+Z7Zz6Nu+c1aesGH6QG9VdQYhP+9vczcCiDlNxNi1+OeyeJ8VECN/iv
EnxLbcpmsLY6OzLIpaZ2KNI7cPzhwyDxARJPqJy8U1+mhtdI++lHguAi6fsIu4oXGxILnXBUznfy
FevbNjuJiXDv6JV0I14BTqtTFIC3VhV79+ejAZOlOKs6oTwm8T9GIBAOwvfU3Z+jsvZtyrwr7qtD
mXOzmcIHHWawqIu13cXC6YOKk8AcZTlBe+84sXQEPo5Ej7w7T2redfnkp6VSz1MNHEUE5NYYYlTR
1a/Qep6AALpjKfLkizvcWeUCWFGa5fYauCAtNTmJHsIKeOCMWkfYi/0uqZC+/gWJz3NUWnU6xZ6/
URje7VWYCyUHTBR1gTLei+v0N2ZTHJFpUbTOAv2kwb1BcQTZO8QVIl/LtMOvlLAm73YxrEbeJgUZ
e6mTWjgtRMq7Mowhkv5MqB3kFu18YXLLCJOhhpNS8J4SqGAYksGMxooPIHatMQGeQUhlSx+bnQ7q
P0rh+eg1bNoYQA8o5RSQi5WOFlAkcMfLUnroMkvP+foAvOGxFZuyQ8XacJwzH5Uxz7ZRDF+IpnKM
ODAt1ShtKgYbIuJevpgG7hHywHJkXjIk/6if7QnUGf17rBil3iATuFjswC/M63b40U5EtfipL076
MPIfAM6YfI08CxELQuJ/1+w0UlukFtHq8U8XcX7HafLWO+GMGvWnWBD2BBq5UY3SCkP0IFisqyld
KmnnXVhepyKx4mpnANjA2JRgzBK+FFZgUB8R/RMzIGO5AHa/GGQHSvyG4j9afHU9Lgym2LHqcApV
Gi6q2mniX9ba+5CTsTTEYO3LwlySf4bpmCYgkggGFusFxIkQ3JbmNkXnDNrFuRNeLPMkHhgOPeRG
NjgOYAgTdf8shKER8NtWg8SX0V7WEwczSpHD+KXnlxXIMmn1gGz5FoVWCeqUupkDrRPO0PWqvBWu
O+egBICg/OCYpifAn1F32ucTEZxObs5//IPma8FB1G+UtPeAnl3RnML8PgrdImrQnEOrehFNui43
pKlKhm/F7YC/IYv/niVyiyCwWM5eIaeEQzXyQzo+K+B7SAmxg+bIpVp6AelLjDjOmT6cwUeRZNgj
QwNvaLz5Z4vdaZWu3r14NDfCHyMRueN5LEtI38OXHqmzwynFheEbzxedIUMkrBjKfN6A8BX08K9r
dvJWuodGh67m6YXkj1lefCOsSGofmLV2KWuqCOcVrdZx72iX5dllkIKDMH644a0hj+jX5DJw5zuo
2rnjVW1zpVNRuZvoDXS3+QiNBz9CN3cEshlj9xLHieLkDkXKHd9UHJCFUfCyrmo3omR2kjfw+SI9
dc7fWlWPJQ9nX6Vl2kRfwpdW7wx/PkuNUd1NCP+1KEL7+JjwfgHEl9ItmgxCMnsOy2gLQMrYHZfp
FYNOoFxp8nVpY0oHco+rEhwmsfBdAxkxnAsExGdqJ/wVCybUOd7ljASMDTdAovC+S69VnaRbqQ/m
2ky0hdssCth2U5XkHd7TOHG+6SGwgTXN6VbX3C+F5FaGy1uPE2SltX3k1h5vCuL3s6CyvjtSflWB
HJGPyAOO1X/yHhldw4UupJx457lvlE1SkcDAANMA/UZkxRbe/D970dVf4KGwA5KL6qPcdaT91HQa
KJks0XDcwvnb9pBXYsU08pgk68wD0/2cpeexfzW63JJiN2KX1zzo1BXFEVfMvLJhDVPL93Q7hzcT
tsBcx3mlsmQaBq1takvCjPZ8hNB4UkaxcUwt+x5PGCv8WGVx1wfSDjAESZe605KfWRjxPfM2AnKA
FGzb9keA00uXuc8Y2pMoC8fhYnNgM7G9hOHnAyVUbDG808T8cq9EiYVo9sQmW1XzWp3Q4lULsDS1
pDnsUst9371afBjTY17MZQXaEYXi6dmY1y2qtn/kUlE8RXl2ugc00Mdmit94Ty+gvwo6id4ww72K
qsj06tkV5ZZr66w/cFzIi0uoOGDBlJndU0vXzVk+DHKDHP3NXJRm8IrKhO/m7ozRbKwMIX1ED8fa
ybrXJrR61mtSVGF5sBXTTdX/SbdgH3hLyjGP3sJL5uGSuZ+Doe+4jHfDPdfoUZxEUwzowA2jcLyw
urA51HY0YVpVPj+XPJh6Vw58l6SfLrZ/SigNebi9wBNvL8WVMfYpQf1O+kLvX8/RyspmD6biaKia
sIXrkzSPtg2LLZ98+9ykRgW7W8m8UM8VMyOllVjeVvoKPx1fYsBLJnQFYXPYx+FHpawZc69n8I22
n/C5GKBM3rwVz7+1K0BQxBGxdSNm5V2vBGseSr7TSYRb5s01/3w3oNc0s/yETtnee5nF5fQVttvr
ftGVphrmgia5KrI7XOHA5/ylDv9gurNQG7l4PYjExuI9DnpmBtxjNZKR1Da3gdN+EDp6d4Pr4aSU
Yb33E9ERUoufvY6A23woa+fG0VCgq7ii88uq6H2UdK1iCZvhhCiizqPpwmcLy4ejbleXI8GQASUU
F8lRc27JMNu84zV3naE4z/hKMJsCZ+7Wv/HyKCjCRQuSZIfsgPjKiwpLg/yz3NOItf/riIN8g7qx
o+kaFKLWgDLVjw0xBJQ1qQ7O5XL7TstAfvyynlZNLyBQFwTXFUle9uXQjizYb2D5ceRaa2nMUoer
wwyxErE0P1RVGOqJ+/LT3UZljo+fVNOSLMwRGYcfj8bR8VVA9X8osvPEMnnzk7PENrN3T5VU4Wgu
/UN6WgA8kZOcRCOqxD+SdxGbWD2LmB24sKGAcWfegFs7eJ09EX5uYM1o7xpHmwxIbCvARy5YDEGl
NzDAPvNsk1f9K9dSiR+APUTht7RzJJrm1RxANCVXnKTKlj2afudbje/iyrjScZ3kaKwurwwwS1Yt
Su9JTQ9T/abef4hosOLsYCVAOdqWwTIKrx+sGbjqGhUSx0UQjvYvovQmdpY0jjcj+kpD574zY1CO
i5GdLoU6Bwi8Up9QiqW159qOsM/rSgllW+rAWslskdly/Mr8wt7MNhlHEhKZ0rPgZ/qZKNuHYDs3
vXeKIBXbwi70B/xScxjffVESKgK8seMPM7DrOxwixPUpZDcbYS95p5vFR5mz31/76BdJTLe+B1Kx
61+DMDksOnsXBgjE2J5iJyEpSVOEh2rH5uI9NfltawZLzAAN55dJ7rzeCh6N7xmPjVZlN5oOJ6lT
/AXMh77xsepGAmHn230jAx44eQiZtR9NOagiEaKQXxDcgU/sO3Gfk5n7x4yd80hjETJMn7bcXoGx
EQrWfKKo27tZGDC46DnnJoOcsLw8PUeg1NKzvQX5fq1zttHOXrqjPQ3knNQ6+ims6+icJADQyKXX
avI0j75lz3ICjnlSPqTupFIy0/HervvL5RaAXwqHuF5ucvZW4L1JaNaVPzAQUipvRmsoxrw3nSd3
4qxRIziZRYQ05WjKXJRIRJaeH55wl3mgzDGuI/pdklI9BcGTMirskp4unfmdssRFm7JJK1OsDtLb
aY3UJs5CnGv29DKgdbaxqNAQgsin0QortP/1kEqxMxlDI7vUtjPbbQMl0uJcuuv/SUMCgVSsJ74U
eGIL4OyBpdpoIyOshADAIba0qQtuewtpT6dON52v1grnB9c5KVIz7bDi91cDx1c48R8BVQjCIGEp
W4r3MGmzV/wKMVLnq7if7OKLcQlqnHPVPS+kiW0RAAQ6ntlpRf55B8r4EDY06IPlbz4gp4u7DDE5
AZ+nU24skaRqO8SbjWVSwhcUsBrC2eJ95Ma2ZBUVWvEvfpywWwqf15JWHZFnJjq4StOoh4pdGsGH
+MNDbXtC/oBH+7HXbvx+Q3Jc9e+7DdClYSCe49r2MMI4Wzbgvcg9qfLqe8Fq9YyrEE2wG+qVmEAx
u4A2yug2CEGVn7lMsrVWrhD+0wC/QeDuzhJWh0IVLwBZzch8HGZggzaV59fn6ctpgG/0gGWoTDOK
aZUXmKWV6eR/kYmoiZdkIEnJb7w6CHtClSoonhbRyggHR3c30FIPgmjfO+w7v6UBAMI4vvWNJ20r
xyA0Ufb7YWzLRH8nBpQJHtnj+OWjB7Vrsr871oYzYy65WGazDLC+PxkpCsrJXRPkgRr5vZfRGbkG
0UcaY6rcbeT9CtkrROgE8WpnTvLzKROLNUlrVgo8dwA8cx8SfyLHMA5zOG4SMPlwPhTl8gNNSlou
T60PVuzf4TRazUgEjU6g97fqwc+WbDZCe7/WwtunV78HszBq3YIWWcW5E5jy0F+vXeB1FLqxzY0m
S/I0bAAwXemcsJWCzPe9Pnp/g+UFYV4PMlt2tEKgsdmuw9OZdExtiLvT8VeoxUh+qPlDPFndSq3A
oC2dcmOVcGN4ms/L36ezvg+I0KFYmbSz4iuHD5anIrI8gKmnDNe7qWNP68vvK6UtwgQPLY+wqhnV
3StYtN2Hr5trsTGf/QmqgSke265yCBLaKPlgoyZmNhuFVdglZ+WecGHE36CNZ7x9rSWbSWKX6Vrv
hhjIL4iNoqvd6N/d361vUc+LnVtUZUYVj0IvHr8Tf2DlbhvAFXS7WxQu37Dev7rIw6B9p7ZVR8IV
YiDWv2sYcJ6CX4vpNLSFnPSVkg5531Ekq5CZwaI+/k0crZXy0IXJ20DI23dk06fHRcNlr9ZnbLMi
8G05yFzUh08oF3aSOh5pWGCMaANEen48ddH9f3AEE8BHQuxgWumXvazcXUNv7vpXT63BtcJq7ur5
ebTCKOKaN1+HxDgDco20xfHqRt4PW7tDfyjDNTm8A5Ovv7Qjpqz6jGvt96z0cASRRDDvLZwQhj+c
CE7MqVvjtjE29jV5HGOjAhkxDsFpM7Qz0A78b/xv+BLcfDGLyY7mt82gjoxzQW2Kf3Q53C/tjIu9
I0302NJoF3x5Mpl5AszspVpaTvBXBU1YLcblWqn/DSh9RN331G/kOcvSJYCR9tt+1pam/j/szPxc
TjUEir9XDx0Ge+o5QNKZk2o0sPetLt8NIl7p3sM5TxhU8aqyTyW7p1hiw1k7ecJO9ZQyWz72GF4P
/oBsS1CgmgLrzRDXDsTDin2Pv3QUJYHpKxlCCeBN+K7RDFqTPORiKzdm4IXVCl3j5LcFoubwoDIW
MJZeXCFEuhgvkE+Rl2fAzwg/S3LKtf28Zou11Nefmf5ROUy0iAx1MVNRmWffMRRaW0R/1YAkI2Lt
Vpy1oc4JCoR8a2HsjUnVjym3bb7I5b403hfsEq8LhqapTzGA42TZI0fN8/p7QdFpEQfBUdsvAyPA
SXWGV8bfqztjuNy+dD7H6hO7psTL+aH3gSyUe/D/BsaF1wD8EKXd2E0g/PMntkyxO0jFHpjOUpFb
dvytnKprwp2tMIPHegQ7IdfgfxnuT1XM27bRGhqCXgy9UecbtxvQ24rwMeKIXwBc1BwrKeqyQFj2
IpNmVGvZu/Cpx9tuWJMJPD1/8lpNpyjaT/YCIKLtMCtUtLG8IseWdb2v6A1cJIN0SEQnC3yImbBh
6ZWAYDQMdSxKrYZsLeDdRZRBtKh1T+RR9suwDYzyHB8gdQG8P3FJt2OzqAdU77c1eYatQfdbs66W
NssVAh2kRFX0gWyLIZGO9MrGefKbYgJ1Cafrwy1c/FptfoLlyWv11EzMVARaAd+O+MV/ODltMA/3
ui5Nme0aV70ykL8AzlUFo8a55JTqAOK0T+BCf2h29ETFe9b1bG2QzCViF9PFLL3cJgYzPUTm3aBs
1si+ynBNu5SSkAPRqFjhpSb5YG6gmOyQMRcCvvBptdGNGbjAJv1XsiA7IxddO1mZNP0ItAKcSXub
XcTAmi5C/RL8hZD9H0XeCUYQTLZUjv1MHCuuJnYLHC0FQlC/Mj7Mj/i57SBnSFG14XZgHLkFul2e
C/8BTptPzkt+A7HBVEJKPklJDcd2/VuJT3/Ny7RilIobfZW/lgJXe9JxdEPqt2+xMpmJWElckD1c
B/cBX5s1M6qCWf0FkOsFi2t872h2/XEOohvHkzrT9qE2hO6DwAyGxptNv2gbxyWZWrydnw8+zO3d
dWn0orwbCuf8Rg+7phLvS+BVtaln8Fwrx/luFMdkKrf0RwS6cFoFctmz81t+A4h3Wsl7nx2JPAFP
Jg+lbl2BaFsiAh4rIPvuo0JanM4/jSW1vMopJbKQ9k0+YQoRiydLNcjXyQUkpCHdBMK2EP+D7VLH
GjdL/cRE/nlkDnIMXxV6s5zPRoxR0SOgrfNIaT73vyF0dyVYa66qTtDMurSWTnS39x7C8/Wtixig
2cRxLtgOkA2yMFSmkM0el9vevYCqIJ5BrL296iFm1LQCWBhpEer5JXc7zPRwLnChqAjHis8tbTUM
S8l2PkYKYZwT/BMKrrfMDoTcnwGWMyNCRQWN2Qyf72kYCeUtJIitoHkqzUG8lmauc0Z1kBM5ll+4
67YboPtLuD4zWFewXjT1XTiOC3Cw7YLvD+9CERjdbuR1rfc6HY3IeJJW2U7leRfpMp/g9Vp7d8nV
+LsBlCz5n+NkIcuQRjs1BIrta9TUTyUWgNC93VJK5By/u7zHboEwptvriBAe7eKcXJf/OzJzUaFr
E0rwqHG9MsviTbnTuVmwqpgWZHghIxWpFUaCjpRb+1bmB6ek2I0iad+xpwb5DkL6/AIk1md2rOdx
7GPJ1Fyuq1EN/dPkKy1G2cmmS7JLBjKicKiKyUc55iD7HU4RiQOLbOagnh3gWZphDrGzsYvVmxlF
BUgvJWBgF4D1d+OekeAbr+svzxPBTWBLPI69+N4v3xUdysQZBRFO+QDXD63iGB0LLXW42yP5dL/U
gwRClSpRJdfq7TKOa6vk3QV69sd/BPL9IL/LQdwEB6HicBO2DwawP7Jg86pl2QmIuzrATWmzxrc8
4qWeK6PaDmqMBiNjqRZl3W7j1TJH72OslD5C+foMQEjvGlj++6STe+eptJ6TeuReWiVG1Kx18KPN
FkmvAR4MJBPvzT6xqf1lscKZGQ3U+RS8F8Q8c1+hXZOLDX1QxiwC3ovfMMl+FP06nu2Y17ede5Gz
yFRo0G/ePy0b5mFP+XXKxFf3f5TtRo4K1QT7JaCwn3i06R8PS+sblGwIXawshzQIwqZ6MZwjhohh
iGED6ZXHcl170EF5uA+nNgqZH9kiyObh9FSG6CEWBv2dZqLTtoJOwYNYUmLOsg5Jm2hffNRyG9y3
B8XgJseXcAGgavu5Mx96FYS9/H1GJ8mPzd/Kza7Ox56tW/nMbu4o3kQPuExvjDPaQ3DA/rBC+3ln
Rz1/4ZlqEHY75ZC028+idmuzWcgfjKl1OgB1N2/XvllKm0jx9D1t8cUgb4EFTcolskF9Q9/kj7dF
01DeBj2jVNIwfgvRpqc5wDgLT71kF7MOSjyVE4gxWHg/wCIntxvF9LY+TttDOe+a+TkWuNiAF/+P
whCzyOuh0UuRUbGUpNy2wWuNxJgVe0JkBoCd1ZeW4JbKtFWJV/ytSebsGBzNbFPO4BBuux2lh+kF
tm56KG/LwMKUW1H7UOAyhzcBrtJ4fw6HJQ4V+vEeyCsdhvlMnw9stU4pmHMdQiuf3Xg6m7Go/A6Q
e94Ypxg/ry2oZFNn3iePlJ8pRaUgDmh6D0Ip45qJqPHg35phw26D9iQzthlt7LPyu0PCv4aiSMXO
juV6iU+PtlEuo4EiK3Ku+vRsXN1Wbrv8vkjDrrkaccPw9SuqfY7Q68YDNmGcSiTTwhm75BZaIP+O
xgpudzphbEP8rUchCzj3+8gLOeRH7LWepRB2vx2kpqS0yHAMAmkUrVA9YtdfnZLaEWQ+H9+wv6hr
JREU/Qm/S0HQnKhmjicSiHFrUJsQkOnYNJuJboFIyD6LnzPGnrke9HPNCZHllOfH+eMWFcg/Kcx2
jnZopf5n1gnmBFUT
`protect end_protected
