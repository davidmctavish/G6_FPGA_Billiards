`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dbKZS9DYc8Ip9WWTccTbJfLKzOrKFJ6Qe5yYxu/5SgHRguY7wr3/n4FJDxW7XzvHyqbnC017DaHC
87e8KZKz3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A0+nTRbFluMLOYzw6AEuwq/n2ylLfv8j6xs6yMwsVWfL6tCVTtCtKRxCyYM7lo5CCwaMZkKGM4Ol
lLudJCv5y38QTr/3dS1AwS7O4l8mYhdvH++4tgt62IUKjKiB7prznlZGwvB8liguR7kuxodBwxy8
P3pWSYDo2ieleulkwJ0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fX00ZuYwqTeXTX765rXcJSZP/WM5GFJvd9IeOiO6uKAHgVhChAWJToCurH5u+K3S5deMgbVPwZAS
xDx3fS8PN010n1LaFT524J1T3ktjKlLpBJylAO7jgmxSEAPJbU2LIK9y15OTicrn6on9T33WDfdi
2aOOQFwqG+abjYmNS3S4+Waad9n2J2yJ9bAJNmDg0nohWc66x61Qo0HQRSrQXaV74dkPddPqXVXi
RJI149vGSjm2Rn+kSgeeng2PGK9YTwthfClOsm4o5GBMfY/6TvnG6kiKQ1cz/p+WHBeWrr/7es+S
VBRZrAzAog3PVQJ8awFQBqwoMF1OKyijq+TPFQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mCUKgVNN/Oij1fqDMgbsBFPSgofHl7bP4UJfEx5D8nBdjUUppTFQ+3qxjDEeE9R84/1uAt7Swm1x
Zk3tOFz64v3Zb27EE6x1LVBPp5OkcOddMcOiorW2OGEFpx22hhkklVTti3gRyhya29k4QISwqicK
VzLRyIngy4UEl+orPaE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NLSrCFiYNq9jCJBuaaXO1NaBBjEFwY7z0OCNa10EEPCu+gMIY3OsvgAwR62RDs3UWgY8Rsww2oYN
BqIDdq1WdwAT/0YdQhyDFzJehAT1UkC3H44mOMVQs/Q0jm3VTVH/Arw6nyeVBaBwjS2Dg5aZmIei
RDN+7/DPTuVX+VLKAL1lMD89w8mjrPhWQ8E8AN/vj1ET+kkzrk92Q4fD6HUA+4Ompp+gb74DXp3v
GkgHg3J8VckWbaBrRuJzoaw/Td+N4NJO5BOhY2MD2tyZcq9cLezYFqc4kFY/wPC5lkEzjDO7CZn0
AytmhavbYZZ6bpwWyoLP7OFGSR29XjN6v6v8Ow==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23312)
`protect data_block
rOinUinkj8YW9gTdKG1QsKmn/xtOS4yOGkPldzrBWCA3yNgahCDqMocpldmlp7kNE6IOGiMq0hKW
7xKlxHCfXoXnzRsgEIYcSHNeXIbTlC4rH1cdrbdhz3rdaCxqEkj24Nyj1Eaa/Uesb6gst8n7mRgf
cQJxWipkHn+thscFAwbWYJneSkxtD9zAWC0ihd7+0P5jKvKICjt2P6+zfwaDyp726VQxsIDmoiam
jbkqVsm8xn5sadwhjukczHzu9QqTTyv0y/9nMcQXKYvYudomfO4oJ55X4G/voVW31kx+BedaGRzQ
8qQkOtDYXsQMYlYMVvG5VC1hTzO5kzgVaA5c91K8i95KYTfLrLCs+7HJWl9l/2qoRIqS0DvtKHE/
qNCW2/VOlamqB1QzhQYsUJ6jDGVehDG719euQy8WZmuf7Y96bGmgV5srAma1PQvDaHn6+AnuX1ip
wZhvsxrdGRKqIAscHdd1X0OYGVOGXuqIaAdvTPsC7pZR7kuDu+D70MhOBEpxl3fKH3y+6qXBnySk
f314b0zjcroIDca9hbPBEOwjZu+4WIAofYDiMIWBM3sCgd+wWrAMEbKrGKpx6K18ZdD0txgqgTRo
sL53ehTQ1/wevP2hGAVJ9QTweyYsPuHNF9k3aBiae1fcJ1LVIETM7/f7Wf62/VpdZoK+b0ecsRH0
O9XM78ZXGd5CtdBiM98MywYuY0mGlMlmtZICjYktcSpYzs19z7pfBqE8Mq4Ouv+Wvg8nQ9LdDkaI
Rdi0kUFeTFBRi0QUho3DDZvmGbcLHML/8j0cP3zjUiz/y5N6lWFHk2Ox8pJ6NKOto7/6xkc7qIXI
VjZcYE6m38z9sraUZJUtHJL0ROUtJtey6hNtjJmTBGIiORM0cS9Z13j8TlJMo9qkzU5ICTF/H7Ay
AEXgfofUbeBhwHwiV8a45UktrPXJxRyhYf9yRGuMwhBlOPM1nNrtatMVb6Xy99PFJelcoMZy9GSV
8eXMx7hBaX9YS5zCnP4cgLUK1bRYZag/RfPh76HGfDzYUHZdlFU8FCVel5jiqNqAh6OrVfjP+5X6
yP3pCDyOHXR2rpY3ODlNx17LQF0vDJplghZEoobmo1spyiDTMJi8AuNYFQ5pGvJ5baHeObuB5VZ0
pKJiep4msb+8zFTMnl1/gTaql56ytMqFZ05r63mrHydljnBJndbDWy9Q4nQC+eMBhwrj4ZGZWQ1k
Pqo2wCVV2Hs2JG39gYuAun5fiBGw1GddU4bgy4gTmhl9KYfu4soEzXfqRt99Rdr6sETUcUFweb+M
x4Rw3csfZ6QVXe5KaiD3/GxyAEi0Sb4qIB266tpwHontUoqIwfRV0CrzKdNkXUKO/JTWhbN1JOjO
jGeT5h4ZHoFwS29AbbyTN3rOgMS4G31frWzUQgKUsp3sm3jR2pxCT13qy6KSjo9BGHl9sr4ReN7I
dcsWF3qzm0WOocmTR+wZaAjxFnmxqV39IUrBDBnTSR/+GyzswZvBlBmE5M+50jqPeJT8U/JwzRV2
VZd3ruInlRI6+mx+AyxwsVkdwlINgI8Xd+tWEY3PRL8d6PxTE/s9hVf3bwIPktmuQ+qH6Z6a/Kkv
eb2Wb9aMOZzqh/GCRhOySPhifXYIGOHZ8ikx6wq+arbI3+Dm5+W2XMZxXjH+zhZJh5ACCR/So13w
uDA1TbdtIKnI48Nkk0h2jmaCStNvydEq7fr3I1vLYV+siYm1ph37O9SErGf70Lao8LGxQVEQ2p/1
zR9Ar+cyoYdgWNSsYJjLfO1D2GHBUVNRHqDL++ngOtz8cXNnPIBabfuTcq+24UUPP4WxyfbdrbZs
OHizzqfYZCRP8NgQca5qbrI35U2zcbvMV6UicoVHKN3xmjAESRvnP347r3UTKRpHGZVq5hutACIF
oM9TfCq4cmQ3E/sAT3o01fy4d7r4/Ptu21H91S+WIxP9WmDEyp8EpRgXz6uDb2VA4BA+p7C4ANFV
4TTOCKDOTokFsa+6zjC/HwbmLr2ZVhbgwgUjnX+XjsSluWt3JyWsFb7qDScBxOnCUQ9V0zwf0gqx
K0TjevEkgx92KY67EA4GqoNOWIXCm/gC9UAk5IGVdCvS/iRz7zsINvrm7BUW4/Ypsgi0CPLMBFdB
3kpz8rLoPGYc2YJsE3vKfWrQ4DsY9XCsqFAeFDeJWLFW3viyhmV5s6oZ9+bY5mMNF2J6DpMYf2Jz
wDD/32uVtd+eTlfDFwxjuJGMSuChV6MZ2smuBDRvDRUd1xRx11hD7V1h1aUOssng7VXfU8EmNH89
nDj/QRLWKttMLKSOzw/zD0JatetTSA2mcI3VaTtIsWEJNAD3LhJix1a0f0ii3+lEvhspMKkRQvTN
FVfE8dNeg8ObyrTuTN6M8sO4IZaP5ygqs+3O/3rd463Ick2hxP2A6GcKpju8siQrOJp16JH43pYQ
tXguWgU53d52/9He0k3jK6URxTMiXsZaVgcytVQpZ+nwyzuLPKEst/za/CDZavUYH0Rt48pBdg3C
IXzxEl/srZn5Uc3/dtbgieqV0vaKb+adkkQTFdWQ9DkOHIeE6/74yCVWacjPWx0cQodGDAjSNDHp
gzblc5oNx20XEMJYDAdM3DnW0X3AOMWv60vR1EPWlGQjsm377dpgzvMzikl7CuOSporP65qZKcoL
jbX3GgqKKCV5NW6i5mOt7cAJDeRsm0qbMDeEa9yg0euIpRaq+WD3PoqiMciK/6LHA0m3LySS4cXC
ddqWw99qy8ygAUtHaidDE4cHl9o2EefvgKWdjCKH4QuS53t7Jz/9gRKRFc1jT5iE6ZVjaK0EIwXh
jOsOBmBzpQoTwGWDg1SpG4kYax82kriIxA1LwRdMjLbCNogjSHwV/+m0UD7dh9RHxhCIpEd74MJp
b7ullzoF6vFosLaeThqgwDadyNXuF5r4W4pVjGJ4kf0ynrHO4YY2xJqgX47nUPs8AbdGdqON64QF
RzFPHtMGg9b9MEklaHVi5rVU2lKhIBo2Ls0mpRh4pjFaruhsgNMMr6mMeeMsqV3iWNLph58EBLCk
N/XpMyV0S5qC+0ZrePV9IgzDo3UsXiXrbuMqpN2+XjumeU4OmY7Nel+lEj4BJV8Jxqz+ILHJb5Xn
hC7Ka0MaIKg6qWzeuEPFgGZOoKnQJjkNc8HF1YLIfha3X6XRqfQypBqqRUghjYhU+JQ9AJFvK5A5
xivPYOlYjDNulpAbYl9C8FlEH8ts0xKcTYUZD0BV1aBOHnwKSBZ1S6Zl4iBs0OWutON3XY6gWSF6
9jtsiG/h9uGahQD7QYBQcinK5d5TFX1NJ1vhiIIJRxvq7b7Atx6IxH59ML4Nau1TTitTlYCuZBa2
jcNX1L8frulMwLYzqO/R3znbll6wFYun+23OX7YvSjG65WVTGESi7OJEgURsIm6svNG2BXcv2bn1
8FBXu+yv8E2ooHqkUuIvxngNizwQ8FU0xQVTLWzcWqSZhGWg+NctAF+a/wOCbH2VGYs2IoF3xMel
Rxzeq4xJWKI3BtxIJHKvR05rp0ysLmXKoZZTC2GEwOuE42F2ruSANJP2jRQwZ9SjF+v5IALzM2JC
/mq010fMd5Iswkj1ORIWBx843XNpjdSiqFjuqMcu8YsZhKG281OaitKNKhmnDMmZG0s3pUxI83Sp
yqLgYLA7wMTTBH1qPI3ry9NzZ5VG+tyRFLkmYWrce7k9Rxm/Mx+kyg0RbSPPKUzFnV3A1w+GSyOE
oM8CAhaX+e50xN7Ksp3nm1EN1Eqm6vX65nw97OI6YFgioN7ya56n5MpLKpQTMpXju3W5yFL3lJnT
goA4DaAj0qbttSf6pCUUsJ+9/Eb6+pVM0uWCPs5S8fkRTqtha5BStB8uDb5NXGECuIYA7+lT7KK4
OvC9JDCELcH0KlEyTL7UJANoJ7xwXLR4Gd4NsPYtDxSSrEFYhtn0ijTpgVQ9PlwxVqSyQ6+0Jg8K
Z1C2/C3qSTR9y3PNQeuCr1pdsPN9KO0f397n1sMJ73mOj0BmL7sFXzcZbExfTCFerg6JLbjz2flY
k0cW52t+lDaxnE44YaqBGsb3zBUf7RlSSJj1QAflxOpFvcK+ylQAl95aiM0cpuVgI1rQJpGlkXJW
041FAw/xZ0oEYx5+Y1jHiWQXlCPk2r8QIbgGhIScnXZAUsLYC50C9At59sYcYqjOf+86Sz671v+W
FlWmkKbnbyT9CyhWn+/S+ZURwm4bugdLN7eWPkvIcBrPXqvou2P1HT9lHMJ1RCtGFYH1Nby8tPMm
y8O0aVs7+5LYGeNfkqIRoFqMZNbtGoNGnqjxPiKkcWiuB228LD/MllusL0/s7Oly4Dcrncea91BI
9gX6EwRTH4oK4Ov9r3m9+9+RnnP8C4szlfnSCsrle6G9HV5Hg6MAwlsDx/+eRW2DghZGnNTNNBEd
7GKbO5NFdpA0fPUvtGh6502lKhneVkYNbuzCt0PgfIJLGc1eFOq7NKkAV74VSQ+qMNG0MSW9Q9VN
dyV09JiLd0EJOTACAtK/vnkI7orI5PB2hCRDFVvpN9IMcNFQ0LukcwqWiiIWZLPEKNgggNIJUgTt
Ok5eIgnfbN0e3iv+4sBx2nG+LilWEuqzujWIkd7rOZdLqCE/CiabKEB7re1CGoW9x0H4Fr5ZAQrk
Z9CQcMNDQhTaJ5GceP/BtAqiLOO88wcCMPZw7lEWlAe8GPIjCIFEVhoDJfssrXS4saVhBtel/TlO
dXNolnHT8NTTGV1/USEby50WcztW2STpO5WaTcyEETMkktPBYWG8u71D7W3yW8QxDBxyxM0X9xqC
GbPiL7FhGSGAVZTee+2dF+Cl1Os1OuO2gU5alx4yYbK3AJYZDfUcSi+hPAh130QA0ifQC4TK69Jb
nMq6s2zB7fT4tOeGreZ66/XiSrO/IKqxMB0fHmhFmwTvkiWtUQxyU1e620EnlC+xMWUcnCVM+2tz
jyj++ftay4+BLFL0FZC/UqKc4zlHF9q2EHiP6mwNdaZct4VDgHaNYDw1QEwfaYzIcG2YSvsCgPWK
oI4gZJckWcTy8+t0sMIg4NJeOIoRNWGYh43SuQPsCOn1I0hN/agbnE9zMSxLI0mJVeIiU0xV3tMx
5r6jdnr1u7z+MiJFOIrT8Rz9X2GnDTIwMSRnsUt52uEL2Cf6Bvq/1z6u4a+3CWwYF5aDPhb5fYRi
TSSVOmv8bimtUf1gPTd4j1DQyJdb/2nXju9kyJrXLTGkd98ByINQpGWHpVbYuyQIadhydyAaFp78
U8pbvt/9m7lFbHZmQpYsDeZqrJuVtrt+f37A8hxmAD5weARK/MlmQfm6eH4KoSZCP4IKmXFSmfHj
Kan9nkD2s+w2vJUNMZAZV/1TiYxEpf28ZserD+HkGylhLY0QIvL99nzp5katWSgG96RJgrm9+BX5
T/T6WBwuq0NjeWCudVg3MyJxfpYbD3iNWGnLH5JIrP2gaxun1Hqxo4jh/w23f4Axf+tf4jbQBQBr
6qd5vyGVNS/PH0ZgWW77Atuuxu+c5wPIVeOVF97z94LexjolgHbnW7IZbfGtQIyCadvafghLzBdA
B19K0NNfxwav+X+8oyMql8TsJrFzvn++muGrkiDd54fD8fx9TZ4vBU9Nhib0KXI4meEM8IuoYP8z
EgX3QPNFNrRO7H5dYvWtu/z5XJ/CPUXxl0yhF1juAhwcc0W0VFErjB3OcvLURYc3IipVfnBps+ep
xT1UAyF2DgMK2hxEE4iTfN7OiAtXuqMZlRE479gLmY0VTtX/N1rMe+iWnQ5BQmEACgG1Bv/JN2aa
wmgPMnXWAIhgROnxZ2EyvA04LmMmRvYijb39SBgJAAAtpIVsxPUKCnw1e1Yb2vQM3c4cw+U3bHKa
a+pmBDvl5ODOb5BJ1TqGBI6WPDOT6bJ30kdSgCtwAt7wMZbG4KtPvlt5cZFziamBmRhXcKkcJpWp
edXuk1GmWWJLC4MsHppWF7Cyorxwvs8AGA//DSor6BE1sJteWnic9bYu0UR2bZ7Ysf1gd9ooIpXT
HqJQS+gVqlounKKOeS2HZrJoxzcvg19GG8uocqZVc8b+/7qqm0zsEtg0BzfHsOpDnNIZgBDrdRVA
Oee3kCUPzc58X/jnBXi0eL9WYiX+JTC6aXVjjhzo4whxoPQ8zb3wBnh/EcCKEyV09SxO4q6+WqOd
eiGlfEdo4G7nPwagaoYK1Hsjf57KQ2tyNZ1Q5eWzmVMO+zVsdm0BXtNqZ83zkdYNf9VvZd35IET3
SEPtZLOfh3xJ2LeH/pu97Sas8R9g4jRK9lr8U/PDzlV/O28lRntVodWD8k72p2w2aoVMxRIr4Wm/
y2b7+mKbuyrlggDmicA/qFb4D4wtACjKHCsNsoNSTWbHuXXB2bkQLmdSYEySiAx7j6D+9vNLpb1C
CqXOCSAK0l8rkiR4rZ6/Ozat2Fr9J4t518/1sGWX9z5UoHz1baAzeCS9YSk6mL/Bdoity+f4S23w
8fFCTrcz/uA0MrHpl2GlGXn8HmDzKE/QucKdCvgn87W0dtIazPzjSegvsCU/rkzD51Qt5poeyogR
MJO/G8nBQmB4Ct/YdsbRjCKeqBgn+FnLAUJh6hqzrSSEN/mNVJFgjkmUq3RjlK9HCBS70kdtIqpv
gZE9JoujTU2PZZanlpR7o1QEm1LX7tdLrTOuXLq0SIN0ciX6ibkGmh451aZ4MYFcKatolik3ni4j
tpvcMTEUX7eewLAAO47s7IwRQSMLc/OJUYsRVFf8F+7+jE543c1bg+MpnETNlWpTEWp8VxdVG35c
5l6qXxwUuJ+mHsuFyxUXud0mO40evtkyttNxf7Qn8MhZb7sNjGeDtgBnei4XFuvZac5C0clAPRnd
N8RBRcYk30rDCMXlQ+gHnUIKCuUH8atkh+M9QZfqHawEKbDiMAGeYN32aFR7R843OVN+moqQtHtF
ERPnUBaVSkAOuzJfsu4ttCKN5VndIBgLkN7eObNdLzNhbP/SlT/Q7bpKe/0QzLn23mB/6QyC7bzG
odEEOigE0bha/hgB4Bfv8dMq3JE1B2+OG4lx/mEayieNsNS9XhBk408SdRXXSYL2W+iWxS7K65cg
S9TiW+sxOy3o8/pid82JAIruEPDixBNGpAPSs0AnTj5zCMB9aJvETBCxVZkJzkSu4ULRz52m3Bya
15fgjgfz3wuualUcgvLml5M84Pq1K56uRh/QZ8oSPGlIqSzUOq7tNMKasRKNmgOTmAg6pjnNpvcC
+0q2SyBWDcs4DIidj3wK6KXG/Rt/7Y2lw2BI1xNP9WkQ4AOU/vHKfJozdwxEX8hK5xslQn7JEQIB
aN/5ZFmhkeTw9OdKNi0nSrkOj69bM1XOD3SliM1PhyoBwknliuKaF46Gl2CNc1bwqRsxWlJDIv14
Cp43bt3d+rUroJ6quPjSDR2d9vvUFWoNSUorVmd6Ud+LsbesUZQF3/1b0OEzJX91FgzsBqyZiWHF
IZ3EOt7UOUSzVyx9Xmmcd/d5Kbxw4BS0QknhpLbtuWnyWjKq58m0k8qhuafLTMr6Ec75+obA4wrH
DeFgid2w7FDyMcDv0iR1oW9/8gjghLoLV+kLHnL0MaYolGdH7I8PugkqZt7KTr1KTyhzpmp/+XYQ
hXdqbmetjJxVOYijeHv+abNbrpj6tH4YWF1T64ZJc9KquWiw7LxWtrN+qOqJYuSuD1of8hOaOVGO
g5OAhiXJwaQ3tFA3uVEblA8Fd9NvvPgrMHQpCZ6UX6bUEmrEuY3upcNOVDz8DOJZ+04aBQa76bT5
DPU04kTYPjaj6RstJ59YA8K1ssVa7GOFQvyzIzywXAShuQATBd1TjzFkcC1z1xSk9R0kqlhLs6ss
rVOf9gT3jQcNXcJ2/qxH7RXi7OJS9LYvrnbxe1iNA9/SK6YKJSsf47t/a+jGtiZ/8zTB94GnbAUN
eH0GyfyxCCYd3tcWyYtYNxzKr9kM9eYIOgGTzo1Jq5i1iPi1byee1jBKuKXpGBVWRAt89q/OyUP6
owVhz/w+vgdM15cqu6J0JJrD+PKXi23SWKX+ufK+98HiryJ/rj3aCpiuI6DlhdiIN2vttZDPqUEs
ZIiD2gx7mpbssEz8bcgkZckHyreySeIJ4U2v12wegPmYW4exc+qpZRIsPx9hcP/QI94wLJ4eA3bn
VrzyWsY37UCc8HHp34b8e9gdarIw+coT1ukFu4WbMz3vNZ1qdfUjid9VXOickMV4+jrBTEkTkYVk
k/vVaKK7koMKwgUAPDpnYbLFnx7RhNpkcvMlBC1Z24FSPfaYu1Up+EqUbUroRTB9rqSItL3dlhx+
2beSgE1wMUVNPoG8wN/yg4atwD777KNBRjhjcKAWC4FdtJPKHD6sjxQ16ro5dNFF4ZTACNWraatr
8JjL/jNvk2d6WVjDsP26OegDOdNLB4CSp6ML443/L+2CuuQA5FZA4NZvpbWenayx3QcRaMH8F/YM
p6oRkcKzwC3CkYFDWUw253L+CT/EPguMGSlj+LzEOxyZJWAkA0yvHXy075MD3iIhZfZ0FHj0XfVv
tLS47Uds0YpMuLgNdMYjuEYTY7av/6Jm0kcb/ROkGsIYJKpcbs2BLd4LE/Ssc78jHdfu/l1MBHGG
D/DU6jnWcxJeWHdJ92qILUxIbgvFu3SNlJ1RsgtbQpvq+3dPsdf6740G74pe0TTD8Yug9f9t1qw4
hGMr1hcw++QcJ+qAmw0mazQ+WrkSzyBgz0jhn1+jrKgxw8NoL4s3IKbJhqvsB2NDNU9fgPRfLffH
u+Xl/e9YAXvy6dtz4z2F1XZBj35oJQVQjLux6drgpiQi/UxEP0nl9sd7we6APm6G3PkICdnjnuhk
45astj4cox929//BMWBaXjZbmmwQt+z0xdlffl9HIrUbmT+0JdmLKicU9sHig99UQG1jyaKx+rPM
kXttWdScQ31ln71R3OeOBe/MkgjF28GLqKkgDNot40YMQiV84o6tOB/3Lwm71A82jq6i4NW+EYvQ
B6OKZz8mB1jXO4SnB7RMWOigXeqQqyPVgB7ok2MZVdponFFs6cy8M4g8hjkPcqSZNrAldbAOJMIo
ZsaDJRfQQYzWm9nuOm/j+e4Vv7mY3ULfVfJUgr1sOFltQ2JeKZ6r7UANZoH6QBNvsINCroPV0yJH
Anp0MirmDFFjZzkDD5s3tItXfz1Z/XRajjdLpMjI7Uv2Hhb3Lp9vEnfGTkNLZKon3Wj2VFJzlsKx
W0FL9ZX6WBoR6NsaS9yBecVNYMfFaGrv70H79ngGe8ExW/8x9xfMohg70Az7HEKdlqnF45RI+ywC
PG0aD8DXUoWgvkHhdMVDrX/FU5Bwty54jxB27qmPwRlgT5qMKnezOzPVhm3RWBrL7ggOuPYlhJlc
VGj2afHse1ot2/DrED+jLNChcx4707yItCVm9MLXXC9vzjPBgR/1RMvOM36EPJCjvB0cCyO3nnIh
1aN+2lpddCHbdORXr6RuKBcjGD5Ux2knsjy2+BXMCcCuKhcC7ZesgM0/uWwcPP+qWLtAe0z1Up17
OCwX2kekYFUQE84h+FhFdZ6hZq8tlEmYrN7AxE42X345+IaqiwQCwy/SWUKpbwCjcPQ5KMHZ6vkd
6YS/+SIndGaF6fJ13AMylPe5k+rZVlVXgH0QCygUEqdIGTT/eZCFqNa8v66cMyfHaN93bEZeQKUz
r4/cqZs+NKJnoBIDk0qmfhFvpGBf23xGM/X+KtI5+VacdKyH6ZxXY5VksL6PD7wHQjQ4HuEY17Gl
G113GVgsbe3OCUEWv0QRWB5KpzWFAOgtY1+jMxBRUh5TzJ/S0Zn6J1gJvpuNJaOmAk+3e/5jM5kg
/iGtwcGhX1lK7ldApSzJFiLHxUXIJY4cW4lwCXl9pp0nyx2wvDbeZxDoyuG4S8eiLBr3RNoiJv/i
BQzxmnaSk7D7rDi9DAhD5CxSc3Pjok5w7o0ExHVhkJDXyRMpZYXHqucNyq8u00m2w8VlK6ys0A2A
fPq5Ag8OBLKZlvOZQ+wM1MqVDNDMVg2TkTJqNsCzxH+RM3M0PyCWBen7wIxEtQIghoG0U04+rrDy
8lvIuA38v0yO919lruVHwdGmlHjDX+K2mU3lP+eafo9ch42UvE3P5K2CJX3jRKbNGUTtikszydz+
VmCqRJVX6aGDtB2THD6IIhEdqVkSTnE7X1yGn0XiORNOoVKRDWa3C3e7zlxfIpyyL0cC8p5isIa9
wzdwH5bn/p7IBtR1WczdW17k72i3+DNvB/B8hY088ii0AMJPD4uIfeuFwuLUwCiALQmqlLvJ6lW8
wkhYrAps7eRphx7utkyrQbUPHrz1rGLhNPzBSXmZu/rSPOBYEuSoYQffKKAB9W2mMLXlSefGBLvl
DsG+pW5D7n2332OC+LrLpODkfMsppUg/J4aAhbdFs0sCeGppEDZKL+fp7QHjNjCIhEZcFlMIxWgT
4vPajnRMVLAJ2adew8R2cMyWcj/fu8PMhbpclYn4rlCRkzeu9A+ueK7mQc6/sBoaZpA2+DYfgL1n
KcIApBu59++Z/XErXs8+J/wL0CTmIhOPVyGcT9YefCLrHZOYxQhGntPh7AHeV3DdVpXC7yWnbVBQ
qAu+PPbvYSySeOHe9XXcqSrj5DOvG4Q0Ji9yoR//sR1PjeUu4dFx/UKRd7P53sY1hJlMNdRNPKM1
3YQf/rUVCej6Eqv0h0PJ73PWxz0ylp+2+WVjMpHZ/T2iDHzpHL0cJT64eaE8RPfr35eWYZLubPIh
ro5uSlFczDOCMSLsaiGM3WSiAMYHIMJSkKSpDvngPOMar4gi1QB/K74jmMpfz63ErtunsUesl0e4
h+k5y5WH30utnStZJaIDEFTAdhFq/VqnavMNteeVfkF1oENHPGbgfH0pTkxzG3pmcc4hduTWXh47
J3wSRV0jtrksxXJYi/8pw0EoaKBSV6OwulHnFnW4bET+wQDOKy6rOTfMtjmSffmgSn1GxXnSKMUU
tkaB+irZxAXod7TJ3xsAy1RTDGmlGkX7YIf8wQEQjAZkaPB9IlnaBoGXHmJJGcaXehOsRporP+sZ
nJlVQSD3m8c3h9D/y2LRAi1Dwb9uIXymjzUXEcd2h9r2kAaKRgIZ5FVyOkU5MquSrpgsfEpJez/z
dqS4So4bU880Ywy1naw+v446+mPp1YnX4xWJrgfbQhUlD+s/T4E2pMVeefbqFn0YuMwWZcF+RRXb
S/BBWuRMAx/GCDT0QIKc3OcdBiUYWGYzCnCA0BcJvCY9WioG+uwS6JPCcTftU7f9xUrv2wMAdJO0
O+fE6z2YoLzhYar+S9VQYsfpho01hJ78x+G0L3CJVb42Cj6WmFJf5eLSs6Y6gns9wgSdry+dzpMh
8GsmdA03KaiF3Z/sy0aQDnPRqJnrOwBNAa8p8g72Eer7h2jJeA5qnJvhLh4BZUd7SSvaBP9SXpMJ
iW1o4CQHJbIVXOHSvcXR2xB7zjK/W3mx9sn3koan8uJWkDpMaFGob7NWSWKci6YWA+SPgGuA5waC
ayRbtmiy3WObthpBBxU7n+LJru9yqzpxup2PIDndtWjwJgIQ0QNLyDrQKuviD0LJadTwDgIfKIDy
/pPcoo6Px9EKEQRU47IQwnTjty6jq3JRe3pFja2IFCrI2fWHwGNE8aI5hxhwhCtNzGMfxqbLKq0V
t/kABj3CBs/XqZv0nd/ZdTsqjy783tC9GaNrOicD1Ce8W/1CiCPIJT6y78wJzHTNOzSdN2o1cVyo
oaQgrsLM7aYoNeOzvZ3N9IQoauzqtHqbcHcb2kj1qvW6ZyhgyoDa0CUCglGJDzN+v3jnNMKyuLTT
mEkduwAtM1qmPo1E23bzZVMiR/I5yZ/3bQ6ZfONyO6RJJh2RC2kfPR48RWNIfns+Eq3rgdfJ3+qq
k5NMkzVxjEtfEl2MHDxJakpCougvGBCm6ZxdPp4BmF0cUe6JpNGrInri05ABW2VzDdlYhAoKFXan
lpBEzCtNAl1Rt0KHNMpYq3QNIJL9p4Ikm7zEbqBGMqa1sCc9V3NndLJ6xXZC52CfujJpb1+/JzAr
VkfII/Mg8owv1nvR04FWLJJWE+Jr2Bdg2UkaYqyoJr5Faxojhx5pqbDqf3YekKMn9BEPbzWCaV8J
qpMEqw/FJ0Wom6L6rdfNit6Cl8ydRy963JHZkXk+wowSszT3ercGCnawYyrmWQT1FRBWY1Z4gPxK
couIwHIQxYQA7VrXHZlMoUlE6IEihkhuFC8MSE1eH7izkWlII4MWEkCRh+QngiJZrBzhPzrliPUY
QZMF8EdpjCOVn6nqNREzT9kj3h9u2RwrI0eW+Y759PuL4ejDTrOIFLY8WknKkmbHcrTWEW2OtG2x
ZuktadsSHXL0YHdLzzhN1z7xKXUNitYp1mD3Z5iUpRsMX48AckX/T3mnftZiCaR9hXkhZyxLFq2w
AytU8rUr/8kRUIn295AQilOzrZZCbmkyGlw0O1+efV+iX5cMLYlD+ShFxnWzjv7h7V8Y0skjoN/N
iZWiZwxDKyVY+oDruweJgxVWgTWzeqvm1ZGMvxDNvfouk1Jlpcl/TX1U+zugTWT5JQj7ES2epf4k
2Z5FopHXC39+0TPOWVMzXPypFhh3Gwaihyapg+OatlAvGZgrsKzgvR6aAtcNb9SSTugeFP8BoEPN
6xjxTSWwyMxEHJYnsQ864E0LTevIPbCnbOBKwkHu2Cf4MkTCqPQZmQXaF6vfcNiRQjoFYIZXSfId
r244zV38eDJqipwgQKmt9McfXbNjQWEKrDMBPsIIoMo8BuMyqsJyb8aRP4PdCuOeUTVHe271Xom8
xnmA03UF4ZtDjpun3zV2beTQ9Bwe8NKoyBdA2eR6IO48jwb41RVERLB7pEJjtz58xuHOfDjSni7p
wbIeK5Ct6s/J3UF4djNXRD5qSuUznde4xrlip/mR+UwgG2vX2B9WvfBSsnpXLOhBiATBa2eSAY4Y
8tx91CaOj9LnZ/6g2f5zQf8V23FudIA85UvyOOMLtM+KSHNaQOY8tSXEUMP86Cyl3APjKM9zTQ8M
4W4xYu7G6aVIAtpbMDpBnnDAmqrpPzXfXPOH28SgXVBKhy9Sv0wLbzz0tsMo4KUauAzZqxRVw/VW
HM96Bxz46it6wtkkUY+ky1jrDwjEBh59WmUiVWq5c2eo+2Ma0dqHcZgcvGi9KZD0Qzn2uerZMnML
MuT1K2NE119s2KLLCR7H4nVGAVJ70LOFoCqiPLNbXRFM4AM8Of2S5/NZLaa2CwlKzKpQWq4DDPze
Tlyf1UomJWT10bHz4V+MR6MyUuFePqNbWcIk4TOiudUHRZOEB1nfdDbNxHfsWB8xQAyByyG2tvCd
9Nogy4+G9o/vZefNMcd+1zM3IPaUo7EgeLlP3rqkLadpd32oQHeFi2P4azlmkkpDX/jM/C8OZVlB
0vPBbTAIhhFrYxkpuq+Q5XEgARtsP79aTnIEJj7SM7TBRbCoaoL4k7HuOn7/PEkPO5haMKpMeM34
nZSas5jeNIfe3TF0FI+FaX5otyGogSyDsouYNkdnNftvvIWCoWhSJQPzfpFKmA9gSmFN4y9aT9gG
AxTS9f17jCfm3uEFn42FPF22daIEHzB/WxS0ibrAvEIgf76wDa5BAhIpKnfAKxEVPVOfRACz/eVR
Ea3n9jCZQxdYZql9PvQ8kq1AF980ZFu+j/G75oj/dd6jIa18/9MG67XWMWMnIcwYoP80/9uwqEVC
DxytZ8cekVnMtZJWSCv4v6j9yXJ7tAxO3xOEIPQap7l11N/1UYhFDsmKmGDWZrWON5HZ4MBzhixx
3Byp7MArBTYiIeZ6jozvpjaL0lj3CA6rmVtTZMlUj6t+WmAjvyyQdurWEOl7c8YjuMQt66YTgCmv
o7JZRs7x+sVtKYRhbp2n4Y3nam193rmX/8XfozlC1/14nLngRs9IFgmMLm12bnhqBCXSMRTpIspo
kIk4onnaXgHyXhPv/wkP2VIMiEqbzO50uibk7blDaAN99MHUTz8SbLhWhnN2CwIwfZz2oRzVCxAR
BGfRyu0XW+DZMPHGGzdW9T8NQ6fPHfWmj5xGOkAIfPz7AAxT29pih0QFQuMnOLaytcX0me167BM3
b5EQmfOo5DMVGIqlpHtOV/AKYquDebc18ZMKljweXEg3zRz383GuRaIXTnH6chB7Dgs6Tm7jwxx5
WimHmoK3XnE+N2MP3AYmGrQsW1xtr8UmLssWKQV9yMv8HVZRG/PlggcUal614aEMFZjUdQxL5dFo
ySYiBxr8+162Y7w2WMhb3NUs9By4q7Hozwu7c1bgvB1VRryyrsQa8fGmFgT5HtoLxZTONLg5MM1V
Pg9l+DnE/ovhWsAVsONWvlwWMhofXj/QqVN+FcWfFTVWQMgEAyczEYqkSStaGcDXl0Flquhp4XmI
7tlGZjPOVUXsQE0IIF3s1LLGPgv658IpUIrTznHzMwxNzRQ0ugjpQQaaWziAco4RKcSCAwjRWu2R
Cq8aAnrhBSDRjYSXco1+7Bs0ktG5vFJzwJwPsjS3JNoFLDmvUbniGzVZWKQgUYSmeKsjK1+Rb/mV
cSTCaGFioQQHp2mz/SnthcN6Rr9vaWzMYKVwuZ4iQ9ibZg4XRqKc6WSGrB0JkZExyVEC4j3h/a2M
94aol0oebCmNimfcnNcjn0Y8/erPlPMKpTC3v8hmOAnVL+i3Alvag/6BhUhFPGuoDExG2XrhJfI2
+A1gDSv0Ng1SrI/HnEWc0toFAvoDsbroXQRyRnRyQZr1OzrMZEXB/aVt2iV+/5ebaUTyuxo3PUMo
Lg5l7d7r47B2Q4IATsmKLdpEUl5rXTor/lPSbNbdyslOoyDCPs05YXGX2F0Q/Wfs2DdalWqKAaOd
e5NCU4fH1YiFcOCA7FMwWnvixHAWVAG/en4GeLcELT7h1KigMZfsZaX5XKxCIqI9RYfnizyxoWYL
SlN0ixNLkPLriXFrPREjQexyr/ih9CbCJ+abR4q91SpgYWF5jYyE2fvJn/V3sOzbZ9rMmX6khXAs
vL6Rq53Xcow/ij6wDaMlqx9pCOVDXZWrfDXLSU0f4et/Q9y+5CINv9UcO6c7H05FCxYTBevJ3Y0x
nUSFCx2QhTrxjGwNtAMmlzfzLZWVhhrgWE7ay6ItJZoE9Ofwrz+Tnt3YGfg2arsEYj6XwxDPrrnD
r2imVyxWnl/q+5qMbCxpj7lRayROp6n7CUt3r91G3SgTvAGxSn9VWWleMiSFg9FCKl2Ih+GixeKH
4j0LRXk435g+AnJpnDYpPNTPBChyrJ8U943DB4OfukDYqAmgCMzEnBDJMHloBWAqCDU2bW0efDzG
su4AZJSYnqDQDwcr++kvx+yZIGaeO0px9feV/7Og/XcYxJXYvpUr4R/0ScYKdMDgxh9x4pvGXopI
0zG+wuBjH//LG19gneEIp05eM3Lo6syGEzY0k8eS7tP8fu1ObYINfvj4vcTSpYBb4+F/9byAM0dP
JT4WK8KPFTaIDNlv83UfDinBsQZrqLVg1JDYACeuvSWzzocwMfXzJZcmW0Pm9+qvSP6cfUUG7Ot2
hxi63aOuDKnUnIZcB5+PFiW8JLl2CuAoOr7+ziOswu2t2D8UdqooG+85P3l9emJdi+Dr40Rh77nW
Z7s/a8HYG9q2mdeEOnuMiem3vn18NH5cw3SXuMUjTHxr940zYs4o2NIF04k28PW3QPP0DnsDJ+E1
xS/ZQe2v6PkCMth/OVg/PsU+xD1WVk8/tIVtfSdI4Ygs2HoCr5qQyeAR7Gdlxb7CoBSygvS9FshD
TJ+9aY4qu8xn1BvZv5LurKCuhmhyKNfO6NGh3PTWwiJL+/cLuPP14RXWuHWeE8SqxRXGQ7sv5eK3
cfQAdcsRQYfa6Iv4ArJ7rl0wHJH25c09jWXf9J2RFWernVGDEY2zzY9tejyejai5qFQvhuryUHcs
BZu9Hg1C5xW3HOtFRpprduZculVrzt+E1SVSh6JxqLM5b24WsfG2fJxrwoGDh/ophRQ9zL9xtY3U
eKed7KpRV7KH64vcZ0oam2/kxSrP7z/yzMxByJsdpxnLjGEg0nve39Bg2Lp/TiG/lyguQfosySfD
O4Ypby7cfywRYyhjwVqnzIzzG4qXmZzW/7OfCTobB/cc8E+917iOaZgNqYpJ/ImSZRpJlx71LARU
ggyykzb2REIPwK2NeiLrfdus+FvweJXFlDB7K8LzhdeIb1g/ay6bYrZHkJ3FrsMZ2GwfXctoQ5RK
yos0J+DZERA9olFBhlPiPB5KNYVNRGlLFz4EDNIQBIdoLCioi3ib54QvGg8oEMAm0udMoPaY9KwX
n/0N8SiD4vupnfr7QZy37/aFzdgn4R3ugTQoZTz7qsjoVexy5Ux8oaXGbShDXoFX96MbVLS4860V
uT0k9tojKxNWr8MLi/pcbp1I5kwmcGjDUWEVZe7TmTtFf12aTstWWsca1Ky9+B5Paw3+Xjq+guQ3
geyGJpE2SCI8MOMCQTfDmmwOqPAqCiO+h2t1BIKJuKtqSqzymbPjsZRPP2T8J2uSHKuSy08gF6Cg
o6mBrQI61nG1vdJlblY77muVPNm3kSLq4y1oOR48OOPzoK7+gkV55neoxOm0GVzS7XZYP3mW9Xvy
EClTXHerk+aGeKd/00pi7Xb/BLKuwXDNjFGbrBpvyn+lwcNWokjzYYKLjOuy1ZJ8HeXm8/VhiSoD
9nct/AVxMHrbMNqiSBfU6u7nm6fNvvO12SXlCQQ0czgZlcBFM2qVedkBhytzsC0VSYoLDVbH4I90
czSK1kIjAiM3CpzTLV4+t4IAoZCi1DyAgbSikZOwwSsl02vc9pTkfhMXZQsZenkjahiYzP/g2Nsw
jf4bH7stb67HQeMoP0fs+Ew+QdChX4rDBRG+0iF2sDTWE2Udsq7kp441dlfVxE14jwoqg/mY3mKT
WEN0y4Ch2hjxU+fk4s1Dyv2iig4jSW2oc/4Q2/Qo4wY/DR1nDxA+KVy18ubDWcAILwvIqcRFx7ei
5Xvt387Vgl+1sgPsIgILB3AvCJY/OWn3FRYmTLGnUyDhQWmKsr9xlPEKscd7Y4qAr7RXHxDKxrlD
OTsTpK/eOEJHc94S0EcJ3Xfegn6U2gsyZdTqz8sXtAW+VgmObCTB48kB7eHCf0kISzvEJKyYKLSd
VKdDztX7ZUjJEkR3pQQ7Q90Jkseta5kU0CY0gkVBd5U/xSCgAHAdrmMb0Mu5lJX1YhEKXmjoeUnL
2VA7QGvqrmrv8dyR2Yz70nsucfiPI605GBf/N4v/SqozL8WpIWqU6y6VbPmrxOULGq0hXvof8QtM
WreyNJKk94WXHiLOY5+BLb0GyRHnJEO0UR8UV9nqdctxIjBFOWRZX0Kc6gfLFREXe1q3ycEef7l2
ZN22WomTU2V1h0ABdOpTfaf15UNRp7X4JSBRwgy0bpiHyUYpEoSLM3amlYlFOHkR0QBpRZWftsWR
FbHnV0cvEvUMfuzVvgkLfanOVqhYxO4q6+PWTmvje7J4qAM97tR26XInPExmMRPt7QPwunxHpqA5
vI58Vx05O8grVdn0maypyx9Umscgv4XbrtPNVtSzz/b8/se0zasPXL4idTVLHimKnYnyKAjVbQXT
bVU7adQYlwCt+JnIrmDUlxrsRGKpU8Q+oYnfUCZ8IsZ+I/0jqs4A8EpCHh6mLDAgc0HTmz4eeiKV
Y6UgWnD4rPg5eey2+3YlMklfx7nyvSYe86RuTLFQU6RLm242nAwH63P5xnWi20IZUYAYw6cnGPNR
5GZZ6otBXg23fpCSFnT6lMBKa5Vkl/K+MexaaYLFd1uS7+UHICoz3nbHN3iUTq2w3VFdmu7nKk1N
XtG9u2HK41YcTD8g4GJNud1dnWOAsCdnJGhpdqZMf1o+2K1LkoP9BRr4q6Adb6AAzKI+OpXs9T7U
7yxsVHxUoj6/7yj+Swk5hkwk01QO0ODCsagwbxgeIntVvepCiGDXAQ3c/1Zef+DB4xRrE6/YCg+N
4ljIbeOkiBnAPZQk9nOl4bJwFRmd0IfHg7DG30Jv44HecTET3Zxs6nuJgqWM+RQ0zqW6rIEJES5T
fr+Oorm9RJGc6/TCWFE4MKrZCODUsoHgWEO8/0tCclJIIMCpJHmAEj1fSWHtIggbOITTHBT4twGn
DMejm+Mpi+++2VHwmU11C7usCmnQf+dNnOSSFe6wZiKDttt5y7pBGL4vGTYJkaZqa1BXsB480Vmd
fnJ5RAZiNGxiMaT4No+WkOU9yyvm9suwqxyJ4lE6i+bm5VeJw48nkNqhIzywLytj7R1p2MxuWn2h
ccgRAO+ThRNWUKV8gmpWwPioFMhLoly+4xMyikZ31RvHpznpNxKRnfjPqMkX1EPFcpBWMdC7+2Vt
4Lt+NnD/BcuQErxDecipPsMcRnoMPqbtb313IDQhefXH65TjRmvadePcQBdJx442UzM1wiUotApN
fFwh1Pv/1fn0VZB1rWKvL4ZA4fa6qnrI+R6MoH1ImHiSwgRt75oJ4i7uSj8RXUofsDv+qlnRpkpn
3TK6sabxDKJKgNCDRhxVgRtwk3boGrObnZkrUyeAvP8bPFugcXG78zEp+AABvD1Rd0X0Lk/ry386
sp8DoNHuqhmGCxanQbdxO0dGXsKmcBwbSQJNdF63LYHoRclyGsNn/XRxWzayRt+CYf/Y8HkwpWQc
mCuqIfrXrcc51hiCVckTsFPmFFzQ9+iNmakToo3aI7DQcsBzvcLQ54eOwMlihzeZFPGsnzBrgusb
nIc0cVtV0EzT71gWeWA3/XgCI5BDqRdZCcSvREb1RZnWDAzV9zYDoCX1o3RRiqxdtT/5FG+w+BSn
tguWV5Cf8IAUS3IWgqvINXDRIqkxQCf2PLvto2FqkJr8VuLV3BExZBXNpwuJx84OrYQSMk3d25rI
aDVlrv2VfTL0icfSlIsBvbWz2GxJEMXiNiaZtvsgaUeWDyClA/9srKz2nRoyinOBBd756kQQeAp1
OKpAZke9QOQEEN6GxWfzRIW8Cu4XlFzAETjIL+vBuDkYN6IaTpSdJtVV+msbIuoNjAbpHB0PauYZ
uCTNNhu/5O1ArRGyIMZcYMyIsmNZMWrr/vudHJCBjouaVwg8hXcN5Kj/PDydL8JvtX0VG1LtStBt
HGAvEpL5Omy5CSu3uGzQ79qhIF+kK72y1Eqj/VMvk2C+yrbvmzmexxhUt7Bohz1SfrEH7K/dylpr
hQSmcolCCtEOdkEoUw9SWAQ7hD5nbghB5Ma10KR+f5K+3bMkpW5KoqYWquU+k/rDnjh2woxI+oWO
F1ZWSMXXIHpR7mTkL5SvNocLWPtWztDAErLkWTxXO2iMpwqn+MjqiAEjhtziRtS0hYR6Bc/lPCyF
x6rSxP0KndKqkzjBm9/c1Mo7AuNP9c1c1ZDsgvjjlx2wUku76WJESwk2qqnGtZeYWMB+plE/ZUR4
YgX/gn63OGAhc/yUfcixUWHn3teb9mCug30g42VzUooO2t4r18E9MQCYPDW4PwROEU89zCNfRJ9+
P999qrKuxKZh6bQrN8mPnfBfEqjALE7Id0Ik+Eb/AanjZJQRKXqfQ4y8YFZ2xcNnag7KLFillAj5
dMANX7o9PLuTLpnVdaF0CtryqCfue5XX+rQ6vVpQCEoyd0qzXpISIM1oT544+2tZeINWDDyyWWxY
woHgWlpqyB9w52b03swirxbD7zHuSxPHUCPbAIBjYQRhg0rnws2J0bE6apdXHIXLjSwaXPIf15a6
p3sOTiyv6jKulJt+T3H/O+9a1qIjz+Z6JLMx4BruZHz+Ao723unrS9LtRzFYkOQsVZU8rlXjGJrY
FNyS3Bln2Mz99vmjn6PNT8nlNCmfUOqbqrQZD7t3bEbmiqGFMXIe34i9DDTPbhlCbFjf69LdanmO
ZfmBJ81W9QZ+kF4Gz7xc8vG9rrs+HZj2kaN8CAUdan0WNKwdPeTkt2u4KUwmNJD5uYGnnV1cMMtm
gJ4UP0bsJ41TiVm9mTL6Jw7PSekx7vJCf9Jr6cklF8bnaBhrSgB5MUG8HANhR7M3s0uO5Ixlcqrl
aeaHBZX7JBj79Fc6Rs0LC+0U7x/mSAVJWpw2SwfQSMR1lWHMVrppCdzSAjyVfD09KEvav3pROIqA
KrAgQcZOVZVcxiBFzrvAcHthgOZjtHqBO6LQQx5b/Wdnmoy4OS5YrKhrFJC/XRbR0v4deIl9rcS8
P3zHyT0Lsf374IpL5Pg/X7lgU9CFDriWl3FA4KO9to620S5UE69ObinonZhxew9H+U9JhA7nt7BE
29rY4eheF6MZ8lzOkYYmBY4fZYrJh1K5+m7axantOgGnES65i0EcOWHURt9Zgfn9KZOsB8eNnNBg
QAehNl60UjDkpzJiPV8GX/6VZWcDAtAEq6JcDRaMdlMtT+2rQ4b4ffHgfT70LgQkq8OemY84drSK
TUXYDu9VXqh95ucib2/ebA0w2Ppds0I95GOa3AmP7znBJ/jYQxgNuVEKSSMLtaTej6V+zUhNAZbn
7nwwZQ7aqePeeRjCIdMKBQb82nJn6xfIYdNfNsKCpes0BNnlKpU1BQ9pFc3F+RELe0kXm/cNAhTW
bbqxTSFWPB1ssSvZJGUKh0ooNS59ljwPDBd3EJgpdg/XAYG/cBtN8ZeI48drOJ/PBJQpFPrGhxfW
jR7jXH9277zM+BQv59hnc575vLLPrdT590G29rEuOZYpPbNIejFPRVSj3KelcGyNJWS2yI9pKMPg
Jst+Gw48pK6P/ZwbgjCKRboJ13H+sfcsTZ1ocq/T78MiVsDAA9mwU4MlvcvXjsqjbM6+f4ARgld+
iEOT9vtX0qAup0ueCNJxkV8s1wa8xIYuUvWlyafW4Ozjb91IKIbQNxFHqYSMOw1jCohZQrYiiaoo
Og+98E+R/WPxIrOP35HNmCFFgTO5o/jpDvBpXNjB0U7I9v9l6FyvJ2pIjgKfss4NwS1ZR5sXXmVN
qcaObCR1puN3mqQYEakv4v1mqADnIwZpSWvrzLWp4pip7WCTBtBHRHhsYrVKPiw5be2rGljy6DeA
Y8lYkGTcGAuLjWHhYYzr9UaPL/KW8Zr8DVfc3mJzz8yUbqDLyxF/qGEf7OEEp08gzgwfAChgIbf2
02p/xEAWlYL0SVpyb6U+wmRbeobdy5Bdb80ANcpHeI1JiYWntQ5skb4D2hBd42vLuAQqnd6W8wHk
Z9kXVF/rUHuba5UU9VDQklFL7EmydCOxC0e/NgGWKQW6lupZv9ZbFdH0rZyXyPVoYFDXe2rOQCeO
fN8Rp8HYfPJ+xJ7D69hvA66r2j9gGMEJ9RoB4LiCsn/R91fdfcWIRnzGCC3HJnjNcK4cduCw+V2m
B0KFAh7GNF3FRiDkBBPO8J4R1/9++MxJR3CpewGEoVooxV3aCxLDY11oU3cucKnwBmrKQPnxZI8g
uC7usj7gmCF2iL6m4RiCmDSMu6caVVqN4pmG4fjaeEny49wwCLEd65A/Cb+3W/t7sudTJ+Vcq14K
CG0t5cKuwZDwXGd0Aog97e+62m9x7OWz+PrC/y+39M7jQCc6ot1WNIuGdHzyQmylVC67warT65GW
++jtas4PKUa7Z4nkeb4+gigAK40N5+dZ88jmUbxnvfy9wTyI72uuc2Jjqyqda01bVNHZe+2tcXYx
SRGZWv06tNoTg0psOnRwoywnNhjxKB+jQMg8Lmo6ctbvodQ79LQBitK3jM4uOc5WTcyE/A3vGJwS
RYNdCRwufctAcqtr60Svt1GlBN8IIbWPxclMccfERdbe3HHX6ptjLqvkivKPBIMGceIxAHJcqA+Y
AT8LIlDLHVQPD1+e7ESapp9n+/q/ND6GuV8p08hdt6bXOoZmwxRCz0w1sSGQNd3E8Wbt24CEPav3
0sIWqMgvlCgpnWLXrUv6VZYb4NRMaLWckkyIEpiBEQ32ZOYCGhO1drSiFpQPBHoggGWab29UusXD
7198s+VYWhSDkB9vl2xiGdxMJMWkuTzxbvZ2L7bkgg8V1LXu5M8u4Sdu5eLRM/Q/RhC0FvCR9Ils
3UyAlPMJ5nKPvZXWkM7m3cAKXDtYSYN1Xw/8SpRpJsklOoMJIq5wq9nsTnYidbjuBAOQrROROsA8
ZyzS+VQ9IirGL+vwUdrVLTENBuEB2xxxpJfOs+/9nfOAEOFmfTOpS7Jl6g49m0XStX7m5f5nT8xf
tU1whzDdUnQimkwf6XwgrBOjeIuGQNpK8foS7DxiHwpnJQ+L64XvUuIGNLh+tdd37iEyR0rfW0UV
pztBvMRlkoj3ozJ6QWouq1I4uptACoyiVqPakFebsnaw/sm1E6UHU3XQlQLPDEBf37ZPOoRYTFhj
44V2VMALmQqoxaEDuIAped2g7qYVN7sNOJTL8fGb6N5Soin6rD/U/0oVJ5btCfCjlEztD3c9wXri
B7jkF7lFbUKBOBdPVN8Fcw18QsG/i+ugQB+uVspo8wdWNf8Orr/CYYWZcX41TJcoPuHgQUZCKA1R
Gao8DfIJLymUqnHL1yJdyDi9F2q3lgC9IZTFUHaCmPgGQrkFhGRFLROKB7yzy4CGzCZ+/ALqVRpn
heKXyJyl2HQ3WqA/DDCGtNEonzpF8Fdn0f4glPBP5RZl3ZxV0wLbfETfvhhh6fCttJE9m/jE4Qtk
bot7eecnq+n0qLWHlI7H/31brW9JFNwGPD3l0ErTUKqAQJzx1D63rqa9WJ5azkRnjTYStSJUHcPm
H9vCt4Jn79yAZ0MaU3FAFWgozblxkLCOxa0MhmI79Bqxh3FetrfFVZzSDv631o4SDzgAmcAoyY3J
E3bDEt2jYNEM5fdS6/4uGtyZ5sqVN2O8o4dUZH/BVQCB46q67Z4tn0epnrp39NwBSOS/J8BkHoRU
60iswhumQALfZG8pHvFDDA4v03RgpYtBXJAKY71iloLmTP2ziTegPyAVJpdvuiIeI5d4Ry5rLX9/
1WcHEfL7TkYbKbJkoDwND3fhrEahJm/i5I7Put3rR4dlWCmaFR9zddnTt/Not9odJ7SvkyuZgby5
nRnFee9MAadwKBqkmbCOb5bwCGPZLhqcchHRbeCXrb1T4yJuz8jb38g4E2c62Pp/teSbKJ4UK+LR
CkNf5y8pucNHnThNfKY+tqt3rKPzLelK2IVvLf0v0jcrs4H3c/tKHQpmJyO/aS4LWAS1GT31yExC
VbF2PQgrYCO18nfE06HSee0fcT6GtZMPbi4ztkmYpUpmTUhafCTEdc10Pc0CaUPLWBF9OZ9DQ+Bt
jfGzvNgTZSNZbgqMjkjplKUkx7oyN95KdTOJsrI8ZznzzhHjE5vNFxFC2lZ0UUnSVWytasXfHldH
U3X3wcR06LDjF/jnvHrtcDzqfz5LIwuImh2VcadoX/yNEMXoA29X2i4N2mMV4Ih91eQC3DVATKH1
LlQphyiM7FuMGQfOFpQzIqMqzwaLHA2pa0JwtDRfqiO4e7W9VepTcKhlS6w0ZODU7vFd4k1clNgQ
pdOqc1TcNF3t6w8rsTePk+EBZp+t+HuMrHKdCRcZe3M+/D762bjjNBjUnR5T9DBRGxDh/MMFluQz
KvHu22o0M7DcoYCZouBsAJVnYoQUBVpMlJSqcPfrHvsYAwK7HcjnDTrPa65025QCrkAqZO4RA8Mb
VXLUNIJPpO636YIWJyKeVCDIkQ+nOpn9CUrg9Cm1sYqQZOsgxp6fgYUoIWbuFvIRR4t4CWhv6xO0
XzvKgxOVSYSsChu6StO+J3AiBxFzibuUMsb2CbqkOLnEClFgsCVP/YpFvbw405vUoE1jDU3LW++I
yVLLedOcme3+hzrj+rDI0CyFtPoffY7501LnAIbSBYe9TRFIMziGFJL5x9E6w7fXqaxBUaJ5sjcA
mXuTyCaIUnMS5unbbYg5vIGih0Z93YV8aywHMnV9wIuptnpZ+jWjHOkgrCComsNNisIgdBqigPNr
PYaVxl066P+/1IGMoBdgS02jEgRS2rNQWk/G0B7Pb06nbqdjjjV5FSIeCVaKb0bsRYMqexrA3Gn1
XO2GoXZQMypLGONkFqqh3CZj+2FyI3tIIOj699Updvxk4WyhpdMvDeJXCaWW3KjO31qxqpTT+NKc
JQLxebkaRkK8tg3lvwjhxaMJQhmpHUfFtWkMPTsIRfzYqXYZR0SjMRYNFFm0PZ7taSYp8mSDeLkG
DFl4zClVcWYdQ9iNmJSb99DZpTEhMxNh71nb8Wc/6uFKuxKi0syzJk4DilTlwlGPRDbrQe9O4Kax
sI9q+CDXl0+QvECsE3HwGeZwhJQFMJ0jxP+BNVQP6hblCKDwlrQEDZ5GhLuAGMPtaPApLs5pyIQo
99yDDD/mIuWRvHdDrjkSMKAbkDY23hr/I7ILckwsvx1F+3Rl1Vmjv8nB5HYwwqiDkwXkCVV7EnFS
boZUqelxpPfHWtAp06YOUhl9bdl6aTQSQDusBw6lUm3a93Fh4n44T4Ydm3YQvQfZ5fuTh2t/H0K5
QS/rbqgo9CLxSBhKMkg195ReVpcRjvNZYVczpOn7fi2g41jF+Mxe/gbBXdReX3zRgZhm7ndehoFs
o58G/aI3SVLhsR7Ama4NFG+KkvZyhKrFq0MeflsS932OuRZ/vo1VPnRID5A/pLFMUfk3gNgQoCr/
I6XFkiXbPTLYcUpwrW1GxkkKsvQdjhbT7kxsO2jZ6NGRqgB+S24toxp1MFHBMani7hkSJRLDXtqM
oDUiUSdxx3JL4d5AIVsObLt+5RuYZOxFJkYWiBVBZCrn2l8ZnVBsrRZv7tivQdwT4M+jO9xtu4VC
rbczUt49H7sX4NenVU68TNUXgXoobJnl7DRMmUBa1sPgGw6/NBduByoQrBodY0xsXydwimmbk+BH
XF7W7W5DL3FdHqGLqRih8zGexNo2ahZYaNmh2QWsbocPEoBpHi7qISlCNfCDxSNFhLCBe9rSoFVX
XVBF2nux96NoTuQldUJWlFM38W5LpBCC6xk88mqo9iejJDppnyUhlZKkoq8LvrwO22qkaYUordaK
3Gi9FF7KUCn6VqwlcdKUcxSRGOo1YMmXWk4YKis6iackV1+xlOKZYLTC5Dn7jUsQfW1XQtXzkp3R
VhD7XV+Grv/5aqDDZrU9rsMKsBr1L+oiZ1ogZB30IEg2sUoUdxcp7q5Lisj0ZJHI1UvaYIRZzX7j
rslatrXAx9zbwPfwna9UZSwGz9BafHFEPKDiQu1Uzh500cxZQ8U1U6YjGYK9iKoGQx/bHko80nSM
6KzuzafIL0GHjPs/G+oa2QAMCieeji7pFeZ4O9r0Wz+rfDEipLeRL44cZEepAxd74GkH4FAjd80r
dVZ8Z4pJanEdj4O79cl9IPuCY4y6UPORShc4vK6LlIxW8UFVRfzgur0B1633l7gC+sXpU54vmk4M
sEH+Zonddww17HYde5rRYD8LgVs9ARrV42lZFg2lRZBw/Bk04Hu+dwdZSt253LRWklwaCR8yTo8K
waIWg/k0wpz79PupX3Le+2plfQ9XTNAfAecbA9cFBOG+ASzGvPugtNYNoOTCsaJkDulUbGaLm8aa
gaF5ofm+NQpukG1dlzaMGBCRD2rY+NFxs+FfAdgDW0OrBfgytY0aEfA0dW4HhdtGX2stf4+fFOwh
HjoAiBPMkGn00iQnFUbB4RloluVLpqC+fQciXIvN4Da1w+VJuGuEtQ8+ScZaC2tiVAEAJg00p7c6
KiR7Kvo9keZPunfZvJvHud2JpjKc6KHJoDaMEVsL9rqfGXH7TwezVJ/j83GRnxB+xFHfNseFNz8w
SPwl7Gp7qVAwHvC4cZmFL5GiohAmQ5351tFmOOXmZ01TBJOa3rIFkKZh75hK3LIB+pRXPOOPOXtT
RtRuvhXTdLzwS8zjoVumWboO1cphzNbFnF53J0eRQtqZS7KQu40nEEiGCreIdxshGDKQRF2WgTW/
DFWOaOxsp+Lk8sD1wQMRLYWjwEhCeOyFDgSIc1oFwRnSnGFkkIuxQjFLZL6Tv9wTwFb/tu0jL9nj
0+O18+yZibo6q2xxFSP2/Wl/SMYGb2Bx09ruEOE1/8nSRxCW6AtWo0n5FhOOoau9xiRE1iNx+Xsw
2N7Av7mxmDHuleS/chag1wdkJXKmNxfLAid8MELZLkjpO9UJYtO+EjHp+6tpjqDM4BRzLYOHIrkg
yxHWGei+xrKdhoPKSNEbuPb8o4c12tFPO/ajyqHY2gKWgyLte7eDlQEqeYI1aDBfL8h3bNKK0q+i
RxT12nBTH9Vj3z8K/yLL7h9e6umV7uWiQdYIhb9GacXtH20C/BWRkCWA4Q0WoeW/ZD7kpv+mPVzf
TGXpCsWV6VYr/3ypFOvClE5zIe0N+VYD5g4q1P2Vd9aKqFHkOLRdt4ggLmF3mrL3GpuHTvICO1iB
8F+6j0gpn0MioMVHxQdOGS3oeuOgE2kP4bKZiN8ctXc8sZqHWA5pYbExtTXRxcAI5aQrF6nNWvD1
VrFRCvuBZHmN2Uvg2A4IDSFRzoO9pj2dwsfsU6LfI1RGpFiZeKRHBChGTD4ApZqzYTFS38Uo/WpS
dKjuIqDFDTxowAYig5tcoyVKJLWaG4lm3K8h/fQN26Ed1JL7Klhv4yFld0uJzvT4tjIWI3h6pvAd
5muQSBPx1dwAMGHw5Ku3Jb5fR1ROW4l0HHEc/3sLKk4iNpTtQmP8RVJhJaKxxc253Tjf3K5OI7Xc
vqeA8QdYCKTE0p/kCWFWUo6nGyHWPOgoaF5/myZUtToh28xZZ1+vHoPhQXwwMU9eEE5CtJQdZ1LG
6ozwnObqoN9uPh9vSaCr/w4eJr6nzrAaY0/YQUC20fGZ/BLNFiyzO2ZNqI3nFmRw6OMTWVnBE93P
WQHkV1pvno7AGxtl2zFycpOOaV48ohtQfh5OpgMqvNwTQ9FLdt92oiHB4BJZg/dz4BTkJqtuiIbc
XY713GUJQyKFH1UnfSMnsmg4XmcHbbqBEXhWBsMu1DuEz7A5hVYojM6YPra5SybWiJkvGAzQpZTG
juPtnkkqIgok/Aw7iWWw69HMPHF1wiKCCdMCdXdhx4mTDeUd0nKZ0GhbZJlrkOOaN62g52lEBh7E
NClxlsRHL/tAD+jIaNCG61cuqrWuAMG3rJZNrzlz0MbI/ZV1aAgfEVTp5QI19SDOu8+7F/WxENhJ
Q8vx6NpRPRhMi6INGhaIwhrFS+01BDjx0gEZjRxH6EH56qa3AMdMsrRYX8IHll4rXs5tDjwvLbhY
yTrWM4/ntNcAka3hTipAOPDYKGg7vHZHYc5d++RE+HMSDKbU0KSEvnAAwD4iztts0BiP6H2zQe8B
iPFEZE0w6VAkl9q8WRX4OUsH7eaXKQiTV8nB0j6SfKlUBaAkMftUOxWKpQZFXFg55SoYPZD4pAvR
V3HDsB4pXT67/eFYs0imXWy4TYf1f2T1qckKcjhyfctBJlfeQ4m6nB0MEzmbtU8urNRT3O32pqC7
xKz/RO/CZa7m1HXbZTYPQgi492+QhkshKSGtRPeoVY+Up7g4G7xOZPDW8Q4DFvhhtuKxQ993cPxL
qpS0KHkntAVKcQQytPIIctiqFqom7JJumoNmJpuYWI3AL9s/NNP9RRIkSQWHRI1uG8D5PrDj+MPK
zs8NwAfSWkMdxv9WAMvf9FTTYfl5PF0pJfaTyjwT4DT0dY/mJi6FVNdS5NrbpfpLqVM/+WcALgb7
VatLW891hYECjy8snyXt/ENsNac86SufvQ5bn8r/Sp5mDgEusGwI3Fq0kZSMIwwsilmHgS1KP4uC
a9fVthJwDjkT8ZZB7JUWmuNI4ZYoO8AedCkZg5nvMzCrMNzdpL0cWH9PEGxghCgAwsg70rvicQwn
BT2U9ifHezvQJnrqyepIhUciA+43uYbXnZvOCJ88tUY+yix1H0rlbs6Q6DYSq+lpmB/jTTFBr3vs
bex3KYiXqWR86Gy39JVomKMrnJH/GbUUbwm+3nL9qCs3a+FDPQ6FY2K8o2GQKITHOFU0NsGwJg9d
nQQutphv3aH8Mg62p555ky/VPLC8h+ljggeT3/ZvNhCcbTB+lZCG6s35ICrE7Rnzo/aVa6x5JhxH
HUHtF3OAKQyqeimPZqsQxmIb7pGh4XSHQURhhnyR9F4yW0GxQFwQTGS/AHPAYPzaD4qOcelqKFje
6vjHDPl5945j/sgTj4RfS1NK03PHbYAr3AGfH3N8Mpfv7V/e1APHNl6INHrYZFlibZCELIIbiat4
HqJu8fxNMwE1rLNvaNXfjevJ2GRP+sR9kUvfa2uqrCPzfIWtRA5xWwNs72LmMeGsiYSkxF5eWRqB
0xQGHJreAudJgKlNyZqi8b3DEk6/GfXPqyBLb2Xoi8vMcyNx4nO/mH6QhAqb3mEXiSTIuWAFCr7Z
+LEbgiTaG6zobh1HaCu+4itUFRjmjNlXEAhLkibwUbnECLiAmt3qyPPr8CyIHDnOfiSzljhovuCT
VPZhfWdr1KDXWMvGu2tHQjB/aWt4yWtHhpay4PkxdRdv9Jqo/bf74Uf/K//p6o6Mv0ZQqUFCW5XD
StXhelrh8oYqdjVz7dZaVWnzMlurOUOuRcqVxLgpQwXqJv7QRyoq2xrCpsRvs8ix4nj6XkaAzN8V
6CG+54StIh7Ix3QYJUIFiGujpFDiOpweAQ+TXI7/WsIeu6+RvF7QZ5atrAoslj4kNnidfgjTpplK
2+5rTidPY3mI9jEf3Xme+jHhZvF9ZmyhNsav8glNBxBqfSVriniuCXuS/aEgPUzsIQok47h2n3Hb
o6aki9fgw38Z3WUMBZ9xcpfdLJZtdbnOBG31DMRpsfxXL6CXGCwsQ1MVIJ3fFADCZCP5+MKuEVfS
Vf2/Rc9HvTjEITyy83pfTXvvHXYAn3IN4AZz0Gc1P7WKweTXT1Dh7ov98hGoDyM3vB0Mduv/zYZi
RUmGpQY0lhJB93kyUfa/dgbq+zKLPCpx3nFS/SnMsEcb/E4sX7yhnU2auKM4fRfiLf7jA6Qjbgvh
u7u6KpYJX0oQPonp67dblvWBu4CYUicxTNNDynTS6l33R1HeX2+5tiuXkWbk2vgqXRfTA4c7fGda
YCu6S3LFF1hPKqgb7CmuY/Jm9eyYSO7tIYNL1hCMXLtYG6RVp97eLQCF+dzisbxRhtkrrdqIfWP9
vqr0rsmesIMha41v0S1ZycpglT9TLGR7/T/HFGp8n8Pkvm7VXhCUdcwSwuAQORj3T5dfP6ViJTHn
CHHKS5770ydzWsqwD2vbCrm8re1V8MgFmGQxnsSi1GK4nzQwj77mYhrNtpp9i2ifOniaX45qk5Pp
s92enUuaI0PHhEcLwgiZGIve1/Qd3h82xWpssJmRUiAaziOuU8zSNoGGep2xs1k7Zp6yDCHE3gjY
RMHdlaS0p0+kBuAv3vHdnJY+Rc1+Ap6bJgswU+htUpHqA6DlsisWdFai5Kox9nZeA2KWzhnlDYgV
fTCuXlv3Ht42IGbGCUBf2waV3ZC94TQGAwqCKVVmKy/o5dDrQAIn6gu2g5CW7czAxFkroce6hh/J
ogiQoEg3NUR+uBLq/Czuy75O2ysFRqM1W1xvi5jv+CUldJKMH+3BFUk2Y7KqW265X97wj/NbzMts
mC9gjmB3Qo7amL5yJF081hGMqH0q1rZWZTHFf9prIPQC45a5WgGo6OW+KfCpcZtcGkGSu2kEMy7k
jhautdmswGgKr8zv2wWxTw7ORvfYJ9jODU4fA/QdyNOGEkaF/DcaX50cRdGhvWLwbZj1lRE5df2x
+F9kFUh9j8dyvJipciYbuYxRr/5VSYs2mQug8MHJc+WdZbc6ozHVjTiJj+NRnnYjiVmV6QS65+bY
MEEtqGgywwrqa8f0HJ8wXkBCH+t3I4RB72N9fvJ/Zo5M/sD5FlHSSQPhAmEz8aWMYn7aViCkIYxr
aaQTCmVLuubne1WLm/1xTNHwgblOYdVULziyrgoEc2HxVplkgEYqZIMWL+ffKT7WPNoYHHmAttyg
cAivAySeSLSmvdNYvi3poPgz/HdzbYMJncH79OCZ+TiCv6jcjxGm4QUYg6DejR17glwZBmJp73o3
/Oax30druJtVouysgvsJS7QBqjNXalzH7CnI1NcHupgVzmMblDy0oYCO5bkKN+lFVliqSNkbMRzD
FT3LevJiawNaaEmE1I9htIXiLBXFhSrG3ToDz3hh5xlPk9ZxIEHJjJvD/Xx6M4Q2q7PiB2MkArpT
75KN6x3vFeGsNZ4qk8MvVFf6XDWLo0iLzL7H9M6JnBMxL5UAc5kG3G4YIkgnrnoBT2IeLBMtLfL3
2S+n0TFCPeuPobvDcI7O4eFpKtCFypHhFcV1tscLhPBEWUtklAoFsROUp7u6OqMUO8JSAwt5JV7P
K07FHaZAuwuuyDBboisnCgNwvtKJz/f9tV2ojhCSqr5kRXNsCpuNaa4rusjMJ8hg/UFYuUM0LIjv
lLeeJYsH9bplAN+HaDBip7mF8x5/1r+CmQ37Nwrgci1uLLmsw6eN/MmXcirYmNxg8EGEGDyYmaNB
a6NNRcXDc/Ui2mkCvlZDD5T+5/RGLSu1aU7bmGBOFR3gfsXC9SYZC2WRCiq4GF77Q2u8fxsnCWUW
uIIN12Da8h4R/CNL2BrZ/7k+psMUYyjDZ3xIEmkZDLaSPLnECG9f+XFfqHMev441yFkuq154IDlr
p+WEK1JbZv8lyvOtXe4qIgKM7D78ywYETBsypumjERVY9CYbmwV33eAiY3cRlMrdmvmGEhkKrjiP
eMOpWna+ToyWVuIuUJGQJ0apwtJJHxPd6e4fsfMtYOzIWXWVNCTkX7Pis9A/OyPH6wPprmyfEJs7
h89kcsktygN4NZQutdHmiqz9z10uuK34y73KNR1jC2+49edCQXCwliV9+OO3dQk/aAmNjJJM96nl
Uq+YhAQAAVcmZGA8exoqtDzTnCLIEHmBPuHMcglW+bS8ehA3s0xC63OmWFrHG8yxcPBUSg9FWqDo
4iNZXd1WUGbF/52/ItU+U0rIqHpnS29xud91vfrcehymvs3LJRMWoBmH4Ded7/wiz+6XAOrwjSOX
cOmL+6uCNc8GYtv2BpS3PbKAkXl2kdg1Ca/sceGAcgMGgQ3z4uSQcu4c6clatVZF2Ju2on9wBRe/
cHv/vLIw+AhFx7ZF8dpd+dPlvwzcTQJz72XRSqNwYvmxOuyvIGBOzQrAZZ0J2kaSCBqzUp5YHw0=
`protect end_protected
