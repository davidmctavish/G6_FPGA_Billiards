`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kfNvsHwfdPI9pRX84ihhLCtzZoQko0X6Uwj3k1FCWoJKCkUzfBogCTgJOnXKX/v/GJ0Q21aSxG7H
tOEVQkd5Ng==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XvDh2uNCTVj/706cSVsNkIGfESfIpeSJsLc9RIn3b9Q+fKUldLkrsRSF0qJ2CKnxoObuyibhTpdh
9Z/zY+tixhPuFKyM7tYYxE06kYEwg7cd18PWhxlsbfSBfiFz1xUaZNgXawDF3REF6gNQoQpFkayP
25HqpGHvk3HvU5mzz6c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Far50RAuu2Q7CNCpC5vTXktKhEj6VikmvHdQqP7QJilvRs7qkLt8O9nbi0yjVEmeJsge5r8NuW+g
E43NNgzLOKlMcyXV8I2QJVzZB3/bbUMRDN0iv3tw+Svar/a5YjFCsxZ+qwiwxbg8Pjrt6DWzDK1t
94HoORgfVsedNqD+D/SrVX3Zj0EkmdfjujYuIP9wVNWj1hCooq31A5A1/pv28k3tA1Sj+bpB34VU
EABH7NXhbwow6RzQ/SaHlVr+6oksBMwyexjG4uVH0g28h+Hml5oldrXZ2yq24FeaoWmLvr0PUjlI
6QdoPJhE9+FZImCXbP2HfaCWli5ekwJWKANreg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BHx7pGqIIGczOSc2CzfGUpuDSkh30+MDD/PzvXWOguJlR1e2ViWvmBYM+7rmMMOCqfXY9A3264WS
dBVtKXNUXsrvpG8+ry23iA3M0dGNpegYW9JiuwMZtir3TrDkk3xiF8VN6OsNLjjv4waVLlqX3hwY
FXXk8fR2x+Mw/3S1AGY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H2eVkfiC9y+hRb8sKexUwT/5syWkkdtB23TSqo6RSYzWgt98e+dVSvXIYaDXfn37rjoBtnUoXLO8
wKNrVdP3phU0aU09Yj1P4D3Yu29w5kJxGXJFYw2RpqeaFFQz+y3YIbWwHawwo3WPqCmvtAYDVmBE
31wSas2+HEqwi/wS8MFDil2Ud1p4uW1/g5SgAP4LGYhThNHRxpuNvEQF+PbHjc1xBUx1x8xUrxdW
wwXVZEG9NlrKd0YNEx9droz+8dRJ+6/fAUrJD98acVmTd+GkPuhkyeruwcUxw2NdXcFQoZY75Lkl
VOqQqvulKVZEBuJ6Gp3qEpwVfyJG4kYnNJvNJQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6080)
`protect data_block
RgAATJWG4edSqRrZGmUp+P51RnaL2K3a96ssewx/m/YUPMO3ANg4yXQuhKhO0OVOn9XLcdC/NMRE
onozUFN/9psNw7IyGQwh4mfP+2/tFpTRKwAOz6ELnwnnQ0QzAvqscAOqfXIcgR6VDVoB33YXF3tn
o7gYqbqNc1+3sTA801YjZ07+Hzu2FIfEhMsIlnF9FHmrfTBbioCS50OSZgfWqfQjjcdadxsUI9xR
pQakHWcX7KzcXGH9ANJ17TdZUcKmNrLPvxqBl67uOq0qtYJnTtyVTrf7q+sSIaPMiCSMUhFbY8I5
qYKa7qQ1vr+/QMfIHj7/oCNFXXuxB4DAjQKjNa2JDTSz238i0uPdTlZ0uB1kmBhWzhZmAz9g3biq
ephxjwvl+Sv05cKPZweJAYB8oefWUO0+mSE6NzfTg70bB05l6IFgxUVwXalvp/MyRwVobBGTpsjm
IL5AWySpKbeXX56ycxEyJT/S8akHLSesMFRBa6GR/cdv7XC4qHacdsIKDi/0NrIJitiNoBAiT3nU
nJSUXubfi+op7oechTf0KHo+DEuu60E7vwzitiPIbttzNfHA+HCQCNzAm6SW47ng5kUjqObITCj8
af+4M2bb/BDcLeLgCIH+BhOOEZn7e/ixCuKuT8gNSB1Gg4Jp1yvlvqOHEdgycVc5/R/kfP8PdSKq
2Jwe3IpeB5YKIWWOT7H9vjbUyw6yNTHMxZZnlnM6dzR+ur9jclWMTVYGLzapemfHekhHt30zh7PR
rVURH2ZQoQ0Q4mX3Y0mhFMMYl76YqVTFZ2Bw9xbZ8kU42F+pwmmjD5aVSva5y6jlzWze1/i/hMGP
hkEPDnB1RF9zURS4W6i+MWytJ2BcjGyyw/B3cMyF/ZqVknDiypzSYQo+4hTOwE9kGb2BbmOeNd3Z
tiyj5yQAecPNGTc6oAa64rzZ4yhgOD9HnaAeAYONByL/oPsIKJYmxOPmvfD03wgjR1HgDNOTYTDI
/qRJsCJKPivW0lm/+IUfDWHdrWz8WjHs9I85y52V5BcVOhZqvwgWsunsS/k2Y+Hg365z77Sz5AMJ
bQQPYaDUIf8LZ0n3ADZ1F4R55t5vh1UnfPTyd+m5V10GsvKezf89h9QR2KlxrihMhVOREdfqIUxE
Ox+oIG8t0dMs+dc7fW0550G75Dlmld+Vs0Vpq4Z2zva0THPkAlM6Xpp3tazGt4QfnZ5GQ/SP5ue8
FwJEJn5PPCOI0KCJgu6X9HhSqx6mx8uj2p+sffiuILu5ogATDyfpWZ4PrCuFdQyKTvIAR8zYrD56
hIeyUPZMtWzEgP53SHheurHLC1C4MaBU9pOIiFEb9gMiSF9JJaG1HjeG1rzo66wQqM3JGQcpXZ8m
EsWdjimsrBRJ38SqoSUTzhF5OQQXDcszddbshDmx12nFwisL0p3cXyOl0MC9DNZYFOB0Z9eJGWyG
HlWw1cjGf123ifN/mGYl7RoSfHho7hvdXRQeHFiOg9vj4kfsE74WiCbpEscfxDQZf+YcdRsgDZdR
CfqZFU9I/vgtBwcWqo9ZXxKMK6X9dzKMBosQpUlwKTNo1aj+J6RxUM3ABA8mr77OQJ5MrPENGr4j
i5hyEGwgwFsU65PkuD3Dq7ByB9PpNcfhTq8v+/2YEITwOqRFHd+GOqv1y3YomXRkAETATt7/m5uX
vxdrwX8U3YWFSx2Um/GpYzRyHozUya1JnBKB/qYCogEvi8VfayT8Zfzh4ko4LEE8R/cRGCRYXuBu
KYmuJX7/DqvD/PC641Jddwvbr/FA5Up0Ovn3RPd/+VegykH6pBmTv/yFT/9xMYu+pPXwvpwq8c9u
KwpFnefaAvIM93bEWmVUfgTjKqCsS36UKLfRK8HqEn9uU+1gxWYdc//i0+AZenEXBljotMYRznLG
AhIul4tyzrSjdMkLayqXlmAKg195ePDfi7iT5ghcCMj1hSnsB6vpKSME1b5UIosSAYBY5QfFMta5
P/j4wVPDvVE7jlUHdHfdC+3PI230kIl5LXdV63qZ7djzFPAGLJbeDYryZadyI5u7hNyT1EnLIOe1
8RdUBf5wR9HRhHs7rTIF79AqSvMkv8/6CHcQt3c5RIu09XsXpgrn6H5ne5fQ80Znuxu98/8uKvrj
9I5ykxCWPeaEmeFqMWMa3YgxSfg3wBST6WGesfkbldUSbq0lELL3ipC0jZ+EGrG9PisTl3Xs/vv9
TK+tRwsqZu9oVp7P9zUzUdm1Hm57hAkOGVTv8lF7+BbjJHeQciuuKpqFtuX6hXT+f1g/sap0j/Zm
W+qHL8MrwCfF8ksVqEADOO/i8fVJZapr8LpyO4bv9cwVZe/sFyj3eKTi8lOx+Z9FrRIWucjlqwWf
OdIcW53JH0FC5b7fjXYwJxEITKzvvW3Zg57vwjnwv6zxNvi4Ia/VBfKCcksIFYAeqg9ww1s4ljFG
MpV2UhcqfWoLxRCiREhtMkXVmdzZ966LAwadyzKon8NhkBHzDldpEZmap7kAfdiUg4ikM68Eg56L
CZYAoe672MdwFS2XkbaZ2eMyeiad5aMkNPvyZtahILOeCMAeTy41+CC1cv5IkrwCMaKKQoh19DHk
+fPRXxGbpSN/HyI62D9akeqPFkMfHB5u36YH0bBiUTTlk/D8OcMaLbwLDJZ4NCP6EHIjIKBxzUtm
mEpWV64KFpW/c875RMldOFUyZ7TrgX5+aZxx23GlmKdGL9JXI8irJoQhLwKsrAJru47Hn/vvc8jm
BDdRpIx5QoBs5C6Bi90ixdcQLaf5FBbeV40WRWPig12P9+HLHxy3CnoTRYiHcWbJRraCaKqzZ5Id
3PmoVwpdpZYgTpyXcnjxcLq/WgWmRvfI9M1t2rfhEBVEEa7e3k4AFhJUcT6sN/mDNdBZuPwhpZgp
IQ5ULEiANeWMAcqx1PIkK9STiU1eHmNOz106A6vf9irNwxou2iXSJQ9dDrsf2MFP4tFOM/zDXicW
/Fe/vm7cfHnFdTd83ijX/+4a2Q/tjCTQiZuTn06QJernCqss5J3uIDy6dQ86jWv3OjtvlnS4Tb0O
fit1tK0SvqlI/9Sf+xIxPPoBPf1tQq4a5lpuuixgUSWjnDMFRfw8g9MHORPYOSghs2jQtTjvOgu9
pwYUf4VeDcET5XYuXobv0u2PZTR+p4SVIO3/0vRlIVktnEDZ+LVG1Vp+OHnpQKR/xClFFdC2xDi0
LBqtxU3cwFqk7upjkmb/wrpEl/caFSqcP4uG1vmGMvbosPTMLU3KubJp7UOgtKmdATp5QobgZZHS
0sx2ZzFeajyrbP/PN8q9LWmKRcVdsxYbsFxI+BwH+wMgye7vaolCVu+YjjiVW7v3pPxuGAKsoNDM
KrD61G/Oj8zBr4LjTI0Ss1FkEXpLnw69Q8O7JwZ0evNPGs3ReaFJ3VtYfQr6Qa3KKOvbltzh57j9
MEh5BVAj86nHyOycNuQ7xisOhg6XkvGlS1KJGN9jKvf2SfxgmhVhCXYM02SX0hghmST1f3zrRfIJ
Mh6e4xg3ZyYNWWPHVk8LHbCpyH8h4bvUi/dq6HvfdxQs4noOWkm5lcbja/f7B19lbSCWF+ZnVNYC
F+yEkmNdfckluF8yupzqOH49BKLztcVdbbjFWcAO0Bf1HfRdo9jXARthwovTyBgFGh7BXgoNeB0w
Z+vkWtnHHTi1OIJer9rDXHCrxDt9cVw0mB2H7N9eQQZuvtTJGj4+cY3Nc2FcpVXyPS6NsqAhjcUK
IDeZ+/x8BhM23iEYmxIxh+LfbpC/y7dKarThsCMAH7NNxJxJDEH8r4e+60d9bmPUTFQrCHpSsRCp
xBY9wZ7p3QVWqCsjrqI2ee6yYk34u/3mr+ytfhGImrLE2jdOS6pac6dpzFQOxQgMI9HC6oWvrKJk
IQdNpOle7u7vjjXSWb2wtx02GmlEYdouzDLKwgr+DIkOb2EO6D6XjXNAy95TPLvyE4vj4nCxejeu
q6g5QTnYm+TNGRobmC2WG/eiM9j0gHXn1jYbALnC5SsFXv7iiAA8b+cAkcVuYzyZwDl4lFFkCDQq
NN/vVrpJ/XSF7Qbr/3yfMUnfk8q413HnqV+Uc0VXqwN1JHX/iJ0hE8PkzCDwclmfOugVVdetPAiw
udP35e9VfDH9q8d3DbT5MzhA76KZTpO/CXyr98j4iJyisUtWBuRH3IMOMRpuAVFDXMr0Q53CguMN
gsedECO3mdYIKp8EExafmXfAuCH9NjtwfBzwccu9RWg9CBWKanWS1QIxNX8cOwfqk4rh9zKeHdUE
e4g+yg5E8VMc7jXHv5mohNDql0V7Vp7NqM3JEQmdxO4mYAddXFE99VXiVYRY3d54cGmBwv1dA8NG
luirLlqupsP3TlfDSMrN24zeWHZmd0jGr4KsQYzDQLr2g/4OPfv+xZDeDHzoJ92n3flEl9MYJj2L
r3O5IY/tLi+7VWy1Wy+FhrcF85Va550rlZRMW/cHXUDhwi3zqqurDtJrvVHEke4ymMNtIxTLuILm
iMQXF//XRfB278BKaEPZwe6CifVA1/aKnGlm+LkXyzLYBmr1Mz3XsHdNmmvVzzXOy6BP+pO6ulq0
b9jr4/LGAFgttOuMAhmFJiXb8wjMu1FWdRtlMmOwk7ev/Aihc79tSK4odimYlkj4mzzaGr06zWM5
qYQF2irDkDEb0QAH6JV1aEXKjB5X9eBXw9BQ/rOzRvx57Wng2SaEk4utIbMja3SRPEuslTJwdOeL
3ivkUCyJy7W4qYq5wTU8KT693/nRhB/Yws+lUNonnMQCnhs/p4+vCUgU/wJAGv/LMD/TsWfXIT21
9CuD0GiYtQsErMxwdptgeeCmMHR8RX7GA0GUnGUKoXXa5X3mchMuPokc6Nd9C6Pb6UKcv6j4vymC
vSrtOb4bkJ9XpSMnGmvDnSnJHT9Rb7Ps150QOmTadHfgy8fa9iV7vBQnl/efmiIwC28pOwgmPeDZ
fPziXtM+761VlCqJKGQ2VhcDwxN0DjRJLdiWjMIDtN0X+wcMLzCGofsz3rA7GES8zf8llkfDHZly
TR7KMTCvhlm2IINsr/P5BtahNviF7Qq2dJBQdLe73aaMx+J/xwy/dy5DCgRrtTTcParolwzXoB/r
A2r7NjQqJvA08lQn6ZQT7JtiohrLPU/UP0Xcof/1LlLSrqyxl8VfyCTMdQaJROvO8L4I8qjIOOOq
rXyIqjxaOc3mV+yccGqjvCYqsIDuQ6kKkSLtRDBV7tI7wZx7tH/OOj4PlodrE8Ym01uUDfj6va1L
SkKwwUXOFozmKVENedyNktC9QPWwQe4EiXfJp3JNA5+JsNlhTeMsn4F4zuIrS2wwdm0dC9Wxsi/b
KSzoPcLXCeUpuEStlLKE2gqryGvZ6SRUyW0evW3YWTN2mh5/vNmUE31lBzuj23GNCRC6wpdmUt8A
y9ab8AwIs6sNsP2uR2UzEuQzVy5wHZy5ROtb4Z4wT1MC/ezugNaPMl+HD9Y4CDL5Jhq4t3pYdbPe
dB+HarSdw7+ZPOgYrxCCNslA7fFy7M9Q1xouhza1trdB09Sz9bG0b0/s6BMltP5OYdTtds4GB/y8
Geif8aN+Z/1+K46hizbWNBfkkhuHkZSXF+vQhO3UlkC0eAkdExHZM7KunEgcvtMNYTJYYM7kgOHD
qr1tLJ09roR9eNhsW+jP/zpPboLeN36Aqfqq+2lyAvLjN5gflw8UOtcmxzNjV/V2icith81w5w+2
PHhOLC92zs6DKExL7IM3CJSY+pmp+09eubX6QMa+ijHAGI0a8oq8+ytZq7FmlIS8p3rEanCqICQC
VcBAmjgYGEiaaW0Gz/WBbtmRs9TqoN9DDd3iPQql7t3ES3+6Z+Ba3UkBuW9vTeC+8ONpYBB0lHxj
4HlgVzSTT+Td3YZWjWA9S6ypPPtvQ/5odHliCfGHGwbu51ApKgQ4WMR7LsynSf/Ybi78DrWagiHN
I5nZgQuY69mEGejSikI70OpeFxY12Udu1q2V6GSN1tk1QQmG6kV3J7CHshHJdhprdoAg7ag5mWmB
AY98pnJxRLuZ/QX0QIgCArKx3R+oY3HlepjEV9DJQWpSARyqSoojeV7PzLCdNIxF3k/d++pwiJJ0
PU2C/o7WNzyr9/3RGKrW9EpX+vogqO6q2gvxo7MZWl5vhqhiMZPc57a4+xXHxA6csPloPlUfUBmE
A4TFHfJ7o5UUUdtRD290/+jLDowwTKX1CP1EJ3YsW9CWIAQW3qRea8l7QuOvCtHbx5zHcdc8MpO6
CpQBBMME7NDhoLgmVWjmYIBeqUHfRwlc/ElXzdCBDhe/b4sY7r+rbHzJ/8iuS2k92OCMcTPDPpC0
9Iuj41DjKfPAKvYAYda5wE2j5P8zn8li6pIiqqNGiJofWMOyxShZDe6/eM8HUrpvdfHh7v/r+6nd
SoBNDimWafQwNRMHTG++/NTBQuv2RbT19VqjfnZyelVPUCtTs2lzV79DM49vPWtvZE9jK+UQ5L8u
wvC1G5rFMM0T5jcH9jX/wbUbtoCycGJttG6Z78TAnUhEwjc8R2e1RbsGPZnihzJOLEY/ki1XvMHy
0dBC64rKLtejamI/tKqXjplfthMkEYAxK8JAkxBVgz7oZic6DoT9FW+RCGoGZzshJ8HXUeBg8Mhs
sNdaRAsB4C3XHZn/rzXvA85UwDldcCOMH6YGCV8UHtGpJeNYGx9cyp9UvMO7DanPYvjUoZelEL7S
aMAMjle/SgHrVzwdyRPKM+RNjxjveC0XSexjcbv2RLyFOXcbRsNqzlMIHPvdPEliozUBLdij9tUn
o9NBN/1hYkS7p4ZhehvfjSdSPHzZPGwA5g4fdsLOKa9plYUd5KUfmusLcmHU8wgYjfMVKoUSybgH
4RCyLEH8oyuJQohDh4q8oiCeldXL1iXtHcoTnccTosDXakevJnAcsX1pnBvS6fXVTRQi2tmn5VqI
W/0dF+MbfwtJj4VptXAWhAeT70W7zxCJjO46BsZf22dczx2FlBCpTLCWhHAiitv9V/0HYV5sg83T
vm6gjsDwzN5y3SX/f2SJHqxWUp7VlEKSStpHJ3QULOlYJpbWV0GcNt0YDEWWHtEmTknx5s38+FKM
aY+sTZmZ6Q9bqupAF2NVlFJmOfmveZi5hg1RkhioQMlCYAmmP+BsiDKBRqH/CiRPxQvpy21NPkza
1EB8vKmclSweuHchHH+eNMXy4Ob0XXs0yOzcczgfyD0YsZvBq55TP9cWqpQpYcN91RRu2x1LRwnf
taoTCtsVhba356XwdXYaRSgW77tTJp8KgHMDNpEQNyYO8EfbuAEX3yKSWHmSfllefSZvxolF/DQK
nX0NOvhqf9RFm5LS2YDnL0X2m3EQUOmUu1VYqtBB1uKmf8wy59QwdkzUl3KPetfMbszehyaYTaCD
rE+PAinSc5X/cix6r4GXDuypDhMX0JSTW1h2VzzaDWtA52hYUKTOO5vqLVJx8m2qdoQ326vkU4+Z
QQRMUcfHsZCnflxzqiJ6uhbJOi3HsS2x2NzPMvr8AHJUBlv2MtUGyfvm6/7gaCAhbz6qkQlTSHe6
hJRBI92eZ5RfA1zSEQBXa/RMqUN/G/S2PWawBE/XsXrQHpWvM/zK72ECE8q+H11LRiOl36Kzo1aw
g3Y5MBaFifo3x+E+ZskrwJxWZzW83DZGwI+hk2aVcdx83Zij2hQl/pr7PDdDf8jpdEi023BaQsUO
XrQNF1FSJJ/+V5lAg9VAI3U9asM2OL8tBtCI6/gpLC0Vrgd5twVrV+AzYe6I6DaW6eXE1zV4Dlt+
I4aoz9LsQWWzGVru8SlUtvFJH/5vNm0DRM0f/9qDASpPXvvrMxxksj7qWHjhY3GCdRvcHI0XF4Mq
KVo00BoKsBZXRbsI8OAPqDaomJmtjhEn1FZOoFCtsWUwUYYQVIEyMV39qNmyaDcHMo8/R21IfLTr
hHK+LmWpLQmB37qo7EOv2fIoZ49PSYxtLsdiPpz/v06Igau22VyOOi7Ey2KXY/ENVdhJM3CUXffI
bNbEwa7mUkJibPzAg/W1ZOqV4YLWBAnxWyk0CdpKUm3q+FihkupZ/cOlQ2Lsw6efuCftlvJXlacn
8AfcCtHS6IoIvNMUk0fcvPVVYmY2R7Turq0sDXafLTz4zY8ytUA=
`protect end_protected
