`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
G8f1gqSMQCnQAMasovp609G+Xtml3VQEkPOLMPqVhr1MIayxmJvmZ4o3wKbACMMSFBE4+TcLKolU
Lw320DyaNQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ug2hg9EpJHXCwIW/al+lR0FQjskKd87pvEXs/ZrL+skznkgUSgLQmC7SJ1oq3QiIqqkep7bUmCVy
we8veKFtu8UfykilTmrnjhTRdAyMYPoc3U6Xbx5Lq7rKnI/dAU/tITqfnX/1RQy97jQ/SOLgi6Dx
Yo7ZJsrm1WJdM+ksPHo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WHtDk6ccWwa0v84+eT11XdXj5G/EYMvPkJ4c5ahUoFGrSqd4gCHCAiolaFpA/e9DhneCRB1la9T/
pcL5IfFfIGM3uNKFFSit1QvzldlM9fpLEMG1OdKNnCRVWp69DgncRuK0JLBlQrlzmwFPjSPfCkyT
SEkKYrcZY2nTdIQ5SLbgqmjNzBcF93ZKwLjze8ccIl9IKNsMpuM1vjvfRM1mgbHdq3Ml+paIzHV0
xzVAzQV7PIanAnzCPVohQpY7U6lCMXZhdciaVjLnPU5sGZdsbkX6VOlL2+/1RPeyueXcWdtS++rj
2qxFe0Bc7E82KYYoGLqRi7Kb8S75TETIsjFkDw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hN3ysJNjoyNBp70dJlaVUOhqqcr2mzYQ/HE9e1MilSDPcz/jN0bqHs9I5KLnIRDQVc/IjMTf1Hvs
CXBTyaSSTFYhpbstaj7kuVfj+BSQj315KjRV1WRKrqyjaqC3oomV+UaFLj2hd/eYIDHnlBcZI0Xf
jKHWzWg0zMrOnchT9Co=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UsVeqgYjuMLz0rai2LA/hZgwQYWVqJGgjFEXQzv9Y+00hP0ur0N5wKZ9COZQf5vaZTwTyOuPtLrX
SZ1NivgvLjstd7l/BODfmRL2canlzh9O8ND44uYj8try0D9PZpZwdkT2+zPnuHOxwOFn6VpPXRDB
8FQLsnOO9RcGzwbgafC0XYO0L5v9yMpxHheu0CqhuQIESPCXp9hByn29OUbPWz+JzoxZM9/hX70F
Rt4HIj6Pw8i0zqLHF3yApqbjUxE3z9pw9XF12lIjbLj5J13qY7Nvp8M071o7YEVT56vnb1d2sbU4
7FN2+vPsLWjaWsmIWAB5eBk4jEavWlXcqmKlbw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10688)
`protect data_block
HHsQld+/7Dz+EiOmk7gLHdNnjCBw31fY64ZvJOKWIqDx/80No14YTTrE1li9v7pnl+KQvGfUcjW2
KQ3j8+Z+QrBfcojaRRbqgsCEN3VXRR8tvvJg3gcd4+Y2du3PNsza9nEQm5fgWLCRAPrEQtqCAfaf
1RcYBqDQ4CVO87+eW/usEHoDNO35oggBpqLI8bAWJHDvhbRedL2vHU7SFbYM7TLBwgo7oxWIX0Pw
wpE/ONYAPpOEAiSlWIfWQLpzZcEEESBsuJNhcl5suVc5wloVCby/5SKhpwpeJOHFCWoKuHhz5dwC
Vqk3GomybRHbEMPIpg9px+tMBZSIFHTq0nmcsUOJbjE0MUh1xpQfWq6UbIvdtz3SUzWz39h4gmP+
zdCGa+3TmEI1GILj9hgg2eDoRuVcg9ZnMvKkf4UU8Vwu9s3hSxdTbt0AbKo0tCsVSUDRAkOkSGZP
Otgd9r9Q2foNREaPP528cIf6ZTPBiqjZ9NsgoFY4bqcBRYACy7YPzQiIniRKFa+mGsU4oWzbmbZ2
WFhIhRE6ugan4H1fxkfxLoSYLzTx/az2dPiI1hfRt1OdDuPDdisrSt0kPcvTQwZWLcchem2WcDTy
G1qrLH7Z3hx5I5UJ1bTgb2NWq8c807i9U3t6vawpfKHA45/WXrxJkuK4Bse7GGYJKiOgin4O1nlr
Grjw6zqc65NzRwwKG4C6DYtBYVg5muz6wmTqTSrOT5OQFX+I3ozS/jUNfhgd1zbF/ojhvdgr2k98
OhMngpmBlOvXPU/CWBqR4MEeMzUd+GsXhqV7W5kdEruzBx7x6nFj0I8optuwkG/HdW+Au6trrqm0
TZljCLVx9FCtbMVnfkVTN2nBr+d1GaZnLeXCb55HvgYJxlqsbcG399YHChCBKBny0KPB6uikWVl6
4f+r+6H+MBkywYQ6/tFr1dPPBW6bOAnXeA6W8xYv+VCVdE5y6rlGkBVoXaZnqxzrNRi0IVb5QoE8
gYygUxtz4QTVM40Is6HUF5lR2o/rcDgQZrmfNHu51W28mbOkob6ehToUPcDhhUsdgCmJt6C9oqC/
2XkfBG931GBN13y+k8P1XEgnczCqOftH/JFfdqqA4h6Ysc1dk4FtRXe+jHmYdKQ5nmTcVL5GqLQo
2AkYkLh/RXXGKiyRgOVX4JLM/J7mbWQsK/SwzzBdPF8jLrOZMHA7fF3J6OsjhxMSmAwvg5BjS1Kr
yw1mfi/ooPuf9FFmxjOoiubyr2JTdIJOcCzSpmpZg/RxmaIyRfdWv2DZvPfxjrkuc/1JO/QAjfzo
qnyb4Dk8tIpik+BXtjejsYh2xm+f2BK9O0V7ta031oDhhcdcSI/8CxF8qY5Wub9Vg4hJyUZp/xS8
+ORO1s63FdHiWGNBI1vJzn2uDXY4EKTvJfZk69nh3AgIk2n95FSP+0O3oFnQTGWNGzGRbAsqUF2C
mmBgF/Y+eZgjn4fwQ5+KOcyOYHiQL732ic6FSfzN/+xOBNrgPsfsuL16FOe861RgKLhKx2wl+c2t
IW0OzFWCgV6SbZorsG9A/c++IEGwK/10qU8GVKdtKoLSDNVmWLikF4OaV7B0SryF3DGRgJuDHnWH
m1RE7rvqbwRLbO6KLN+Y4cEpmuO10GP0iHRaeKK7G5p0t/gGgpahlS5PafntE6wfKyra1i32EleC
oui5JjAZ/3dLcnimzsOcPMRSBKeMOrpa8av8moMymiKoej+dsYDbnjJhrEdGYitbn20a7QW0RvC9
SDVpFC9GgOenhWqV6IxHbhMq2zJa+hj9Xa7qO25ib3MZmBDoGQVeZsHbBsvK/ByijQ9n2KxvTAsH
No39PfE3AaUrWp3PdsVWniex3CBP/aJEsZuvoIXeFnAwWkZwDhDVPxwkpl+S90DYFKY3vBpnj35U
mGXAkLV44VEejrb+biDE1g6x+o6/2eeLqwmouew4U9em7PxtMDdoljLI7LprDQ+sC24tQgFxNGeV
XE/qHr3G0ieGUkuAZvkMiy0TvE+HHedYXSJHVkJlVDNr3pUQaFk0TKiK0oBlQzd0pBZdeFr8MywW
LQQDQuv5Nzh1DHWIksd7kxCS133eBDipjVh92XKOJ1Yj/W+LcRUYdc+UHKynjhA/HV2vNY8kBCco
M5pgFvQfDd7JB1zOiwM7C2x3aG9uVg2zp1MTjPLI6myzF4d4xaAz8a+P4uONLXMVlAmQcGIswTql
V+z7CbOGcmmZmsR4EJsIes0YkOjrWA/LhOESA2WYhGKwbFUmkQVbKxIZ/qZrqR2prKaDxsJpB/Q1
KJZ+CvUaNHAu8xO+z91Ftki4V26PIfswL5BERN+e4ry1eHJzhPOfC3eC2wvK8oR1elwE7Fwi6SZk
COAR4nz0A13YPWN5YTQffnrYQ8K7qkjSAtBB0Qo9Ob9lp8GjfH8ytzegEbfFCBFJT/y+wbBQeKcb
/1qQd90Rfr7MuFzjkY2K8+HAHIKcuScMask2qu4HybSYKyDePNXq3As0oJsuMeDlxJ9+YrqeRzgR
angHRgBFfH1ZqIW2sRCMQ+flUQwdw9e098Nv9ZYm9uYsTVP221YzNnbOP8lNWPAqFzJRgYiC4pvy
S+AMqD1GdELfeN47XNZKN35ndSDY+09TUx0Oeup0Fk687Z5NhaP1zXfTSpwwyIvJth/eVSx80UFw
kOSHuOCdYxF2HX7KCqWx994AgZowW8pv0Xh03fyXSlY0lFY9lAVh+amnI+CHbcb8zm4EQS3HrHMy
eo8HWSsiemYl1zp6KTaLa2XeJuA8JcJs2A7Qh5eqRkPXT7fIOQTzGFd/k8sE8d2gNdEIK1iY5TCz
Bqg6mJIAnwYNXx59zrG5G1cjnHWFMgRpfB9beck8WrwNqZBLFLeIiDgw31/E2btD1KiMmTJNUUeT
xzlCM3vcF7NTJMt5SaadnBnN5TBoQj2xT15Ki7Ymv5LDVR52AnjPL05CWfg5oIYLPWKyLD+Vl7Gd
YnBOJvOeGdyb2ih6GZXCCbQ9wxVm/Hh5m9jQHqf0/5WX5ry1UdVsdXchvIyYxAjrCiLMI6X1nEOu
3ikYftBeavMC8+eQS44Qlab1OHnUJhVPJtWnekoguEU9eAW+ufNp2OP1Nd8ruS4lgP82MVIcSwdx
LP+Df2ue4ZPNIzbrjAaAusH6lfqVCGOmTz7Po8HVkVL7Ga+pDjoc3M6iQR1Scg0z0E5Hqh9r7oJ2
UOhwaOmFir/2icNfukLXM8EAkIuDg6BWUMzMDIdIZ+f58XMXLSPPl7q4ao9kHa1U7+3rZW4q+E+Y
ws8LOLOqRwiNiH3ySWZcmYaI6zf83bZzceWXSs5CvbCELMc0k3y2eHewGEmvnT2LETxAudBfGK0w
JZN0JKDP4TvyZChWQ19QDTtClEBui9XGzOD59E2LzrbCBc9Aa+pqHOPkaZnSdeXBpNiplW2P7bJh
eSKXh/jziCq5zpnmeZzj5jjA4YOJ5eMgg879NJV6NEsncTIP7dOI66TwQz3Cjgz4U7WVrRBbM24B
vcPNCUmNDtt2hcvOisb3nc80duTpF+oImp6zv4wOHBO0lnzMUd2kDXPG6k97U6hhFUULH8E9udKm
ZOg7zSEP+xCrHOKuNTGk1v1AkWOwWrR+HgZwEmJITNjWEf+UdGJe0Buk3PfOpkQK2KySUXgZSXzy
HWsdgtgd3KL0TqYiVNQN1iHd9qz/0dRQuCafEv4WCYjsGGMj49x43AZo2xXkb9cD7qb9skTpImfd
vijnHdQv91OeCf5eLsTrgYDXXSJCNezjj7Z0OZPoaQ6bXjXZUOGvTabvjtIOtAgN3MpKk5Xd7/Is
eIscc5WQGucIB1Q2BFAUCluSn9gUEoF4n1hoHi6wp2OnRj7clMngp+DCx73Zqw2p6PvB3WHnaeXm
83zjmC2FDFgnGKq9UWLzl0G1Q/UnvKo8R0kOnWGmatITK2scMuqJDdaTrOesL15lRz20yJiBadjp
glS6sd6FDhz9d9UBmc4Pv5XqJRjGh9Mtpie4NIqP6d1mOuJTlinbrwO9yXAYEXM8hxfaRvrfTlb/
3ljiUYy89RK215fu2cx/GshPKeWcC7eTwI4H2PpZOeoDo3X0fVvPfluN1lUUuDDPUG7YBPxKZtyz
L+JCTeuPQs8J0GcCBGYcL0wDBAiMR3Nzg3jBw0rcjgX0ryOEhjfPaOEYEYXcjbKJ/2kinfKVL8CO
cdLaMEH36jZr99T4Ar0ClQtsb+vn6SEKzMqYk7g/GFU6EFkZdyz3vV71R3o8QXSjXBHz0+8sxA6h
wVDgGdSAyFKv8nIB9Qm7fXH03pCasLPmVFI2+4hLMDWIfjRVWLNv8Su5U0LOPHC644os3xx+PkB+
U7ofxyw1tI2pTNDNBthYN94jG0eanF9Dtxa6mQ4oR3gHrvv5cUKxXiX/Ch/PbZIqeiWMtFQyjDC4
OtmvJA0fP03MztghfxIadCj/PCCu1G+82ZR7CWggOUtnvvpjylnz3n1R2c2dbfeg06pjbzNDOHAD
/iuoYb9BC6S88/bg1g6rPGKpsou8OJXFSG27W7c9HnXSqQmoEmIkg/jnkpy3GuygoYGquk/2kgn2
3n1dgnbVvRVtTjyETGX0iGczsgf1gRvWRWH2V/3lsjL3com2CPAv9e9g5AIvGQg5/CIgu1z1IuF4
yS/Zjlczyll4r7aCMnSpH1I55ihjR+GC4ucsjY8eWnNDOsKl0UrlH+jJGzdXwWe81nLI4jnJKMhg
dCwjKoj1THQbYcopJ+RmCiRkME0kkNRUv2ukTupaseZGuVutuhaU8ZfN4eCHRmKcAuvkcwbJFPeQ
fgguHzqOkXRT6XgZxULbJHWQf3axMRFidtT60vzLHsZNaN92Da8rKY/QuYyLWqucFWfhvnG9md5V
ohtp3z8phCpctlL4rHLaFJDq40uIXNPenMRTc7Vt8fs3nBZeM9wasSJRVEpl37repcohGFkhRNeh
GjHSyPcRw7xlWjdaNBsXWvqyZjaC6qKyuNr0vk+LAKTFvw0QH72oQoPzU7v9TA8ORp8OLMLbUGan
84kUQGvkIoUDNi/FYyaS8lb3vLM/V+wAnsz7oTlplNPS756CrllM9C3lOl97OLgYTuyQntDv7dzD
CGC2t8cbinUzbvJVH4vD5mJRz/NUTBAROloZx75citPsagIRItOPbTvAlMVxEeIUOmvFA5/drE/E
vxXqnCEka5CWUKb9h9SGCGvAmw3+VIWxWPTpNWJfgwek9LcamkDu2ggs6W98nbwGFWliv7ouI1D0
YSF5r7/PHvN3Tg+n3ogB/FWMfA3mvngHfZSbl68JffQconu/FllpZ2TDP4TpmiIjBZ7T3BZPK/uK
y3qi8vQFUqZp8sAXdJI+aTUIJVsTIhaA0HrX+aV7wnyyFpqm321j/chz4ZJmcDip984JrazzDqaS
uGcJBwO6FVzcWmPeKyJngUEw/h5yxhYxc3f/rqggA8fdtBm5zbDgODxDbdGXBs7PKCeHexxKAD42
LSSIMyAaF3x2oQ85yuhRaNkhCdh4juBvbc0XwMxn30xonLnyya84Q8iQOLcLy6t9bs7fJiktVt5Z
Tdj30otHoALZY6giZEdZRX9t5lKjZrKI5aq4z5F7+42L7afbaCAeTei6a1zRjkAslI/TkVh4zsAh
9yxj2Pffw2PhwSq+TV7KEBwa9Oc9xJi/kTKzx1avHwMgPS1DTYqZkpYwecb1okUbEggYvMYfQEe9
FlwytVY9KatFYiaRSB5XjwY9FpueU+ooQFY7cPg2qDc0nYLDsgjnaIzysuYDL585OJLboQ3/KpGQ
hNpZ7SbPmnKrZyZG8L01K46/W1XmbDOj5jBqbhMAnn/o8lE0xlkNd0qJ5NuH0UQOKQnkMiWdslkT
0giPAPhfB4lU5OqXy+3taRmiv//4iCHD7faJQ7/cda2rTLuhsIAQ0rRmBzTrKat6mh8d95jDLm0E
4I93ewdCNryCNQD4n4vmUhLcoZfiUJJe/iSfuLi19bcseWILvYiKOR2/xsP+3FoSZNpxY0R+zuEV
SCUSjB2ECT1+oOZm2qtlJB5dk/kBxveu1ZkynQnjfJdX/7WUfzZNRPifcUuyST2XB2cERLO0HXZ7
Go00HdYx4uhs8cgzJMxQxedMN/lXOEwgWle8daVh4Go7W0QfhmSuqKTEHwtJc3qqkHgYMcJr3DjL
eEWKN6BRCJ4zI3m7gT7FFqxkR8kOXnVPmwcdt7ZR541FQAw7a4z5Vatd5MHQcZo1T/xrYh6Jx0IN
vvQzgo14jdajuuPvvm3bWwAi0/xZ+USx+56AQWwlbLwpEqB078bm2zxl1hpEhOkloaQI71Il74Nz
a4GUAF70h70pS+ncf5zbbSvwaS5Xl+reIVx5lDuBtTwXvZOgg86mOmYdeupIuzDz+w28V8WenOk5
eiUtEAd+FgP/RL5qzNSgD2GmFm3tJEb+pFdt3Zq+eCz8u6+Z82Ke2t7lKVfNbjCIRFXu2D09v35A
Swhc8qzq/m6c1TMoUlzGjr3Tnkd5uy6v5aPmXryAqR7ZC4UeT81r7/4TWzs06Q0Yx0jLowT3MzdH
3ZXLKyjJ7A33MW5niLN38EvJBUIObmlnl5f/Awpox5Q1h+j55hxrJHYVaXsjMmhyHeuPasCBm1pV
PFMtK0yCtiPOpt8VJNapPwoonrxiVU76RmgGBPguok0ty521tmizYDpePdBX53lteoqJLLvVrMcK
KxSgsvkiUEqneAUkuwQxglTAAoUT6PpJ/XEybBF4Vqq4KyVjnzTufwIfG2e+8f/fAzg+ix5bJCtv
lgYdly10w1VpMGuQOxGBHZ7ArwJIjig4w4Ne1A/shsKShXD1tLHEXqk0aA3BEWYnicFswUI34os1
H+pcFk+2IUja6etA51BgJe4OS35zWAuAQ1mXTq70WI38ZCoEaB74UhcLuWCN1omLrEQ+KKK6FQbf
TdsxkxrJFkWdosE7TXFzbq0v+pNjVDZ0orL3F25yJZqKxZhxl4gOevy7HdJaPWWSWNyZmaitybEr
nDIpOk9axeQAo1e6/py3gG1pyAEroFks1gzh/BEzkIGjY5JdIdZfT2bkQY9cW0CKcbgis/0yYXg9
w/sAykvQrWSOihxeBkcPI3cfStuilJwuXh1OJegSH9Kz4owt0xikAU2YWjPoyXaHVB8guzAUueet
h8qfOOLo9kMzlD0IfAHhxCNdx5Cz/3CII9SFfUitRYG35lHjHa0vPwU2LQIXhOkhgxAmRL+v7M9E
RwbPUH3G4o2AIO6Z1UGcAModkNT+nwkjQdoo5hDKMJ40+bgev0nbIShWpygcNKRxv1RwCxCwuFJd
J+WL+GYepcyazEObMSDjZDW5YlvA6snzeuNugX90mc6T6LrpJuoDQD8CLW68zQQHfxJ3q6PbfIBd
dfmgBjWoeGcBudkmBNiJc8GBz07zsnnSxnsRptzvUWcVsVGP+r4ztrSS88/jihRLMd4w0XhILyWx
noj50BgGfeqEU+smkEEotXypMT63Qzra61LRuxPn/TCYpW213ulwDuDq2cxdjZxFaqI+6BJBrcV+
Ov3xekwinpgHPxDkWdTP8vn0NVhDUjn/0dZSzbXaA3vtNAB93OP2RdLOZKcxJ2RghGWI8uC6t7i/
0hu8DXAvuaI5UEwfDOcaEbrnmAKakC689EJftOk06d3CuT5ktLiN1GL2lfOLfnpN8aW2zbJ7EZnf
RXyviVtqeE906KBJKLXcS5wbMzhMBFh5+dXH8uw2L92fO0EU2uETpVH9hVKcqw2Me3phPOfF520o
Cy335DklPeqQCTskxdsnI6LT8TDpdO94KTivj8l9Nad2jsXlvlEc2deWQYYp/4OLAuFYq7uvB4PM
HjadFs09qoPJu+/sxvrudAoDabChblb+XL2llJY4nadZpwfCMqns3OEARaSwBsLCMYXxmJHjhTYC
S8m0+vYDSe8T76teQsc7OO61HI4bckpz5Eystv5h/mz0PgSEIR8wbqX/dfZ5NWG7Q6+sHssb82hl
t0UG6dFrwnu3CVzIJgeE2qKjSj1h4useak1sR1DsfiYemC6XesXvnR90Q3SzwxHvbwm/SqiGp5M+
8+5dLQbZhkeZufU8Z58EbGRJ8x0iJCGvHmv0srLa1L0rnXmol7idvs+k9SroK5pJ3GsIgZdTEacv
pqqhD4gjZns2Zrv0bKnpmQg8EIyur6Gc4eINkC8GGvdpwKYmym1v+P9dPAQwW5Gq7L483aEJ8HEG
FCXe0yAHoSTOQWznLazhqsOjAtodxnquxUekNFaguOLXEwJMelShtQRzcXOUPgAqx2D1of9daS/F
mbPQrqE516iMbyqv2pSgfiyFB8a+4RiU8aRZR5qR7rwkpAjXoeGx+CgXV8FjDGm91ofJL49yC8nr
NNiuQ/zf5ueWp87J4tHjvhQexGpBdr8NcAD79kFswWmfrpnL6uNpE71zXyHr7XHoQ/FLiqgDcixo
kuoP+LN+T8Ljh7Qist8+e9KFx0NJsoKLBMMF7zuuEVtd4KylD/ZxKk48kTUKioLPAM4ZaFvx6jfn
NKmpa3kuQCWurVa5N/X2TFQGOkvuB9cLKnWKTyIT6fmfgwBYCPDaBVkavmL0jl//tNn0vPc06d5q
N9Hd3nTPVX6++RqBn71skXzTNRm5+qYsGD97yU2rFl2n8NQXY5pUFOvv1oW3mQdzFfgybRL0CwQm
CPA50NoYXEnUWyOQkkpkMg2U9TyS9G+FH2XnH9Os+eZJcpVm7QFgeRyNFmYUP7G7jrMFmhbLlm/M
8gmC0yffvsfraxYjrcxFmn8mP3fnQPkQMPcEs+yuPiKq8UjEZD5qaIkjgbT8ytDryz33qY/JPC4Z
VRMTyGPt0drMu+3eKjdiILe0hIv6BpfOp6fCjpDKhDGzhipPSC76R6h/RFRfaUZKl0VwmTGLzfyy
6VpRKQoUqmFBHALJk1BnLSfmNXC/7ERjU1DMUpRDTUUHfAgHpZt7MhQscA4mSkMecSuOhkDx85hi
wABQreKszs41eGS2Ew/vTaExdx3DEsWSVQAwaraildDpMtalkD1vkb+qU46BHYlobN87dLVaFd+v
SaYDJxZbcSyRIP12Yj6t3ZewxIYIt15QDq2XsmKlnz4q2N0bvjAs/RSXmUzZqdZ/pGD3TzvEYoa2
/NDpoFSwnhDoWFeyPqOpcoWjiLcHBwsEy+UClZZrbDJiw6StvwJPhShiD2dLG1pt7Z6UmV8Cfms2
AgY1bWG2hAyagYIN1eqwcspiqQMMP5rWG7ytC/5FsWtokjJ434hNvwYf/m3h13eBxTrQbqm91keu
TiKnE4RK/EpbFycuUiG+2qXLAVPY6OdS/ov1X82YkDe79h3JHK3Z2oXRQyAnrLyZHx6lXDc4C7+u
UzqZPZf4dypc/P9PbJEhF55CewglWQUFVel6ZheeWKm4oNGRLfXBDX2XXKE8Ldy575Mu9nNSZRUw
/qjCHdPaihG/yUGwlB2Qz2tcI6nfsVIZAHTl+8cpo7r2Q5jOoAHcHqqDoilhhT01/BvL7q53vxin
tuFlWkqqs9xuyqGpRlyRKnBF6240el1l5Odgw9tIAQCiMGc7TSsVbOU4lQZ6nd+49OoV3feopIhq
i36XivIeU+BbMu2elLYnO4HPf+mxbDVuv06GoKuARByy3jZOaBeyLSy+Oyum3PrKPUbh2v0GT68F
LU8FFcRuJ7v4jFbfPc0PYEvL6TbVYFj55v0ytT0Ix4OKZfRfwnNcjqJvklQYeG89ZQPXCnhhit4E
lbnpMwg42M8zMNRvXOt6f+e5VkeHMSKpMyYSmhn3hbuzRfR40xpQ8WH3zHbpxV6mr2BRT7wdZCmX
vg7FrACRksoYyBLvPm98L2wSZX9ViuTH8Qq+IyHwhACUTV7YoBDTUjEn4xCHhCxc9oTOFfC5GtLO
R258pqElU8irbs2Uz5yD71F8TeHl9d53aWCRBpGnqgDXeBzb1gGtdm+YSNUL2UwEGqXGc8feYUM/
O6pJmEw7BTatiNscDRK4D3LSIXW4Nt4uPb+Q8rpuxkE2yId+xXyl6hJ07z6gZB18Iq19NzeFxelE
BjXZVfSvXM37fReR2VYFzOxxAL0HGJ1ANRblqUZ4sH/iWISimXc3wDttMw3PCLg/Ub3NRsVBrT2A
VLL3oShJirCLYvfD5COg1C3hYXmyclC41KWIkr3SRRv/W5J08yA4ozI8PWFu8821ur8mljyyRmrI
/AWXGDI2CnW4s+p9qFSqgKAziHf/v7d+EQMQKqIMVpIV/5JmnOOjqm5V80asUepNOO6z+FWOhmKn
H+X5cO2JkazfT7aHMdSu14RMZxk9+B2UPz7k3UmtNeRZY6trDh67o0xSHEXxQ1kyXzS/CYNWljHc
tHoJb16rwZBIN2zsPQYDju8a3tmA9BmNigKg0JIhtUi9XbieMKmOV9S/476dZx7FvqcVSbes0wMI
apd7JErGefoS6JPiBemIX/DtR7Wq0XfaLxXKrK2Ssk0JGIzaUxeIGk2KJsMIDVslzcK1l9jrsXrX
7+EGlW/9K5xWqLWWOwo9Dl3XqSN2+W8UfAKrdsbE47iHqKdfPwXfbQgoyEfjn0YLwRbk/EOF/wys
nQ6o1BwuLDXOHpmELONs+KQl2J/wcuMMeSLUBI5z5WP6vXNpwUPvzt6o5Cq0qlzfd5696DXCxxTz
w8ATZLfWcl36JgoEINTGQYd8qbIW3LKZ7Q33YFCVQw4hGq+lqmUzwnwYQJzChd3pA6ANde31I9zx
Rrxil/DKEqEqkS2uuZMpLWu5cIUyOH2jvNGSObN+iK4ywjscZmY4KP8NSNQ6hNPDJ4qtY9ETWNsv
jA75dunBGl7p0jlGI03xyxP2Ldj7NbevgZ3OUmaZ2Lm54uP3LBpsUXv929XzLz0yRwdZed1TW4CN
2V/WzNjyq3Cw4P27RnGskUlrpIZqDiow3oYhTMIXcG81hnF2sxDFNS0+vk+UUYjYb3uAFINR39X3
TGDf8N0qBSgi3qNWIW4BesQbjcP+Xyv6KbuINFEvFgicshW1WBXxSl7q5zm98ZKnPOntZjnG0Jhg
8WE11GQ2+ASDS3HO1vbsHEJVkn4blANVmOlltZNoVwdCgS41xG/unhP4uiRVRC2m1vjyB6zFS8Ad
J+ek0AYfgbyqnhJI6I112VbQzjG+Qj32+ykpF6hIkV6xZs/xgoRzhxB3KHn7f+MUVE7+/VFmx45z
p1L67GAGmWASJY+qTvILhI0GLqmac02hI75WR9vbq1OguYqC39OiNTHfiTJPodXWgPJTzKHnGepv
stwzEb5YKI4uCLL8e2niu+qE01DAAYh0EDDQG9R4V03MvRu0N2L/bY9TCeBor0W4phwuAOZQTNeJ
kPFtJmjCc4eCeBsH2RsA6xM3m91Isx7DsG7L0mscBfMM3Kxw2I75o0gBNrwo87A9jNacbUPcU55q
wg2aQqPDgp4gBhgxnr5FHYETFlH/Un30k1f1vYyXjTXJZVDH65L2R3gapNn2Ca35uGWMYpj3hQb6
uHJ3ffkWjf6Y7MkWMQTEGyDZrvApuUwJMN+5fu1TN7hkEHWyFzdQTlMB2IvhKlWhoE2IzQydzTu/
+veiqHWZjnr8hPgS/Y7G6iHrvpMN4W48R4Ytr9NkJdGDym2OwdTWVDJ+Ss7Oq7qcLKRvsJSx7s2Q
kFM/P3TUnQTwToj6KDxl3iXnmcV3EOEyY06X3a0y8rYpKxh2VShcD3jSpEhF2hLcU4wbzruwaKjm
st+Te3dYaFRFaVdxqVyeMbD2AM9vMySy68+av5m5VtvFg2NkIAYzIKK3W2cu3910Plj7GeeL/GjW
Tn/J7+XOxHpK8ocrjsrWi//JDc0J0mWPPYQ88KWdAy+zSeJrwMRPYp0k6+rMIrz+ZTavA46fX9ir
L5uFv3gSYe3/8pTDgwqrrQNvn0HvK3BJ5B1/kLATnM9l1jsDlRYiCOr/F90Y+GfDN+nmsIqBZ1s6
xrOa3PkqEqPVwMHyWy5BUWvOtmxs7MFvKnAIrTDGId4BxKalgZAtNrTnyYrKLYMgnt1hULbkyutE
sriaMjYxUuToduWTle6aAVM4qXDgED7yJLz2Ia3sgaFt/XNBg3rmS+mBSalB/ABjnXQemUkizrac
AqgNz7UGPAzurOqnK1Wk8N3fA+1Hrr7/R3ImKKVhS+yX9xMJ3tBRe2mRz6EFRmopyAijExjXJGCa
+TaYlqMtmP3DiZvaLJRPLS4dyxomOV6OmFyNIya4RRozE6QuY/jsHLDu2DXbLIvSMoCtMpGcYYYH
46vp01XxdL2S4wrw6zVy8oVL0fNGeakDZLqxmMu921Y5DPw6S+O8Nmnn+OUiYi3F4yK6/8zu+ymB
2ayZUUAxYpdCkNeQ3qVauAITCaWI5rLzvLUIlkwqTwttpBXkZkK66Eo6aSCb+P79TvburZjpf4qL
Li6FkE8xmi0fJH4bBkl5mClNJ4rCmDrPdpjqYTHKdidpm10uTWX9z6Mw1hOcpl0i81E4tbbkbtsp
SuNDf03hJUYUoUir/iLFrYwSuLHSVGyABKD9lbliTK/mfbQJIzBw/HkMg3LakEfR7i4OYn1/6XiQ
Qpx5MUR6HwShZFhTBsjIod6ICEzJ0cufm9azvZ5MdUcLu9g2pkhQqr8T7XIfjmznXbwrCXIXSJL0
0QRRin8RfMgymnyp6DbkbuNCHlh8RU+IqfgCO+v9hH8YNxc6H90I71BtD3MjVruaG4+nzTD/hdsC
kmadIjnD8yFljLWzHLw2g54JQA1eax/w+cOxz20yLvvQ0af2G5yZ0Kwb4mIJsWkQTKoBVobdP2H3
2/F2zXLsgzTql6IRq87YfgKcwgqrYmjVE8gWfoyBFikLJ26wD0F9xG4gRx5zxAZuI4yhbv8relVX
hn2D1ld5eNEv3jJjeaUcLlbpSTvL9xizAtIz23TT1EB9i/tjcuIXA6CErkopzS9dl2Udxnsa3ilK
rFqv7oFFca3zIZmVjuS+3x3bhFp34nLcKOdQf0iT1ZJ171ITpWduSoIOmMthCKfurw2ccNRfRfWt
U4Ae7f/VfhBNx+/Nnw7dgQQGK2Jb4i71uuAFSWiklh0ulmzhb8KRrZFYBaIg1/kTuDrrgAJm0PKV
CNPFLO6KbW3ZOO9XEvIkrCsRlSU06xtTYEWrKJbhGKOiq3HxASLTH0Tu45MFCEGjRs1tBVLRq9Po
AmbhOSWsI6SPiFoCd0e1h4WbchZ0cuA8OhJRvQ/1zGd7/VEAG/yeK6yQrCR+VjdkSTPb5vTG39yl
SUEKUSY1yvC5tKoiZIcUJGCH221B7/SPlcyXtUeJjoZ6/l39Oc4xoBTxhW3K57rVuqGYRWfMHugN
IyWdKqiXtqQufQGmZTSyBaV/xzNp81fDA0loOrXbDI1+prBh++A+3WwI8dlDeaQpAxQas1g0YPZt
PuLxStvD8gebyEoNYjugE14bV1ePW1QoNZJFJp1gxu8BXVZIUHUob6iwN0FcUAw7E3cxuoSDvP9P
V5uB9wX0qHQGGymnWo3O6M4Xv4qiayzxO47piQAd2F2gxz355gUzIx0rll6qX5Anz3MIv5cujHPt
guPeJOTijlRfjurUklv3oC0vK1N/WRXHX9aOjDUHepfbclW35k93fcTTqvbfgdh7mGvTlz3q7M7q
BlFSTNcnr8O/YrwWNkYeIoO/eJoVvXza+Cm8zxGbDUOjSTJC8NqpJqUh9saKEv1xWX5q0craSzBu
Vw7pzqqLDzCOVh5P2iXvHkD9pzQr2uOZ836wM2S028rD9A2Fgb0Bc6lXpHk9eVBUr5Y8rRk+Wil2
BFEtipon0BBf3R34nLWEngnD7xeR4U6HtJZL/zf9C8hfkROlsRrxLcKfe0byKO/MP28d3+jjyfOw
q//2DRpgxeJUFDoJGmA0tcwzUuPJO50ooTOvkhAXf+LK6KHKtsgJ2W8nEJ+J4r386AA23lsyVSYk
flKLJ8qhQx6T0mr09KTDbVAAP2bc9Nim2CN0Xg/5Gki459r63EGfFS7pdpKR8ewGjPVwAZEHvr/P
g9y6PwdhJyHAPY7IeFbxMoQeAaOjGRjtEQ9Ro9tfO7tAjfrzmSwFO395j72lnU4yii4vUAU3sTmL
KQuE5uLzStluKJZOsWy8sib4f1GDY1r8RhQVRZSuRZITwf5KGeYXsCoAF1DggrkvUDsOAmacjgP0
WsNj08QoZTAy67YBJoZH7B5wEtxwjweI+NAtJv8UPxfZjI/2dEX2CwFBjlvXMFBFbk+fy2dtGSzt
cygR9Ou2G6PM2sKsYGbOcz/pZgdlh9KGmchRBVA=
`protect end_protected
