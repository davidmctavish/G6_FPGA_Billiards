`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Un7ltTYolB8Jdpc1piMiqB9fjB21NuT52z4yiw/yh43AqN2BcvpsokG2fSNL91M563lXE9uzCsAq
I7BjQLEnyg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XWwowkgAz73aMkoOXpWBzHVDot+mz0DG7FuErhIZAph/JWP21ARe/7Kvhm8tjiC+s/wgMLuC+Sy2
8Q0oMU++rCzzKrJrdDzQv0h8qQXeiQ5msl6vFaKOW+GynXijiu+mW8Cp+n6PiVjcjDBntx/HmbVE
9qBTwUsq2aGG6IMNf+8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j6vNxB4JkqdKS8RrcDH1x4abPaQRb09AemthIR9Lygv2sWLiXpks+tPlgx5gkdGwNdstflq1ohP0
/wXT7qR7aeUBp50eJUaghrlho77TBpOO8f7SH9iX76VHkW3Rnp186gXE7+nP5ZOarzPIDVyw+RPG
S8LN354iZeSaBMc/Ns1s0GI0Die5KmIqIPPj6CorfrPr0+uO5VJnjEZt10iyRGzeVtTnBIY3cVos
LAqdSmcp6XEEE3n8TujPRAiCcIk/FQGw0w5Pr7/6VKnhJpSYeiabA8RxKvSMolMi5sziA5AwyoTi
dlgipu/7lfuYrxy167bGNjqLQlt5SxYFF0IeuA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wiu5GUPsCm86ya6CgVqvvD/1rNqe8ObDlN6xn+25ucL5qYqiRTYWFgABnLsQswJqyS3xR9fTQA26
MeKMPHTF1R6iGJUpAFU/rI/SHumIND1goGmAOanmgTpHZ1Fs5+9/Ele5yewHd57wgC136ucEOyJL
fOY4CBRX69VqCXJ+/Wk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
niiSrzUUQn6rnOgRNOUFnKgRXi2qhBj2P3FfeRenr+sOg4CBPDkVVsuWYDRKClfA9o8XuG5jI900
uWWP+d9QEzt1sJeMW7PDqi+3Sxu/6P+sBsaHylQcBHMeAGwWOjdGjQHqOPtYzU+hsdhyTh9KNjSZ
SSeZ+o7p9Kw8ZDomeRFR+T6wMZLoXiCTBiPCdzha7KA8Cz2P/15ger+Ssu0L0BNYjeFzWZVTYdfP
7iY/AdoE73Sd4/fys278OJTbRmqEQqWwHIgUW2YHzEN9GuUT96yfBT7STFmCLdZem6oTO+uex3mv
nmXvuG9TlegDWW9BAj8xx+Qml+MhALambjNsUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19440)
`protect data_block
KuoGa1AvyDt57v9cR0rcl0OIYxpaUvNFaJeSbTcYhCGQbaPrR2nrxJhSusolYT5BMuFciqDEhfg6
72PsfNNuw0yih11sPo92gR8+hPs64i5Myaxj2XEYWHOIqzDtgxmBiyBDGgiOY6oKYe6qIoH55/dI
DBpoRfFBQnNFLCguVaC/QDmGIknWSScCh/tChLrpdomIibALJnDXzZYfoBO/WNg8bzrwHC33iJKX
WH8GbKjGiXdNKwf7mzrh43a2WZbD8K8x86UEPuyCVTdTeghKUlKiGwXQyGa2CHvHGW/wRAxcBsXC
kA+p4ZRymYkBZ9SyHx08req0ZhDbPsgxw4OY0U2amLem+E0etRTX4t+njd8ojDC3GoGW5qB/eBmn
k9U4fVfKxt8Dv9V/ZTY1NYx2n1CjayWUwyeM6LCBvM3i+M8/7ASQ4nRlngd89R42pXM7xxXvduFJ
+Wv2+QZ1f4cdaZexKK5VYSaEfm6Cayu7yEtjLpYx90J8ahDpLyPRfSqX0dkH0lFGoZBz30uuFfSl
P5pHm81mgOr4lZxFxpu943YUB8Nyx/UAnU7ez2nbLAP09HJxyHJXBZcK+vsSjCRwIqnsvmPZbCvi
bfD9wTLO4Qo8r2/8CybdqQzY9puWMuKc7SoBwrVrkrfzEM2banEyafuGyZVAyvj8zTxYyPiKxSGF
RxzbH2/LBV/AmKF2ykxxJK/bXTE3fn2TJ3ceDV+55/TmCfebVVKHUku5unKf7ClWWWxoCrYQLk7T
26cBqE9Ioc2aiwXB416ilOo6+uZj+uXERYTitVUjMNRlAvtq09fNPAbmAtAFvohZxyzWwUYh21xZ
EpQ5LE/2fzYHElESPJ0QNHE7sLI9gTKgABmmjpX9+eTHvU9lJ8uv8E1WC0pVmjASq/6fN15mhmkB
PxN1qJO4Uv7pDFgcN/RamcLlgicsILlKBUvocPmEFnyt+WtHbB7cUDWwErbEaJMb5j8KVxuTSZNR
C4sYs7r9td+y07pvAmmlk5+kZMyUeYD7UryOFHNMZYm6REILcUP39IzmQGWXx29f87IbeGsdKAJq
ML8I7Zvd/oyFavwvLuQRSSp0GZJgiPGCYDm3Uk1OTt8QPF0DSeQ4hzjK09WjLNpxPuH5axCjm/R0
TMMF21R4AL0ZLV22dR3I5ucSC2Z27OPwytW2hzpC4ntFS331P04a1YbTSf4Xybfjbgys4yMl8X4K
uQ9mF5rHn0z0BJB7IiyeWk7UNmQnm4UVp2U9g9aZFZVq0J74Z8VBGGzEMqV2+oQN0jEV9xQUFKob
CH1jTU3rZ+80Yax4fVwAAk3NjeBnVjfv3mQtedk7qmyue+uJsTb2x6pgLzyp4k7TVpfKDgDo9Q6a
DtS/NZEUQl4J48WKXVgcH8heQZpZCa6KVB1goq0zXNRCBVNvSaUm8xTfp5suStrqjeoU01eeVvsb
dXIR0J1FcmvjMd99yVSqQgacFEmCfk4lehFpX7uRsaktTNKkNrX03/eAJ0zyI8l6bjqQgWJjc/5Y
JCuEEowY7JI6gv8gaWsQRAuQfsBdi7lLcECdJgzxmOTrVeb0ipg1VJrX34QzoK1W571eaMDI4BQV
9HHCNG15u2zBvr2ejqaxbI4jQ3aBkvhfPsFVwpUTy/gfvQMiEtDyzk0zcTnOE0/Gcn4sctkwxrPt
yIwtTX2uU4gcm1zaQboxeLLHoJnW8ExId1QCv+R/rZ03Ddgxs+9LTaN97WyZQSt1YXZyweRiHF8M
o7NYdpjuLNgixuMShP/jDldyXf0sJz4G/5rYVEQDstfBP5V6OPg/hGmJzL9U2vWIA5UtCRfWqY+E
jqDbbLy8lcWJpz+Ex3hp0yUfq4rrAn8xZo6b9+2qFCOH+jnKSrivSr98aHWCrxKuEMTuCylWAkzn
QzRLMMFEc1N+5xaH9XnIlCMXPfuoT2mhwm+J4AgDTPEsvHXNl4EESpgrBHwa+ajoIszXd1Xp192H
d15garBSwsmV5pkFW5N8oOfagCHXDn6qqm85tyyyzXCe6tB3lui6sOfrcCxRZNMlc2LCkzwYtoi7
t8bfolZBLYy277jIEyusbzoHLuk+IQKBK/qnXEtr4K0isIV8eY3HwGVqT/ZsnQKg1PO5uVM+I8AN
xq6VtFjXfZqQ5LMbxSnaA3G4ZRcpw3tZHU37o8maOPcb/lXAmum6MpV06TswUmR+dCQ2FF7//YOt
IWCH068UTS0OoArjrbbZBi7qd1uBOCIC6nDhHAobIa6vRd44I2SNbFAU/CIGCXCoC9mi8tD/w+JD
Cr2ZSUKsvwqxbYo6aX6RdHh2ydTJBCOcgisOfJu7nALWhP0oHCHlZqaiGRlSS1BdFvWJx92ycrcL
yjWa+Qniv2P7DnzwlIg1mcB2CWF3VIIHL+M5Wdv2/v1a/x9kkriyyOCFLggRMQOZ6/bNDA8tQQ6a
rSey8Yn9oMkVhChyw+P4qEnAvsKATRFDMSBaqju1mbq1qwbpc4oSO/u2w0t6RsLUGKfdKQiC55Ea
cOxZ3ZllwS7pMBPjjMGKzq6PZbjcjGvZwmlcJFGDkxAq9mstK0Hhe/zRgv67IBfj7gTejfmZ0mvp
eiByZxj7S8dmmAS4JtydReYPUVJeA/aT+NjKuKHo4uvk9RfTQsxtPY6diNJ1xWJQtJp07MP0pVwm
ZrA8hvJj/PS9nK0s1naoJqfFtNmFDRC6adv67NFmyI53uV6P2DcXHbAKS+Zhs/ZZQfE5usuuuaJP
wHnFUyyCLx9Xls+aWjDySeYCtH42XUDgbVXaFGNmbeAk8GY+Gaj/lyOUQfrskUudpqwcXWY9XVen
H/2tpGGEGU1Nd7MRBRXx8zuJemAICD0Qxvm1cJ2GozwQMtXcsS1ZUAy1OFQDDHrCyMnKLvyaO6nv
ZlqkjrJg2x+bxH0XB0MwRsEkNxuyvkSTQjSvmh7TusA3mYAOz3lnZc8tE/NVvjstsIdA+hB2Yj2b
QQp5urdiShzis9KgeIuKeY/wivn7r8gOusuJClq+El/1NyNNnzAOyjPyseBSzL4esiYNPTwJMePb
b0kSgM1OrwSJSoJPhnym/v7bJpVol3ogPcVeiisedw8Pi507TdpEDnKZXw/3n+hjEQTUQ3szu7kx
Q+Y4yHKrk0ZABEbDhSGyoeqFbNUMGhIaflRrafwFa0owqrg+xw/2Nt55EHtl6dDNpKC9JORgbbQQ
d+MQa9MePEsOonAK96gVpq7fDSJQ7fAJZYNgw4dbkn8gycvGtfXnxts36Tldc2x6PsX/90z+LJNF
OvjB40te1liKtPBh1BP48kFi5lqtNp2GBxfZZHdeUKmViHsfsOu9EgOkACD+1Bte3fo3TfAk/6BU
XApPCchDFMLSovj+u1vH9e8v3YCcuw5NucV062Npb357TnSVOVS/wAb+KY/2H04J7eP4MHON1G0x
h7P1oYnGyf62cq0j1jDqRtcdMN4OAVUQbrlEvDWkF8B4q4dR7t8Giuoi8rUCKSuZpIPU0bClVPyx
HKKTaUOi79YvtlKdhlx7/lQar1sRnUYcFOcUo0GINHvNUi6eQ/SswbC0JKwsNlh2cMKTli1DSHNg
vyr9t6mdqPrG7+KNgfg7m86SiUSIy3+JbaJAAbu+kN3QAhuB6VXbTBFXTL5yFJCJgNv7ASVcEMXV
fMTCmlHLX3qnDiLwMAAfw1TfqxE0HOuvRguX14A9gBIM2cytTloqSZ8qvchucwMEuKoSWSys4N/4
u7n7b3YW11XFj6uyQVEY8LY4H7Zz2sEYkfkOtU5qJE4i5es3onthbvg/u/LtgpEOOHeurN8qv2KU
8v3yjfrUwVRYTuvk7/ghbiBtzM+V9ZklyxSHeaVthooch5Cg7rLevIYPZZce5Njzjpeq0Q6QJax4
ygxIYpXbJcZw5rG7Mf/mVSz8yWd3cJo9v5qdGSv+tFGgOi4uZ2yn5TAaNC54Kq3BlU3hR9R46Zh8
f+WIDve642NA1PiUQDpUGXCO2AoAdWwIrlzb2OUVHxS166bv0PKXyR9sCrVssDKJpwn+jCm6tv22
+TDbtf8qteDuw/Y5D2nQoC+6fNm9J1+6Lky2nCboeIhm/SoRz0INYbLAKy1yvOm0TzQC0xbH/hKT
W8iOrOFlu3HUAvdLGYZ2PZp0wm/WGwQ+BhscE5x7fbez86NLQ4YMVo0LURXXABrlP/4Jny6J+sVT
+4CJ5JVsAQr6T++vaOV5BYH28DnEIiNQRxhnPjxwJBisiiMETA+n+hu4fgtGLzigfU4bhzwb9GUP
JdepRnZZFgErm7koRtBpBFLcboNDU1ub4O6dJQdRVHH283XjCB/nKTFFIB4YRv0BUPRxyG06FMs4
9IsZvlUqGD/JpDpIUz4fxMALeJMjaJucBRPDPTQ72hF/TyyIAaXTth3DqkFTbGjXZmSF2jn7b7DQ
QE3Yfzr7GuTMlC/96Xwj+snQu55Aju+DegMvhZdcDxNCEW9EhqOpGpkUJH1HgQkJOPyIyJNpukWz
cGtYk4vS3r44V+y1SCmK7yKKBpBDXa3U4ExRC8fTin5BjAwf/Hs+OfEtM3i4wbxmWESWpgSNnMwj
nBlI9TcXP+LiEP6SMfCqQ40DzO0IMif8WpW3XU4ViliuNhWts+SYtU+rCkaop8QrceKcCx2gzY1u
lIRRQss7jm7DMIH1q++ooD0aHAePN1xJh9FdMov2SXxSVa9Y47FlZGCoCYT9u8oQfkU9NxS/QJ8Q
EqEaJ5m5Eg4Kj0McrKxM5q0yiAiYoNCov2aSKMICqMW1ZhLJ/EbRAwCNFt1qNjoAmFSAYF8PpSq9
Q/GoOzsRrx8DMvkhTpF9+Mj6YOEimQOOV64pQndiW86PoBZOBtPDO+UO4KDAJp1s+vULkHHXoLdk
gxyEXQZ3To1afQygLi3kXC9xDo9p/X8RANaMIQPE8pMjG+Wa6a0nORHkhn8yGB6omstyKkESfIHS
voSeQ4lgC8dWecPDiUVz2nOXW2apDBiI+EUF4mOPtbrmSDWH7aS3DRDx6ekSHoqtHDsdJcePxFpB
tUSy3UVL+ukL4flRarUpvy7HldTL7FQFEjZgekwed6wpPq+AXBRZj2IlX7ppVuaN29M5QhZj0UUn
XwdTOcF/tm8iDq2ru+QTr/IEw/dA56EkZYYSbPEfCvBAndgz1t8hdQlHTe4OcqFgvOylUnrEvr0r
7WkURalplfTbT22UbmALIpEZWtAV0fP+DL/rttB3WSct0Txjmzc54UOhHrdtxwBNBIBMi+fYn9Tb
w1eTEdEtaucOxDFmLEjMZ3HHFuTUjhcbldvCeE3PRBO+p5Pguh/plPzBzOhL3VR8M1tYLrD/6sKH
/H9aKbeEpfgcjXwvHZsxQaFVDcWEYyIOxCYXje0U2lQlF8ICP3mmuF4idiAW/lHcaS7bbkBUDesx
XfFVtd38EJRULAJUC8dKtLOz4S7+iTUPPgyldKDjJht3ooHBpJgsOFSOQqTFkwAk7wHkVdzHOrvT
77POyC62VzOfdyt6LBM2O9dug5/8aJaC/n2b6YQSOkPL7YcNWtJR7DKb6xCtc5DRCIkfFf+EnXew
0oSFvlDP3t0jWDJ1goX5ukGRESdf9q2DBvJjO8VxuQ3sII6OlIeEWZYKbIsdfd2sUcTiiRWsxO8N
sw+aZy3AczGrMwuV0Z/VycAA4PX0AOHeJ52nouTJ13ZGIpmIIBZiWBYS/vgyvgOCtoDpoz7E/4Cs
Eux5L5t0KLK0lLd7k32Sqv6gb+z0IooIchs+SCPAPrBjIaIyk+BMVGAieXlOwcGwsUGoJvHHMS+Z
5Gqmtc6hEL/3HKMgp1F4rp7WKXLC/Taj9DkLOVmwZZHsokMO+io926uDwVYONEVMEOsFKjYwufdm
orNjHA5SI+i1njvVTmWjjJiGyGLX05r4Q7qmS/e7tY/ZpI4+IC2XizVm3cYrslduc9zbvPmRgJL8
S8EF48/PsDXte4rbNh4/CQwypHegHyQr8l7XH2W2CyL6lc3FU+DJkW2/clwYf3Z2tqTz0j4m5I0z
Kf5BW3GyFIi3TDSxrWuCZFmCHTmGsLVQh+NDmdQ0V3LQAjHyJuY49O2Lw1nasaVqx2stXv7EnPzt
XQq7YtaSWDaWzXlebEuNg0Ae2aSzMWeAg3nBK2CudeS3M2XukdkJBT/wbMmH8NGg1ghbXBH1WnX+
frJoezTXoXFFuQ4dfnVvIvo4kiOJ0O9ELv+s8weD5bR1JFGsQLCUZolGThM72JUvKTUD8SSwYJ5i
gMPSPMt70LoW2BTE5iG975fQaOTXo3WsdRX+g8RCEKllLCsLEbPxr3l+BcpOLLuw8udpfq6iY256
RBD2fy5hqGrCZtVl5NiitqZ5qoZJbvraBaM+5BnBgaUDXOPPMGarsrFPhsfVXIfCG/VpQs1xz+lY
75vIdLjw19rRDOnzOQGbgL4UYGCxHMY49nIqkxXOpSF85lC3GkBs24cwnWP7jTX6HSU3a9IoD3nF
Q6dlwU898i+G6ZrJ4dNnibfVnfeVuHSo8o5Qp78uwoFhtK0i3Ng/g4GlTM5wXoAlJDGHn3407Cyi
kytGaRJAlQRQG9+N4/x2hGRq8YFzubUyWovt8X/hNrbC+pPF5/9Rstw+zfDana2y2HBNV1SBOame
ruYmOUUrxFTQAiIRnqK4dBy2UDmSrnbFXVEuesanr4W5hOGOzOoR1/C2KpKG2G7Z6T7duLnT0qNQ
g601IWIKOGon+c4K/95rV6c16IfNm6EL7nJPKkZrKV75ieNAwKzUC4cFAnvMAVi5Zh0oAJaDoiD6
uuR/aqpIjq0TMtV016IBV+IHHaS3jZ0Yzxabrmp/QiByCM5reZx72R3HJR3epwHCLTy8EWcrVsm5
FobIOPltxW4OwD7ci5wwcm0i1yYN7rkSXAO/aDA276iTU+OpAAxXkClup59XZrDfey3jtRW4vMzl
W7lko8vrKyW4uUJEV3Qem0k3Xkb3SS1dD9MdAbD+KgmlBmyyh5yI2q3fYi9Jh/UyzdoVhVagzD0e
EfUPpNLZRS4oIXX3USShRpTTQMJjWlxQr9K8A/yAMwtCTCpdNEpejogLF0Ibcz9yiur3Ke0l6sLu
3IaMuR7rld0LPk+eFpYgGtOVMWuguup+CkeK87lcAGrpsUoJG7LdytIjpeTBMgwRp59sG8+3reQo
hxR+TmWMUb8yKbY1bGc3ZhzVTNgwYuZK7NvT+aFDJ8tshQ06kGa4UQ9SZ+NL+UWFwW9pj6maZHhR
Y5jfgfZo/feG+rjK2giU49kX9zqR5NVbkZbcfbwDKUSMa/4y1ej/7fjAUkr5kgJte9Vy/ELhNdkq
vN6ZSMEEn0vNLlqY9PacWf8GyguYhQHUgerPdQT6PU38/jwtaUNeF3CPkKF5t2e4FAGeWGaiHV8U
QgN9KwkeU51H+ZuRqX0hTwsHo3Zu4My7QAExw++pxfSwY4ybs3HUsE7LLLyLlT8lItpRLWsKJ6QM
V2iSse/BSkE+s0SGCNf+lQ9RUc1xHhnpp1KQMRHfGg1BqFzsmT9hK0CKIkZNvK8gNT5ok0TQKyjm
D2pIVc8XbrzvL88jqI3UmCMfCUCj0o0z8JpzVP2cO4ntRjyGJr505ctEgmKjHyLP8Cir/qMR3fqd
U7fzQDJnHS1PpVqlx4tdomCL1RyOz8EN6apdA9SEKAv2AJOZkbOWbfMtDBEcE2T/9ty6ZZOOOKA2
zz7Aq5GGkv0h65r8tu/eGy05XNcAf9RpbC2pTSvYHySyOnleEZ5jIQqAvnUqPdvZ6LOlUqlgreCj
u3W/LRfEY90KnZcNqsXwkbv2OMYpTPBQfMtWI7MCXTp+DX154SnPU6wX0uOJ16XCb78EVvsP7rLC
K/c5T3a9O5CE8s2M4ShFSp49E24hR2aFPs1mKR77XMyEdjFPk/e0xQu7Zz/6Qxb86nt0JyNKVFff
X0I/K09nL72w0HI5wkNEWWSQl+K+wBdO5hy8jTNyAkbUqRNB+t9PRp+KHwa/VJVOIhoKE+eO05DI
16DRIIT/TpV7nJViSgq7NhrnB7w4HJ/IE5+0fP60PtYRGgeaV+MGMA4rh+siRIa4lrZoxl25kaCF
/6O3xHaB6Kn12RgnKjRSU0cHygbn3Zyni592JoHkdJb08nxZ7glpYqdNK4US6fGXpKjoxkarCwCA
NjZKqOt+pH349uLUtxC7hRtnzGSf7BBfmZZyMTnzZ3+MAPYUKxbUCOPHLJTTVXbJDvYSmSdXkx/k
Rf87mhJGkszUrNWD6u/hpRJx7070j1fmheLguzB773BBlNnCpTYu+nO64MGoNsUqO3n+hbTl/GDR
XT2m7ibatgze9knKHcsiWAmkBe9b8HUEZdB9yfFc9Wi4x1GPPM+PQ5iYzGS8twIjirqgJE+cRzIM
5knLhuPM+HQpO3NIM7UXCMg27QELmLsSXtvnLF7O6/Fq0odg2U5ZYIMHLXoRMGDA1YM/vcDEDhUW
2Fd2Ym9jrr7N9w1kRsT7B0N5YNZ7uGqpmxLaSAu+A77rUXpxho2yF/iysc9ljXerWg3L4N/S/OH+
RB0XktnYJTjCoTMHNnS3kuPEF1E8JgoYdDbAnydsz/0HCrJxiWTdYclMZETpV+y0Q6WUNIc8sp34
7jJcHGG1G1saEqo1behnyRz/1E1UmVuafWMGHKqi/5CAX0iz2Q5adOvp5uGOtD5/9XkQGbLOVUxc
av1jKPW71XWHdCouaHROhLoufTTM+RvwmYnZ1/PV1c4vPiqH1dmQz7EARB8juUX1hJ+o9CFm60lI
lMHSZ2DpD66/UG05Y6BXosRWYH1DzBRS0ih8D81VBcgyLUi0M17a2PojntNCwkO7Td/ijKP+fZiC
aI1nyi+crOTmaJUKV+G7qfMRUHjXIpMIneLMKpsLOHyseX3Rzf1Udur647m4I/oJ4M6v3qXEamDt
hHg4D/VvQu2mt89K/buZAnrVXZVzJa0QzFVhYaKHd7FL6r+kF4KT6obTieOO4VekRL1pRC+IIjKZ
roaBo6/oPWM23RirSM5LwPubcN1Uv5ESNCpQNNCrYUjHen6hejQt7iI+wKZbWVLV93tVHbZoF4gN
uCSlP62dzzkyK0wLfqyw9v+N+4U+8EqihyGDQpstem1kBMVnDoNuxemiFh8jvGSt6WFXPdumg8HH
K84uVZ/SJIm667qZWamzqjJrDEeXfRZHbF0hF8GjRKSS4SKOQ2IwbyHIrnLzgqlutDKWTFYxx6qU
iz9Lnxsw83CRiJkBNQFfi3DhzjqH1uSjoPjRu2vX/NYKJaB7DtHDjWQeq6VyjNOcDcHnIg9scIdi
tsp7WhG+zTado11f2+RcHr2jPkpaN17TlsBJpDnx5tvETPw3I2uHvk53bz6fxFT11rgauhDFc8X8
YeszDjl80S9OAM9hp6kp1gAZ+Qokl46tkHR+8lpcXF6KAa5b8QlWpEgXyBLSCDmlh7ziR8Khnnq1
bMTjQh9fNoK26yrxiwYOnne4Eb8TF6jLPQslCobsyiBHLhWPobk5jCiXM6klWm3ebSluOZg0MzzR
TKrNmWBtWc0XPL1tagiph8JXeQ01kmyQVBpuAH+pR/IzV8WRzNfr+KHleL6gF7IyWpLSil7cPz98
sXTKy4jSwhzEXM2pliusvx5Mgqjlxr3mnA41QUmAeHMnOtLp/q092Vd8ZSPF1FxFpfqYLXVr6KW9
OE3FoubrmIZ8y8qMcscWXSZGURHNfPwPEkQqcRO776Nu3pl+NdhbNaWYtgTLs2HAQG2SxIe7eQ6A
S+mT2HUdemuaJuaT61bzQR5L623uQtI164lIZG/hZYYtrXuDZqPcAgXY6fq/YZsvo+oI1kMS8KI7
BYWF5+Fr6Ygii5DpKMlrKbyOQ8gQngyWYeSIn7HaiNbY0ZtMIia4didqj8JBR0qtvYPfwBNxquc+
2J8FCRtMr1Ghg5h3V1UJnjtvl5JvcgY+YpuGdG4WK9HV253jd4bFqEUgUjsfD1d0oCtGqBDTodmj
EFr89HWMi3o0PVNqYzdE+MTZbK6HTdF1Ou3sxVaV2tepLT2nSmpzX+/aTfRV5GWV1POVNxyTdxhd
3gqLYz/ikXvuHus+KKR6XFjfWQOowGax5qWAWDC9PYaKXvton3LzKeYtgbzsXP3klBRG0eyS8yvN
Carjv7dA/ZTJ1XByCckuJTGzrWiO6it+fkd++32UgThReIQ2B8wgGAolOGIsFMGv+o7ODEcZoqVU
Xa+J0JmjaHzidTM6OqIZxP6Rl2QfjLWNms3biePNmSFt1yh7oHXbUWygBvEPAJChY63OyGbCvZwE
/RzMBn1tTbO5fvgffkRqv0yKKlQ4DYgYOa/aHuZ807vx1f83dyIYqX5EHNoEcF2EccQg+g1UGkEC
mqt7JlwRdBrX3Ic1DTJjcmtPU0rEp1Wp+Q9VgG4w/LWi9FgdecnFT++izxNOx7TIqPsK4LouVEU4
Y9s3DYq3oSAEMSV/5xRcrGvEppL4FNiNUJYQvERuyAJQfMiU1O2giGlkz/PD4yMdh9VW+JHP6vZy
kj6uHfNFoTTRWA1UXL5XIn3Z/XKQ7xVJx6BNBPXdOv8ZVQe6f/n2qjohaT4vSmjprVgEUyBXEEEo
G4orrkb8rcIxncXprPW2ZYq8uxdYAH2lfOOAhNH3DxBGIsJnpbL7MA+WomAigbkD7PXE4KSHRXrp
hfc3neq+dutOLwxlOA4bHRo48LoHDr2UisgniZfv3D+Ocel+V3thezjKAl0iM/TCMkbd8zNRN+sX
yaqo/jhTktGvd2d/BPObrU4u1M6/PpmFp4sDD3FjdyGA/x5R89iBujbIORwHh89io6YHsAFse1IC
HgXRa6UeHORW5Ot4iCh+KLVbTAcsgCg8kI3tHUhOe7kVyiZT/3k/UQgWWwEinEh5+yh1TyChPIpm
zjTPSiM0X2D3rXy5qlzWHH0tveJLgEsFsr3NDggLcLfnt96ddX3hAMD2qAITHBxkDq3b3IqP2FDh
8KNk2zF9ab2/85rMoss96eJyFx7FiKhPzPhK54dMXcZ9PQfHAi2p6epNGPGWf24tfWKK5zo3iXqv
pzGCGkAtwEqmD6Vse4eXQ3tKe1M3YnG5t4tCskA/cwavyizhvAs1bXaGTsr48gMsyNwNYHid/0NS
pyigbgdp4hKXb3E8/22jSxu9nBB8aDO8hMMe+Xprs/kkbiNBo9OSUeU9KjndiGqguzWb7RBvpQ8a
APMA7cTdm398PJ2Lu7QyI74ueVwobJee/2NrBDsLs3okx+5I86RzfJmQcZp4elAAM5DHhG8b2Up1
KtOLpjDWaaEbVzYM6616u+gRRyBsK/SwK7NAAp/p4JPfoMsBN/qSZsrjz2PM2Agk/Lr50VqKKZys
T2TMm3hC8yHbYhwPr5REpEK0eUqtDuPAXGOfWu8HOQZwJxkLcUUoV+VMUpNKhn/alnXTDETnqhvi
hQg/tv82uvg3B28IGuUcyh3ch2bqx2QYtjsdClvuFBK3nD5bDClsfVS3j5XuSNHUUCLVXeEa2S7U
Uq0Xd5iBRI5CrfBH91WOIo8tfoB7OkY4gVk2YaHSgoYAhctRsGULD6KJdItlyCW0uYXntU4uY0GU
I+mMByjfy3KJ0WYVBvwXqFiDIrKPD7IYZn3Jpm41q2/nUXbV80QqG0PpqeRlJMr6wi/Llh2FbvJV
wz0aLa8ROkBryv/sCbfub42m3K/W++SteiXPo8ZgouVJAlF0HArEM1fEjJxJK5cBEU+WPvm1oebj
euuw+LWL5Q6DbTaO1OrAr9PdqRnCCcdegMVlGYbKvcVbuXna6Kop0iQ2TdRMNUr/D5DKHDaMQcve
90B1d3J9Qtl5pZvQ2+6vIjCF4ItM46g9E7rburj7liXKYU1mV05+yxu9QRP3bUkTuK0QRYRwhAVl
j1GezGuTqrgSD/DTkXJT36j9TidNg/vwMIWmjcirSW31T7FSj1HVE2nzY1QecR73aijbylLiDbYW
VbUYR8IY2w0IWbDB/jhS0B3VhAs9fT4paziSX3vaZYb36lA3nHa+S7lYOe9YaskHe4zmDdzB/6gT
OUalcZg4VMUIkweM91SJIQBrq3hmlBJflBEiCVvbY7Ha0kh7ZVzSrI56melp3rRkkhI0H2KF9zWm
eFuXGmCXA5l8H2CQITjSKuXTue8gST2aRf+XiCGQU5c+Td1vKzWyYenW0xaBN4YtHn3KcCjkjTMo
+toUxjZ1qFJEIliRL0trenediGxAZZXqSBa4f6DNRV8i8K0Ehuo2KASZDtbgOaU1PkX2K31ydOWN
vAwUERXNJbEnIrlddtb1kxHR0GEw42n9wL5K6fnLCdA/5EGa6SEgAvWmyW/HtVlv8ERUBpajP8U+
JNAMiIXPyLCl07P1wpHwsGfX7G30aPZzEOsFvfozJST/sPwUccQicm6l3A+VMVKdoMdWpPHxADPa
IA8Y+nzZQUyUZ6cK6huBhwsFSerBIR8pwlYYLoByxUAQA5zED8lYTCs/CBoPqzEfPGq6Vk14E4Ef
nx2SKJ2kukZKLj8ZiNoGGwWSPkoU0CaqrhN6pW7QBh50JuZVEybgqVpnctbE8DsyabTbBPjsGfo3
NxzzQlGZw37lUA0pDV5lvT2Lfd+i+++hKmXY0O024kdH0gARPuTshY6GQ67GGWPF3ruqF/cGosbe
KF9VCon3xnYs6ovtShgUdiawQaF0FlO+0pWNTSJGzYra/BYXlBjTy70fPSgfv17TR7FLer5Ut46n
5/Q/J65kzNKu0HyNLz/uT7TPmkRW3Ego/R8oB1Vy9ASAgPSVJ5jSYVDuWjevDL+0IzbVJ4/rnGy0
8hRn/a3O/dhcYUzaRVW47uOHJPhRp7gKf0NEUOFvsKsjydV/ooPyJyK3768YtWCkvdCD0stoJX+u
ccdmrq4psf7u6y8Z/QxgB+rGkGvpnPJK61stUQyRAPFggfWmZRlcpAdzy+7vItyNPd0uBa3nX23t
l8p8/iN19qxzPhJKP5rAnE7qXId1cWYo+f74HarDw+of9SfaUtx4BEPd243T1rHFLrGoRGx6QMdd
MaBkLATP4Vd4J0V1QKzH/2aQyQ79u6cbdtwG1fC0JMUL4VL2+7rqQWOyauLqt+f3w7M5lBU8u/Mi
RtXCX7CB0q8wZiekPdt48ERPACACndeA2gFLZgIibPzKg+YO+y0hVbgoSg4XMWF9fIQYguuscdXm
uZ768Y1cwcUT4PSw3izLbIejSaqYar/cNAMbnHHlj9WPEmifgUm8nGCMqAoqcMq4G/t5Kog78bEY
zIS2ZBAkbHMjYRQc1untVy2CyCAkqEiDIkXoSwAOXQf2hSh65Ot2OdvfxU/6dLFuC8UQw28/0Izq
evdAkefI7z/arWj7nLcy6PyqatrClDjVtLMZ9Wwrfi+QBK7FnWc0iyIMzuxNYI4dCewUkg88GkML
gdkVyDvJSR1YC2auKUcHIJMgixKuNCO2SG8PUUyg1mY2FB8CKMv5tbrMxhYqTToLHDNk/simgtvB
qFBgqnRnjThDUAFl9mQt9w3sRKIo2qS2XhcLX+2Q0n+voE4wjGXOejIw60zTL/jD+dz1x8SFkXJn
DW/vqHfLyiHHd9VypqQOoj81w+nDdsWZEwtMNchMSdoHRrVd9BOzLB/HkREG5kJUpN0+7RgE6KZc
IAcCFanuR6SJXL3TeIiz/dcyjYQTmy59qSMHMll/LKjyUDBGjrnLpBPrtvyAqeTfUsqcOEmz5Xg2
Md1IdS+0vpbXUkdP43l++shJfcr0U+Bpulyww4RFEjlc6jJj69ZzhVdGDDlqjGdE1I1sHx+7suwh
0DU2Yc0BbSnpOnPPqHSkCpuFi+yqm1FjvXacNGFJNqlev2Bg8GjE1AchaTcg0laTzpJrI0UqilH/
T+Tronm96FoOkTTTkn1uVfSHtnAzbusx35ar9YnxeS/Z3hQke6yW7ASd5fhdmNx2yXY2c25V4AI9
t454tLgLV+SC/0BVxqFjwZ5WFZwWAPhFcjlcl3mkR/ow745PlPRredPUzPRzJQpVIUuimJGVF+5n
oMe5ZDxPkmj+M9tUEJ6F2BVnVaqZvZ9F8Jr7KL3DStLX/uqL18uOVlp01H4HaFiLZ4rw1vAij+Yw
wCpPYMgfsDz+Xsn6d+9Pxdqufj57LzKz3s1BmZ+ULlM8817+rKLWGjgcvZ5bjCJsqGgIe84S5bZT
YYSPEBF1h8H/+RWqDM8R3yOdbz5j/KpBmb/8H/MwPC6icHO2XmbZJULWuyGHZ6g3qBbDzT58jTDC
2LDtMH4Mm1f3GEbPtD4M/WNMjORY6fMMutZorOsTofKxshDccC9wcJ2qjIOop9iB35VGmAw3sXxr
zrTyYzXioPdlJNBxV6wmKGi2dG4eNv+KWIuiCfUipueMHBEm4VaOI5435Oa+nM0n8530+NpSNI01
jZ8H3u64uuJQE6zKeOJVpLMJW/R913HH4O7/IEgatshE0aoLgaKn9XkheoIKFgKWk4FpWmFnQCQ9
L0OyxBfB/FLo3eyBEOBNfnk4UPOxAQVl5PMfH3mvilF1FFbG+ANZtkhM/0ILCrXc0n1H6X3OMxv2
jnp1QP4iSTSPKBMRLW2/aoH31ul3w3OBjwvFazflKZR7Vii2pg/VxzAo0FtjSxR0VII4+UqLgTzN
SvtiBoYeBJI5jOYFUsBF0cwdFEOhANXcdVBs4cJcKOE4cHLaQwPLgbV+4HfPzYST9jSMsitGsPch
glqUwNdQyAt+rNBI7Zz8lc4mCrKUeRIqnc9uA+WDRay31XsRzfb+SiIxSq3h3coiNUqEutqA8Koj
KsYQLDmGrTwssK3Q1Tg5h+AZybSv9tdRKJ2P+TSdZH19tE9x7w4K7SWcwhUTYA/oXYXBjk8YoI1+
N12ZltpJCCI4nlbO55t58RqFPofulgftl2eLMSEsT2qkJWFa7HANtjNtpuDzBo+xA9K/+HL0dboL
jo3/tyjYkT/3HaxXcvPOUeYuphNyrUZ4vGBmwR419fVfcBzKBgjJvj9IkJWvz/UpA81q6BTEkEC3
O96rKPNzIX1ajuCgT9brCd/p8Bl+Efege9MqFpt3lN7i90ARy2InBuwNjIUvmPisUf1GlAKB177a
oWVaKL7TCngxTyG5WeatbXePBR4wKmWNRHyZr5e5s45y75AOQBCHk0TPpSKIOMimf9Blo924ZTY8
btd+6V3Qcnr+LhLTreXeM405d3i1d+iQwjMH2JKkXU/rXOVFpA1gr4yQPBhGHNpBmHBK/1ouZgMY
SvEZOFORPb5yp9ul6wugYsowcZaDPrvvCGFPKEZyMVVLkzHTTk4GVvr1NM0RK11c2fSX3KdFeJqG
UyT/elrhSPlMf5DylXFXKmy62RgYx7p6l5FYVr1kMfuFwoOjBTb6Raeq0/hSltqTu2Qp+lMFcC6N
A2K9tBAi5t+/vLjW6Yh1dLtpJY0aLmqgb/Xa+r9vFvbLo8GtqIYzYfeBn6WXVZsjWnTIMPvqhlom
DPfH8Ao684FAeBk6CbJvnZLJBpmmJ0TzccJ2XRHMm7e7+jgOror4i+UzCPh8a+bB9YquWEptLgoL
DB4e62DVjtiLtXUKd6XOzODCCrl8pAUUAK2DEiCurRtle6m7WirgRZvdlpkaeZMv6Jf4YoQxQ28g
AxAi40t1o2Y/LcAfbdWyBQ53NkVsWUf508DRycEo6d/BSFwx7l77uAcDo6VhuvGEHqSG2qzuVcb6
/9hbKVtE3UFJ4bdGMmM7OoRcAfo4gtYBNlniAN6yWe6Aj0WhVzUTVMAV8lfHw5jt0OUWz/DKSHfB
kqjUtUKH0Q2Oj2j2cLZUx6To4eyZYE4l5dVonK2ikcCMg3gEKi30PJmb3h3n0oRgOLiG73AH1Iqd
x9MrnuCBBii57/hGdVwhiBsYF0RwTf58ZmRyQxksXK3oPGqKX0CyUirDgwpCF67seoTPajA55Fzk
bnx/+FPakaIflmCc3yZszxxFZMhHCtW9eDe9jfsLoywXS+7Q0nbPnswwsP443KHDrk2qjJrB1iBr
ifn1iS/kXUp7BTmpmwc+Cs6z4aHJyNHyNMbk1HLBwGAshaoBuTtkkbu0n9yIO0JgichFgTLA4H89
VqeF8iPl5TxrGqHv3Cnkf9Hu8K7lHlZdHj+Qi9X2iCt7aU3VEN0bNGWqr6o5LrbtIdjs6TJkTBpw
55aygyh7DS/jSRQszDrNXxzct2zVvxOuA0o2H2ib7w804UP1PsR68JrdTUpg9qUGr/wp/eUQpEdi
7SM1cLHcZ0J3jSywHjTdq4DZw+vHb/hhNr+aEFHO1IZHuu82hQfT1l5q2u/l2k5K7FYnM/pUuJjD
NE02scgz0vAXJZuFprbvEdiZYBR8A6udWpMmFFEmNoIdoEdt2Fd8ypiqrp0guA5o7MZIBSKkCemx
2uEYTYp5zNw7sbGsEd2zfD/7M8wPzI+OyYiGym3TK8t4nXAyGUTn4+5FbZVPqnGmYHKKpgPKMdah
03Aurg4HaArFZkOc4ACJJhAa5mJkCYbQGmMGsizXcGPMq4j78JqJ3ypCdWd+5DMkYU27LbUPCAjv
pc8iH0gaJB68PB123XorLu3gAizPZBqt29ZCSRz4EaqlPeKqmLBCWxONgZtCm1CaxAdCv0BzDo3G
/yOaG/vbPexw+FP1btbl5XbdpnW7+SAacWKwLzVZFkRChP6r9J+IeP+YoAXi0b4uO2mhGl5k9Pas
vMR6C3RQD+Ew3Pj3Ioe2aSo732dwucR51sn5xiFAMwLqf5U2dmhSzRBgbJmIiIRbr3yqmIl93Va3
Fyu05smfTDPlm1WnhDc+f56izD/dvKyA17XL4zQywUsiVfpCUbolJLxTZc+b4Ate9oPp8xkDdchc
OyDuWp3M5pZFP/qhnLnsC+pPv2oSDjIvIgEdqwpqFPoVVlSbJtnicapr3ZH+E5V9CUMj4uU7v4Qm
vkXitjUBqAE8mkTEBVxzBdhwEPjr8XsZTYMRaQM9Ee4uj7ONTLiYK6h/eVfQ0azC1JbhflOdBkCQ
NgImoZx2+cfwbMxOo4YW66WHcPbTZ6kK7msiQniXVDswlbDlfL2jfLiBJFWAltR5AFObVAXbUw4u
H0dwHAD8BZO+oyjxfo3+Xu2xJB830TVdoe11A4tzKM5h46Bhr455lKZZhKfP8E88o2jQLggsun72
Xz3Y6COkFHhSrZyjasrjhqFyZHCIvs6JYbVdGPVeBhCQPJryN8fCUPn1/Eu11u3BOWHE90zrDk70
qZzDIcF5LiqqEaJtzBr9vMk/g7JSQcr/yNLfqXGqn489WJPJHTyxOckeW6ji1bCAJEWDPutpVUOC
unlkD79jmSnCCrVX29enCAeub7Jbvz9cB274uIUsSleqEvXQcWE/gMTYUf/se0CDuBwVWMECw1NA
dYJQGPe9gszucRbMSHRqP/Z8sX2iwkEjBRF+2yKn7wtq1EBee4xb0bs7239YwYsuF/QIQM88rKUZ
SMiNQQJmJrLZRo1+R6SMfQDy1Tcsx/NSoHeM8OjwW1I4HkUKQsI3/uywi8KmYcOvxYU2Up3De0Zf
BbwT7vOym01ETf3uddyfmIZ64mPak+j+/lAdkXLuvtZ4cUoZrrIRBKiUUkKFj4aXEfzPZojJvUj8
0Hfq+imfSCNMogjetxWlihonSsQZrehFCoFavZX5O2Jk9/MLmxQ/Gb3v9IIHhQbUc1Ek4UhXDJXC
osJcgL0qYPzNKR5m3xPLdiQ6rVLgpXWu7JG0s1oinLrjbOXG2SnjZXQOoQ9WCOhB6SgkLt1CGFIt
8dJUzHtiTwjXg45EgvRy0a9zkcWBQgpgMr0rU94kWnZxo+2kXBzF6F9juVylKzrzO7qTge9HLEwI
dpwZko9BklGyo2T1SxDkv75whXBWFu3rlOdmdDvtvot8erHqL14jeotgJXnVskOV7PehSUZ4dzC5
GoNAFwoWkEyPvNg3BUg0Vo5mOXE0g/PJPhLNjdazXC2atuPJFwrEcBSBfAlkdNjNWSTpawizdwSQ
Q7MVK8n80wg2n3ECPnFBsn+dDqWG0WGlr0wEGHqTu2DEL2knX3TDfl7fgG2K5P7jnIgM3sYvDYo6
ulkhonXIc94pJkoquDrk5ArxfmaLWbU7KSaEArk5b+hBDsuR1TkG6aFqzmime/ItA/0pSptWmq8s
DRoowP5F2car9g3d+XJPQ1jaic8LEvlHKeEMg/yV/kcWW0vAKWmLyzb2gUStcmU1+TTppQppr8jU
8k/NlAtORsPqmtqDWlr5z0PjoNbnNbc5M+8f20nidxPdDF1zNJPET4D750ugR2++EZGKHGptL3w8
ctO9YyxTpZ5guqkwBc/arC6ZuL4D4bg+Y+24+kTm3P3moHxSdf2w1BzIJ8KP+DcuQHHoIYyM4AMY
PeZN0lwyf9ei8JC9aWh/MsPWmXViThJxAQbpbeWjBi6SaDct2m0AucxR60C7+PmczfehaKtchJOv
fu6zgyTNFyFjOz0GBKGERDqhDsErxhJhFQeMgmdHY4yccRvgLkot8ZMbRZ2yLo3TsPLOEtuKYpVl
my3AEBELCwpEn0JWpR8LxV/wedNrOfXazO3/KMIswMAnKs7eH3RyayLuVtaDadi/xnkAnNc2lYwx
oqqLAL0QEYT67rxU/rdyGjwiO65iCyL9uyaJfaNaNGlH601VScCV6Zx2EHZjZ1tSyhVgAH6hwu1c
VQRjaBckaC6+5aHSsKjxg1KlQ85mwdRMLdFp/S135G1JNQePMRBkeP+cKuMpCADg8722a+mZty26
Kg/CGhZ8GWBUrsA9mea1OJaRQBoc0JQPNkdFG5kLUYh13s4PWSoXcPvQIpi0pUi2sS8anfiZz30i
2ZMTK2uHbdmbbWHoJTyRVZuCItsa9YDmzrqHiWuplKsBZdZRKuUG/7GEMy51HeC1gHHbk+RzL+2G
Jw7eFJFYia30l3movTr4EAn6RwUGVcv5rd+O5kL7Tmy6yKkrkiqgC33FjDkNBo/ialSrRx7i77pr
rRyZtVNYIvvsTC4lMdZjcuyU1NpctuAQDlxUIF4Jf1lc/SEKOyUiBnnBQ4w/NL1h+ClV6faeRpYl
IXXN4yYnge8wA/PsPG1DSJIyi0SuN+1x8Kxf+h+UUYton1iNSoPLb00NRvVvDPPmg++lxMqGW4J0
hfh+KW4wagh+gjfWmWB48ffmpqBbrRozXmP87Yp8+lAiXGT77u27i6LnWfifyvmmcJrsSC3bJfld
kqO+t0dSjAYyVFMfj99ej9zCY/nTfDxUeXO4kR/yS22AjA/W5/QYdXfvgmvB6fXdjYv4uFK+Uk+u
vIKVV00jahjAmfvQ0R5ijOEY0cnYug7J7cTanLtqdQP+Ue1PPpV1zEH0c0rMW4pYk836VJN8vQ0n
rOIHZEL5sMksbOEEmf97aY9j89/9YpdZg4VAMldbDhlrjTzINJFsdakSGeE4xcseRpvPDKKrHwWv
k2fOUYP4lVGYWmKHaB0cml68IHsZO8HT8D/8l0SViYfzUtlWhZhAjv/wFNd7ntWKgNkQetbIDrNI
KbYc0AACbrlxLyNeabnqd3tB26wZRtyLi5DxamzuL6aQUTOrCHdHVeId/nWRu1s82v1QkzAo+c3n
ndZKUaaQ5b8qIfyD3aFfa7l7doT6I3OEQDPMYxjaVSTed+rwIFvUy6Eta2yzJcfeD5rt9vwIIByi
f/pTng8OFmP/tuNFkAXSDasSfwJppr2bxpVVdpjTMChG8iHEZO8OpEn97xNRJ8Gfd6Eem21lYy7t
BXaDI9dtYIj1mYJr2mIpz1MNlLNeLC4Y/DGckSr4w76kMrqEOsiiJNOn3VmP50B1ow09XkPIde6I
VN1WtrQ2la4UCwT7UWj/VH3BB6BI/KoekkYc3ervSNOc3Sl7vVFjZn57BTreEqD+Z3/thN+iYnw/
rpOdipLeEzTDL74tXbmREeT7rOxJJQeaT1LGAYYpQIdPXLJZjJFwAYbcOTTOlyzlmP6dtWL8Dt55
099crpI24v8r79f6nz6xXvuKXeLA6Tufa7mWMDJfGt5vZRA7njhHG5v9RwF+jxcuJ6xyzkqEmdqt
q6wssbHTZR0fMLoETZqKcpa8hpAdXbw84tbjvYWjGoeD2UDaFHq0BPMntylKqfTRoKiWxMs8wkf3
BHp+6PmqlkrLHAubF7hS6aX1TgE5nbqnwilVj1tyM1sqAPiTO6dUHGqBuS4ACr1TTPwfmIQiNW68
8yIePWyNo5azzt4LOsGLOVEWdO1yIx0zhOXYVqPJ8RtbtjL7FP3CfHdvirH1PdvXS0e0RmvIKIG7
htHlyQ20jGkURJwqa2Jerg9CbZyw1ue6VeNw5Gz/ckMFTYba1xtgH73iKq6qf0V0ihYCHkuvLRCK
jYH55LxpGPECp79aYGsStfBXFZhIcaov8WYr65KN4vD3rt2QPR0neQ2gOaYWoF3Z1ohX69VBXK6L
1jD8sYpzY3TUQjCe/kEh1e9AqAmzAPwugdS7tjCygW9kIvmL6f1NZMLV+JGQ59AMeiRe6nDyMvdC
nvjEuMePHTq86u0fUAD7S2SEvWh7j2iUSA5F5YA9AF2Fo53hcopHZFOBBabmBkuHO9CxnC9W6h1Y
uPhsslpdV3ftDChfjx9RPbetq72vttrFIdT7TwVi/iRQ5HFXkSReBxkq0fDB6zK+ZWPSKPznxTYs
X8J9Twta+5VmcMlMb5h6DcsIDVsx4dzOsGiexxcw2DTfDVnrDAu62bZ82/uTA5E7pmWtelLLYNlJ
sGd1z7qO4XSDqHZqg/dosszWBYHG7MbymKYCqZKoRDilcXsau5OUNm1zpYUZIP30A16c4V9ZoUbG
a7NgKlfDIxoQfGRNlnn9fd3SQI8DxGnnzoNTA1ijhl+/FoB8FwixbzZrSKiXc7s1g2XEHDNbyevK
2mBWDIAiqo1RN3GvcveDwc5ZBta4RyCMF0ELk30cHG3/Xk4i3BazvK4ZAyRWVPD5d8cjjC2NfDMW
k+fb3xI/V3NLNKUtp/rtbjlCAgssR7FsTzpv3T0uFRy5dGaYcYnFITkC78J5pM3JPBnnxEzPJ8c5
pHXNYsuwxch6yZMukfwSK3QFuQakNPGsDl8gI6vRwyLBqcoeN+DjZPmoKVIdMDs9wBOaVOEwkmEj
wpgtmRWh+Ld1Erby11+aHA7GRd/3D1Nl4Jcwz5lvGleyK0xPP3cSLh75BTXwImfwogTdMrM1bzXM
Rq9NX4WYFNtATZj2pwL99o0tks1DX6AqgRMdHBfS3kHDDzG5AWupaiWVNSppISr6HoPdEmpEpSgT
k3bxFsSWArvq+zUFyvPRTm3PVZRs9QauHC/l7KAZj6wfPt642rae2CBRCm3ZbjW8IsmktB1o4HVB
cvKMqNkR4/az2e1SubPXAOvYKLvXXO1Dzcux0VMpHZiWej+xmHRpJXYNMhWC3FsQLmwgklQMEoz1
6fsYkS71lMXaILIYVcpUMNU2LCblyV+nvC9zMHaTL01DwIdaLdkO4oVfNQ8WQ+VM9uldDieN24gH
CZ9kXZfSjfsnoPUfZ1T2UDU3u7LOsTdcYvxv4+0fvwJ8hriCKTr9xnWWtewvqnq1xfEFs4AoLVwx
A9EFnydG3vRW33FlvFiN1csDNqRIV4EtaUfFJ/egwU2cU3hEfb6dnBchILdEzZ2nINM5v3hw8ZEd
UzKV87bwQ8h2yzum3UJqUPhDZ4MpJVkDFXZ6+VykRQf87tm4W5RqG56X+kpnmxhctcY5suPiwogy
G5dobur0Xj8D1M7ZC4/u8rq+ZxZ6NDHu0uMP5Wsk+JDq8QTAs+7t2Zf8/XEUJhRjRXCZy41zPPX3
J10Ax0Z9RzAO0XQk9A/TohiB/73ukh3LhYS1vZIsV2y4bBhCh9zSCsahNGzYd1v1QgRQskVUb3B4
3fo+ZR06koEhfBL9LVpWX+sMNixO0lU3L2Ae0asUVr7dS5+u5R4gGAl3FfIRKNCIv5HgmUCwRqh0
u1ewsyHGLzYNXau2/JsxKyTnZn35zPZ3b7EUxCjaLSXqgy1itNCTxDLY8tIMOQjaBDKRz4Bn7T/s
mYdvWadbuQmvXCItbdY+COc5iGrIek11BOgiPP6U79Rdo0v/6FPJUAI03E4NtBYwCzD443SHGZLW
wlFc8JavqbQ6laIofnTJJlJbcDgkCByMh8EjzQ/R92Rp9+wSNSYQDY6L2QT3s7rTeDZZWXVOM9OK
qkYy4Fpfn7BcSkWfcAhomrVZrNl2SxlHysnJTh4brxhz8uUPbv4TSNhDCMQRLnKGabypURehMn1m
zgn+OtXCV7vkAAxSgmKXCdZ+veUTTp4xSb5tYOaeF8dOynosTBO85VReer91zm6bRIn+APpRWXoh
w8jHpUXm2FcuG97fl4GoMS+m7jm3vtOcv5zg/G6sRJLqQ59PC/SQr4tlulLSP99PPno0TeEEbzNO
jQvszgQATzggEJtabAXEI1h6jf/QHEvalcD2OoWrKXdM9EKU1brnefPZc/RK9qikj3rFC1PlH6LW
alE1v0BGQg7KWiyQA3SY9iFtBWGcuCNJYnHChmdwMv/yN1tIanW7SbkNrc9CmxxmBkUfC9vwlb40
vlW+3gkG4iZaQqiRmnzm5GZ2Rv5hZWfepctpeB1IKr5X3fT59IJGTwxJ6t6Ca1YcOncvExcKpN2B
VSqVxzNCE2P35w1JnlhndBDntwF0ssqfpCb800gQ2pEH61YMGE3g70NWySNoop1LCAl7EdRxju1q
7WViY7AIQ5MVd4EasiOzFBe5DZIwQ7eltV25K7UdwC+GjYycISJHaM0kBycq8zCy/f8D6IZ1L9Bw
CI76Ul5VPmsSGzOps/gUf59qSMI7dD4U1UJmHjmbWEnu/sPn9O2LqgRvirsjbUC7WgAp8AcM5Xj7
gOfDScdZNs0oaQ2JTHE+i90JHQVTJQS6PMrfn35wxGp1m1+IzVukdBZUCtA3gjQhn/Q/L1JDLwA+
VNSyvOs1UYAYEmdReZSCW9/F7PzN6hB7CXvBhvSiq6PH+qVAmNUVo1g/gSRtc62PI7I8bCvX7K2O
4StXI/ZebMhyakp+IR7N4Rf9uAN9IRXEA37I442n/xlvZXjpx0suCUZi5XUhx22UIzuA444s6P2N
FOpHrw656waxSXvBQhl8RErI5NJFbRfELH0iQ+H0vfK9GRli9ta1G47k6caPylJPK8wAanVJq3F5
RkjXrDvFdErSpYtQHECzUxPN6Oq4wMan/0aM4mvqjWWMckbRwcaPsTU6iAA7cTpmKtQ4G6H0GdMC
1aNSVJaFx7ZVrPOXi1AGHLfsqsogFuThZC73fJVyoM3v1RzkrzoKJ5Fxl9Hbhx77jxpXrvk9vjS7
fo1EFKsEkwOGIv3gptZaokCY07/qFOjqha2PirTgYeCEL4b9Uwgw2bwYEG8qfXLLdTjjgMd+PLIt
PSolUVGZA3mQF1RjrVwsVLm7j+i+lVArQoCWUVUi4PocoxtC6k3HpqvSy1hCwMEd/M3oeslWJt1A
7zJx5uGgq7fnTlYKbN4tD5YLxro4XT6yRIFH40sJxdBbHx1ezLaW2YDBh85o+FNMfj+fcLPcTpq/
EBHT53LJZAmq50LttYGpXiE/73U7zNV0BnfvT3lCzxrYvYXg/DfnOoadXVzLIR0xi27/30vVzsTc
hIATS8CcfPylK/c0h20hPqRtpPpK3w30cHzK6FSQqLeER6jLDnU1ycY0zOgayVfujB8hGuzGWA3d
8W/Dt6wxi1h+vXfPvfEjzwxtoUGThpjVK1yYwRXqzJN/DktcZCI+jmel8fsXwMNjD1FqA8JzhK/R
p3RfCymxGG8mIXJFNTZaiwljiRjIQ6X1NMmUNLr6ha9Xp8+ZRFDiAu4+LTOWv2r19e3xan4cREkm
ODOPtWVUX8/scODNl0fA2uYXYPyLUzhjkIO/4iZQXyaFh8TWn3nL51txL8FyNVVx8iFp4G9Wb7ZR
2EwU6qOlRKAK+5flFKeAqm4TacE3zQIk7T5spflrdNdL1sG2nPF7OKdcdd6etHMmKoE43ny8+ov/
OPJfiECQVOwomNc2LTwbOsqvH3pEk8GvhFw+vdm13Sle3pRUMiNquXh4WHOV5DwWhy0z+ZuCysRQ
xxnN54Ql4MKN5RXn4wC+hwVdWOVRE1D3qUWW8IUig0WOtIUJlirbc1IBYy/Tapipd4MFmkRd2HEg
rzerYObM+4dFtryp11A92i5UE2HdOv0xMdRQLXAU4KkEYdvFNfyPwF1dJM4fcMczrWtJtgUWcaBi
mJH2x9BbMsp/RQhr7ZYvAOkF4AkXcQCroIkQzF7HOg80d7GjTjPC+dpLXJOTPnzcfgjbhjraLrWU
kA72yJKGkE+TCYgrTcTDmNjbv6Hi9TxyRuhDTJdQjeVmo+4cGyeNStspl5F8C9Mb3Mn+WXrmGAJ4
K46L6IMNqiNrzdtJPhdAhhXX0xPqxUH6JtBgqZHUwMgB2htbUnwXCByDixTvnSlapgBhZqDfTEol
CBmgzZeerTodxnAmvcriRcXOfEvpLUNAp+zuEGV7RHwWTpZSJLwuw/JyPCcZcTeO62a6NFUrmdkk
j3A4GhDj2qxREicxAm9i1OKmo2gCWpVBz0VkobMFNbAXuzyx7lURL9zsseh73MtXYT4CxvHBufo/
rRa0Pn/XpbBPm4G1PpUanOMyo3MP0QSX7I9yfbS++8bjGx8QzHT6OtUeiTvQtxIkbpQrksb3/Vg1
yaWCXKkv+W/dQZMZ8b2yxA+HLr5KAuUAXYc9VEqyWBnJpnLwk0Fum0g0NeKznxeNPWy+UKc5hVN7
LC0k7EoHsQaHRqi4WSU710ycKai7kUMstkaGojZ1BPD2yyA4fncNwsht5RuC7YJOc4ce2ls9aFP1
0uWBC2Fwznr52U7wVRmC1KOjzCfxteJo9qcQcnWJhlOYecvPn6feEMNhX9mgJRF/+cINq/Ghe7AQ
gna0R+PR/tpYC3aucRoQELmhWLFKv8MXA3DrL51+9nnDz5XRjdjf5/3n0+Bnq6aeQCTC47D2Glxv
4qVN9VQGg5WDXgc/O4kG9E4+X7/4GJhgeOx7WQki/iuRLRR12z3IIkCv474FNGAjVCaY+E7T7aQZ
VY2AHHjAm46sMjt7s1CR0RZh1LqbGJLIeQ+UwlA/maU/y8PWVk583cteax9cSLPJcJ23W84WutC0
E9IiQ1u21HYOs/y1uzprFEImpcTIyFzCSR7KB07kciEFUNoklUjcTpNquj+TZZir8QXSy89Tzda3
LBE5+RyPgMTtMYU/txWviykC731VmZxCqEqZhMkBVPZaKmPKdBxQzsOuG5tBXy2by/1meRSbAcoa
DZv66FMr9nIQa60C8G26dfwk/24L5B0oiARnvfv/1c+sqjIOYPIDxV3Z8yNg3cHussqpFCxbmeD6
R3I+smsjvEBK3YoPlx92Wi8DDeiaQXKkJmw8GT1BaErl7WFjf6Hnl7hMmiugmXBwd+nzjj6gj5fs
gwNPMH4IWZ7aA0Av8aWfWJ9wB9vX0xOSMC81km2z4uNqg0fWSoCFkpTV75QDVL3TgporUKtFXXGn
cF4ETbbarv7hQQKkvOKF6zCKHYiGmaFJbuB2y/gOfFXjdpqkjFbHL3GsJixEEAB5RDhSPgNR+tOi
J2PSa5IQ8NLXHXmEaQhMHSLBQEpDs7ToSw5O8eW4MrCFl2SVWGDFNaOGAqFB/OFrIaU75EObAkkP
/c5A01cDjlY8JXngzNXRDSEithGJEiXvyJfAcaRGQiHKZym1/6uuRwx01CKb5PhNryxtM4qgGr1k
d2og6FXY34TV8rDNGnLKuBbK1q6sAqe/1OIKONupOnYW8wFS0KP2YJGShgZHBYUZwla8p2zAl9h2
viCuAUnQs2kN67KHg3QNix9W/Dr7p1ZcPcTenSN4Nu7ubsyFZGOdXmX8bE9Q1wpuGgQRP+nNDrRn
IvisF3+csik4w1L/efUWQcRSPu+i/BSQjiUn71H3Q0YbTYtBB4HHdTQ2unaGDAtDES85BxZfzwm4
N6wI
`protect end_protected
