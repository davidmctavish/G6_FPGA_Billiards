`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FKDT+ocEOnXfz9klY+zJEgZZySw6ckSFdXs12C2iTIDLc0xq9mJuWLGQcHQF+FuP+e4PuVWNRdbc
De7MiQTkaw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JB+vP1M2n1HPUp54AJ51dEeEfzN6d8Rl12nao5OOV57kMZzidmoZdOcivg0oiYNFri844tYYe9RF
wIQ2PN25pl5XcWJWMYt98OowShtfHwUKq/Hd9lYlQkPV98dYuB4MzVUiBnvdvPyXOcPzccsKbl25
gkJBs0n55VEATsAv+FA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sVSG20XoQPYSqhpTWkGyxfStqficsjrB33v+rasb3UDbIBprr7UIYNKCfHPb4vgLl0V6LE6p1hwk
Nr4oXVhjyEDXP6ihCsqdDbcSWuM1ix8WCofb0muLmPBeiC67JKuM+vPD0YAhAqt3VfqrvNsGGrm6
r6hjP+9N5/a7EmCKbrcOR58tsiITemaGx7DeZSiEgSDlnE8s16jh3YBeRmdkrCXu8XL/2pAAZQyh
CvdVftmEXkgziToFBQrNuKOaHC8UQ6ej21guVs8unNOkRvM2z9qYBkCJCqhOuKP5Af+kLOetl60h
837jS5yB/mdV9fsxcdBKCr14dyEO6Yly6IyI7g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KsOF4o8LshVzzZmK/h0pVmJBJ+bqDWufyWN/tStzrbU9iUFXkJqaS0lsvbiwYFfNJCVAmtCiC1Mo
IHW35kb5N0Rsvf+a0HaYZZSZWxzzcmwpxStFpJGhKudtxJdqZ69vflFflvEzgmEJv10raRXDTIpC
M1ve6ugr1SltnemF6Uw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OmorJ0rQ1RYDmFtHk4mVm3oNblQQxYVIdu87RUjKtaKVDBEKpK812nwutt8yCPl9+XTYt3n9cfNT
U3r/+5fzyZbZPRQsq7GJ1wzxIyiNDiB+X/U/Ta2YmW1K/dhz8sAt3z5Fw4mkeVF0NtbbCW46miUC
pCDHaRpHzf7KMdDWzX7sp+Riond+bZOrOOYgm2Ox3yGpBFSYZJvMzwwAn5yoGoGKh/wD/Jl7XdMF
yaB7SAk8tcuaYsXSFqFpPYJlKDB3tpe+yTHmgZfkPveKvM5oWtJhvOHFggo+8fnKv7nT4pUGnfPP
0+QVSD0dU0HKiByRmFEoTnXVuipj5+1H5qNn7A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34496)
`protect data_block
THvaMDtxxHD6n5pOYf6clS9hHtAAw95hnghs4CcYtju2cs7H8Dms9KmCUltlwJFPFGNfcXbfNV4h
D8052MCxBsrfCtPmk8JS40xSRtZeRiCtHDA1MvzY7fBTG3rg4vGFVnCIP3akwE5FRpTmbZcYTGh4
MvXl8Aafnb8Q2mR1bVtor5bD3bVb/CJTxKI4L1ZlhzQIJevI6QspbfE3tnMI6MdDfvaM5x3jzaJx
vw4kD9wXE/gM5hZU1NAhjo50yjaIdAhMzGbR2R8zqbdiIQI0xaxoeDh87Xd9s0Hpkr9tNehUiRFz
pXzAR47PoPIE3czDfdTi3SViO4IBz3PdhiyThP48fqYQGABwiJIIG9K4l0Idg+CkraAjg81M0LsO
t2CyIPlKCNErAhUwhACYDQ+XGGnf26QVK7rEf3C1U44YzfGx5a02fzR5Ik3Mlu/1c+tD5HRLl5rR
yBgBahj41UWc71tAW3shkjUpEAgARR0dLg4YA1HIUuqfgUQSfd4w74//J85XQkDqoi0ki1LiIsQd
0pktmHyYAH/2WmXKy8Etc95WJwkFc3UclvFADhd3pMCRY0+TZRMISZqULJidKFv0JK39Bo/0bTMK
NIKG8mFlJ0VjJJ2ZJ64W9edO3zM1cU9Z0M0//KfFr5ZxD/MdXf1i7/ZI8DbqBcqLp5XshWG+5j0o
QKFHVH1IRH92o6JyTuR0cQMgGYAJ1hBAgBNQVaarRQlOQW/N+1Ta05/1qQq9LH3Bc51oYUZpZr8c
rCYDKsJy6xDso8HXV64w8LaMT9TiWKyXpuIREO/BenQuHkmlr5csfplFX5zbOcr3bODBLv5jL2eh
sBIDacKR0i6cklAsw7Lcv0W9MeV5N3lTeL1h4WRp5CT5K0qab0BsTq+Bro/CRyVoad1oT0CuHV0V
wHPmtVOzmV6i/J8wR+Qpdub9UMjwlvhqdbG7fjXDAnh360oXEGzzYLZATnQp2U8R+4gxSgea4+pg
f63dzEvDlgPnxOABdJ3SY2PgVyECn9bvPOxsN6Ur+REuTpPV0n/iQEVxshV99uUJ4hbMbJnsvZJL
F6lz1hKEO1jXr9/FxGtS8u4aG0lWQEw/IaHQk6IafLA3oseJFoZk8Rhbk6VFhHZri3kgQc8HW7px
M6B8FSHjgy6BfoP/TZlu9H6mwiuNz2ZniQfE48ZxQcqRFHWv7j+0UKHHQK/uHMuTjo1aLCN+XDxo
Jw/9AP9i/OrWiaoio6P2gWzyc7G9l26e4yk/F1cwcmawjYnIXMwbgIih/nTqFrtb4+7GsAuVHFrh
q8W8VRxj4u9Oo4ZBi2LX/mkRCjtbb3s4Wxg0zIkaMK9POXhz0J6UYRpUOB6TPlTfCC0hYb/8FVR+
7G7rOJiiJKs8qq3PHABjZs8vceIhHddMpxlGRxWXr4glrRV8aH3gkoHDxQkMnl2KaBtJYW2cQpGD
FNnlMXBjtV1sUgbOHwdjFK1bKZr528RfaCvUQDcmPeJuSa4BF4xf7LyJcHfbQC96LAAoChaUT2OL
aCcfha3NWAD8jibWtLGglWPpDni2hsq+jVbt7qysDzzDLVZpuOSlnZxVfDkFYY1e/MUx1PqP8kGc
Ejpf2XLxMdZoB42HyBL9NbeMd4epUhLWiFTCfMo3AHfHmXe/acFfXLw0CJt35Ear8EWurdme0kly
91JsN+AkVvWKolJWJIQquMiDZeeYOkjzeKB+cVRqU/wQcyC8zFdx93ZUTRoj/R6kdpWb+6saeLUY
/Ai6H6kbybvhoft6BXE9dOXZUJcJjQZfxbcNFjPshne16hRoKAC+CErUyHpROLhCiPhsBi9P3hwy
Gl82Tbqu4eDzjai2Zx9WwdbEnSzt4YP4tajclqa7HGJ/IcXRAOJusAK10DQeRFruupUFWzSAR9zN
ZHlwmFcejKbI5AVTCX8sHzsfPdoy7WkrDT99T3Qc3JRBnfgTrjgiTUuW052+oT7ENE6LymquBN0X
Cet015nwlA8H845HesybLTnWcjYIK6Hd4TTjbmhyaimDNJsgfX9NJQ+m40zGTg/3VkeyIlkcp56t
aa2h3OLD3Uf6CT2XubcLYvGtxsceg0tGuhtM6mfWILK3bZ1HNJ5jN4cvabbqqUHX1Wms0z5Tn29I
ZcDH1i0t0xTFgjm37qagTN4zh4RUl5V9j7ozeLHAlcC6kFPsVbFCNyvqdH378uWfjqJhW/74HRfr
AylERle+XgsVKgkG4xQDJ9qF/mpDR3oigLH38ZW4vfLHtocxUApVupx4IjgR8HZw0hJzYU27s/J5
riUtEZATG1/5x9RQqdkgysvEdaZE/QIiRUIF54E0VoHv6ILZSzMiYmiYnNcDySnPcVrtKRmlGBsE
hoMzTBIJ60CyDhkSco0sTLZPlrz1vFdg9paKT9Uw/vNFAbVym2mb88LS2VASe0xnwYBVBLOVLuJs
HgM5I/uDewr/qGdOkVtXkJkbCDZJU2v9DA7iDjoPW154Kz1RMBD0XCSZfdxYiNjmfbru+zJodz4A
0kZw2iNlSxS1NPztj8b+NlxWhiqpunFru2QFCq2TRQmGuSGt9skj/BVc4TJfCbfwxn2Zuo5mqqo9
622cgF5/yhnIWyrAjNc3sTABMZzML2FufL6hI0JMKQCrNphYdED55jrUF9nyKA0GVoAlF9syoYC/
aSHo5sWqEHMK2xxwWVcQMf2wROefyVRfQ0OkIv2HAx8MnoIsnYLNZ8ed3v86ZTsUjzPzeT18clH2
OllbzmNJ1n1tavuyftBEgQG5Op90UPATKRjavY4mTjjiovXTzn8ugl6bQ4U5CbN7GRMZ/hAoNwdt
VXvCzypooFvlFlnS5vrKIHv9+K8YxhOZUOQmxoTdCpiUwQ6w6fItaETPIXJ1T/qkVb6+Hu6x5lrD
XZ3Z4CPez/4UxhV8loFe5D4KstsOQuFOAm826V/ZEahf4MEicu2oNYlT+u8mg+D5Uv1cZ7FkqXai
zhsQ064Jomd/pWCheMz65b7ooAUU/LXdQvC9YWaatSLzK27hCGpNRMw70DLWZ9nlkJG3lcoViZIa
vx6MGTnb8x2HmAljZuvTL+LUKKcxdom5wZ/oBYZvrCslyrnALrMaQAETdm+oHKqDPq8pNSyu396S
B4c3DHDlwKhQ7Q9Fh4VxI7E5boSCuB7SDiDXxc7/ZkkYxX7adUdgPKa/wcnlE+NFDn8EoRoQR26E
b4pXKEamedBARwTEq9eDEdh05PjdxF1tWP5nWCKeA/Ynyc/HjglWEx/VYkRqsDjS08HvI7aP5Rg2
2JnXDHIj9ZGOrAZEDYqiKZgQoUKApg5YKNU7NG90G3AF71Sau+idOqCSX/lHsUoYxRMlF/XjsmYM
gia9jPFbvafkTNJ0yt/dGYoVSIRIOwNel4yxwUtDXNap2cpZi5KuyFZ4BZhBlOWUq+IcLRacMM6s
45N/O7At9IvLO1DdNCiFTa7AxIrGMRq0Mfs8BSrHE03M6zhjXOvMTQYZg608nH4lXMmJCJV7GKln
4FLS5Pw+TU9Yh8P4wfv9gXLUS7iYJ4VIrowhH0i4GRYgFTPkoq93vFICmZtmN4mBv1VzTMC2FJyW
RfY5YReX06XTW76uYLhxrNZl8UTus2jc8eretzP8UQPRrj23CCROBMceBtwMb03uohVtBOipy6Az
PcDwBDI8FXZLfaemSa88/Yc8hoTutnlDvObX0MysEtJ8XHqMvoA/6o/8pkVZVZiatsPThhv8nxbW
QFq1VRvnqZcFRlNuKEqIn/9G5EZLtsYCSW2+3B335xNfM3qT8+ME2GbTL+rSGhJWvduNHqSzMguR
q3qeXKW31MVNllThCZ9wCP7AQHHQV1vkwnU3UxjW+jeE6z0UGd2z/RMWKWu6dHt0V0FlbkGgaA4H
S8tih0jAaevRhLgqld70YUmCdA1nccN6qmbmU07NvUuY9uf7UaQXBOefIc3xVsEXYCQOWsSXxFn8
4q6rJvy9IP27I8BiGkNdYODE9/AcAsv58jVoZb1DWocukWxTJWH+0iDsTj+l8m7KuFPyW94fQL12
tu9Yh8uUeV0bbKogY94DYtoBcsMI/yC8AQ+kV6UQLSMI9ZeWcLTD4WZgnznUC95pxXO3OoTnMYbu
MBq3xHpeb3/FRnsjHHyrkNqx7snPbHNNDzdNZ7XK46ZUe+ZILDz0dkK4AtJnYr4oG9iw43wwJ04n
HQvhnaLVos9vEnJYte2qpeDXWprhOmsQBfMtq/AXT3StXPDcdSkh35iVrVOU3BEdotdm0DOVkE3d
wLeyeDr+AENCXVkTIvg5My0LfangowJ77MpJFKyO4HjVtRP7CdYT9oZVadylKGgv7heQ+G/K8xWn
EgplOOAnUetyROrJ5v4r+KKTPrc9PwaSKmJ2b9w2UiPmYDoXi4H1MLSL5jBRRnoxzcTINH4DrDb9
Jw5Sy2QVfjtX8WYgHtqAsxTvavhHewlH0KeweM+D4MZ3hMM1YvX9rn6NUCSEwDUd3cbpEPo231sS
nARXn41o1/+OEbbhSOTeCrObDO6MG4p16xNa1piNxCcU7L+pnS2/puBgsuGDjt5vvH6LLf9L+qn/
Imp9nBFoGea2ugqoEItTIEG2d9BzQm1srNFBtk/rxlQenzTs53ZO1uvqsIQlkX/gzVoyPS6VPaXi
OULSYRYxLMyfQ4KlrG8Q5dc/BH6cQsALHMJ0FsMe9Dt6vxTeSjddhvug7YB0cM9EencukWLXTek2
ufANIE+iExM1lOy7JIk9e7wuUGbd4fuUAvhWOR8U8vbPpzGd0Luf/ReFaKcFBxtJva8aFdJg2DiG
QhV9lWJ4nJIX+jg6kjG5qZcQQoY8Vb0SvzevptqQdBolcb56UrYCAdrfQz2jrXLRIvVOqpdiY8wY
boQzbAwS9WhLSHKc/d2fjYxQD9oR0Z3WghDaWpTyB4aMAkcQx1k649iNsIbSLP3W40CkDBES/W36
eH17DavvtVyc4joLP0cZUYyc9zgHpMTot1jIcu2fZ3wza2wmCLqewNz1w6LP2QhZB5cgMhGUDg4i
4GfdpZpTRnlFOI1HF5wTlto4N84pFna8+GREcl7VFz7DUAxkIKW8sCTx2uCXsmYzChN2oJljBTIB
qEDH+gGkZdC0VbfBAvhDDy1kV24kxm9vEhiAU1eBT0AwpJva4NffkEFWfjlRwEyyhssqmdq5ceBp
s0uHeQyuyfGZwP2tQgLfpkVuEFR0VqZQk158OP0WgSBY21vaxkVTVkj4Wd+BMIYC+sIZqRiLSeP0
ih4BAkp+Jhh0bzjfFsJVjQDF0zDEr3B0s8MoKyTtAgFmr5kYklDqBJ9397Ow7eHibqM4gIWcgcJt
/r82Y44uANX6i6KvS2abtFvQBDLQcy8b79/FGGAay7wYpXDh6asYS3Nl7NnN4cnOjpsz3ryXUH1z
THUkOWuoFvjpvKiLZB2YJz2w4VyXLOLdwQKJxAUFOuM3475Xz3NMQT4AgVDhpRygbSSeAMcpgvTC
2NxPf6mkiPGpySdrGwatKlLbUa0F2eNUzWfoZ1W1QNvt2zm7HuhaQvA5vfWiC8YDwZUkDa0Mr7Am
qkDo24eVXcj9BYChru6H96FyXg9Ma2TTQQAVYfAFVAHBZ6EpVulsR3kIDrHLxRqzMdUJwwgL60tk
GIKV3znAVZ6r+J17wGuPKuOH84cU+UgAnC7ZYN+KabhP7alh7Cvuk0Ht20nbAPZxwnuQBieEkb93
G4tqmGoOAGcA6gNK27RGjPWi3DsamGmC9C62wjSuaLwJIpIJ+U2VCOtcxLQZkxEm2oY3C0OapUg5
GiPOFzfZAm4C6gPbyKDy8EV5rY/WnqjAlxj4FLYYymU8mYOEJ7zKD5yEEwjiHlZU7rgDUD9h3xm8
p1SrJLRvya1bhz86zvqHe11AYyDY6gB61pj792d2wmNIxXUIEChTqabHGUoDLc+p0oAsFi/6nCNG
2/i/j508tFlg+H4FClpGGpZ7TTBWUdNswJpIPLuR5VNegRjwBJPCu4Z+NQJ8HbNFewuG4gcpHHsz
gpx9rZMBm0CJ12KBoGTOagWbxgBwawS6348c2RMdd+QIcG/1UQ3rgLFTBOzvsV/qXpyRqRNEZKpa
yS2HCaelNyBYOAhwIxUPLoJxwD7J6TMa4GCXDQAji5ErPn34REbramjuP645FK3fKMBHR1Qi5QPi
Qp39x7Fw5GZyiYiGXoqd5GtAFVrICWm37fuqeIystQ4A73QMWMKAp/O/54RQ7wkxOCeOrAO8+Mrl
ToSpHbkHOXIZglftkQpVeMaTUqnkRbGMQLvsxnnVzCnFSS3akpXpTG+98nBQMh+iLdgNVrZaJSp4
GFuCKw8eFotFz8avlFpW4p8kk+jGaB0nffGBbEYODOHKTVst6Jv+2L0Bm4S/tGkYmC/xCWo2Szy/
BLSiPg0CM2/n70QJIQszr7itY+w2V05+YjCvGfkc1AeJki0xikktGM2TrQeETfLwSPJPHXFqrDfB
yETttDTZ6BLxHy+ktA3h2p59p2LbNBiCnvEUQgeVVRiNiABY4GkVAUMRNSBzUhFCV+gcmagNFJSP
QB464TAnJn7FriYHnGwzxvUshl5yxBUqlWBARWLphVUn1d3VRHCvX5I8KYccMpVTsIs3XoI9DiPh
i3P1BZiqEaiw1Slo7xCiIaCoymBLmM/2HN83TCm4ZkI3RbwZzXhZNe+aeKgI8xXSTb5O69uZ+3ki
QwKxEWL6N0OFVZF17F1TCUflTGGKMlTpFXxkWGAImnjbt87c0HJGhCWDh3lCJb96b144aL+B1/Mm
r0qsVl9dNSPGIvKf7J2pS6HrqhukbT1R/WuLIWRWmIOyjiAMH9pU6qieUoYeOwOJg5ot4JlJZyQH
Dqxu185JpKRlqGyXeBvwnxoC+o93C470qc7TSXzVhSQNSA4WjK7lCdfNVXA5GBjLQYqEJYPDU9c9
Uu62rZouKIiIJBH7XYtM6o8ZOVKpRQKG37lwnLhIi4gRw8YUWDoiqMuVrSllSJBEgXuP3aKkICqr
hg0gNs9QtHjbYXSi9xcbzlr/YkmG0/YT3NBzeT9HJla2IEM/vUk1rIuuj64Pae9EjXn8S7NYyDeL
XJ4EMhyOo8AimmQK3mclKtPng/LBFLCxzfk6ICWnJZKhJbO+kY+TbwDr7V2k+iA9wT//qECi7XDk
xfdxtwzocMehzmfkJUcWPYeQCvKvbXVq2eDrRgUbTnQcPCluOZMuz+NGEsMPTXW0PrP5NN06jIIg
BS37ImePpCgY5oDDO6z5zOEyl3xNAAXCXGc+DSoOIdxMDQfihQZSY/6Sthktg5+/qeR8PK+66lbm
HN8hJt8KCiAAypnRZc+Vr6G+qE73kkkRf/kDwRfANqLRFmHHu+bQuOyVhvMkyV2LoYNf14H9kHVB
OWuU5tJMLkxO4XSyJ9/pyYGY6WkrxmiUSDYlavuy4RBqXI7zJ5uVobOXRedpx2dM+gzIX2gEZSlN
kbqG1l4LFo1wpY07GP8gIB4Gd2KVeWnc1NQNRmr+2Yyuqzcx3/z94qOdhxZfmmBed43dWu3/Gqy6
ZpqujCE5M34WzuKPd0YhUemhlQyfXpBpRqakBk3LOsMhy5QtND0bJBd3PfXv97vAeqgT6N6rQyrY
RVkehL2K368a5WtbNA9+bm/pYE6gvAWV4jDfiIbT9WSb03w5dFo4wSwn79g8QtzUlV0ZcO5KDxdQ
n52cO/lEBkFRijfgy8Yhya/YYZlReNMFi+JrDbOl+2wohjGBvGy8+x2wAP5TixTb3zCevWN35V7h
dc93cttqg7IWrAh19V7VUnNBmCsoA9TnXeWI+PH//+NBRoxRxyEwqOzWtEcRGgE0JaKljEQoKHL5
bAq99Wcv387qV9YQ+9+HreCB48vucj8JNpfx95ocuXT8KgV0vMawSPHMh2tE9dgVxoWxbAYubmEk
1y9Bl8M2yhIQ043he5rmnVjQIClOytcnG0n4dsCUBXYKYE22NElP8YxNX+WlKauIUKpmBzddpV+u
oKOU85Vy7LEQQBn1ovsCpnLh+m6FCgSWpe4xI7UMpxo2idk4BVQofJg66hGjqE6fhfQ+w4HACdjp
8P0dC0o1Iuc4jUV+DWB7bsLd8p6ltbEtMMJ59+OwBfltvcIyqQmmMqkl3Y1VXTN2G1cn+/PmW9/j
pgK3e8JaLm9VGFxYzPbMr7OWhxHI8cMO3+JwVKqo25DXAm28VSYhI/jOnI6BnTeV6x8bKOKyVgPa
cSudI8vpNFyGVJG9pRlvqfZ1tz50d/0Vf23xkeSZw/mF/YJkoNVlMRurqf2HXV9Kgh1oYo0Q8koN
A8KF8/MjnuZOZ9nJggeu0wEJJI3ftsVUiDxz581cDKDJQSRe69qaCPx7mHmEzaZ0rpvvJa/xrVRz
htnEQYmRQ+9JCJaCh+BlST9vnqwTUo+Bg5dALbMREsqhkVUCAMWlPSpmI1iB5a9qDDhij9pVGNRZ
cIRSolp4eLpLjLOCKkmTMe91HB1o9lEPA1zjeH1ImcqQUR1DOiRagA703j+Ng5mJcHkDYMrULNEl
F3jbPSEqFcRySzV40bX72ApgmRnn0teejDwMFwmrUdaC0k1RIAdnkZGc1Utq9EcE6QmdM75jd9g/
NOnG8w+70nMLxFTwqzeG2fzfyIIPrYhojEb0qO7yT8m0OoE/RvH5mFHJDy8/rv1UIkGuyp2uipGP
KxoqKUv1I6AaT1TEW/qkHqvR8E88Lph3Xnebqogg6yB7Ry9CPulNPSkI3atI+7dnQ3kACBlnX6kc
uW+KSUdaVWd0aBDWjaaEhOGIYCNU7VUlhZTn30NS6Sc100sv3HJqUBiIQla7vi44OcQn8dTTiJ7b
4sC6wr0Y1GrcLLJ3utt+Fu01/BxhSsCgK8qX7K90l+kYK6hX3elW9PLXGkuPI+PsUOi5nINXIXGx
exSmLjg8bBrDsGlA3ixQKaRK1o+aobWZzt/ErdX/b0GVYIAmOLX0n3inDKFD0hbma0uN6PETJEhQ
smiZZjSv+sUGuaFOEjahBz34L3S2xA+y10b7ZKUDiJ1B+AhyHtuuDtyJMmsiM8fFnx6lAG6arnM1
w2cy6ZFcFwts7aIrnmnIbic/A1PpoHP2gm2zySL7bnhIwaNhzBwyXGLMG1tBZV1dm3wBBlFKaMJk
E+0mmfeEMDc0elN42rebkxMJQQs4Dcwok0UGu/T26WKd7DCKA9EvLdMvf+FKfhJ/o2SWEfhMeThd
ykWDIwtxyu9aGprQjomYRjhOrdUvZX5tG8+dBeyb/zkMZvCn9ndZ9ArFL4tByctxPvIXis37j6NE
loEbba00BTjKDTPuqLGZuiXtmx+YAlMx+mtltkTJLqrplJWCTOsyT9C4Cg2TDMnjWM7AkV3ayUmi
8g+0tDJbx9ma6Pt46rgwB/BSX4Udg/JhEXK8EOQ9cYNVnVhu8ngrxxLUxxMYunwlEQOccmQw/3gt
koDdDB9MeKzd7r7wocsm/Zmedmdfvi0/UeWelIhy4FQOG0QULqsqeQDTp0ecKwFm4v2Dm8mdiRXo
Eus1IZKcBamTysNjUi85Px9zutQQZ4jwHLgd5Iq9E5sVP66SMmKV5s9BZUuh2BMqgwraYLOOpsfd
wE1ZngVQJ1V72PvdQQoMtlRqnEQChW9Eq+pKIddP7Z2+hLnZHVnk/Ng2XYQvl8T7+54rCgpNS8Eu
M8DEKdD0NvbCNnvT7hVnCw+/rwSax5yXpBiBWL++MAYKRSdCqdu6RsyBGNftFbfnhF88caQBxEF4
ZDzx6PZuO3jHSvXpCwALDUVR1ttoI1+dvienjqip69sFbvjtTlNWPHXfw1PazTqfH152fcX7/dQl
6ZY4yBwBRV5ZELlLSjdAMbspMcF/i5LhGWQr9kl6UAn6vY+kFHzzy7QMzCNevdsKVYUc1cpL0oxv
TrfjNeLmmPYNcTqInuUPji2sc80l3d7lN73Pgg++hDjK/E5tuX1KpfykewNRIn9cXzkqZLYqgdtt
LxS9pdQ8C56d2pMUEV6IqJkBrQZxUnqoiVy6tuy3Y5GNJbpB1gCpUJEWgvlQP+1ZTJ5BzUVvBjs1
8biVoqsqjVoXX5odaMgEYiYuihoKA4/tPF6+jw0rQqWJmt8KtWwZTJ5dz68PpqqFjUPDsLSmr01l
l//3NkXzS+jbOe51LDTnbCySH7Y2I6PNb4f0TvWNSalrcgZ9wZfQOQwKEjhmcU6aLJlTBBIUS2RS
Xbm26HevA+GcTvkKENO2zcuO66O0K48S755o6xvlG3v1EbWC/8raxhuREwFrM7t7wdYrGLdfv6h8
1hC/NKX+qR1KaK8zp+1FkRqdSPu2p2Xi2eG5wM+40zNWRiu3TTI0+1GV1+GTHtm8hH6jHyFdGm2a
i0d0LFIFLonDaZmYuar6m7zHZNWqFPCj9baqVVxz+oGuO6ajVjrc3mSxptXDpdd//ggVRKnCJQIB
5FjpgBmVc1avnsD/e1byDhNNDqY3Vm3PR2XaKy/eMNIUzMX2KCjuWsLak7uS0/OC/LF/TUMc84wH
PhUuAIx/W+0XgoFOwAf+j1UC468zDOL+DacuVlq35J0+K9v54s9uwmhNDxghHDpAbNKeiOhp+Dd5
E/dj11gRJ7yZK4SqM+c23/XVngRPVrnPq5DUymxWknRH4NQzLe7nAoRA8GLC8NvKLzbaOgWzhTD7
YDefpwJ0eTQj7ar2yfdr/WUtRtg/b3W8C12ar63vwSOc1cVCMvZdWASqzW6SMYDnj6zc5+cyup7L
C+2RKDtYaNMnkd5v31l/GSlAAi0HygZKZn9cTsddgBvd7BPpV+3tA6gtzW/wvZ/C0AgA09DrMDib
R1y6wwsh5/+DmqYn6uHOo6MJPxj3SS6B55Z22L4p6KhvKzQn0HibJZ3xo08EW8TE+o0wgZEu848y
MVdOSejXu3alKInCFjivJPCPGjbojsn4uJwD8E4N0aofyT7tTc1owrX2i4VAmFcD1R7zAdr9Qbno
mARGip/gprX+kYZhMMbm8eHthyYfZ/QZ90xmMyARvxVpPnBKQeLZU6943r9NsKMtJSpkusknt4VY
4GveC3sGGEp1SobfsBHqxS9/tBZrl1N5o1hDsnK7IGxWjKzn+m9Xcm7/LoCwvTzqMGXKtgTXVTsv
+1A4cNJ6LoD47f6OvmYVe7gTosNliFGcaR7eg+HVmGY2dfDNOIOrHt/FqYretn2CXS2Vo/Cw49zK
6XdZZU0lTHhV2ybnxzx9BZ3Sr2x9chyrQqt78wXZVgr+pqbA4+Hz5kfhGYMRCw06VoixFi518hKm
PWc/r5J1SOOweyoAtC2KpPTwN7q0Ij1LyAZ6DGkeuZ5hNrdoHcmO5u/Vuvxcuw7Sa7g/WSEtHDDx
R9dRg/JebtyBe72FOHtfQqSTLeltUa11D/3Nr8r3Bqt+C8qKyd4d18uewM26/1GGy4K6wRactsNg
DNputIJI6hAGgzQsWK/5dKqdxIgnYKI0/5XjHNraknVocA9+GwPLuERZqyMqud0eFeVNuPwSHHzv
L4CiVuji6NxTPRP54so0HaEecq/vFbrQ89KALBWxYZGcuTOOVs2sfTdfwh8K1riU23mo8OxyyGTD
SPZMDs71UEnui8K7m4FSe8o1NAu6j/cd9mUqo/k8byCeP5wBSPDgU9xKgYLliuUrN+NzloPEBrT4
+6eJvvE9Ldz0M7siZcys5yZwdXwVOhoQjV0YEXfnqWaxUS49cvwr5EanlI2LIxELLp9SzggPDM+P
HrEzxQmX5xcoMnGnLJaZ40QusTMLaagCLm/lUmBkRx8eI5UNtP4+CR8bHAV0hL2LYUsUdMoOHcja
0ffm/w1xw+HyvgR/7L5G3QCFasuI9OmRw3o6KiPO9YrVPWfY1HmcHam1lPLG3jJSZEgMZhdsysSX
UWtLBdtRfcVCHv8rDjt7rGMquCGZ811AJsgoXnKKlzW1sV7qKq7SaGqBf7hewBhwIKRfMRqtdBXk
sX0FuqW/WBlH7RJpE+lI4aUlsb/HjBNDDmxc74Stx+ncBB7Fr/AkCc+reyNnI6PWrg84ZXRsMx6b
H5Aous/P+VpNG4W+sdIIBjD1yqkMP9xGHAye+Z8GeODIgYXGyeBS/7p+Ev5892hCljTgfSDPoNNb
h6TzL8Q3fsYYovwGshkFLvAOtAJAC+vti37dgsYJRN0dAXNfheuBZ5GU1JYqKT8hHMWQJD5Twir+
yxDlA3PPkK/mxDjg1IlvrOzSVeR1HyHSkn52Kh5eH6mA5IrHGwqFUD/iXn+5lwEGPGdXawFBSQWT
lwgnGKiCiqLsJ136vIu+VCTkIOW+MvLCtUMb7mCynmLJNKDQYFQdBSkgSmg7F/Y6Ap/2S38mUbdf
TkQ1K001ocELOjtxXBTGppKAX3RoozfUtUoyxV3e/0ifUtaCdyn84W2nMni0jsJr1G3P/jXvLqxT
w2gaau/OsHASYpPFYxXmlMxiLfPy/yknKJlzuUMURzqpuimcakckT8lHAtVqCYlBf8LYQ/emLBy8
W47f7Ng9EQc91rKJfcoCJEo2JJpGxeyfVOKu8e8RxS0xt3Gql96dXEJVPnx42421QmpM2YAnpiVF
+/h/5RlIrTflIEOdaU4pMBfhefFOYpx46uRxwETHEg9GDhGsCNYusjTXf0P5cAMoJ7Qfi9VtN0zn
2sPTUMhKsCyFfJdfyoDBE8nNTnAlEkVEcKHx7ct5liaq+OExm1mAA7PZAzJqcGVtEivfZXiPTvhl
vfgvHPEAlGuj+FerpabNejr/pN3g80uYQsXpOthShXg0M4YzpgD4Zx7Bhe7d6jxhfpvWv7GCwjYm
KbV69SpiN+/uLxsrfAsFKDcxwAW8TCMYSq4E+FIk5wtD2T5CO+dU+amJpaDQuU03DQ9gJQSpfrTH
gp+/lFK3VcMYjgNnA8quR3W4TpQPUl11haIBFMki8x+xUdDU9v8WpHH+B52l8wr7OVqYQqtjtz07
GflAivA6N1SjFc3exDAVrag5xjYBCpWgbKtjew/QKjUqzIo/PT679DNDEBzyiyEXj4CV6jB5rvah
dR8I7mPb+mIYEZGQmsei8CBzQ3YSyZ836ypK4qHECHl/5FiM8mKa8E7q6tvFy5pze2QRisYQaEmy
BE5aZ+/FFc90GZDi9jNnjYfZmZV64QP3sGw0fJmnWRDMNCY8DEi4kTtZHlznXnhAXkL9dRovPikJ
/fj9S+2RdeEL29xD7tEBLUEcAKJ83ZHoaxxHkuoqsSiMDW7TwYL7eRt1ClxUlKTyhu/V2caGnYB7
3XxHLZ1aCB1ahhjHNoFDYxZJ0JqpvjcUmrMKGNvFh0Wu8JoQqscDXcmm1WLi/DVZdN/R3G+3a2Wo
GjPmYPtbxsWZxc1ekDbsRqjPQ58A+xHI/Qv9dmMALWV2/a6xeSCdMzKBmwc9MLA/bfWMZClp/+0H
qCrJS0kvzf/lCf7QvMQdbwVvGx27Q4fE3AteJA0NzoMCVDhRagI/ExorsWjsdHPFwh/1WqxPmHm7
ZuagYQMQI5YWLdwWiZtD30G45EWX8CPvgAVOvasPznz4LHk1j45S4eiil+b5pzWLq72/qNJT7ess
yMlibtdHtG4QezcC5ALgMeloSx4zVXY8wAoeBNMuRmW035L8kqfjXDdTa3zGB1cG0uh0oZYtrhxH
uvA4CT+2zqgSNrY1aVNndpR6diYrGYZqlne7Ju4GcGumXo8MIVRoA64vWVID0VY3ZsbP1QlFa24o
uVaW5Dvq3+h3KCHWdGn1gJ0ELMNNYTZcjpGyUDX5QY5c5jioL3p1s/BeqG8piDY2NxbWGU9NH1Mr
bOAbNQG9tvG+b4bRCrTdpJQS9reYc+F2nnt1Z7agc4d30Vlp8yaiXtHvlNeHhX4yU7ZMIeSxXlnA
V7+js7VOEU80MobNJU7r8LY6J6aAB5wBfoN1Ou+Q27oZlpcSJNZC9haYAqLy1+sHOrUUMmOTDOCC
b74GrgRk5AE7vRUNxz1YedoDfrnvv02+Aow9bdXQ3bVe4aU4WOciHwYbuqlLoy0Wcm2a/sw2f90k
GUedfo7eJFNZd77x7yrxHRcUFxay5En4qhlejkEG1KIkWR2hOy+nLQvmY7wOUQxd98OeRkQooN6T
pWCnChINf1d/Hb09bcMDIdziqYioJ9MekVhYyQieci9hWj3DkYalAmpJTQqUnx8pN97IxZ3a34tz
2ZkEiS5zaFdBgYD2Gfk8Tlcr2NEhHSWJylKSANm621DiiMwHUITYvf2lOV7B8+xn+CXVUYNEC0gp
CQMKgaEFDfjo2qtCYh8ROjm4gGypkvTI5BPhyAsYbsLCsEiUJ6mMJ2ti04byaBuk2j0hV8ZBBkmm
9YOv/u+q4PS++xmSJnrcOsnTNIvFjPog/tt3rJllCLPYHj4YdO+8kD+OoIHvD9pCVLtMGvuZ5iKU
l7ulH+DGY+NOd8elqeH63X4D1IdNCrf7icR4rRkNnw72xXLw6zH73DgtU7qYceeEs0IBTOSSgdic
r0FOxv2lcPWGHEkZrye8SftruZuamifCgE11W3FzatmQ9WXjoanWkAFOKMY9TPMCa2WwXheWNKyE
vDLNeqNJF9NAUV362w5gXzWguJIlhZHBNdx9pP9tDWX3ci4TN/khXhuT8/bggbK6gmTeAPoMUhzP
EbPRyqhdAxHVyEp/fhDYUudnok3Mb733jCfN04uRKPzWpVpWuNZlV9UTcqg8RD2r9peX/bCWQaW4
JHndHYS096sn/Tq4Mj6We5XZNoX1gdCSzdoUXHFQ8OKe8w7E52JTCBShdOM4/NeFn1nxBWZygyFX
CPesuBxvxQX8hOd7V7eQDW/266TnznXRi2CaJl9okP6P1RrYuKMRotHDRqI5Nq/EGORyyGj642Hr
1H3CqrZ1rYT6Wmqy7Na/WSuJ4hnOBaDk077yJdexuzVezjipvHI2SzRS1SKyGLz/sF8AqYzVQK6m
6xAfPxtVn00+VTLpG1pPkKFj6WGqr5I2F9YXHOoZBMC462b942ft2FD9FNILlbVhg5LmjBk+yfgq
+BM3WRulhIBpByO5CwaIhn0ME6B2yqSB9gG+eQ2km2RvIK7NcfM1N+hnb66tTS9t1S131oN7zkWr
iGrjWgGJZ3Td9jvEEvP6WNu2fc9/+BD5WanEDDhbdvafIHakvPQ1/yWXdTCMtDZgOOlrMO/o7QWv
5qK36zbWtt7HVmecWV81u78nuoRQHiWciL9yVXmtNzOUkeqJrhPkoyYs1/QwX3Lqv+7M+TrZlShM
oSQXMQOISutepX0F44NeP3KbZHOIJ4GYou4uDlCOO0R1sRT8aT2fpmxggzLcjAeyxwh4rmJbX9Hc
GLNOQJPMfB7Kt8FPEZlzjWXAJy77NpvrRqSNzrpQvaW7f5ZZCrTJXlO6But56SNdwwQzoYGIXRDm
cB+Ac0GADlehCt7TeVR7+bHxhOFbgH9auBQqyPbV0F+imFOvmUzhBpJKUSqByqarC1SHObeUm/1r
q+Ofse3L/oO0mt9CW8wNhKUycwozaoYwarw0WmijY0DlK9SOuhuhXD41Hyqr0xkLUW6Q1gUbx/6/
gwK1UUHhQhE5RvspVuWwz2GIpUU0t18awSoTilfJkU/J8Fp422YY4jjR6uGBwplJFsJbFCttFudT
3kcFTKwIHwtzSxbqPNpmj7xOa763+Q8YbrWW638p+0A4FLEo3sKqvv8aV+QpIaH9WkzWcoCG/gI5
t0VKflUfs6I1MjJLGtGo6PIbRthtSfngFsBy64WPNVLNidEb+EE4jk01xf5DsSj0ydHRSdxhVzIt
WUps7JGxG/cDLjkbBjaGtwhElR72XyWzFxBXUye7TYbnhkP6cP3Fdm6ZPgQOMwbkNdPDgPq/c7fa
DfGQVoY4i2aH3Hy2fYkGn3tz1Gyp4E16Gc/RJxmWmzuRl3E5f9KBOFTjlRhzdkFZHLGdKxJ+1iCM
oNVye1fES4ViZYeXh7+tV+z/pfE5bwv5BWk7B9xfSkzGBbI+kuBT0ZKEoGkUIGSsZTI5Vjb4jEJ+
LPt6dhFT3F3omFy5YJCWuEhqAOL3ldhbiFBNV08wWt5PINpHDdUVvKXp41NFzHvvxB5DzikUIsy2
s1On01wtIHQ1Mj0yz65qi2Vk88jWeSvn6QTQqzVOI3LJkO6KiCYzAMCHFlZdYgzr4oJJWSRP2T7r
BiYqq3LDy7AMjsiuhgGAfOZxB2lN9P87zFrJjK7fLQNtQ7mF2RNU8WXkGg3GZcnUwzCI57Gm0bgL
HE26clK3WM4EVEDg0YpR5w/rTOC3MY/khVTSZh0KBGXuFejELbVY+GRc+Mzk71dX7+0NDvWvNdrJ
9OKSTH+3pTrDo/lJj76ORqC7YvnxKl0Ob8Ocm/Y7hYLl7OoJl8aKUycRgVHex29K8CKBaaudM/fh
AP58tI7uZX6Kh9npO0tbDmfwYvGeZqqEuVRl9HqfT+eWApbxG28JjVQuhrGEGvrbvfwduwXp3HYz
H/vNvJ3+ukj5EezOCoBpOjReeLyccaMcU6/l7kmbdSiKQ5g4fRlQFm+fdt15p0WcTwH9mHRLmLTl
S/5sLvQPRXxMX+P5qGYDUj8x2AN2UUGo6Q1w4G7x8jf6lJK0xwn1UzEPfm1xIFhMaQZu47Eo+A/R
eclHwt6mcNk0RxETiTBN/xSKgxlw4NfqhD5ff5a2DPwbL0NCNKnCP3X3EQVNcaSKd2hoAYtUHvbq
pHjwdLgNFrXmQssoZm2O7Pitd6z2JLl4CvxCg32zRDyHc7MnVe1AaC0U70oKFAZSc4XkK3IlyNkk
ctW61/tLIp+WY8bm2AkJeN8rDoykolIrU3YV7d1UhMRT4E7tV5HvFhrFeeAE5ixb/hX3z/6b9rbQ
gNuIm1E9MbwAKzuv7fnBjMFkEwWwn1xO2BHgZZf5vQbM4PooQBfjz4lTN9luv14FqNUeaQkSABF+
ADzCBnn+DYlOkXsUHCAIaDrDaJYW/KqtMeHXEf8gnZlkuUdnCikADpd6qc80dUASjIl50kOPuIdT
Bn3StVHPQiV0UAuLA8SMoOgA9ILnZJPDxkQ4k0HSGzHOoT60+Tb/rETyWZTH9zABB8B1lUjthP1X
Nu98K8CHKomq7EU9VJNo0WJFpFnX3Dc3SOymmBZoQcGBXEY46lNgbLwZMXfBFMqj7WxnMSKxx8UV
ngn5j8U4Z4n8uwuUhPG3Vkh9e3Drk/ATeud/iCT+oYdsyaWt8ycm3IllKkFI07Mb42U7lbeY8bff
x7+Xm0OychNJotAcsI/flLLTqZwl8sMiK/Vf0uF2LczjZIYLoEnT+3v9WmDC9FksvLY2GsoEDtSg
QQPvdmJ6iOepGBLyncKI3PV+F9lmajcqvPIECjtWbvFur8/81+IjeI7GHjm1KUUpTgwSh1iRzvhz
rrn6y29FAJqu9MoWGKOkfylWutKtG/eDkvXq4KEfgOhwu++h8MmilJyIr/TvvHgnU3k96xCKKd2Z
ofiiauAMTm01hk08GxHVOHdH5sA7+fkDSOVy6x1acz+CW8sKmLmoSDiVWsNMvyGuLJz7qHYjkPvK
33YUy0vh0qqT52O2n0dzVq3EVXg024lnzmYI60k0dARlxQziKPtffv1yoLv6rFMVQpUqNrdl+Hmq
aIlZ1/f/oM3OlAyTNdwYeFAYYNcrKI/92DKiSjjFlxl+JsSOo02K1C8jUm8Ao+IDmuu8z50PB8nt
2fv4rRvA2z7YaULgtfyPNCaRGxDnmFeXvyEagIhXXxWgQ9fs/Ipovlkmg1A6YZOehlspABYEt345
EIlTkWfkKFH3tUFee7UDtKSS7aj5cpgjGP87p9TQdwHMkGu+CXYEzlP/kN/JPRXsCh2I187XtYr0
2JLvUW/Gv+er3sSHCmLivxwP+qep5dl9cosfaAlyUO9Tg7yF8dBLc4W3tTNrQ9KFeeFntpYiVH5m
JW5l30HL8Sz8A2OHa99pw8eddlC7K8fQWNl4OYqFiYy0s3J4oHWdYnQ65X/OPv/Szdlp7ZrQJqPF
CZLiTXIBUWDLJfuOElNUvCEY6HFQLIehcWKsdZT2XKgcHqXglLpe/HvZfjpBbn6wf+BFsTeZjH+j
5cMR0xraaCV2972gpdHsWiuEq8Gq5V8EHoJy9sLOtsVES3CCa5VJxi0rrNZNZ2yw8tHuJqYmOl+d
wxdV/69LGnJ59fUhelFULYyy6z5nQ7Bk5fZFm5hTcyl7bsVP3mgwHPFC6D3lXgktCW10/4iPg3Ni
iImeFqmS2Klt3tiii3NWyRjkmzurd4pf8s9+s8FNhwTGu6B+NByuSORlLBrmsdebZtYrM6RhtPhf
eozoJSaDkaA28EVUaVZTiah33dHnJ7fOMFOnmzd+7kCH6ri6Og2vIur3gS8aEcJIOAEwlfmKJVH+
gV6zTnrwRX/emtYiJRXaEdXUGWlBtYOFqjJIpg6HS6wTGctCpGmKJkRi7IPkKGuL7kju5JqQ21dw
mIrC/TzvH3qCanVQVHn075hpZZvVSgMe5XNB1z5rc47hydj3/KiYE4iRzwDfHXjhRUpq9sbbKstH
64pqo0ZkDSAUNSVrNTYTptSgGIIWiZ8Eey2aRKnaaFrQKmDEtxJ9jw+e4fRVgnzm96ETaCABr2wH
n8VFhMBVZNe/HEzC86fc2HxmIWRQlgc+sVxvPMTwLUDjrhhy9HNrycTFoTmPGDC7GRvI2bS4Ea45
dJ1gNl6w/kzRCKlI9MC42ZL0uWU6h9qwIb7J86ZC88tq4IglVffzqvkpRZ409Juuu4DkZgUGCAFc
WdrJn/ikNDlaC2Qg1OBMDr9zgPCUHc0iRQ+OlCTePYaJfDuh7vjFzebHbTjtI6vm4SCbqZRX/UqC
jXdxxCc7UUFmHcR2hazdH8SjthEUI8R4LyOaz0v/TmwQf3iqPKO93/IE7QLH7rk4qDEGkjJALYMp
pKOJuE+pXh9XmPrLKvX8uYOQ9lL9nlBMpnbVDmFZVO5hRwvz4a409Kvng2PkONRwQvSjMphLPsBC
oaqRiRCllVDnCFSnbbiz9XLMsHcn7lsw8JCGIB8+CpwsPD+AAxi6DtqqvvhC4yHrl4r9Pd6arlqg
UIi0xLikgW+GGnIAL6ceNP3Uddd+xEiiUKICFH9a3rP8MGHWxUBhkAn6dXwmV8aa6ZdH5BiYxqhE
VvKznbR4nGb5wzzl7aAjA+dt3Wqzgs1MElJbj1W7A/+lhYI3bJIV2zFAdrgbvzOQrbvOtav23HC1
0QRZXb+B3kOuQlN/8j2oO9P+t1uuZ89FPduUK0kwUTrOJuRARf4CKlKt6fzwRPwFdZHXlXoFTXIy
jHic8VgkcoT0z7dVmvdbean6Qsi7SZ98AVMp8Hnhbw4z+rvob+reDePWkZp9C8uqUZwRS2GUku7t
vnjWeNMpbACgoWBYsSA5wy0DLdbhe2Uc3v3IUpaCuEN0JFUf7/gv7KAiGDJJC8otUHXlfz0Fapcl
l3HPTJ9U7F8wr0yThS6PxTp7NzG0Wui7GdP7qWtFqtuE/by9ux2vM72o24m7IRvdAfFuiK/9dxc/
upXZjt832XU3sAFg9e7gphaaksAqWDOqgWHRT7rFWUyYCk6KXr1FRpnpACouaPg/9gACFEXPDbXa
r0vPn2U3V5qPVP3VRadvrPD6eHvFkZTxR/VadtLTx/Ggd6RWfHLstwRbgP6OsUjkpUuagUsAOpqQ
nFXW36bpxQDR/REPWZD8lrBkPPG/PZoaZ55IELDz+uD5CPxTXSfs2Qa/7Qbv5civUv8Cg/ZO4ZFk
CwqJNDUvCZOBjTzKywIw1rCxqHLyc0u1y3Q1zDWMldKkVQUxY0FhtVNQQ3yt8jfSzFTVn2at2GvW
6yu3p2E2e2BkOaUoIuf3OEdJYNzZrflJ2kR9svVwUnWAQ2AYA/wsU8fdqMYNiXA2ilq3bO/RXxWL
byUaNqsCMeyVYagAEr5C2BgAvFwvQxi+Z7l+jhUDL+Vqu6zU3hlcV2KMbgX/BtsiXXdLkYKwS4EA
Z5ncbmaZBzxFCNxBEthP+Q5y1wvm3/9QqHLJxz5pZqlOSMpAF/8y286T8wZIYRb+weN9xDOOvKDX
ecJQG3xrYdltXrUyfb8oONIhv9I1x3osJCL6Hkp7MCiv2quRv2IC58R0pwlZ6BiGLkFMSscUgXlJ
IuYHxymIdhoxTkSIjptlBOugV0vhLl9NLBrFLT1Ud3m/LU2GaSPiY9X6/sCQcgbgHiBXCtE19mWs
h29/NJzWz1UM0lDNlEoxn7nvO5djM1yDbPYcWtn5iRkmws3OFZc2Oqqx9mkkLwpDxLcAwJRcryVI
aXmgPwGu7FcSO2ins+JWJWheG4zWk9Za7eK+45jXdAULVyeEO9BmNVpFAsIMg/pPQk6oGtQmYJIQ
Qh3RXDr+ASO2+YqxImtuPExNhfzI2St8ZoLCpISFRGvQiEI1f9t917N8BGyZ/UF9lj513jKIkLkX
umOFrod4EEs+h1E7cauCOq2Vp+8L0aXzVeyWZYb9rjnVFjYQRelj2bsLtZrO81+20mTIuFZgqRCZ
KKzeq4NVDBtTykJo6FNeRMX78iHXxb1Dn9OZ15kZTFXmGfdCGZb60C5yE3ZwfH74N7Ws/OS3vdtO
pDYy6qhEEi+yALbPfqd2es4CREcZq8vK5HQEgjPjBP8gGSMH+lP575l2FajYWjS11wM0h9EOBww3
SsOOEk/XhGTeXNah8un3I8nIqVYLrTpJGVjBU/gXeWvWwwbQ2dlR35LkJxzAjDG5KblzBSUMbYHz
316ryHQDp+SaM95IwkpYSAgiH3nDd4TC25JIGiUUhBkLktNEoaVHRH7xRsg4ygg39Ov65Uzyf+gL
WX1vF36W9l9H5n4Q+qH4XcX2uziPqFbSBhRHSXLkNM0J0PQqdCOi2zrY+ww+7+hlOC35t2JWbvKm
Hl4t959gpxdRpuW6YkOsaZGaSlZeasQj1N/yhil6GP+A3gzhfZW+9tu5juFJUla7gk/iKkAZvVgY
Kq839q2VSQbTsr9BNzG1l9+WcoZpToqFNnylE4DaJkZk465jra/uQesuq6XeXxOsxPxvZFqAkBw1
rDUyB+1A8deB7snlZfNvsYramqOMzy6pjM+Z7nuq0hEuQzCV3Th9bV0Iqyej69cCIQQMf1yB63C8
fm05S7jn8KILjI/ul8Togy6Dxm5kpO6XONDeumEIHHD+Hu9pIDLE3/HtB2cjgEKGahkkElc7iRTI
P8h9KDZBm9dkDOWza7oIQjFbkKwIM/v0V1p0XJJ0Be59c0P6B/2Cm0oFNPbnw3rC2qygzhhI9s4y
BpdYzqxukVPi7BIkjZvKXsS2pJBBNV1jvceNSKUD7zOFV1zpBNcjuJYDJBslnMERtpk+YHIGsH3+
ADTxUSwCZ9Q3y35LoVWQk5Tyx3vYvQ8t9ipwNAywVer9Bhs/W9awmpOb+nxvPGkOsc7Ia1QeBe/6
3bPf6H3C3lIBy14d/9JPMyPcajDr5QmcTUcoL7SoUp6/2g89LFh64gDfPnJSuS6kOpco3GIoVzkj
nJuBJz3qBOakE/jqCZy5agMKUy5IKoyZnTBEtEErJ6RU2vxrdLYCv+C3lgHHv+80Hv1xDg9X9MDM
H9dKdhBk8vUWM2zsSm2fislpXDcr6VgolSaDEu4Q7zkIJ5G201VUwNVlWK5TBc/vp1tYhDzIqyaK
OGe9j5ZtNZsHW/8IcFoh7WL27BOUiuog+DlqMJ33Rbg7iFu8oFj+2ibUzbPbMU7xDHkVdPrn+Lp6
LNe5ANj23QgagN4LVdJcHJRimx6roKX2pzo6d/PORHgg9y9RX0hlEBSTYWPHE6sXrJoYW9pks1KA
/86OixuaB7jd/PdBHaf0msFC9aedJdQ/VhCpxeqJj9fKOzdCTSXkNEVYFIGs0nJwiKvewxD3/iqM
jLAKq4GVJtDvVxnBQUUC47pwjkN1jCIDfgvud1c6qp4xpu1EzHC0YgE80iIjKxJDAGuuVe24Evun
m7ke6GULx+ggQm+g8t7sxUeQzLUGpbOG+e8nQhynIcYkwY6rJm3h+mzLLiYlDQoid9XK02QpdZ7r
xJX/HlrDZBSgO6DmT1DWhN7rE6VXJFL8NDlop/tcBPVJ5ZQ+L2zpsGVrQFTibba7O6hRX8+ZY4qL
cPWWOySQX8Xf6Za+p7Zad4Qs7xLkuviDD+OFqdegGTJQvB7tEn41LBzR/nsBqWt6gXN+7k1Byots
AtKOs536hW3963lnuaG+QIw/iDn+vcDlrneblXbIPfAxJXb3Ylbret8kPT+2J+vcCHHkxfvMi0R4
dB+rErqH9NMYwrqzZOOv/9VS0YtFXfKMUawWuuhtosS1Z0nCDJZ1WbS7tbEI1V6um/MDpd+Ko/1s
E613s8BRiYOeTGGabtQQyWmWbDY7RQCsAr7hgHk/xmNkDMRFQzuaioPIhRzH+HTlwp9czi1/TNv9
Yfr2zxS4FjvBHW+koKkutdYyd33eoembi123ef4N3njMwB49Voqu4Euk4+Jso5o68YzZGuK9li/s
VneUlTP/8O7kYSivPeBtBrgXOLz8/cp9V5Z5li7sV1nHZDn7nDTKbzXDcfMjH+8G3GGhQzbhLQvC
xlfdlUXGOTl6/377MljDGeWXoDCmfJdJy5gwvSjnwy8umvvtEKL+MatHMljsbwL7klL2GLWdGlte
FmbvfNKsiRMeIpDDhyW8ib3UUy7kEijy64IAAnx6rpZ8HxIzw3LxVYU3rwU6XwO77/hyORXCAp1/
IgRupA3nPiakYJWx+ses0GDhs/RDbDRTrZj+bnyCtHstN/tt5mnMgYJ/dOO/QZup+0pl8kwbEGap
dzY3hv55CAL9eF9sSpNe5p08hLhvlvBXP6/jwcPBSGuqV32ymNImr+Ci+J3+7UIsEfM4UY4GbPtV
UhDCaQJy/+ewI5iyaGBDtysGk9d61PcstZ+P5sHvrrXo1TkMCv/b7uwD5SVoRW+CHPWbqN4ROjp5
/YJRxSeg5FGJMV5y/fbJz3762yLAXln5WlnPcO/vfp4yxsyL4JjXknVJcGo683Nk5rzZfohcfO0z
Pc1N+zfUpThoBEkXn223GHF7xwWaVZWGPPtQDJ4TWxyrxDN9wG5g33y1RpfOQqY9h7IaVGLEeC4D
lzhAk0c+kelD8Feuvh2ue9R8xY3D6hvIrAH7AaUts01Mmw+t6iY3ujhmFQSpZdH2Ttg3lIGlDBKj
tuCpFtgslsMCG9ZLxRn08+OYhZxQcx+XpndsnaDAcx/9Dq9tqVZyDncgxkdyShQOvOyXp9Cg2zGA
u0Ow0MlkSHgcONVidzE4eamXrXGomIASpPrgsU+RcuzJDU/ny+bkJUA0V94cBn4XmN7IgSPi8Goj
7e1m8NQ6VJjDMIhthPyxgzdEw3kCrCkVTgAs7TRXd7VjrfUaU5LpHViSjS0d1ajW7fsaXrpJ6v90
WmjHAaJpFUd53eVyHBIPoTTsdXfzrf6BW1SKs80ArUNxrDn2CSAD7zWBg0NRjBEb6fiFib3j9fSL
r2+vD/b87m6ejt9tU8zniFF8CbueUT//A1p02tAL0bwZeDrAej/qGREBixcgcVD5z49YnifFi3ga
o2CJTZQ+DBO+p5/Gqj8I18sTyji6dvFUfj/McVe1pHxPqJnVAE1NLA8vLWzpIXDnTj8as77xxz3P
8zt3qFKN+j7h3KfIqitND58IdsdE1XZeu2rKOEk67J9fwa1jAi57AYMIH5xEIXxsiAMQPh0/EwI0
VboxgrNzlagWUWBDTcFuzOTFlu+1VZOEXMKmq/5sQ8+t1QCgVscQK72llVSZewtaJ8BC6OXNEkpq
RfNJRG/9ZAArORrLAx4KXa9SNYiDol8GzhrFGYe9qsxhghtHXIq6MfnIg/11lxs1s560qd96qYmk
a3XnxgaBtRk47gWRv0z4JRYMNZRfmLIvHgCJAi8YgsYcTn/uVQkAk8K9JJT45RVFc/9nXnPljaP+
dhcuqzn2t19F0o2IKmz3lgp0NfelvitD+UwxFULBfatJZ87o1IggV3mpItWHYzbUoHDLj/+8y4+v
+qd0ZmiENQDJ0c5zFKS5hceHd8fmBRjA2Qxktao3aJBFxPmuw2igY5wcsjnM3gIAWA1YrLH6uA73
iQomGwT6sfcy8CUFLfWu8e9qjqelkqlfNJphaNQThmMlCwy4MlMMmTcZCtPszUdxddSXFqW6KY6+
L3xkaT9w1UVS/DYMfDZtYdnPcCdq5+lgRKBzABVRWdBjOLSOvD45/OZzNfGgd3dMneAcuv3jkIvM
aAHbYC3t31tY8ryse+N9daLBP9l2h6KHzceozBIGXlt8KsAbeODrhWOmn2mjENh81m4axN5Vt81e
bpvCrSrdnVLHo2NI3Areh5l7KheYoAokZOhvloaX0yUiEr4wn5bbQ9bYuohJLmaq7pb3rcR0umBB
uz0O2D1aIL99own4c8MOx2r+Nj4uTfcJNdLGI/uphAfw8xffC3lsc5bswM/fiPEgYy1yxZ345GMo
PmqzZmCUWkaVcGZTqpPJoccePprjrk052XAScq4HiiEupBSxVio5UA9OyJMu1jYFdxCWBhcL8J62
lMmnD1uCb9W0Oa41UMASkfkMcDUkIQcC0w4CXO4/i9KgftHkh8C2j5EiQnuv4SeQM7wvpxLQAcHI
KAU48O+1h3SY5/8LUJTPVSzhuPi47Ak3ZktE5keEUmSXiZVR1QdTrGkIA1vVkC6VQ6PRDfPAWEeK
cfFS/oRLMH+O9bZJXRbiPfWmgtMlfDZnUwoFvrNrGNqFi6gBDV/dtC39xfAwlzbt7SGv3ZIhHUNu
IeWSifBhGty/wTJ8ZsGi9/U5CtsxNSRGQ2oCZJq68Wl5bp+Azc3+lXIwaxNfutGG0NbyRiET5Y8P
5cSO8ZWzSTch2SodkeszWKUR2P3dwUZo98m5QDbhZkLrd0nsyVCAZKIZ76Lt9pNiCPbazHNzI+NL
PQ1HLUJ/kdQbZPk6unW1lA8Emp1v46G6Y0JjzuYKLet4KeOOtzmhC5s+S84VdCSeTaaJ/d2sHnjG
EATijhrBkjnh317hdtnTA29IG/krzgWtZ3l5U7Bm0BpPBn/4mUYCQgWv/yTtY7wZCpM2KiU67ub9
SuJsLe1umT171fUuWdN+jyMGqVE1rcfmrg21swvpmL5JGuElG04z/e9G/2NZBagxWFYYYJFo3n66
k0lTkEjXdZWr7MIa2ZTrB57CksKMoR947T/isRGi9e3lyubuvd/kPaufn/4wmV8J/A/WFuKjLiXt
cjzeDbU9szit5WPX0CjhodidEQRzhNK5+zBuIndDMEb8PlHQsqKR1Efq4z+B64uUuPdc8BTqL5L7
0MTca3BL29+lrRgCCQjpLJbGUlUT91qP8H7H2f1uAjjvwcNyIH8R8A2XbaPRjEOpV4a/DBr1OdUA
KoABnZDDDcUqZxsSRiUvQ9mYShj/Q+KGvGNKeoXdEdiSGhJXys/4zOAXvVtE4IEr8l9y+zWa1DtU
shvqtCdKXdMM1vWfmMG3lRPlKpNnxDiZMCLKRD5Nxh7mlg6TfbwmbMZVHCCpm2B1XW9ed8Y6d94M
2rbCJLqdTJIZliF6X88PNh/98Yem2xbfXRUshckSIA+7NAEnjiVu5IWHOyN54456KxMAJUxn2nkP
ZMYZi7vm+HeCw6PtyK9M4W45mi+ebUFD4Hko3xc5c+hR3wARn3tCEw5X1hO3BrwFEL7cZbirW2Ug
HP89R2fAD94m/zX/ZHTsbObkV5lx6cslEtFNu8bTPdHMpJffbLX845TtrDAQJHW2w0lkn30dSff0
hKhbFVJX7UJOrjrjuCg70clre6w0fh1YYp/f46rngvr5b6u7LmZBY8lwH1WcrqovkGGhpDIhyWJu
o6MouKsaATIkGY68uVZixrSNLuU8n2uJ0YVN0IP4BIDi+mL88dIko3Ex5b4xZpF1oYc6f043+vBl
1fA+PDMhr40rRvBuWOHICmCDpAJhlbquFM4XQjEBFHRa47UtKi/qfwF0FvXER9k9LnNxblTY0Y/F
UTYrJrAYqlx4Js+rHhGwZiM/vZyu4Vz6seIAoQY4JLm0kRjRd1p6tKJxep36dQfPioo2JXgALJ3j
XvJyM32zcyx5IrQyGtCJ0UHy6pQYKsJVv1hBIGJVAo4+2PMQQFkHf6/dECovv4w+URtdRvNQAdTq
9STIb6DNC+LPYCMVwWN4bqePgeANt5HhuYoHfpmh3TxntCHgVXQI9dCgtZkllVHqL99s6K+1ZcoD
PcwcVncSb4cKluEPHT8O1JwNhYYDUmCUVR4dsc4bC4FiW0Fuq+gd2V1eSTwVBilzOYJaGLXB7+ph
y0ukhIJvLCVf2Gl2Idk5TDXLtNE2AMV1V73dzUT8oCE7a3j/LOzY7vMey8aLf2eIOKUx2hgOvbtm
gwHv80/6eXku5fc9BDR8u9wp6ede1aV47ly+DWHz6E1MhUZfvlKIEKnOrBC5y547ejwKB7+qL4iX
/BEIKkc8GMAwelSvMnOOKTSKgFlN6I7mvl4EA4S0O0ymiYFF8oDsOAJuF4833B5Dd4u/r7V59TSp
Bc1nvKzSiIMjVa6U4/RBZjTovKkNoKf6/DYoZJGl6DBXKDh68d9pIqf/MHQVg2MubcoEZGyxFuK8
Q+RqhUDWS1DShVJzYz68DPu9fGcC/aNaOl7YTgIbjSNaoQ3RwERTrFHXkDDxOZzW9t6h7WHdmPsz
nH25RXX19+pdFGpcSQv1bB/Tbau9+xfB9pZNRl7XnOP4H14hz8OOA8rBQbGF0V+0PJcR+qIMR2oP
jUcOA7Y++2MzcVwrzXbT68ZFx9Ci5arEEgXsZg++tVbb0BdStvl/l8P9i4G5S7p1vVpmXe2W9lyP
FWJjRZcllZ8vIZq3bURk/LwFWacCEoCIf2BvhhML3mqbV1Jxrl8Cx/l74iRR3I+6Wue3vqsPd7a4
2/h+BVSW0m3oxBZk1yuo3gFJvhvH/pJ2XWd3xZciZRaIP96zNHIlyWCHnDmwl1PWzRzQjesoCa6+
ThErfWns+CrzM0JNz8mT4bdMtdTGNI8iIpQ6A6eseYCEoH2lNsiH0sg2epPdwrbZnz6OkvzT6haB
L4+G62QMuDNSwaq216JFF+teU/uLDw4wvp8fhSPJDXPBdRpffw1P6wqqnA/L+7bPI/akaKYTR9xP
cOEVW9EVoxbgVmWX4OVMlwshWiou4OEDINt+FdF6aSHkpqqUYo618DQC+ha8Tpd+pHYHEs6bEE8I
5stkQXl+rF9bL24WBFaEDy7Irqnr6FXgZFp4v4DVodq84iNuxQROPSE7ELQYMyJO9RAU/xynTorQ
3QX6cDH4Us7m/sDfhwBcg5XL1v1c4bphgC++qYeNWiIaUbg7WOAON5JyfJYq49NvXS1LdJUTLUpn
FoBOqoCOdxMzGBOgcq0MEMzUajelO0yL67is2CH2fRsdk2JKHsF21TS9oo/kxULOu3qYwFj1nVgB
bn1TIYm7cukyNKnQ6PyAVFkJQVy8ijfjiUuTOI4nMNFhaFU8XYXdWarMWFZbhLEYoDs0wFbuV97o
UUtt4qsbjqkegCEO+eGzWusfu4n9Zte8Q5Lb2GCjqhb9OGm5ZtpmxdHbyHbu4PPrOJC29ov9iI+e
qRqmRR2UAGcwI/Khk6jnIymwo2z1Zbj47cgoAlXb0uTxNBKadAiDcehB6h38wS+VQgEAkNHwdE8v
FsDfFTLx2Wex/8SDuz7e3lgZ6k4VH+cPeToclbDD7THIU2eKVLFkrDYWqEQlM2uacr8huqbTFj5t
XoxXbVMvI3rS2hmj8DhZpyH2PUcPcxYwMScnsnp9A882YaQtOTloqTc9epVtbDPvgRvBOZkpHR8t
8njOaxoJFgoQTEYuWjsv/fZw9JtTeLr99qNZXwP4NaLoEUEC4wPdIOuO8Bj0NJhtYHvCk5P+dk+9
EsPzHSJOFOCT1dsnYl8h4+njIog95P9us4wCwcFJoEDGOr/nslYzrfytiRtS7nMUxrWEzlcoWHt8
jprVOusw6KPxGlX1PD4OlXI5xIHQY9rHFvMaj5N0WvWXvKcUlORwVmqkCHLn1pBWGeqICah0a/Hb
DleCElWFy6UbKh0c+njogLzQ4LtOT/0LXTfyTdtJvnCD7O3+F3RdO3urStyktqn/ia3aTA1HfZhY
o+RbqZX9swTtKDaah+famnvoNpAG6KMNE5xVNSaeU2KyzzhgdK8QMc/JcnlB2phi55jrvxkvqWfG
1sJSnme5007Z/qvTP5AbuDFTAMFLnipuraWH5dG4Pdiaru5e6q+mA2vNpW6jldu9bA6eGjUJUQgq
rrGvel4AU7N/PwAghoAq9RdjlyhfpJPVAopzsOu0NuF1YS7QPWeEwKjqTTKST1S/5Q26aXx/R3Qx
qd6nNtw0t+l8JktNNJXOb0RL8CGfIrYk1ZBiCH9aDTLT+e4G/TYNEUpDpT2khpaAtSkz6E3X/vDx
3ZLQd2W2Xge+Y+j45+XM9/XZ5iVy/KjEscC/vADmjlHex8JtwI4gP5WcUvLqIYYq1sf6EGF8OKgO
aiSdudtydZPnSnGSOcfTw7s5QmKjEuwnquYNOtCc9H8KoHF5tPuZJEgteqzB4SXfLLNPM5qfqAT+
g+ogZGSzv0kqimkPVRsNbpwMnXJuZ30zjIkyNhBIkGb3paUWj5VQ7p5Zl+zTfHH5C/49M8R/Bx+w
RumWQxE3LXDfzrMoHoDrG9ZL8ke2iTaBEXdOXCNi3OQz5IfTgtpfpFOaqk9TUvxhvc8OU8mEbk+j
d4FG0LkOl8kFDhPKwLOUhFnHr34o2GvHP2Pd6wja9jO/wjjoGfSDFo6itycnabpveIwr8rPUlt3a
VD5LtO6gTh3fJ86j1pFa2VWGkDHrecnVlpfZHcA50U26mSpd4TLQpZPubNo/bXFDYJkDMRbLZKc3
ejn2ts4XNZtaZ9IwfdQnOXn4gY2wazmKK/xfMJlGpfXZcPsRAAGalLn4ZfBcY/Z6ycEW9EweCaGq
p25Mncr1+r9cSfVpdMpikHmvCCiprhAHZqrvGm5tu0P27mqiibUczluBb59VIApTRSDI47c7A+zn
dBrfK/vXU4gOCvjQvPRSogCdol9AHKCpoPPLCedaNjLgh4xy3JdbXkBxejCrIvcmw45bMxNYZLjo
oitco/qeDobWzpawh50cYV+QNRg4uJWBxiInKsw5PcBn6UZ9FhgcO+Wr1PbFazYQoFBALyL8xTt8
nnpa1vIjMgv6XiMUwKGDJQATGFMr9g/94IePmR0imz31osithJttn8qVl7/IsYIgJTcAaDj1ZZd5
TOgne0emGfKxUWVNGKtqvl3U4GvWvrllgYdgJcNDPSnyqlubO5q2/U1cKQcM28mhSVK8pll35PGk
4J44cout4HBznCC++xIQYZZgx6V4Z+bEFGAYD1wxfq/rZIKv5hL+La0l5CeymS8yaIKG2qo4VmeK
NAw+4EXMmApktkv9zzd5YA7X0AEX4w1OT5sM1tixltpJPuQgvcJ8X6P2VCRrixLbrMcn0KD0GNRB
0ip9vYlBTFmdzQZBntGPl+LYvQla615GtM5XUnDb8seoJrU/obdQREpZIF+xaQo49s4hcJWzkmay
O4ZBAusTWWsxFEZTAI1Sx+PyosBX8Plv2hGriyvM5wuCfFZDvqM/H8B944q8GeLso+czzBZ8XrEt
chmPB5TdOYwxKFSAFrHuArxLxtT40cEzLaU9ETe3E1oluJnRg42o/V9AIs949IZ3HRjNXqLQd+5h
cw7lkCDoUaBQsk7u970UohNZLMDgvS75gjpybKAmS8zn6ROSd59nobCMPrh0jOjWXf7xQb6DgLmi
uGA44h3DK26LoUnT9ZXDL881pMaq82QUB35zRlyBRzIecvzigVSVqCEFPealGSnoCbr2IRES35/J
Eo7wDXB1QQMFaWqfbNuzi0ejT6fzr/813i6QNZ+82oLUa+McuSxdARLHR4FEDPSrpQu+1g7DixCz
jOWCDz8B9jYCI6wHNezkcIhcpyJfuMj5fbSFPTQ2OCW7qW3fGQ3u4lEmWTMMMKq+ZDgjeUPkF84e
immYvaB6e6foDbiPs6liOV8RYJwWW5bSTP3WZcR5btazKm7dmmnX9Va3mXEjEgMi5GXB50uP3Z8i
LxrNrbJfyXF7pRO9lox4/WgvcoouInt3aVw9hn/O1O5eSu2HoKG8of+HydTqBhS8Hsgw0AaLtq9M
1hTlv+Ncxillpg7Y5pe2HKbDhlOBV0V4ps6Zzxt9bIn66PMSDFH7ddnzC90TMcbiko9yxcZGNIz2
5yz0eP2UjSZsDpKzz+He2xgnD3OHhv0DyjQvh1671Q9EyLvKCICApeWOJwoNRP6el0rXx8vtPDT1
pq74epgiI7CNNopGO8hApJKxw9dYtbZmKm/YK5cPDyiZ6NzcE1dXmVN68wg5JvQqphSIxR76BZUA
t79H3xdrrtLbhN/ICouRgZCEwt27nIEFACnBiDuFmaxDsHDJT8mLr8AZH4Kn7qfSTuk1NyVkNEHd
hpVCAurWymjhZwZk/cFNisflaj5frhxiguyhfFTGkf9NdxycOVmYAlvKfPF5tjUu2eYjUPCQI/d2
wCLvHhXHzUtVpR4TN6BqdWdoeM6wjQl4BCvJUNHO4nqiUClGAF49oQeHbC03S3AyWcgVUwAfUH9n
jEQZ1f7UCAPMsreq7NGFiDWcs785OWSUn1XlJTBHGHr4FyheRBA4VCzyNaaPHOvVNj7HysxSjUcu
lAr+KsG6FWqnM7JrA93T7EX8Qw2nNC1fS+qAiOEL+CfMuSHlcjLnvNJdCQ/EjwD7QodyZji0C6l5
F4AGf4ZLP4gBGcZp6U9T1fRQae4rN9vByYCtEp7P/LPhPyxRrrQrSIS+b1Kw6d9DaKK9BEqtL1wY
LMj0O7iMvXCLv4As+Dq+6vRDVegvszi4EpVEbFZ9P8RkeUN8u/4wwss5nwzZQRKyWOit/Wz4QUSk
dQAQi6hgMOj01iW3rswZLXmZopX+Rs72RHxlQzQYUB9MxxP4Zt79FAoU3YtQq4tEfimh5FLC8Nhn
p2bLGq8vPC7x/1osieh+A1Yl1W58dgKBD+78ZBbnLlfPgycycS0GxT1eVNcJFkxK2zQNxxFdt3Wi
6lZ6dtNVgt3zyA605Cc6arH9Nhc5JuHs2AOA/1G3qdZ4aShiyHqXZdXg8lTl6wICcSFCqJ3Gbn8M
3/cU29moXUhKPbUEOF4Z93MBn8ZACkj4J9i9SEinn3K6oCljwyb1g+HBN2qbFpwc4c0hC1kCFvkn
sjVDtM7MdKq92/1O+Glyn4rgFEPgKQ9N+HhvVuqbsM4JF4hXc+25FVoz9if5ME0bW3z/XnOleCkK
x32V+M7LE0hg/Vzg2zXg9SdIPQNXCa9qDbIwBcvSu0ZxXZLu3sMKju/mh2uO4lfMFBROIzxlLJiR
LWCY00SwB3DGNxQfserS5sWJUz2N2/1I7URymmn29jAxC1fOs1rhM02Rw/X3arnSZRPoSJ0UkvO+
QOPv9HTEfUxn/Pg0fnm4LMEGVcSlHlbsrbgOyQv7Tc+YPKsaQPBZkpN/xK2xC8Y1Q0Z0qCiaU7Ym
ORfYkVSeZ9QfsnMkBp0dgCdV5OjcaC6t/9rqy3fPKQ+1EoV9wBknc1df8XPjR9pqxcW4tLc81/LR
cVotuK+FhSuR2Ve4Y0VIJgRPVZTjcD9Wb07xFa3Rw4hNy1AHsg4lM5v4aA22vy9DFtk7J97L3NCb
dziX/mPMq7T8oAZeiK8Unyh4bvAJ6Z85G27WiKZ8HTTyrXJ/jvRLEflm1IXb+x4Z4DceyNynykMP
yqM1bWfwAxU8Pbou23ZE5R9QtARsvRvh4B+HcCSQxXKFW+8u9O/zSwKLAdpzzxFZu3XJDdguO0KI
Vgx/eO+MYPjOsN+BguZIRr2Ky1yopBuq4AdkYx+F0akICwfgj3ex6JBL4fSAEjg4uxjLPyf+peQJ
91fH7dlkED3fxQsRMYdLRJ2riddFM+/GoBP5W94vzAD+FyIJG3Pdttz5rJw8Oij0UM8gO7TDSGYq
XsF8V4opX6GzkA1oqG8rSea5L6WNKRCVk27B9x0PNkPclGAiR/LBShW47W1If6NtxvWfOEltWXfD
ZiaL6vzBpkuRT9mG2bFPAztQ68piuJsJ4sk3NCcnIgEpIPOBOnC2Snz9gfUX9CRtGjWujQDSSEje
WNFry1kY6laM9X1DR5CGZhxsnWg4YfKubtifK7wIcK1XcQM4XKuA87Z/+4OthZ7jdQfenrfg3hG8
uKFxV0uBzxbU2QhtCVK9x7NBmWWVojkB6NPCNmhLd4dzkXYZNG3bjQp9pOETXH6za5jlJK7a6kKt
pLe5/LSItIXWG1sikTFMSqP4+sKKXCSnoTAZf4B/zP1dqaSYpkJHzfmGGluxOG8ePnP7/fw1jPk4
JezRA0Y5HoDrYRyN7ITO6R732QjkVzwiK/sF3n6f7Ggx/VYO6a154om8AQQH8ykzyCDWL9m8cXLS
cYce2d98t4opywW6EHpBCrMYgxcAkeEaLpTkR2bvhfY2qBMNML9MKUdsCuRuKDcG3DHH/S8np9bX
i02LcfBgrASeqD7iDbysLZpgabNCmZa5rCJudi3G0BsSEf/CBYcgapf+sddhRDwCCrgaiA8oDfKi
x7VmIO+2cH/VtMd4GqVt5Ag82APX2xXbKp6BzNI8AyYx/5zD0wJHezxYI0wiMJyGZxNKqKSHwuwo
lK8P/Fp4okCaMcXZw1mQkQcK9bEkXqG3H+kkVyYb0kCraEQ3pQS/8aGade841Sq4DDOFoObFTvSv
0ak58htyXV7kWh+O3r+NIuXqKNeUHVBmh74ZMdBv1XZMvdCM+CIRGg5IMbrZEuYrjk3xytKR0WW4
lbdpQkWam3ahScaJVOE25LGgcsiFYE8muIHyqq+twBuulo9tvNw5BNlFpwXCJQ73AxLS3hZ1upMl
ARG+X9axv3OOZVwxItrWZcLdeuOSrXKQvSJ2YyjL2aGCiT546dC95e/IYU5yms6zEUBFgAXJkMyX
N1IoOjj9lTyiCbI+0xdliEe5r7smBC6qEMs8Y0oM/c66QONeSMbWrtwY/A3eahE4FZbe9bEBmest
5VXWbE5GCf5cwCOoqzNZODurg+cYQzviIyaPxHmwEz4KIMb3CXfkK2FMxett1Dqh9CmZVGcapSRC
rS1of5r8yEwZ2zMCikbsXXF/CyhikdhXIbyU8vaDbsBUgoc2Xaz5s22qlhRYvxjFB8JUJJxDU8/c
YEoFg9VgdQlL5T7FxsNm1sUzzDxwMc/d1HjOr8Kvpt9KSgvF9FPROILOlZlGb8g4WCk6Sjq23Vnc
kGKkw9c18peFSYW8yyjxwLnTsTz4tGF1hyeYePrABO+t9oJ6bdWMaCxTgKWoZoJ7u0jmj4QGOWjp
ajCbryUF4Xr1tSDWTtswzyHkn9glzuC9QTqTZxaE88JRFPHWaiCMXSnI+ZYaAzLtZ5+v38GQQtcO
yIlunlseSCzWztYwEKZMNQMGGc7D0OCtP09c0LODd0XA8zENQBxeFcR/P5OU6IECLjwsxO7gzqn+
I3t5FNT3AxzisXmvG8i5+2pWsSMowgYhU90N1+ZsRNUlJ6xHJ7pTLK8fFYve+Mv8/z/qZNSzDppv
88wt6xz3yCyeE4ygJn4TN1MVFVCfzycZqTgu+aF/ZgIjsir2qozmYn/NLFgUIEvSYheLznJQnvUT
L7YtiVuywKDXzoh4rjkRg29x1Z1K8LEdxOutjR11sHWKEaO5rufhlrzIMVAdx+uAL1seV7XACrr2
mIU8ObmCnk5hhu3mRVbgqIOPyoTRbwwi7nmkHFXNSqbxcFI68TFuPJJqOkK6we4HJ6UcuOkOfA8V
SIcBCFue4qQXdciQjYzO326C0z1q9cb+ctQGsLk4HTvBgK9DjJDAg77shPyvUwi5M8RM0AMM4NJc
qhVNUDh/VsqQzDBtrHraPA+ia/SESsNwsVCwdG0wgLijZkeTSglMI1s4SLoM9xWS3rbintC38OwB
APxrSaduLiGhljL9/DTWX6o7or9ZTfAp5ctdRDLyVzMT4DdkABaKWz2oat3NXwI5nbVlFIsu5oca
cSgwpqH6OGw993/z2RadYwiZQpwbHzMNK+z6MsdL7AZc5PF1GgDqYxxDUOYhshqtGqVOaWuNkLOr
AQ2AdSVY2QoTBLZE56cxEHcG6ASkAxCXaPVGmezCzVLuillitGiK4ZWUVtcxL4E6W8mfrFPedOFZ
XNN4xsCxKQTKpiamxJiT/hsJtkpwvJCzMkS5NAopHqvi3wDoqAOakfkPgXDSip/Au9CpCrb3tBR+
WM/Mfjc19ijZ1hvMhtWVSi+j+eRM+LFeXroF4cdqc0pxVm/LF+tXex0o1ShMv7pXb8QWABKfPGIV
iXanCoYPwn+8IVbtcRvkeB+lBg2D0YWtlFSAYHvs2GCxgjVPuvwY3gMUfTeZw88eCvlxwJszx+AL
lyXiv6DHyaLK8v+wRVbHMqdYgEJw30+kkzWMpaErEH5Q4s746Z2A6ot3oUXOhNcwloEyopXFIVkR
FVv8qEs8Vlo4i3yjFxsLk92Jq23ybHc/oDZ8igwyrRwm6kxzGSxqKBlRiD1e1vX7+3z+/vdRq3JW
zlH/mTySkFAknfUFDmFhozQrvIQ2M9+qEr2GvlpVZ0Q15WzDU26JHbDaOZvrQ/BskJQs+8Np2fJO
+yqc8qWVz+QHGABx+kP6Aeu6NVzKuTDJQ67GBNPMBUiucapksZTLMOEugd7UpPI4zQ80HSiaMBcr
RqAGNQwljSwVZhto+yvQp2PPhRwjR8isfK8KzZYwFUd7nmDnDKzoJzGYsFasLIsxztKtwzbilkXs
nn385a/2VkeaT2yrHtpk62ax+/bnUglE/K5VEY02BpRwLoKd7/CQjxu3s5vPcrxmYCpsvX38ZMmy
k6Xs/DP901ypuMrEgEcCHYzWUCGveGzUxzbGXK5BtVjTmGezpSyeb5m0fn2TAQXBGg4nRHPdDyYm
xhZxOJqtPeo7gmp78BozRRIT8k4Nmx8Ta29JwAl3zK5tsbB0Zb2WPNETIHhrRRkDA3uJUWKyZy6d
DQbJ/Kt4AvLICvTGFPNWfX/MT+Vddds0YHoCoDKa30LU29d/PYBCvw/XH3QBHICe7/vidLj1lSHT
Bs+/JWu1caFWfyL5m+9L3J7i2oF8MYbBNrmYL++TR0t5sKxL/jEVIkqbQ1CKrdMVf3Q7KigsDS9H
SHyTwlJafCq/ESKGB5JkfE15LvjJrbJikopbA/90O1M25pVPuFxBTrS3hPUe2hDK0KwqBLIwqFkt
a/clSQ48PPxf1r5eMr/iKjRvamFj6mJNZNO/GogItLRJPHJv9h15/Oe1GAAC+ExrIYcr9AWSqOLi
1YP4YIefKmiZ/LUMrpBCfZSmQWvH89CnayhDMh8QtSVQs9Xi5+3/SwXpnZh8jSScc8qVVhwYOwJp
gEjg5vhzB9Xg9+0ZEVF8P48pyDcGg4xmuGABWPSArX8bafO809Cs9v8aq1zI06mHbN15vaF7WWix
x0A9TocvvGd/CFOJh8bkzDw4agoZALio+K4dYV6gcQFrVX9fEyjJc3ibiGbszpoGQn3r83FPrEOV
AhGql5yJiT9laKTYQWmyKC/+ZJxNoZDV7cHyJAtBzC3TwNyMXnaInWMRxIY/tvJ6FiMoqn52GmTo
Jzz1wpm3mtSh3HSN9WaAnNKBpcjw2UFUhAmt7mx/wAkm+XkZWmAcRqqEpMlGP4S2irAWd+xnAzu0
hwh/safOE34amG/RUwOuRbv9bvKMqT6+pJMuiucF8u0C8W/jRPJUJdI6TlfeU8h1C9no984rAEmi
kNLOccnvfndAjiIWZvOL4K71AHlk4XIFX1aC3Qsf+CjGdzTD2bR5IyZMx6ANRxNFVOxI9MXecQL2
0aQ43Qb8UuqUnZU7RaaulKgMSwtJhkoeaUSQ1Z3eQck/wppmLM2IAkRgxa6DX5ps8obZQLWOdFfp
8VPra6imaSC0giqju39Y+Awa3wSqv8z9jB6pe5uVGZKeBUrxoiK4XGsG4rzI0D9R/S5SV09uF//m
2MlnuSzk7XdUTYS4bxSknICRr46Uiw2qa7wBSowGvpKPq93hWb0e7hg3ry+j9Wq6wEjYW4cQ+I4W
G35HxXI8yG0l1bwOxtk41vYSnkCI1B30x79tiRqZ001Gr5BAJBngEUTrTPjXQytpE5nU6JgBwNc5
OifishDyMWujw8sdKtXNIRAYZ/6uYVLXzquuwtxnzOnMjIRCrXXNDQ0seaJcVa/o735pThTyKU0R
TqosSh3g4jMzkQvTQSzEa5r5+ax55uoxoBNC5Z3MpbJhvKQB56681L7XaOL2HnGZp59pEkLozIZd
GgUyte1UE/L6YylfYRwXSg+MIRkdk/CwbNKraTW/kIikSww9lOEWHEctN5yUmg1zQRIfy2RuDgvO
Gqv7A0ubpQXU13fhJR39wSyESJ9IdwdHlyxbfsUOnfew1Ak7bvRKrWiU6t2IZDfoeQV0V53ETn1p
H7fOeaQK+536g8sEUMi2lzMPSENkGAgloZN6lECozKt/yCKZ7xYV1OxKi3l8eD4ZtFVBBZ6C4KFA
V/ofVFtMZhQCP84c++5UPMa6l6hCI1WV+VsBkFGNr7/hN6kbwPAYLUiT/GA/Sw4G9sbKnAN/nmL+
Zeg7/Ux3LtOr7rBgD94NzSw7E/1vTNP1h6uvbZPmFCfdxT2kNAqTrbBaEyjWUejpLytQycKqHp2q
Bhb7zvNT2q3MPAmyOgBS9FmmUjmFKOlCxDq1ysFwXx0d8Ehv/ue6vC5BlPRyGPp4o+IRHrZoEdAd
CVNy0AIdgKw73M0sUYUqzqoJz7rEgdlTPfy+wApTt2F6wds2T4Q//kWAn3UbUymzFxISrQQgEgmC
2YBUxzFkq45CPZ3vxUPMJe+8S2D4yPhwNsHy93/gsHACBiQIxvBQcs/tV1m3+BsuGUCQ9Ljv3GA0
qxtr2xaCDTay+TqTqFP7nq3bMw7pAojzu+19l46fCFxl2TM+ew6Fgf70OYYAyUkr5QhqGfKEd0/U
QxgTfgn0+8n3OuXHgnCVbNwLPDPvFHFyRBKylvA5k1lq4FByATUl3aIqZnOaE+nSMWeq/0LWIAtq
hP8ibDZz61Iok9XyFA4nGzDnUivc6AEeto/FOEFOvn7HzfttH0l12pG8FUZGKAdxZ4iG1xkarLhB
kqBZANUcBuLfqW35HjroLxm8Z7A8oQORNg21f67ACI6Nwiwfa9tUUwjDd/jtMj/Dy4XE1etYVsi9
ftAeO0bQ5hJWThsXeWbvMQrDTqC+MmBOij6mHeLciLb+PSYUbv0l+tn/pPWgQb5VTxMloNg7V4o/
RSzkMOjoi+2hvRto00JsLQqZXgvVPnWg2ivOtKHLdrwtVg1pCkn96iJFElrAIfTa+CXQTqrKl5jT
IX9dI/7l5Kf79hNkQVjRtRHfSCIirIU+3/8mZS/yFy5CLpPx8wvlWp65Rww1wx0HblD94FUuxfRc
3hYkjCdjSj3yoT66RfqTRG44rtB/gJvDXkKWWDWqxqzKkokSLizxf1wJlzan0PlWLno2xYvcmNk8
Gw2JElbPz+xg+U3ydORzTv24XkZ9xK2x3F6JaqPzjceGD4t5/dxjfo93bt3AsPfH2eTYq0XqkC6i
U/ddUMPpQikrfF5i9FS8cE0TV+alSDpmpGytxiXVkBchcsThnppfaBpj0zK/UNbTQqqhwnnIBZTF
dkET9z+xlZfO3GpdM7XB9IScIzlOTeoiLCnFB4R9EM8+r8BYN+FNzKVaJICUd6GKv5yBqBTFh9n2
BFbCe71DTPSq37Xn8uJ0VM1RlK2q/OFVbFax/ZACuwq+r3NI4WVnegvxDN0H9G3MQ+VuZ43cZpJ0
fxO1SbQxWuMukl3qkg6ERDKyerYTVftZjntZK/7JdNYcg7Gw0MP9FKibNpm/VJKFQMCLIAj9aOBG
/JnFXJZVHViNl60/LOQ3igUDQuHuYz5GIzB2lvyneGuBMM20fShSlRt4u61Pjw+X/8iFrlKGg+pT
9Vmk8b7hsFNMQXuE27UtR9eGXhVXZRl5wMh+O90nmDULfcFKSGIDSFrAAoRDt5AT0fegU8BUPie3
CUat91QKAMWmOvpZ1LLLXS0eIuuXMSK7hC4scJtCNWQYAb9zo4YZ4rq4lYHW1y6AZX+OKdW0E/iJ
6NZsvqWLj5gJ+bJf+FZm5I92VFsNoTec0A21pLTk+8DR9rPv+ZYbqTyIv4sBJhXrUpLKco7+BFa2
M8Oi4MVQlj+zslEuLZ5xeVc0ywArM1Ph3fq8zztvVgpjrOkHDI5T9QBNbwBAGFfAUZHAJas6Dko/
cgRmshK2xnA+0t34mk120Qi8qN2GSX8UVLWIb/mPc0P6bywzbl7U3Tic6UaVt6ejx4suIDi2Neqx
5gxm0gQZS1l4qcswO1pyZro4qSezmlk9Ia6zZu1nm4wOH+9usXfK9iFnPxf16N88U2A6F0MjMmDU
haYaPrKPCqyJa0Ezqewil21oYNVOOJX/7F6J8xyYBei7GxGAyhOoW2Out+8ZH9AQKQAFojgNZ6wG
0ogovPRng0NijOY6euF0HhU6U1yNDPtFzck8nVfELdyvNpi/CsScTwlhrzN+Nt654pB8vN+Am0/c
ddVnxBAbruIsWgV1qxphSH4qV2ejaMaDn8wgY8y5+A+zk1Gx9ku0IAffjTIJmk+lOdOemER/ozju
cfDOXnE9TyAJLtOUsYLIfmtZORfMRpM4BxQkmbifOemSXszTaKcdjTO8ukX+ZjC4fPZo/xanuhbz
0HyUd0jvDc8Ueovm2UhkX21ZQ66pFxA8a3Sh/B8mNU1YjM3fpy1O3ZKtFi6unvq6lOUZmu7KIZh4
n3zq4AkD7RVRN/n/XnSx8zRS0t79MtOs9dCrGBsukugsFym3Jz7JB+8nAmF18XJ6uU1bPSnNMq4n
3tHEtGMuh1xjxW4M2qx2hpOnrn2MpeGWmjBx42Q9UKTtCcIxhaxWDEkyw1faav989SzUC5VXx5NE
BGBHGX0NONzS1kPaiPg6Do1N7mPJ8GLVLmG/V/upT/+di3ZWBTKmsFxzSxlHT36swi7daf/u9Rhn
tCtKU+/MhYEfCZIUeCjMQ5CJT7vXjnk/8U3pkbLH76Df5F2RGqwg72G+KGw25ib1ku49oPIV/nux
jDWA/q8IcQp9OO76YBqt2uBDJSlRpMCQfJcw2oITcfMe+6/C5QiEc07TNBfTM6GM/E1AsQUlywrL
5vd+FvEyBsVVTjhLfqXNgWKJk4DW9w99E2DUmgvREuma2VaqmflwijRigR7rl8LK+P67oKFFqPaa
3Xyxhu5ykOM2spq1GUD6BvORdVVcJrllpHQTi8eE7PUm3mbr2uAigU1FPifO4td79UhKHYlQmZNN
hIQs7bXP1iqBZ9Wk6CC/fALNU5prNHMxI5uAhszwNmuvLa/JGzO6e2d4Sjh0RQzK/t071TiKlsuY
FrSsZ/LaehiBVwlb8Yj7cza5d+Kzg/XRJhMpmOuAk8RzzgZ1f3mZeAPDUl4K9kA1Yc2oCLBfez2V
U5JDvpYH7e1J6YoTkNvPguvdGQleznkGpHqsqrsHZ1MVsrEJr503veUdfpwnx/de04YgW810zIw0
Wbgdl3YQUqQp8kAE6Lhq0ZmqOVZRTKvgcCrSRj09us7QgQnolunS04AmVEkcG/EwQIoCzSjHSkgk
FjsvOo8srvw3DqLJoiNsKPbfdVqTUIXcc3mcxGxivS3g9NVwwcPSlMsidb89HokwgzVyfxWg0l3n
nGSkbwhZYoZPbU5ykCahgDcfbwiDtBeyNJuI2NOGzbIhU5NTX+IXHiZjutmw9hsl+Py+4uy2Mnnh
zPiU7OB6Wysmcw0Rb14z9lvO2NL2K/Fp6zA/5c+a8vCJ1LD330VulHrW+NK9Q9oNAnbjFETXvp3U
qvgDExIeEy3J8fhu4H4+Il4wmndlYCL1BBIvm7iqTSZNXHLNaWlngSG4TPt7HoyU/HmLsTaIDvGp
jEgdhAB7AAWHsce0cveupPeIboJvwnVXY3AiHb7EPscbj3tyGwxAQ0JF9Mn89HlGNYO62A7Mep9H
99jRwjdMHVLErplbAl1XVx48DHF5IG/hLzvZglxjKS2HLQHtpIczlByMkDazVAk3TSvV0qTCfrSm
PW78R1GvYiK3pFnsta/tYvq0LWrdYsubTsWl9z/8Idc9bLZGVmhLbeL3V0Zzc7rF70q5v1cQ0n7p
bpyQ/bk8Tmh5kj73H8NNaUP4+ShJK7fGkFsXv02KLW1FMr3PI8P/LY/xER0wMg0+Z2AwI0CTiVdx
MRsuWZiZ8IJSpSR+3RoZcDwMvdbPq4yUliSsNP+PRu02WDHrZB0q/fZNzMOls3TEghZwhL10zoMJ
P6fjpFBA0osEoG9c5CaYi0qrSQBfZ4MK3WXjeQGXoTfmKMF2bQOiNBkUZF8xZcIREQjlRwRMFaWT
fId77aj1vx6jpTVC0j/+aohMdS8iCKAyly80+zZrrZ3NEeTkgU9tYJSvSVdREw2L5L38X9doyQtV
st/RDSWcNedD5qHdCbBgy7tXv8tbChMQj95hFDKrKsRLLISNr44QxyMClCpbjHBIZApvSW6MNbE3
RaAgO5/LVepLmMxLHFpzAmTARP0WKN1f9XZr8L1yR6ntwaBaQGJr98gsVSqY5YPYKJcjD0xZOr5H
eRJaBcLoAX0tWAcHgj4QB+WTMLj6Dp0LpJcDUagl9ap92+sx0HVC39bD1onKhbt0oKxbdLHNSsej
P11uBsVVznhSzNG1RCQPHDnF21fQAI2cfMFZkYzPtRscNay2s9cXyhGpNBD4vEF5OFUumS11mo2T
fzeWrwKkx4xEMvO5oSV8jRiu9VuuH7UvKJ8txLG107vLWyGpmI2KFBudCGlMnWz4XURAvel1FyBQ
vocQS3kQjpYu6v4qHaWir38t+7f/fnfwYSlR+EvNqTWf0vYJu4Qa95jag4BYO17BTJ3csmS7kWEh
1Xr7Hxm/N2akzNrVksSmlX5gncerrPzqf1TkiFaVRXhBPNtfQyAoOpRydk79d0X5J69O/uDABkns
CucLRC4T5hBapXTv2C24FC8lNdgzE5fFy5XCY20h8XX4RIg+Y8PMAyFB+dv3/kbJHQW5rQynn+On
6NGCmqNaltG3bc36JhwvseEEEQe3Gm3DwPmxCm9ib4P9A+K20ykbV+HiKnNdJjl14PzCACSHlUqw
pPVe2lYHyMfSKZsxcdaFGPHLeKaKSez6ZskZgp2k25EBiv2tVUGE1XqsTp2bSzmhMStKFL/zT/JL
iBkSjr37VaZFDqfzeXFE5GACOB7FZLh6GJ/vGXDLX42l78fRLx7uqhdbelvqtZJCGOtkyBPqj1eK
GaZNQInPduMl9VAQDmlE/b3ODf58hGbzkqgMmTCiVw/6rT3e4DhTH0RXkPHbmgTw4T4wGSkyq6eu
O5XTLNRYEVFd9KngOPTa+naLya1gpi7ZvOwrlni1/bOh2SH6FTKk/BVdYCB76pNYnmtY7stqO+lS
Fjl02SMclqzkDCChFJVmIQrqBpuk05ND0XLdvMAsA/O78WH7zHYXfwB5+hH1hSz+a1JaeHj3CBK3
tk0xCskvee8j8etW6Yiisd70srpywKtyDGcj7g+NinnQQiGQLO0wLNSONT6saj+ZZmUaLvrULuhK
byQP5tUnYWy3YI/U2SpnuXlsHGKNjd5zJYMEwShyhcWA4+W01YjCSH/aLth2HKwAx/I/aVJtcZmQ
3YJqHbVv65lToV5xznkgzFciCbO49lQk26ZtWVXKj538hMLm3CkO0IdFYYvqP2ghxdeBubEweMvn
gAEEuBQ+bVAMemfSGFf6O8UpmV2sG7ekCx+Qpc6bKxud8wUPT6Js4gmgdIX3HJQXKCZ+FtnLm2TB
9S04UpceZW3qDVGBlHGG5e2tMD8W9dzYP4zaAGS1DnWRSaZ6P/1Rm8jH32+lhNbPjCWFX834sL/v
qj87sbInNIaa0z1SzWFWgCA5x6el/3yXEk5Bo+rVURYZecU1uXeGuLB1OUi0vzGzviewM5B/8EPh
4USRNgKT1kTdmBd8Kth0HzxlmoKaD0cc4HHn4CzY3U+UO5ehToFMsltvcj97GkE9E0QUq+4mDxRL
2x/UxMa3HkS5w9YVa197pOCacY1JV0M0jP3zhfC5VLv8clJjIIUdGeOa3rOChQ6BDZBbMDmRJ/vv
M+s+mYkZBAS1SS3UcOblvC5fUi6/9ORuyoWSqSaacbfAeTF2MaftE6+csbBw5RHHA11HBwk9mori
73f3p8E6/nl8bIT5DF+hfMr1rq0kvO+dzam6uMKSYtZ0g4FKBmJjWioVtNAip004UI7taA5dQkKl
Oq2924t6PWrx7/jFc2H6hiBNT0hYj4NPB93I+F+sn8jgHd00/EmDBKD49qmyKIV3hdRv5RMU51EY
VJDy0rJUxxbd7XYXcpKRxk3gkAzKTRnC/w+QFozMki1vqSrdo0SpE0bStq2vtJcVsNiAFvKAWOBr
TJwyjiNc8MIRabWw0QYqANJYAUJcLf5tBpmgFz9aNTqDLV1FjBcEXOJwoFn3HqAngqUpBfjf4bTo
3xAGM/7IRWnnVRMU+DxyIH+JITY+iB9ICZbBuC8Luyv+41QrZNVJ1Ql4vD5kttj3VeSubH5NN1t4
jZhmZevGNCUQ8bOeL7xsc6UqlKrebu8iwWrajIpkIOCdrMuFqKBIoBuI0SsIeJEeqjrFnTNfgoYO
xdssrPDxdeRaoxJqup9TRC+dIxuPspOeQgPok7H7pnfDGZzx2bfc0ZB/u633RNtVb2rFAgVcJGSd
pPMFFaLXhshiHSTMaRtYQ13u7CHzLsY7NbWt/2mFn+iHLufJ6cZhvQGsXDDFguzNaL4ZNvTG/BXw
6VpMrqqBhG3aqsqYdSr3pbZZpYDLlCPb7SLIKTUdHjtTMSQzcLTXWBkIFA2NYo1hnbUhLBT4gFvs
asgv/EQSrjvr1CEY3jHrH7V8z0bgcWbwbpOhDNvsRwCS1p5gtErWT9XhtVUFXaAP2WlXpKZ7RWNl
cbSML6RLsc4JZUfhce+xlZM8Vx1A8RbAl95pSV3p1fYNlS0MyrtUU+C2OEHyXh9T5K2qX7Te2vqp
dtvyM7tNZQOrrUMzTRwWGh3zmaH38Mwb0yEdWkUEQdOhjYB5n5iAsv9jrWPMCVfyfw0y7AX0ajGD
pE9Zuu8si4na8GI/6fMMxVsyqgIzHSGM5NXO61lR4oxxV2AG/B7pDfNlJnDwGFs7GMWzoXooyhHO
BeCCM3m1FMZWWa0MsFjZMNiab9uyPql3WcpQClLcuXa3AXZORUm+ZQEsG4+nw9GAyIsZKaaEtS4/
OVJ91pX4+UQI3d2WJollTyhQT8IqYs4j1OgD+QDlXxZwvhRW6IpseLOJ8HpTKzfLomtX+Qa9SJaA
pNXEccY9FNJn1Q0ceOdBXOgWlap8mOHy0ekabyrAbCstIF8YhwvlGxXq6vm0PEfm3WjUYEe56fHf
ZQa+uj56CeE0uvshKh3lexinszc9J4PBHUInRYE8OYUAyBfaXfcbsfrUrZqZOTbWvWt9PJiJqEDC
qdjJ/3P/2E0QJmSi0uiLkYjGBG6ygc0VaxnEvezShvys033GW4rlZAW9Eb4xjJbwTEekZj0O6qb/
SXjp3O+wUvnvVSbOltbkLNbORqFrY6flJfZBHWBAvNripa2xo8n6ntfOlaPQG22TnYI0ueHb+Bcq
4rEgfgv+S7ovUmLigjbA7Rnm1WCIkROJrGk+YRHgHLmcgJ18up20oQqmUT9qn2LsAbPE3KGmAOqO
8Xnbbq3ru5nm6OsU32dyu8ol1KhphC+JogX62n0H9Ovr/OKI4jeak/Lb3HRDC0aNc6M+BjDiRe3h
1B+dINTV9vr2D/+v7foJEbnewmUQFT0rzlOY1RL7grLQk1CfPysrKjR/KZsDlE4JNgLT7fKGk8k1
rQVcI4+frOX/nRuXkmfRi+e/D4W+YSyB7dc8Kwo9Gd/FJVlmzPWASfEaP9ITxyPRUNbxOXVBLOQV
sB/pq3lhl/1Hdm8JnWwZWVARyPgd9LmPQwUjm+/vIRLJUbWKsxyBOkxUOeY60AUuia4ZZ7b2h+K3
yrlF/0RXfmE9SpuCjyVYHwehaHDNysgjDhHPquyxgv9QomL/SzBELOawR72eiDHBscqn9Qa3WwhK
7ySDaRBUBGZMIOCYhTNlSmm/trE1LDbQ86owNVqOs/k28vdulPx+f7xS+c2oxLfvUhxj+j0IuadI
akj9jigxpD/EubAhAwBG0ZP89A6Dk/0z7L9GeQn6SBxnyI3CEBokQnh5a+5Ub1low65KxPja8cRk
FS2NGAeblzaK5YfnG/8u16MBRPF1tmhT6cTI4Eo6+6n3j/Ny+7LqjiO01JbKsiLRU1qWcsE7lh3r
lwn2/kDNhCeJ7ogoBge6VjXFraLougNKTl83GTO6BhS1di8dVIxpfZrG/cmED7wlMXeop3Do4RtR
DPLa/HSQWsipt8saC+MWGAU5xrLfAoE/+QFfpopWUUjjHIpYe7MsDCpVFYE6TOq6IEw82n08dagb
TxJjnoKZp+2/vjxoowVbd9LZuvHxomQJ5aqBHBg7oPhARHkzYBKlkVeHeQIBWkZk+DbLZ2ID4bQx
zV1slRg/iN8fCfOdiadj5EzAoPjheHjC+tA5F7pE21cnfEa41h6GknWsqOP6MAtEjJ75cZEG3XwR
awkqLPs2oYVk3pVSIScYcdIAjVC0mGi1Mi1QfidFy0RnZppGUtu0f8FoFD08WJYFok45CPzaiwcq
0qgt6XVJWYb9QR8eCECVqajB7y1uCaZheGTfm2UI0lNpZ+wU7I1tU5koU71hYPoV5sw/PUHc9jql
pg71IJG9UcLavl4pgX35eguR6mktqPf0xqtGsVkkGnjiN7ykeVMlcWBGzOnXlqeCHf3rr/v3HQYv
MnZcloP8S38Qv+eR7ga6kS0J0rVn3+ipmpvXBjCow+I0F5sEhjsANJhDq8S6Hi0LK7MihWfRVKFC
aFgcU7IuBfMYkAFqFyNUM/GBq+mMt4qatTX3e4SDbhhzWcWTEG3u1hmMlMLuf8eUhvEf6cpnBjPS
iqrSSkM4rpPRZfsCPAiMc2FXEtAglKN7tcaFSEg+lKHExI2J7CzVWnldkQW79HDZ9BjpC9lPWpzS
g6N2Jfrog+pufNU3BunQJHyddTEMGXSPrajb/RbqkRxPMZ96efm5Fb0bWPxL0WuMZVgIIbO/mayl
+PBGuGm4yk16PhkpEKuZAIWmCNGSo/vwjmfqYOceE0fVxygMACGVfXIc1NVdz54fYRb6hAJ3BGAZ
6+L11XE+t1p9dKYLbQLlBmoQ+0lE1rzZlRXQqJVb7uZCFxBD0msRTaVtWgqmxKDp4q7ZXZ9vNf6i
47LakIwyq56Mj+UK5ET05J45c6F6rP0pooHVPpfKl14bGfb6AKSi2J9oyQBl2JnDXxxBEIZcmsqg
rduITtHQgZv0rZ/AHBK2AFoVT5u6sGiCH4qGN/kG6g3IzxugahPgYSZgY1hPGtphEgVzvqwx1dkv
qewZnyLtkzR0BOm2Df8uSMrVaD6fmjJHATVKMKMT4/Rdy5m+PbH1Yw/03b44f8L+y7kkBzBkRL9A
uCJxCY5RYAXcxF6bAtMhBsRQSYsnYybjMsw6xxROwQ5Nj9mH9OWS2nHAhRxdVYi5hXa4MtKdP1hU
e+oVkQHndqEZlQPKiHQBhJPEgLz+i6M7q8MhSHNfX1NMg9xcr7Z4ZdMtSgpnRmWEb6i3RA63RwOP
4Gq0N9q7r3NFFMK5pJRe1qXn3zfj0NfeYc2R2wLWr/qUpBxv7NrLd7uGfo0KbYZSytflNho96fuc
Z250a9GgNb9PbnLDceTpPoLf7lXmDaVH9YPSnBc8MPxZ347497GtwzHX+pcrrnxVPtHN7if3tS6p
Ghnu6OjcAjHljxwW7l+tUrVlFrQm5aLZ0NduMSVDKfN0HedJprf5ItgJNX8d/AFtGhKpNFo4XBwt
angFEpxgYxYN3uZGdmJWrniQFfIXqXzyvR/UqFzZGrwDEW9+4pwYJA1EN1YKfYtVPp0+46gVkkTp
XlxV7FrIE6BUFB4=
`protect end_protected
