`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PHhkNkpzHyCJ02b/zcKKV4H67KRxpe36QtGSXZ4oANg/Tq5UCNDHZf3jnecctZQreioRQ/cc6TC1
6ycytB0hyQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bWdkQD7iXQyADDoBhEMorxDwaorw5ZE+71aQZ7Jppo6RMyIponN+UMss01BI1N2b3FJS4Zu3aLYO
px6cO+Vs57h+OQYvM5Rj4nWKlm9nBZ41CnWAwleG5eX8bZY42EI0UWD2fk3svZhWuYfYksxWdUez
7k4lE0NIPu9XIkcIeyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o0D8irmB4btVuZMHr7825UqIRFmxWPRwnlzuAQTRAkVGag0/uZxMccyUEuNVjWpjJLtX9sBqvYWy
icHrTQtTi0KfJrS8ikJrBTfSeheDRWxGwQbktHiSZlVIs9ZXDCQSHR9RLWTw+n7qd5CPOqFF2ZBz
CDIGHs3Y2Z49vgia3VU0kO3DEW2bnOB7tyT+k0mbUU9gtzpb2sMIdNXoECla96Il3oPqhOn6wnqG
fxyvNEDXX+9ggv/b3AJ8f7vQxhTiWZRghRRZKvz/tDenZJMI9gW1b+QTVFaCpXETDE3gVUMo+pDT
gkeaydaT0UUCdzbodNgTDg5EzKNdDk7z2pWJpQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZ9fmUhBpgsyORCOIb7xGyx21bVvbIGX22TkOkC4OYVBlblOkFTGwpEfpvP1tBLXeWHsaAsYDaky
+MMNQXyXlzUHdky+SJLxX8DromtiDW0Twg97DXw9QoHET/lH0ZfTOCzNqJMGsxq4/5CuYlwtSt63
Ens5BOQgrG5RRH4Xbgw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fgb81NiSq62dSzr2ywLopRavTEU3BAdPPDhwK9GAYtd64X7TbKUCX2vkWpAUxqNGlnbwV5x+UovV
u/ZXmGRsX+eBE1EPykp4L/3bM3DF2RydBDoHDxeMmK2h+VrqiSaJktj/VTY2xfqO+bNMcU39RNml
fvwPsqHTJOMpNsEG2KsbtSnC9aPwzo5OxbfrsYwLtETkRL+nMXUlixjY6elVH0lotf5n9KrLTEVj
WB4Jxad1k9nwwYOxN3dJ6njufJIBiBpOT8n8lJTiWbAdxhlaZDH8rzWrGbPsBS/2MHuGWVgaznBU
bEpdCIot1kexUpnYXmm6yrI2OYokdfrieezi0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20960)
`protect data_block
AHSHqOoMIa0thf4kqVQotnKCaCeUSG8FahuRKCbb/d+LtUBFiL8HGVeGX+MM/gXFLLFWOrDXS23+
ISZQMoXaI5/hHbaU2R3bID+XdP7Puxr5RfSjoeUIW50/7fTzKmma2XvwEWW1IGDYzAX5wnwonl6t
mavn4M5zm14RHSxh8KWymBM2vqTth0R9w3lN5ycFvKzsS3VykKsn/dXy5nzSiUemGvZ0pR38R+q7
X2KX+cFDgzcfOraZIXKniiajtIaPPhgdqRHZM3ow+4Ba8VSzfjEx7CnnVarwOBxSprvbCZ2/Hwzl
rjpi2VCpIseGSgDJqIbup0RA3FShHZGTloWiDeHgKR8p8KjCLqogPqKJMP20s+TstrlqbAtSRm4q
9ty/rX+4Vb84c+tjBt7swY2oF7XP3xNL2kxvs7S+RRHrEZcDK0FeTiZzBH/lB1dvMIBFR7cnEZhI
QgH8BinkWhW92vN1XjaHZrw64R8xDPZ8X2QS4xnJjwV3OScHRnxklVSugE/CDI15exFo0NQOgKUs
ZaprYTdalEGeOcZ1ajIrTR0EPd1C+lUN5rkfUvXo6AJ58D5JlIhA2rQHd7u8NaCSK+IJbeLhu2hm
P7LuImCG0BN7VRmditV1rKLD9rTGzqi8l7V7pJYyLBc/bEnEXQohcPwVi3MFO2DSQO8p6qhEVbHi
bG3ReliGce6Yw/L/JWclHf63U6A4wBlCPOpPIMLiMYvH9XkzgbOjsMTt8YFSijcz6jVKKUTqdbyw
MFlpc4MdXLsi+P+k0ue7gxeeYoG0KMbQkRh3nUjeXfrAwUm9vyEi4ZjuCgbAV7fH5e4bfl3YMwos
P0+npd0O7JZEZ0LFP9fHIsuRomCZJpl7+T7BRxyH8BTJP1nV4S6ymoT12czcIfXeCi4MQmVOLcoj
OTbcfLEXFJnoLF+TWnpzDk3FcGgIpUafVx1mguSnNnQ/as6tDjm61tOdJtBATzWyhTCrrJFb/fx1
CwHNJlqFuJRABiZueiid8I0jgTLdJkDDDodSAMNB9I+bA7YdwIZ3DScGpRugZWTkhOvZwNF3FfYt
M0ZWV76P59PXK6mXUy9SH85FKWNUWU7OJ7KB8BG9jI2zEVpmJV2ZaMQDJP7Us4goR7YCMAQZm+Lz
zEefScDKjpuhd9kz+Nacrp28wOkK0vfYuPYjbF7jYC1tcyvsi8MwZPZA5RsB8YL8Mu+vAvAFnWBk
M/brwsvuVMw85HPZ6vFmpza1mjEHT9UtS09C7Vh80qyH7ZPQO/gIY+jjIRgLyRe9QgA5dYCMPqZR
i2NZ5UxzHTTxFp/mWZcLA7q9ZD+iCSMoOA4q1fFv0g5DVu+MAT3Jgyx3GVVRX22GzOniDydiiMym
ogxYJiXalzh5x88oDbZ8DW27U1YsWF72Tx5d7HMJIeYvgFB0cCi7aWtAOlRPu9qvj4916bP/tLOJ
9NJX68K1xk2A1wXWv7yGbf0YbmlHIAlv5bCiLjFNF3Hh41L3gvYUldbAOvTfyHpkDSFdrCPkB21J
ZpuQ6dNVf2Ec2vg//d33gqQXK2iIt2GPrv8CYayL9RYPngJK9W8LTJQ5d/gFUcSG1JJ/+A5i5Xmx
cu7tf10iLfHkt9sGRj35XlpaVrWKAO1pXV3zSVJ5TBS0sdkvEV2ElOc61h42glxFu8e58rUC9a7X
MV3xq9FzDHM8GsHDP9EuosllJBsXJaSsbUS1ApCrAV0htWDGB9jzKTVJ0iFEYv7vqFJ1NkkHtyua
6fUU/QQex7DWl52sT4ES/ePHTG3ZfRMx+3S8L5Un842wOWN2naGjWYq/y8TzC70S/dMklblOMccJ
0RZ021o4bxtjcFLn7gOKIsK33LImUi9TKHH55PlC/gSuUr0p8yxrCMVOs5Wtcn+1NEROgwvHMjFr
6iiLeKyQleSR4e/XssHy2Fqf7KIZq67OrtP1SeOWNOURMFRRkTcaDqv4IE5VRfxHVHEJnMqA8VWd
ho2YCGxxdP3fNyVhNnisD50pW5Vn0fJnKcPIjQBKPwBEIPE/34ku0AzfWtgb+1q4DMzGh5n/IgCh
f2Zi4zdvEgqB5miGAposcrYIcFxGIiNBLcoiLHy8QwbYq7SVFUa1LLobpqryUq3zsbUY7C6H2Y+u
K5lkdzUWf5JZW9/HniRe9waQFi1WJFylVschnvPDL+fAa0Y4KnOxRhB171u8hBmxSKM9dscpc5n4
bbg7sy60+2tq2IRF+fXMRuYbZ1XfasgUFcAckVjM+veG+nvZmPhmF8KkHTgLCG8zhPPgJF+JnbyK
SLCNQQfV84QarWJRU/pQE8gLPCwSAVlbIgXefFF9Li1F40c9l51TAYPNeZkpJqYTAM6lz7y4EZB3
9NyfOIEriB6AmbSNHnmRW6hFMJBlII3xUCxE/+K+bOX6R/80OHs4MNgZxumpyFmPLrGjNJIogEQ7
F9nofhW/tugx6AW3XPVXEVUsjmKThwBea5o0A3OKxW8vk38lUXArm+6ZySpMNW2yjn3LnDzVl9gE
4VJvdSoB8muTS7ZJLpYbu1ITHbcU3Yire7u3nfgnDmXl0bwetoYW9b/CXMwWQaDChZptFmhaloth
RdGTlb6ALUyZz9eTzqrlyA4tkDpedVT0Zd0w+U4iE3iphpd4LpHPMmjUc9VqXzrM/nf0/7PkDvXN
Z+AaeUOjGdgUdXYGUO3wSe/IFZaV1kjeTvmlzCw82NNheAXN6uSKAFRCbIMaGhiTv/ONYgogZ+5V
3o1hEsjUaNx7/c4eHfG1atmsx7SYMBwBn1oy+t3Y7DwUmwevriZKgowuN9+p+SbkWUHSTt/LVO+S
5zLYI2mffYTdPhFCkbH9HgDrGsgcRaOWPgxBvvW5W7adQVi70185/3s1OtyICj0H2dGj7Dng8RKC
DSeVL6JQcluvEiVBteGGbzKYVaTp8iIIwdvxF2ZHLPO23/kX1GnIsKM3huhHdriy9UFj6uu3qFsR
fNv165Rb57nB/fVA4ag+Fm19jIntKnXjbc7R4/lOLwI+jE4nGSRp5mdl59ShTJSHAl7DIfXQM4uD
w3lIRZsopHJL8rQGypc04Q0k9a66gf3XHBMICOokLJ9/+94g88siBSRbXCfKaSncR2sGY5+zYHlT
KPywbzkc4M8Vl8b5Dj0Xzd4X4aqycz85oINw+Lspt/w/wRdlcCvrkFBA27Kh4zrjjOoPRqIUt5G4
mDG7o4WjMLQxMGdaJIalNwe/UQiaZKC3IQXRrjl9h1O1JqYx4XFm2lJ0hPe5yqgpocJ9yF3gNFbs
dTag55QPDEZO7QInqwW2nc/e2z8MI9o3nqdsrnmE4Qyj3t8b61hEeL/G6ax5rYCnM5pIMLIiZJex
HEo0zL1dCtHQLLAZORa6J11KRswjjnBBb9ebl37PioznhopK/8BiieL9EuESoJJf2YtAenDSWQG4
ymBXTE2cBJU3mNanS2QcNx6EwbuExunORnzwOSQzk5HAHrq1Zib6/eNlThh20dJhLCCo83vcsbFC
gEiTjbvJ6yJX0bR1M7TDEQV0Wu2oUCf0/vVDZvnFRsuJL3yc+w4uOyGIwh5MyPFVZuMXdoNfMSV0
/6v1dpv4saYXjS14NWM0jlWCAOLfFW2DjgLcSEWvmWtSjjbiT6OVF3uU9qjyJN9yb4VHS1JBeew7
3f09TAOTo+u6+ytUmyK12cgqw4pdj1UZnVIuoCqqsbvYWtU2/V5NxP0NQMicQdiQl1RBT7N1G41Y
6rBq8NgFDD3wxBPj9P4w/m0NG7CHyHKmYf+sjUIg3a2spB7/AitIKjXKBt4ogfIfvAk6b7Xlx2Qm
KR/7m/5ZDdFdIx5BntoMLOQWmOiVg9ZN7f4pKVhBJfyx2tCZdGEZ8bnWgKpEZ99JkdDc4CIhVwWu
3VeIE4jvIpc59ziCuqeBj6Q2lrXrCKWkDGY0M6OPAmDFDwtX11cVsEqJQXirfVedneR5MuGXdKyw
I7PM8jUpvIvGq539WEnTp9RnuVkmRVi0o/BG3TKKANN/F7fP8u7mn6f9EP0fuz03/5GUDPmPob+P
9X2k9WMIbOsbf+5TLaXfkldmt3vv2y179aV37cmtkEAra3gAFtIexMFnwLUjUDEvUedf+0xiGj+p
FQ0F8l2fFrVUD3RBh4GuofKJ6PDSJ7DSL8T8ExphTJkBiD+qHPu1Ov2MfITLyud2KZolqvl90fuo
/c5fF/I4kbTg+PqeLBgis/YvEaxyDaG7ypetNzf8G3V1Ek1q+cMuZgv2I3o18T3Igwiv5WkOgsEy
MVCG/d+AjdQ/MOFU/Rj5niSh3n6mjwMLiTEihfCHnbNMMBNyuFmojPiE4GOAj5KneHt0/g41MUJi
RX8yX+1u2klvDddJbS752eZSb4ydeDoqBB9uQHaGnoWyFLIqR5H4YfGyCwAZ8+VDBPOTtSDspZ6w
4Dil806Qfj99UtWGib4x5rHLSVZ0Dla1nuY5G5rjq8zHd3WHL/svATQFZzLIdXPARelgNwCA+dnf
sjhP6Y6WZZeowcbHEAAFDABZozo8i+5k/u19RQmBHLlocAx25oKGr4J7hw7FkyLLoSvyOlRf46GA
mK1r00N+ogUTQ1mz25MPwcxdSOb7TQB302Qg6RA9cpvZOJMmrcytKg7ZgZs6ilM7AlhNk0pGxyFP
BRyW6VZFPOpjxgaBTzdM3gCD/+0Hkj7ooHXEtomOT+p7N/lS13kjg0x4NRG+fRekt95sIdGXd9XV
+txrJ0GeFbw68zksnl/EtWDRzpyqRf+c32gE6DL+BP+bCDogyK1kp76msDKAG+CXkbNq7OG2Psjp
d1DFDQEu2akPMcnGLDBhQCGMNHA7VCsOmguUs3O71CSzXp+2SocQtvhkgP3vla415DhI5tROdXsT
CYzrdtBxGXw1+ctkvw7wVja/sjj3MM5wkEZ1TZcocO5HepUiIdFg0IijnJIFf+SqBaIK62aVSTFo
R8ZskwWrDwEfPXuydmg1tkM2i88TpB6Ogg449C53o5SpQrkrJDIPcKZGzkCfOwaJhRjQCo1OM9qw
WImAeXqXJEgp5355JhJ2UIaQpEm4li9V9/EI9L3i1dnDKwkv7LkOp0XOOefpT1DIX7AH9e4oe0T6
2Rne0T8FWqZEdxM95/8Q3Uo0AjXq56HMsvGBwbIOPTJuo4Sh4WalkDt+3d2Y4t5GygUH+mIJUfRT
sdmdAcYkjXlxhaAfurA4zx6znS2Bl5F8/LfiGf9ZtCE0QeMuTHnWPKUHf1aAuv/EJTtX3r7vUS6Q
b8CKQwVgxuRbCKyNonU0yWCL0KnILaV8zzXxUGx0VLAJtUeEbNJl5WiqHg137r4kj6lWxm13d8ow
+177d5sKemC/bWf7+4lq7znRAEIUcYQlmkzY8xMLexQ/YIdDX+n4NP2ASo161s5IeE8cBGHZ7IHc
qY9NeWvOHCG0GPGI4ZyIQhH/d7Wqud0eDpMV1uRpl7Y4pqixpvRl/uQU2oOosritknnrvEpsopSy
C1vDn4rW3pPfXX/8TX4RinoDlpoS5aeN4RzzTA/GHOWMIrxVYBt61TWfwhdnNkIRUdUiugb0oJzQ
pxSAeA0krLnufuOTUKBA8+eQuZaBWOphXGRSNpFzq8187XS262zJvweMTKHGyBSJSAKx/smV3gHp
nd38McHxCIyUKqxkxEDdD/WtDTKhGF7N5VPNue+KXM74i+ikHvEbpXZ61ZdrxgmC4acxVlvDxqdZ
cNvDu0xXnIEm2h2w/NUY+bGGqP+DzgHtF1D7/hx18yltXyNmUI3F7yqS4at2D2FoYHcmqxk0uFau
UNe9Pf17HxQmsVAkq2B9U6RctjZIdJO/+LyQDhexpjGBHedDS8YSm5Y4gN/MQE1iC6yFX8G2NWro
bF83cPH1dIhl9xPfa38uAx6ipR8MpvMZofR9Wx0/kocMe/jLhLUnDNnH/2sW+MrlunjHSWbvPfPA
5L6fJ0LRhzsTtJ7i/UwbdarpgdCv75+hAYwnVpufRIIgbdFtPChdzKhSylpC0siCjw+e9wcET9CR
Zaha7qR3kPYhMJFDWNJX+dPp2sicBnoKuBuRN8XFJAEPgW8lhj/PE4FgsVdEzyT1FsiGTOwMxaBi
BkIhBm2UgA3ZjkjepJ8IIBf4s65uQfUHfKjfWycjPh3Y54ol6v74nTM2qrC6Q6gfZaZ6rK/OU2bm
uXXfRbBGfcpsKDwlExyUPsObrAk2Oc73hnCXVQdlCRnSVNP+vRnjGF8Ny9zHn7XwW70LRNS4rgLk
CYX6iMEwkx2sJ+G71zzx3emwa3bGX3XnH5jIqM+n9kidDN+NfzItZEVmrOHpDwLtzlVmDUL3tERp
llM128UNPS+oPtWX5Nz3ePiG2xqs/S2dEYKlpcmp6osqRGRpQqQCP1wF7EDFcxNLrag2XJeGlruL
yJoRtAtRKmOzl4fVZbmhk1+z6zML6Uzt8hYL5NCS0osmWUzF/3iV/FTYXDr46t9exXq2mBnDahkG
4qgtF81Mjfg585q89Z43IC0w0FO2fwfj5fXUtOD2BibYP9bs65zbr5xy8hhzDlUhY68gapkmjQ5v
XWYYTCucJYhHQTXGuJtT35UWx/0q1LQLa43Rtc16XRb91zRLGsh/Hj17xCvbG2HAi2+KiG45D/3N
CID9kMClAauT5BpYpNQELHDddir/bxJpsT0UidZVFstXqbQIoRAc7jrN93+lO6iBTOBQzQYO6bMD
8xutrKaJzWOXRcRooIa9FtGFAS4Ro9Qn+E6m+IH0cioCAJxE+MQhgxXz4PFFpXhcGPDXsnISfOPe
Tat94iRSy8XAUunJhumbD6C6bBgWtNaJmyUEhhFnWsKw2h13vXgAQX6wo3qyA6tDAnFc211sLFG2
og75lx6fNQ+EMbxtoY2C3nIy22hqgib6NRwr7SxrAOMCf5ZEY6Yak3AznrgNlPubw2pt0VeGkqjQ
CDmgjdnxnSfB+lfL+2ZCEBv2spxzIFKxA/9P0Fh6MnFKIZzlxhAFOqCi/2s3a3U2fMx/KPhPGn2+
Gd6BNohXNM3M8lFdgNB4OZuFcNiCQ7XpUEd+cLJMFgGssdiaTMNecSW5GfHRGb9Lz0oWE5uGW/WP
NdolF6/TZ2jW9kFq3w8RTRtmGnKrFLGDBcyYwz22nD3rGgGLPPshqE5ebHmw+t7r09U+zODbsHzQ
MGGJzeCOGNrsDr053ZW+lajs4lA/9P52uz59TY0jx1zdzQkaQ8dbZz4GF9VRzAj+udKBCiygMeF7
+A9pm9LntgO+S94lOXxssjb4Q2Tq1422yWKy5l6deyPvDPAFc/X0u5jd3hkjFdn3DTfdiXyjBWwp
PhTdaDRIFjuf5O1MUPO7fdK5CD9UGSwhvxlNA/OzfTeXKHPmzkoOMGOcAst0/lbw+t5AvQXNsMye
dfD+5V3rKL2+QnD0zPn0nH5h53cAdZtaXzdQRKAGJo+IOWqWcWi1zXhDR/I9lBUBE5Zxq52Z4Vwl
JxdF/ynVcpym4TE9wdrpSygdln/Hn28AI9DiAz0Bdm3LVO3s/hfwOloZGSIy+0oMk6NlFnTrl/Ew
u5Y+43H6uchTuxgMdE19QYO0hM705rRIeEeWX8liidgiFT9avPtJFlAGqqpE/eYl2w2kv1WlBhuR
JnL3Qtk9wCwyYG7/lO1MtI7PAeb7rFPXR6D/ujv517ayvlGzNkLGdoaaRquMcW2RCmTow/mIpbIZ
G49QDE/X6y4rbHDDWEpINjAbDKO2HaiQTbdx0oGXPeRaVRHmGfoVnFXxIHiutF0+UYakIHBNcFuj
Y+ArXIeOjjToKavh456mhgQU8PYF/csfdg7oXieRZYocKa2GK1ktZVqjtA8/bUC1rEfugo6cR31r
PNHD4MYqA42Z0es96FomVAw1AZY51wzGDeWRR7KCpnte4V2UFyZ1ZRf5PVNm8dGdgC4guSzckrhh
er3NXJL6qm3DQTY6PDk2R8uj2WA/CUBxaTdwVLWzFkG4fzLlNw3zWNrhtRhtBlhsO+sozol8Mfns
yC3wELeSeBOasB3ay3UYVnEtGAZ4u0dao0xMbciTCknaQqRr3JKFQJYjUN0VJnfk56HS1Tr3J7o0
XjSDL8yhPh+zpQhW8tf1Ctpe9PtEBEGMhjm/oieviHm1LftSXBOlfnRN+Gh2PrXcCnL35pBGye6M
S4t6uenZ0NQ6L5ecZ09N5nYuYUyZtfkfPopulnfs5dpXEsrePUqsvsw/XqugrIf8xdgbQbLi+0ud
dT7bITo5sxrihbxU+z4HswoW9KMmCcxNc7na4AdqqnrkQhe40B2mJCOCoYb3xDYZoUmkH5cd5Lf/
FhsbZ4riXFD3zKUs75YzCDSMtHbK75N/DoCAB9M9fu7wU7blevOlOhtK90l6KKGxptmc85tA6gY1
M1HwPBKKQdwR+7fsP7rsmRgMcwteCQx5PnmBMlzS273I3aHuhKy7phFJtLy18fR9O57hATMOkGax
hE26vVpNORUQ9nFYrrt8yZ9+bH8+r0ZP4B28EbUgZ1UVvL/m0MMIV11IZBUcB0t/6qHTh68NNHI2
K5WNd05JAZeA3UOAqToEQ9GuTIcsT2tH81BGiSLqSeeTNBI+rMWqlsaPLiWakZR3/0S+8NxOqfqM
I7BpcQ756Xw+7IrrUzay25d+Zob8NZ6lhmXkrQiNraL+Psf0YmtVRtSO6ccQ3Oa4FqZ3AKP3Yj3B
4pO7sSoPJur2TVU+VhITrvf0lE+hJ3C3dTyX/pPt2cxtsFW+92H4OQEGaz8Hj82HSQIx3b12UAdD
wJUrNd6LXqKTG8xKzGB/gJy+kl5cf7wsfpO59XiTuH+TBLnJ+uc8AQEVyv0Yuw1Fv55SrdcF0PJG
nYVcPL54R7n4bpvw1ZpiLnBr0tYv/zZQKxLVCsJfi4SzWa1qtkoEfkayFbFuU9epUgW0S6byhTa6
9FACoQPBChMGfeIdzdBjZeuFdPXRYBijAIR9AEclr2WW7c5k6DqqRhB9F8s8LV7cnvO+NyuHRATT
A6pdqb24IN/iS5Nmf573MbyyXGCAw5fszxJePuBvbdT9ek10jAUSnDDPhaoKkKVlaPdeH/OKc1X1
qvsBF0BNMOywWSHuEwwSedlCAWMpsd7iV1eCIXk9p7KbmFHnB2KcuiTU8Np6h1Rq3U1nRZSfouwp
Vu7nDSViQCHKBy6Cv9cNTEeaUMC1222+Pf1zLHy+A6sgrGKISly47QriCCRBUxWCWa7npnpIHovB
3acQI72VxbwohQB2iPHpQhhBk6cONbhJmhBqa8VpWowN5DVhVvT2kAAmRTrUQQGRRm3rELFavNlU
4i9fPXP48OFDwSXiTnlsXOvYlM0qP6YAWRl/r9BoWYlVZFkyjCyVEUyMEdqV2rynpHBtawRS7mu/
k7J825PrMFL6tYvC/t6q3tbRis2XW6kj8A/zfc8Jb3pRJmfYl8HuaBZjmv9qmqAIqdhOKzgQ7B3o
UWInic3lXWIpV0fTde4zJ5GWsrUf7EWUh1j84NWzFYVsdn3SgRFcEIZUxjLFB+zDyHrrNw5tsZjH
InijZJGaWcJatL8aCcBmYvM0KJVrX7LE87nJ9BcMwPUlzP6ETZT0kGYJlM6zsfmSz7rOfhPz7e4d
u81j41M/dx0HjvwNQ91sd6hHRRpqk3NpAe+mXd0E9tR9FidaYbudKqNUJpv5XzkI6MiL5btn9qEf
M63/XlLL9rrA0AuF6NapyhWx9zhWDoou0k5/GH4SMTh2h6nAOumC+U1u/Qj8P1rgoom4EoUVkNGx
ntckniAYpFYK6gbZpwZINwVYFsCovA8VmdpcAo3y5ehCDrgjQvcLVKLsJy5EXMZ6qG2eiSOhTsv2
K4bVZjcNSL5boMcjmyHscXcM4CIQTXSkQ8iUJtuWgNRvo59z3h2jlX1Qfyt+9M0IX+IWlo8N6UMc
ZPYNbACDdiGMNH9o8L/pVBrnpzzh3VjC+VguAIZ2hdUojtEQmQTDaBBOWoi3Kk+U9K7QOcLT5IZV
gQQusIVqwsqf4EC3hY+lB4QeH3dqfa+mM0Q2g0RJgRnUJQZ9rYJhSBd4Yu4MxRQkUTtwjXrt3/47
+ZOlnBtjIF4oJZkcz/i8W4It69TCi3SjgWIdojna7pDSkf93s9lh7lPgF59Tn04NII0iwiTe8sCb
gYMVSHhyi937qDPBjrrQ+kv0xchqrM7M9ZqaJ7YnhBjTGnrNatCHPi0V+nKInu0QWKLaa1+qmyc9
YCOrj5FLiy0cSXd3qW0yhqEfK4tZe35RwDcuDi1AJpLyuApdtQ7AGcsnsazywbdXUnj14NwdRE2d
ObOkjKYu7MMfM5GtxSoxskq8Ab6rAI4sxLAyOYGvmk+EDSw1eGwzY6k4wfwyE3g8flLOYzZMuQBO
2XtsN+GUHzeaau3K0i8qm6vklm5RAlGtwwZ/hL5cxIsV2IwV15YrASPAK+28tBGUht9ieLYhwBGB
/7Irvx38YavK5p94FkBVfEnHy6MwjOjEteiJ5UdGwg94z5etnHllvvbn73FvIf+e4BD+Y5m+lM3I
699lIVCeElRSfip3Z2ZkkSJ/SKBfWzBy39cniwZU7swqnE1WUBpXkEPhK5wnc7uxa0q3YbZa07f3
ZbsmCAzTF/6CmaviXzlNco2Y1y/zjXVdn29VxQlEJrJfHJuTH8KWtcecI+HYOAv6K/16zZ1Uv9eM
+Jk89c2yierBy2GmasjlhzBDyd1WEgR9YYdE1ybicJBRkmwk28YcEOkf0bZx2zkokDbyTJWX15KC
FvNaZXNsY5UEVTEbWZcLRFsEivZjOj6zqaDDYNNggE51RwasC7m8/v0/yMktUY03mAj6YHnB4yKK
NNhY7+m1BDxVvwLlYeszHCy+ivJMA1iCn3socS/jJ5gNpQOTPjbCw63zpuQ3tXk2+KFlFh/GzJcG
31Pj+RquHEuM+IoVoZLVBOcDky9gCPP2Z2RpFNxyuZ0Uj2TNQDXk8f8/LiqrX9ayTl6EpHYHdyde
WiikB6gp10X+gEm/LaflmQwbBJvgUAcCiSCJtZujH0a8e4ZROu5X9azYuWcxi5QPFPUbBHsqoome
SNU2IQrxgKkGmKqrGqDcnpsOW4ENh7xRm9PWXKSjYB6rHvPlbthJHp9a8r2QBLeL1UKefrg/4ODa
sX7AY0hvqXl2a+fVy+FG/HbWyG+oICgblIRC2kmUlzdmTmzDmTegzCcH1L3xRkG8CxQma6jc7Wxz
GWRRUnXHY+NWhJsvH0XWe5IyD3O4B/bb+zPL+/OThuwSdONbCJ2vmkHflLIs/laz11Kp8n1bfrKT
LJS87koXXvpDjOvidkCk1C1AM4gAaJfwUxHgESNvT7nrLGuR8JOSFTDT9tYfSvDqsWL+VQcaUg2d
ka4WsBMnvxeZ92bHfIbQMe2EIwrVgjLgB4lYUSW9lXorSncAWsThZ3OemiqzERDucgOI2V9pHXjL
DXIRmDxsumFT60v4tsq2c66qizHgvaLLNwHdloLcnCjjabVbZeKhRor45cughv+hI0MBFSWNjijm
q3Xp0ZVZpGS9gHDpqkJc4iou9tqBhZ5Oj3UUtGAw6T6IRHWqNoAvxlEu4meecUWYs9df0FzMKBGz
FOKvKMklxqQOj6peMuHnxoAL2lOph77CpVNCBdutMuAqqYx6dqeCZnvRqSmRrHmG6Q5tGO0q1cS3
kwnlejDnZeZjBw3ytig/JBQ6Klu5hd61EMnD/zFT4vW6wThUZjgg5i4BrCZH4yPMl7bqc6mSzD9t
V2Qo2Iqy686F02qUc/fKuLYsaxSSV0xp75uggpIzdhvzJVHRYviXsMaxCiLaHkL6ptEj9H3A1Vv0
RRpGWKZzsjtUHeXMg2TS7cM2ruuLWzVoW6/VWVn2PkY8UhV6H9OZDkdAcW1fWGpMgh7Z2yEw8kpa
TNYCyy4YplSbpdhRsKKmoaKzK2nqOkbaXhUt+ACc9EFRnyCGwSFbaEMPGcztaao0ixWjHXKS8DfM
tirIQN8M1F2ublcy6d8qZ9PWgaUQb+V6LKva7RLmOd/Uehz/lEw2fWCpw7bFLYxxTnQtpbWyRafw
isOOmXWab5FFfkZwp7xQ+GwjuJyAylbzikHc0Wc8nclct/J62s28FcDROhQVcqi++0ygRye05UVi
1Z4xPvF8rH6zPNFVK2k28wQNJb1GW+0UPXLrvck1qww6hmAcy8IaCgzI9QgQdlwmKvebUT+TigvC
r2Tcwcvmab0vZfjAXU/wMsDqddsONK4TRnCcLDH/Ks8hZm3o02RdNLnZI7+gx/6f28WEz7bJM0Ij
YGxsj0zZfFaG/hlqd+lQItMw/XYNimsy54w0vlIDeLg8vwSfVo+zzg3l/Ms2h0LP5rPuGWExZ0BD
H9ne96ihEBraHIN8ZtUPMD/2mq4m1pUlsq/n1U3AQlBXpbYDFrmIP27lvnSz8qouraDK+XAqNnBe
L5xYjOnr6ALqx4iLpvmn06F4m7kiQK201+tcT5w5dqvtZJwg34z07G09+RczjqUpHm/6ymUc47F/
YQtvC32ty5i4u69xuZLHQJsmR8V5lUbiKq9aOKuZruk8Fzwm/F13ccGC7D9RVoRscsjmzA0k/hUD
4wHnzpx3raPCROsPdwCzL4T8++TzPBRzqzpuzGkU3VuSsUMOOpmnH6eKJ/79X79mvAbNMyiDuyox
pTtYpqPKFSSu8ooRTpqUocklRtPCyQ/JHJP6P4g8njCvj+w2b+u9OOSsQ+ULFoUswSX5ak8vEKlX
VQBeg7J0caQtf17t8GrlGVvz1+SwTehpI+yqttnd8p2XaMzn3BuA9h85wRnlCDIxw2BQJkj9GwUw
szGl4NzkkHOQ7vUQmbD1TTwYGnKpETdlbcaESE1yYvf5VUh2gV9frtqNVBlcngMUvEBN5tHVf0t4
uRtuTEXhZdGNW97FS5JxWjDRUyBiXBFlvlSQa3ZKJGe0/NSu4LH2j2NcdUsaRx9HI5ScpyiNpqz2
VD9bRMyckJVNQZnpV0eKSHpoYfIG6Y/E9gLpCfjciYaW9FKuJ+d9wi0CsJfdy+lSmrRfENBZ5161
ADn33iF6lU88T1i/EYRadRzRdONv1PY29sk2QPunOiulWlBaF9ckrhXeSoi1BhuBDTEQ6xBWVinC
uJH/UIGweQaLwalPCUhuOyvkE6ACIV0GDuM81CxkF/HZ/ngRwpGywkfCVE5wHZSD0Sy/DlVZYJ+J
Mk3dccoUftURz07b9w5ZMYlTbhmh5kp30me9XYodPuM84xC3ksi3zemArmUfmDbhEpbjyPE0ckFY
5a0eh1fRAm+rjjMDazRWEknlG/pYeLJlrw3bro9109wB/y26nKK6bOM8R2uXsVXcVgfbke8QBccY
I+/mV1+uO3yaYy02MRE/XvmCFz7+8nBGXonVj9g4HBFFeL+RyZXdaqSO7qkwLjO3Ln1Pk0l04eua
weC3Zvr2PsNqlfiH0yC/St/A36XYLWtCgSk05DxcUYcHlD+8+Fgjo4WWvqTwvSKIouOvHhnIT94H
tMVIOZk3k0cVnlIcPDcAYEtC4vZc/EsEkhi+1zw3pX4jy1LNCk5OxuJwJi6IlHffQxgODm8kXDBO
Txt8k5RbUYVsm/XkJq9OKXRRObpCeZgSkWYUEf6dBNIIJDO8naYT4djlVY2zg3j21onDnEzqnv/+
mK6WPtpMUdlTbZ8v9udJBR3hczcPBH044BUCan0bmerEiiMVb3wxOnD/UgLICkY8d6ZKyJAH2a37
0L5gkLBd8N5hSJuUMq0e5qLjl4QLnkGW1VXUbXKUmNKCXmCXGyv6nomJLYmfRLWc6hfw/n6wgEaR
HMkSMI2M+rbDzVb+CEdR1o4oSN4a3wFRwxLQ86tDNzolv6xWABlJpF90wvXiuTvxdXlJ35dzGc+r
vzSIGhzvAXyW27Zv61CoQEH2rUE8pOGGBwnC9fEB1A1T9jT+qwvwXU05iSfHICZA8cxQvanSBA1m
QSEGAIINqT8n5gTdwAM/0QMu0zeBQjLnU/TmcfFmnu0LyUucqxCKu3wFm9Q6qFEpueY6zjlddR6+
LgnInGhJzKodhGdexpfIuIdDr2m2c1LJoXNI5USXPgXNiFQGUswdT/PAa2fAD5g0odP3O9b3Gy4A
1ZBvdP6czmNvgLyF3jRuccUpzk+0iX13R+rZ9hxdTTou3lcl321EUyGTsykms4SKZuCorQFuV5Ka
7Ho5YU+7+7+E9LdnOSq0lUvvJapN29IFQQpYJsNGvXfODE9S47QXKhtbUXc6DlNEwtPlH+pyKlXj
oWzoIHO7W1Q0+/bF9ckF8OWAvSvYHjl+45hAa4wUGIEmsonoKVIFfm5cqSGkXHT8xYISJGmublzL
Scpp1ngAxhC7CjdWv3Lh8sKFmkog+2JQine5+a84WiKmdzsDOur/TYqFGsTDicoduOLGBiAX2fEZ
+bZlIbxN5go2xmtR2RYI6LW3/OsTcboyDwQEDo/sAvGN/ghpowGpdLtkJfYAUfB+pE4AMSNa/9WO
hGzPxNk6MZ2Y5D2oW73Qeu7NYy6ODzUBmIF/hrrfSA1jq8kiQ3ayqpS5mRyTlYKz2NN0kOXTm8BU
IU0KEw1inyY7LBDodh57cWUdpZGvccir9X9zSJH/HAjoi5Jyiy6ZUGoRQAGtaivEHmDyYz9zZHgc
C3VL8uuxZISNLt81lKTPS85UwgsV55f+uNlFjpUQZIoP5pBwbjcS28+eyv6kdrZVskCKqFelmo9O
bJthhJuT8/nwZONkQnrE6N0QEJBlQVMUydS3S/m28X5j9fcnRh7GVQ3uzRVHoYFNe4f8R2tnDSHp
nqSbuv6K03ubuCGIxOtYJIDy7iafaCbTZo/IFvsRPH2xm11ypu47o/2kCgWRZu4uPydh3jSnGSLz
4idyUyoki1P3C1T+j1+XEVvxwmZG6V8MR3kqRYdR9OIxxdRjOcPH9vOBY7LX1KXgFGu/uwRoNhF8
Vm5jy4KXih0e13/ig89m8fcU2yZ6Opc3Ce0LSEwGtW+oCfomNyc59bnqK25WfuDN31sUANrTQusq
zyRGkPtkZposR9f6g96ORRW5lKg0GvwPzdOH8Y/ca6mS+lr9TM0gWaqNvmEMLOZRb95S4ZbQ7nMw
M9ti/M3cb2vmdCI7DK+3zlTn7VIb80B4SlZVibckyOh0fOdXQ5pjHZXcaoeadt0Gu9dts/F7b1J/
7jPRbKKCobu78Yrjyr3oBeisXOqbRKg4BptutX+Jv4FKdc5xJjPcY50enV1+vU87UBlfmgCggWtF
2VhiBQIaNMSJGp7Y8nbEAWa7guH7/M+h4VReIdEI3ILTXnv6fJiEfheSBld8yQ0lfp1PsFcEuJVE
UwyZUrxejOv6cgFRNyB9lu7OxiPqCKuQo1/QKJB7zaaSgdVvv24xVWO2nmVvu9sUVgY5BFSFbqDX
+VVeyT1Vb9PAHFJDzeH8wcvdgQQ5ocJv8qbi6eYxy2l+BvcJwRu46VRcaaLZTJIkY1oKsiUITtKh
kuYmAY+eEjBiWxpMvvbj59LSeyHHXhVB/nNir1qz8pqln0de6mLdcXi/5/MicNojyaPlbLuRZ7eR
3KptI7hmXPRDwtbicn7h2MfOXjlTAQpSSnmMikpIVFT+xpz3QCM4xp0It/Im2Ng9FaYX22pQ5kMh
tYqVULjn18QOycSOSZnEVba9yvED4Oio/cMWgoNzydM4lZk15GpI0xxL/tOlgwpBci9Ss/YdpOvu
6d4CCzCyykCoo6L6Hnebb5QQ4ZBU/pRAj4krpWSbeRSq2bevv3fjV4Hgmwki8NpoicyxgUYjJosG
JfcEKA9shdFaUFzKP9K+Yfxk5StJIB1kN1iyW7yko1Fb1iGCzx4MeH04LR/OKb7+35eVTYk77U0X
1kEyEwf/B+HQJ1yk3QOrR6Pt4m/j2ozwzCELIvd3nrkSEuLOkPOr3AuIUWHO+5S56PUeDhW2RW3P
0j42f4bLuQPfKei8AmB/DARGJ5SCzhz/66Ho/TkBs+ttbXRxmNGNrm4lqegcuUQB1H0BQWYpqjPq
95MwyXK36xs+1JjxpKkqKCiN8sAbjXJYg0ag+hjHi1X2R5rb2zqcV+CuTx/6urDxwEJEGyr+vzbc
krquUNtnkzVhi8rZRMFi9cwbSE9Am7ZdEkQudGe+lfakn89/Ar8VCUPTsd6pZvGIKcn+579us488
nKxcuxvk/3Q2bsDlZjkmNLuZ/jinybQJ4aqOVU3BqGTvtEdgPHPwLyIGcjeh6TL+wckV4yWh9bpa
GtlMZvtaR4jNmGm5zg1uXtKOJl5yYxUY8ehGr8FvUWqRnfmeVHFebQEZsW7+SZqee4PQTurix71V
ydLyUuAYvRU88U0bJWPvrZnUNJsPXAXA4FqKL3lZsygDAicOlT7/8/Kgz+x/ISE+HZZ84yehcL2y
p5kVipThI6qGTWrjTtEq91F6ENspSR/lI3SXNpWYC0QFsWvnOkpuKNcPGsE2d/7SJrvg+FHIM2Iu
JJXpvDWXkwx1cUCFyU5MIt1P5u6+qyKgkYaBTajuSaHBcG7IGvzmo6CX2VA3wJZRMOHhR2hhNwcy
jARK/9mvYlrlhITs+R+1oMmF7F4SS3JJAY4gDInocYW+07r3P0CY45csUqK2PkqWviESsngvstzA
HLo8vh/Ls5SV996WO2cFK4z6XzmOnzEGnI4ncH1C35V24Uh+a0+/Yq8WZs37gNrKzMpanHrS6b8r
znF9P6FPkZyXF37lNDhzpMpVcvCq+fKFFQwZS44GIe6QcLBI7MtdoVH5t4gpAYTluxe5DE9YVj1Q
XDGansaFSu8X76ek2TEf1cNS8yvG4/7XD0ZGqd2bdR1tc419BXMzDVQ/g/lYCY0ljZs0jG2Afd7U
Zi75q1mbToo/OqGbKrkF380WPDO+L1Exalmne9YLmgaLZlLNBqI3UqHHk7nF0jqGP6UP8X2cgqVn
ROZi96PlEGC31/5rFdHKdI1+lpGU/rlQABPIm/iZmq6NQjlm7nbAxaTw6mSmovzxEb8CWUBk6V5J
sSPqNmwJ+cypApUTY8NEsxJRsOwVoCNPqlSWnN0mfuBblWMPxRMZPMSlB5t3pDAwebPcny4ho525
AoWk7B8GhS7wZGTZiXf27EXQSn80irREMEVWbkr3zqi+3wtbUUQNnzE9w7ajklTKYnWi8I8AEyvM
KIoP1EoP7926HhFPUP3taCRBuqugb5/ZiP2OtfuV9xrXI3nq9oSP6+knJOx5msOFBnQIE+mtOpxF
goXPKxK3ptZ2w+YCo8Lk5/N6dpwmfJs4B8XvGirt1BCWsIxmE9KHIaEDeuZ3jwX3sJxzJ4NQ9jwV
bdGDEz7GPQAC6BIEL7PDLkfOCoeruVc2UTBjUHO1NR4nBhz6ms7E9Fo997GrUqjGVLyIsKoHMVwW
H5estSdD8oMzKr6wlwl/kkwFICX6U3czrYjqY/I0CEvi5DNU8wHBlrxmwa6cVk7EtNUSpJWa0QVb
i51gDkATO/89+bV+51FDdFNxYFzTYc8kYGK87OlMq+MbthsZ0ETsz16fSqdI6n6wwEP9801eCMHX
urRnHZRCZgkR6aryP0qmJAsPzdGglho4fDdy3HW1qCb+m8AV5mw4SWbF18KbPGk3KTN9yucnObfV
NBjxd3GBlwg6l7lY8wEkd7vjY6JyIThwEgd4Sd690QRiYFfVDux3rojILTav3Yz0N2XvE4iqUxgN
kICAOz8tEdHrIcbjWfZSDSI73f9o85yTRuiZgGHJy0AVx8J3eU/Ry1AnTk3F0XcvZCUcDS3AqDH8
FWbxYjsecee1/fJndbO355A+u5MUWuqZS6Oyb+kaDrIERbBnHRDJpl34HJhAHuiU7nz8GapdkEWB
ytpT0MSvMUsxtr3zDri80RXEqb33QiSfPuW+eyPC5Cq9c6rzxZWkAZcDN/3OVXre82IpeHH3aOLM
e+3VSPzJTGCMWMICRDUAhTjbGnsrkbdL18CBNx8tkXi3M/4IMhLYf/CU+oHGckQ8EEkzkGG9qEig
BgiaQeazcNo3KxtuwH7hxdOI4hPdctCbe4bIDWo8vNr8eV/9x2B+l3erI2lMxRsEeIUg5FQ8hN3z
n7wYc7zWprPd7bO1Vfg0sseJj+mleofErJ2Rdb/VSVrG6JnI9c+kU9snARhJVWjn2WxOO+YaNxrl
Aq/SpSSrNlDkVAVAazy95jh/lbOgpMYphXc2BNDmxnldr3u32xEmd1DKx1JnZF1z5ufwDZ6/YLRw
mNzUDZNRzeVlJgNp853jveCejXirSy3hWZmmVQ1l8jY+Mkbthm5vlWBqytH/Xw53HAunpbwBmEOW
3PoZVqncoWp+rRekSsVWQMdpu3euINd/qeOOIxUM1rkxU8POt6BEYJ6IjZoBfZ/ZTTC2fdiZynNy
DfYumlyQHeS5VOBA9BkMLgVzf/UgiC7cbS47tSeg2u05NagGi2imWYSby0P06hTKVG/LiFUJ1nCy
YLYQspZQHsGzoYgmJucWkexdAFhlGTGvO1ZeE4v0NVsUN0PyNIOtYMxVMA4BjUkBDAfbNRg2gynN
EMd5xHBr8UZbdka+BbYrnonKZauqea8s6KNZlTz146azAM/5O8iLf3QyB2lBwrhmXr2rBUOWOaHf
EwEOEXU4Xkq+wIcgGjENkWRI0N90vle9tmhOdaDLr8MfLd12MvnxoLbpvthNcKIY+ZrSq0oIAngh
olBlBx0Q8OzSp8meNYuQM6lCGkCDVzI1SYAbRTvod7Gvs9M9TWvWC/w1ZKLho/V6An9tMocGQvbi
/l7nH6nJ5cggfFTCor1DpejuX4dUO7ubSy8D9EPu+lwD/gdcJ+j2aTztUriNMtoH/j/Dv4lNLd46
5i/IBmC6e1ovnRs82XJk+nyMESd85Wu2fdRufSYPG0KgrooKzGI/3tOs7e5Pg1eyJisjdHoXhJkp
zOm/oWwR9mGYbqC6ySi8JkZNW8HABxwb2Q9pgbUyXe5XI384UKZ24V8ZMP/zpr6GOwXBFsmM2Oxh
ncoOGqbDIcLSAZKvI3xlVMIn3qyD+iHzFB/DHZdFCmYvBd5h+rD4MdQT3727yklj94ubRfOTCTa/
zn7UcnOikLIoFGlbrV+gpC4G+1K+uSycOY8QTWfmxLzhImdZu8F+DW5Bwckck+IXNXGRs3NR1/gG
zl7CqSfdIW0L/0Hl3fa9Hs8NMpvGPRwgECWyl9UBbgNIS/iisGx60E3NGjxrqk2VwRn47Vbx1aD0
7OyymGDU4qLRaUecAst87mnn2SlYHtPbMd+nDVxYT0O9nQEyT7xFWS1lVWs5JN1NocGI+4OBaeSI
H4niHzdYaCkpgvcySEGxcTmgRyoKQV6H+PfkEuZsU/WCbzSlCstt/It7a2lrsBl8d0YPbjU90P3W
/ApgOLHEo5ljvoDigDaMjeyrA8Q572d6aQ+1NY5VhLozr8zk/L8uBkUwhGG6BHXuUy2sbHVvXjDI
PZmsLfamFKaXSMCmO5o7T+SfOW7hiJHPNbXpBGHHf9IbrKwd5Pr1IkrwuLV6axbYa3TrymKIjYgw
kOxcE4OtVpL/8sR73dKSeTwm3zfiROynZXLVRPcMogLG46du14MPG3UwXxbwQ+KT3ZS6ld4mqNW8
RNsY6wNN7oaS7w0pEv4e1Kv1XfSUb99srbNjH7GDwL/pKWlcQncV6dvp/5f+Cikilkwc/r5Bo0ey
BObZAZCo1ZKBVVrOVS/6MryQIElRssRRGXWkivuKKNiEU4Ut60hUioM2R7tvS4J9hB8BMSOLgnA5
kUllFBzyHCCZSXMvMP/TexgDO+ykB/9rNBQjG3UfUqb5EEdaYBsRB1UKphItlh1BGzFRxQdndItB
6/Q2JMQUyzvnWfT+IpIBOaknm/YbXV6JIjT5TrkbL3NFgl0SKxtZ8f5r4O6KonGpqCcipOYTQCr9
DCjaxWtBMighKIxrn5j8rO4VrbpilV29y/eAj/OwJbxjkthMpvf7PeHMY/NYxiGQoLK0WqaTXA0o
S7kzEGhI3G1fEBoa1V6hh29Zw74BHnaavU2T+97xMvbEZ2MObaqlmMr9nQ3RA+IBa6NgYocwuR2P
+XZ70/Pmd/ohghiEWrSJzxtBAki0FfrXDZtQPbYKsRYYcSNxqT8L6GkCOw6WrBoFZIcnrBm45DDy
YMfsXHTVwcj0GRnJAoYYwx0EiALoLLXQQBw9jp3Q38aKjnqnk0zcfoDnRumIh8TwhTFJzewFGHua
4ehB47Rj3an9AKjS3Shhk+x8WHPn0P8aeViIjEIceBCDLnCmAQTnRwdDqTxEICV03UgoxzLciYZb
v7h8hBIJOCb9+PZSQ0S8aHVv1TSqQV7CAZB8usI+EYWaoFmL+b9qIsTRihSLdFUFOwfS9CRP43io
7+FFUWkBDK6P5i+ZcWNTHxGEcNuO9N3ncPh2v87HmMMcAv5kKdMXe3P4el+nNbbmF8YAhtmVG2R+
0GIBA4GYQixNE7Pfw9hWSJZMdW/ijj5sR3VFTIPeHA6ehtjSyyVbTsfvWWUa9XKnaWiiEo452KxD
YP2FzJTxI6lEErq1pkPHGGiBeDKg2AebNVFqTTg4Q7QNMTvG6Ggr2/VOY02Ly/m9WSd5muyISR3E
nqhNH1Kn1kLyLwFnHClqECvvArrINmp9M2GcW18PCZ9X4t6TsIcAlOn0/KhwwCFsTTFuNJsvDrgR
55FtELS02WbRYg5DiNilV6N0efwLGhXfH6KyKgSFBibf9d300tpOr3kHBxSnK+fBd4e7O8xw6GgI
v3mLimLzjK8qQiehaeAraTc8TRuGtJvkjBXEZzaRhllzB9K0m+m7qVR+ircyYsrt6+Mb1zrEUkvj
PK0Gugr3YRKNbidXl4R8BfAcTpKP9huXNh+ZT+QVpXJpWNvSc1AwgDKY5U06wGkAXCFMBMynkObs
yqBHaIC9iZl8yhhfcFHs8iX2cXEWXeZAX+F+101htGiGQuddGTRSygvai9ULAzdIZSxHBTOClXx7
ForD8gqrTeYiFkhr2aMf3zYF1YQp0Fm5HXoneoL8XgH9ReqUtYbX0+hDFhcRjaYj77kYNiTejOhR
Z+1N0P7J4cnM8SYoc++OrLlAIGC5G9cfEnaSQyW4RRMK1Rh9gXpUJkUPRd9KpR7fOFpc3bH8wn2S
9G9Q7s1v/UJbesJIosMti62igOuI5TUCU7qApOxpFixy6Mc4BTOBA3162qUgtuzsoyxBI0rVVYKK
NokLpPwzajPxAkaOd2iWHTxXzYZdotuuI9dDf4J5EFkF8dNfLyb/JL1165m4S+KOwvi89iqjZuMl
dGl2TWf9jAYQ30Fg52CQWgXGfWdn7/pujHBM6XgiInDZBrrnvIwch/ryvg+Rj49Dvr1JL0Og7UgJ
Gu4SiPrFTelJ1y3p4s0/PeLkun6UkhETzi02HAu+s73pEbfIs/LwYThXgPqXr4uJF8OSJzIqYS/E
LYRxy9E4jkOKYeVYPmNiMRY15TUair7N2ahqy1wAer16LsE2Z/Gs1f5dvvsH2ocrla6C/ObezsSD
IXTTivOpHHLmIqWkyYRDD+Z0oV2XYS4/BYrQ694dXIgwwNmtZZlHoccpH4uw1cdhqioZvXfp+xUn
9myVFu3z5UavCC6lxZPY1mx77Q3WAauouJvdJlIF0ExJCAneWALoDkHUlW1K4B5hHVnn1jwp1NuT
Bzf1Wun6VpZW1lAKLbv4hVgwJCX5Bo9qOWNf69HZ33g7PvodNbWwCEH5RbwMuVA7a0Hr8ByPcR56
bS/jZCHZqdvBk1pLblmKVIud6r8yj10aUUAofscb4e4iyL4FNCPXLqjtRkHY/tqPCXYG7Wc8QP6U
9R1Ky6b+w7rVaIN3RKMJudOui5T7cg7Go2xrpldOLTodbQHhjQg+skQKid3uWR8oJr0Os6K6fot9
kWBjk1z6jta8XQEhUFcnpcjJCnYLVZI8EGViXc/gPNe/lNS9iu9bDpBGTH2j7MU9HO0iVk4DhqrH
/gFDNdh7W9oH29YxZrFD4OFf7yFqlJvVGqR7UvhbHIwOJrspQpAauE7RPA9GMSxLR+crXgm+L7oA
+7keCo/e51SfGvYrmErZy549DkE2y3TmNLM7cVgtKkDRZrkv3nmiJHRxaPgeAQ1kMrplRQH8JiPr
oY8PYvg1wbUqauYcerREKjK7AOtFbs+4OG0spp2L+5FhOSmlLpIuHjS9a+8NPrLwSJlux9/6MQ//
TZqtXIsjFNoLcPpujaQOufpMUyuQ0nZpcGyLOub1JL03TBmEBD0EL7Hi0f4G+JiHmb6YDvlZOt/L
eERhpfYubKD7sP8kl9G776e8aoZ+9MzCJhhis7Y981areisGNGt+5W7pZhu6/N8DM1WVRWjwrpOi
K7YBW7kFzWGufq6pNE+nqb2JP0I7emrTdScfPCAHmLOF71yeu3yr9iS3EcX7SbH7+aXdpoF2P2nO
/CTUpDO520cxKuWBbFOR1Mp4Uag465yd60xWU4Yb/swuBn3DSvOpmOv3cKqMbSpUMNUFJXcOjjFV
ZGHN+nkttAlmGVzELMr+TJcM2cxqJ5ro+Yk6H0SGGfh+kergFa6xFQRWUX67Cdu0zWwi/GSf7dX/
INveVApQkYVLb+dbqEP96bJwWcIyUqZZnPPgfHGiz6ySvfYciGAxeCOVLU88qi5fDD7DUvkgzjy9
apCNjiJWAILN5AEpbtuYmIeXelrxel83taBUemR7Wnz5SJySbj4Lp753efcX/l5GZ8LZCvZcOsa1
SjeRKZws93zBOYDemo9PkbLFxQ3HUebaxaE4DpBR7k/qF6PfQhW68AvAxxnWljFMf/BlYSLe4KjF
To/dOX1BuwMUlsr1nl3pYDcBZDZ1oRDtBVMLoGWWmtKlpBIcjHoq0kREn3iLgUebJXsIlG/ELPqo
CHGyUUxx4425+j3+lnmmB+29h46VboThCkn+61VjL90TtahFmoMFLPf4C6QfMV4x/qJunHNK4EZc
M/gpY8LKQzLnztV57sQVkxk5hs6uj0rktFx8X++x5KhlK82SdN2yQ19G/HPjCfunAYFxIHnnfhbp
MmqZPsDwZ5/7KIU/QCj47b93POzlDtgqmEKVCkbKlD7ShZbUWp3o7L/xsolondzWNWmSeMLex7SF
EfKIsVg+EQCB+dYquTdkhWudOs1SNZRf1W48/GKYK+HMlBtU0mB4yoBQAf1oS0+QdtsvVe+fCfxy
Fv+QO2YTt4DujfNXD08chg5+8ZP/7SnU6d7QvpuTopiTAlDmb3PLcDQ7dNO/XXDoyGH2yjyuMHIT
ra5tf5TmOH3pfo7BmTPampANwZXxoVLIQWRL657zPmfCytFI2K0LKCCFY2Ju742+Afd8RQkgv4hE
qKo2hx1ND4PSAlK0ZBZj3JhJniVmZY04ZVMnzjtsevLKaLHiDnunYaeA4A7S81qY6OG9PRv64BGr
EGBLnmZfCn2y6q5CgE9UkQijhdsL5IIADnCdB4GOGUQhHF+TGh8Gl93rfbhAJlZspwMKJc/akdzs
pNuVfx7TQEc+Nz86S9zziomrmXFAVBt/UjUqpSv/mqNmkZCx2gNw016390QV8BmpNyPR8cJDznBP
DqcerBvvuXAIqSDYsHToh9myJDWzXq6qbkgavL8ouWLGTG7kEVPAnhacHH9TCYRiqlGhDsw+iOaR
H7xPG/H36QbKprq04LyIbEDqHx2M1WShzizvUMZ+q2O8jMCbiE/KoAk2l1LvzNYY+S8BmHQGErxl
sCILvqwoq0YSeGgsExYFDCqqgswTPQV0GFXr74CTIaSIS6W4WYIizzukvNAeRx/h46veu42rnc0d
285mZ+JAMH/VJjXGKFfIQSCUO/kseB5WdfFA9rwK0ffZdKUckiPXAZkT8v/R9VCoFQ9VBf1c4htt
9Qwsk975O4zMOlyjCF+HxhK/bilYdEdwH9hEirZGegjMJRDvqCk7FYwIlQVBDpU7uQ7Du+f/S2Z/
aqtj2u1FqTi8TOs3l85O4MIKlYmGuP9Z1fNbE9Lvg6uePujAFNxZO7sofjWXqvxuTx0ORBlIZ3bl
4q9Cl89jnCGjB5ZR3jBoZYN9rvHrluP6TGeiZpCeNQI8TtyWZRlhGs9Fh++6BNUZARxvd1QeXIS1
CRzSLYAsJxRh7mo5qewP9sSWDpgny146n1dduFMjX7DxAcs0vGax0rz12NBk9vuBGAxnnTddQLRc
OxjMEBJzuG7SSByO7uvmtTJNtnhAgIJyZKbPtecgI+gSuKTq7tKnc7CiOnF4w3YtFjIvo48dt5SO
kcJVf4+bFX0JGW3vChyLmvf5hzFK0txLQIQMMfD/fF38duP9ambbC6aRtVQhchHeyVIOW4p7sZNS
H6Eqhr1Op2JKYUEf2qIWwD+dnSqTtndUvwbcvMo7cokB7spv0yw3KHKj1kS+3fdLZOXnOQwkUDUR
CVM4/2ZeC0GWTSKtLxFB0GXyrH3VJL6ZmtX1ZY8q0peQLj01aV9WbDvNvPjCHQSaQlJy5QCUcRzV
oPoSi96FpGOZ9ATxWMwAeZuD+wJeBrdjNTAiZTjrwt7tkGFN3cYiCCLXuusDX8Kd346FCSxGU3nT
lLqb3hByde/XtU56ypMoyJ94jjtPUvGP9c0Bgf0cxexZRKIrFGGw7FbXgEh+pi1n+DVr2bxTePft
ulXLQk8olIUVLm0JzntQKhBMzO7U/g2JP97X/RlB2qHEBuEt7QqNWiNmQcKryMRdYJB6r+4nZJHb
DlAAOj8+FbLeKTB35KFG1q1uGREFG8KygVkfktNViw9E7fyCsft/JKkXMsn4ANOcHe9g5VAEfGfp
XtEPMl2kFLKsa3nuNlFNHI4oN2WkdPOvuW9ps7oGRb1SrX8bU+5/IWkCYwhg6a74rXqliYKU+2N0
X8KucXR5HCpksRFP47gfoIZPkEaH8UI+NHtdcX2ZX4kpCg4wxdEaSkuG6Me9wVh3monETDYNHLqn
I0C/pSR2DI+G+tn6f7HYXCrmibwZHPjmDNS8AX30Gu/EDq4TJOoKfIfiwjQdV35DFPMHqE2m5Hx2
ByEeA4XACTxHA1C3iFx6Wruu8Iyj4J3xcRo0Q5tqJVOU3YryKZkWyE7RM3/bgM8gAlrt4edasCSj
v2Nifpe8MEGm4YDgVYPFlcr332sEmKaN6jEcL61Ajb4lMeR6RCHNWzLDJhH/V71bFp/bhA6GM9na
YRYT0kZeJQmuGlD2iPAoLO/tVoPA3OUSAv42hEGyjJDusrZi/J7Gb3pB5/kzywVC6kIB8UcSje5f
suiwrUhk0NpW6mi62hrMlAUQgQzBBqzD1oTkUwBehkneRiEGOFLkE609CoJgbRszTUOu9mwAEQYS
wyv07whnf62AaufwZeQQeiZ2iS0dlwmfJOb6jUX0sI7hTG2gu0ONyaLn0RhyZu1LjAKPmW8cN96N
1rYr4vUZ2YK2Gy/JiA/iexlBDcpeVDrmVfIbCP2LDZbbUG8mvMzhR4nmcjxYgsEcJut+DhMFnPHH
Mf+ibhNpFwB2O6VitcCESc08Zfs3QSPo7pcnjXh/QO6nILA29V5JG1a336u7iRv8PAF83yKVHNCy
W17VOvKSU9NzAtYVoELSqgO3ch5W6HL9xrUVKAW6ra6BAL+CUHBfvmwXboEnQcolR5qVIKWWDUBN
jrZA8iyHPivXMlXAWw2bkT//HjVtXMH+DzgBFiiJr9M7jKI1Co6L0QzAzhYzSvumRt0PH88jR/cx
TfYqzInIBO++7/6r9c7847RjdCDu4559Sf5+8V/STe8KvrxqE5accUimGRIsrf6deXLG8NFoMV/U
q0x6kw1QDWGbgGcJNdsw7trfMza3XeVA1Uxw8dre3d+LEnX00NAIO8n91vMVOqAPjFHtXZLfNtkp
YjkL6+SO6LcCEqtULRGNJ25QKM5YASUDgzeUvGYs4zhQd3C3Xl6UkjYNKTGFuzZp1+dH6iLiBo0D
BFN+4VgZUwm9yLvkkZ+vW5umQZQFnzpXyLw25sQSOebKNVWgdaSBQjwjhCLGvJiDboaiBtZOZdZW
jk8L980rads3aXsnaX2Num73dmSxE5/V0Y93Ds4Y1siJC4kTSVAqQHbHHSbiZpmh2LLufD2zK3eO
xWLscV6Rs8Gga/+jvrU01oRiqEyoqujgo1QVOZe7IjOOSvnrqLjNOgAt74DRTrycD6vEKsEm3UH/
ALTcRwXmk5kIenH0GlBJFKLERldGL+dpjhPsajEfOO5zadqB/yzUlFx+cYmrlcm4Nx5muDzeTsCZ
3rUSsfzzzNz2m2y2NMArBGpZhvZ/FPEgl++FnTtpnlpj8FzGD8pIT2zKnbJlB7TY4azYXdjFmOir
xjtTpZniZ9tIt/57XARaTexNnWBZsuWhb34wl6eC5fRAwrxUZCaeu2Cm4R7Sr1LzT8niGy1JNTNu
qxGuRfH/0RwziXMrtTYI+Ol1xAb4/JjSQOh4M1rAYnEgCRdVsq2PCPAkN/ei0G93fkXvtSW28AcK
Vz7aZaQxAQmF5+1opWA2MIZEM77zL6aaprfYyKqDusBVELHqZd6XqKm1V1x59aSjSPNyBoCECu9v
TcPSHFDYvSorh259FSOLPYEE6DFfpn+IOy8w7kNiZonzAsA5FqV1H2JMsmnc4arwoY1Jbom2R9Yf
Wm6UlWtjfVvVAgUx7n39yjVzVW6FeXESJRThrZ1ObeJXpJuWfsIYx6eEjgse6o7+wIiMdyID13ND
29sa3nP4cd0DHiojc6MIgMk5qUCVIVBMYw0VBHwFkqOd45dTwPAhwvnLuj8yQ6FFd/Yhmu2eJzv9
gC3x8SUyrhuQvxhZr5wrn4gbCs+9l6TQSZYHXM6zDdddf1+fk7VFfvGqTp/wUFMTKSKZWMOhHAbS
vX4wPV3PjA1Y2iV0acs72zgnzC0JNlohBHj7jjSs1FVRSyKAIXds9zKuSZptQWWNRaW/BWjSvAuE
jJfsX0R4L6FkeZcH1MyYWbk4IZQC2hjdCswMf+RYpCnBDGbve8eEkgN4esy0gv2K3hzoKTgD8V7c
HsMBLB0X6k73u4XoA030gFi0H9dJAPVz1XlM43UkbUOZy7Kuzum50CXxh8LaZ9WZkGFt0zsMltUO
uFkO59Gz5gxtTXWaMWq9Axhazee0YvRFk0JbjbuB25WWweAG+/bDzX2NRhpNYJshQBp00ABKJBQW
sxq0ftLevQYKMHfqAQqs8VNrjliupr4LqPnEEzl8jBZEVQbQ5/+i+embS7xbw2081NRYjBI1ml5i
uxRLgbWi6pMKJNP9e9uRAw+ZPqKdqIONbWh9wlyY8FwWSUBg3UG4h8QvsFe8yDXOoQ3gMsRuvCCS
Nj9wkCOVBtv8lgh7YdJTr9ooxHROK5qt4EUCafGJFbpLiIYextwR3O6qdDQm3WBIhwG8h36+DCBa
QnQi8vQvuthaZWmDQvWC+Gk3jTGbLLURhL0Wmkf9govVoP+alXe5Q2DT6FFDzyN1XIrMhw4mO8DB
DoUmWWHBdLdYzV7VLzTzTdG5Z3+FkvjnMUXwL9Zu4O2QQQXSoozxtECRp7ZZYodzKS1zZXQKB8g3
4hAFwnflsaGZ9gMVmdyV4V5/yrvtIyYcz3OzINw+9sui4jUqWzquJ+cVEV6gS+SrNemSP71N2gUy
LKfp2pz3XuN7zHw7WVS1ViMg6/6Xuhitj0CfJg5MhyUx6MOhi2LNHtVCd6sRM5A4mxbsdPSejcsL
myLWg88479TkWSty6B1dE8spR8Qe73v7tWq/luqXjtbusBDEMNZggBibrIVf03hc434GP6cPtKfq
2jlklfku1JIKRTKDpBRh2irM00OfxWpBMBTAZghHeMN5AvYXDXNRiBJf4CJE5n/+Pt9ErIBn+KN4
2Ilucj3XEgc8DSMc+woMkEJqTDv9n9l+zKXA6gk805t+A05REOCOgF3gpG10VtBsFRDrOUsmDCFz
9OD9/M2sa8NrvIZpLdKxTayrUQrkr5q9kaEevJdK/2t/CgGLEXVzi1BZJ/Q0+OOprTWjPaU3f9FS
VziXrVaVzHF4vk8NnJeAz3IWa44jpfhGXYv3wcdtpIBhgS33R28e4TE=
`protect end_protected
