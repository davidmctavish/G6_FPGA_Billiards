`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U5fR7Ly6jiSnzpxVpLVxdeAF5t2+COWyOUR8htcQsU4ADoQEM3sR3zhZU5JjWl4RatPYfsbeTYft
wYNUBQTaaA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JcrSoLMVnM1/FW6D3akIb2to9//yc4kk9QHvtUmHBR/geBPupjNJC2ERoNhO+F3zmHiv4HuIEogz
r4Q8RzHSOq8YxlWIgWjTw6TMYbsuTIFEOwo5AgAT1p085bqstd8Dle00LtV/SPqQJtpaicUb+bcf
jKhn3/vwrkAixLxKMrs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WGswdTKoDvzBb0OdTFrc+G8T9pgH1IlCvte2o1yWS6s9T8D/L4lWwasMR/dq/Dr2RXhhmRgHrcAg
8YiyAOOh6JqhOQNiyvzcKKnYiMW3zQfM3RAwS4uFveKnHtiUkiTmv6patQiXXriS8XP5eFuBLtmL
eeHByW9/bblqbgDpbQLXjThT9YwQvMp86KMTG0ibeC3CbD2jHUsDMUFBeq0GSalmibZUJ44lg2JC
GC0CvwFvXEgHRjZUHXTTDhaeEB/Q80/P1rV35NQjlkBnEg9n7RcXjPwGSg5iM1RApbt72XVi10Zp
ISS9lMY+AhlJk/9gVUqxDoISekQ4V3NPK/qDJQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nStovpGU9Go+xari3N8GyyGoDvYVeJB0DthM/29iK2C7jagufawZn7elM3IVigG9PBHoiscywZsL
98Tdj26Yk3GhrzkdbppY8cMejlZrDEqyox08hbdyK8qXUMjaJjAQuWpH3ol2bO0RTh8J77Hwpk3R
iltKLX1a0kqcoYF15ww=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nXo15/AHkpYGC5tcNXbzPzFA+jd2VnvGSS23YFGlpP41iLfXCzX2UaYIOuHkNc3w5VGh8nsjdvMy
8zvKotY9TuTnjqYl8CMwVtmYhudnyfdwmJY7Yr2ftgmS9GzFOel1yvIy5+64uWTbQoN5wa0wEjjn
7X6aBmhyF2p3tXsGO4weXXS18oAoklW/MPedEODCOqnyOPUWgA+TWTb3QWtxaw0yctE16h6PTCxX
UE1JyNqFpyu/mgzWB+0UIFNXnlBlE2z/AU/25Zc9JyejzI2JJGREk0IABbAi/Rs0w3oX8HDTDwoq
jYbFGaTav9s0VEz/ljyptjtGzvv2Nfq9kXoORg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8400)
`protect data_block
8yV4sMIf3/x7+Vos1XIvTk19ai/acqQAfUPgoZyM3e4wIrEPHB+ru3WMBTELZYO/j9C26Y1cvNsW
8pMweth8XZxY6aPwevPdt8TIpaXGMTuVeboIwV9A9rh3oYSrugI3Dne1FmDH4HZ+Bkzb/UOPsBMA
nBW7a0JHkBIKwuB1ltX1XQOWxmWblgMClcNegCSsN8vj9wFFbUcnn0K2NPmHR4N1Q7ZPcHrNtgg7
FnJe0Pt28BBTEJpeIQCM0oTaUaNCjSmlNJr4qZq206AayDFynPV2CLin872CX4XsxqolD08dnwzQ
bDmZQRJNhYrne6t/ssYS9iLOxJJAruYOhNf3pOh9pTrBbzW98lhiAzBeO/uCRbuG2H29MBNXJl3T
7fruG9LYsSolN3f+CQQS4TsAR0b6RqEjofYyHRYhkkJrIzTcbUqWi4qRYzKLvvpv8DzhqusLGdHg
/LYhr6RVbTVNnJWnDPxclJSE+uJNVfzRhXm9SxIsdGUr1xLxnWzCGD6/h4ro8ISKD/9F4vd5KNOx
5lA7k7ZIgoXjHExbIUOZvq0Q/2RbQjz6jrx9SxVdPOodMhcFQBOMif5ciYMb4+lzr8OKTBMYCOzf
XnojaC8fyXNAi0JLF8Y1Q638r8i71He+ElPJz+TS07f8I5tgxFqfeI9ETE9rAVWzFNE+VF0MooKv
Kxf9TQGvWOKRcbbynC1sOcgoOLYXpq7xHgR220nn+yKIy+68GPU3dK5a7o2BwROvhRVe+oyhJ0TJ
Fei6ILAWg/x4oJSitG2WdJbfXsjECWK1PWPxoKvBEPZgFJR7e0U7PNZ1AwKnLgDK+wnVfXvP9YDE
coUa4iz8nExlrTQ7dVLg45wak6h+/jDQxPA454MCPcXvEcfDIbl42wz04vo29NHzMNaRQRPsssIp
T18pNnPc2P/vYC2eKO1rKEhXren2uFrllB569L0C5eZH3ET70Vh72V0I17jtFmF7qOFsiX9nNKHg
NanyB4lhYUf6FBnHnyYzAgPYxFnJ1xrySjSUX2UfJy9mNKshkKctPRvdhg8RAUcUVQGcICrRBeab
AdnFp7Il5vfnXgpnyUGjs3cY+3JzKb8dYuyPspuAtYv1DxSfoIvTUlVy+j1+OYX5qDS39P/eTaVO
QxyGXOCp+TJNCnUvpPYsMQm0fUBz4Vx2O8xpyqo3TvDSKgCjgIfOofzObueiXw7Wz5dkOOEFrWLR
K9pL7Fmb8LpTxpUiKIp+g1YVhGa/mXlqUvg3Wf/f9vFo+lAViKYEiO0ONjLOG4A4X2mY9gzrdB4S
+U35xXkJNW2jmaxaEvsbezD52FdO02DopZiagD/3ErkidWH2pzdXoN0xcnToHqdJAARw2/JIk6ce
2KmtHgiB1kpOj3wqjg2LW656Am5Mm7Jgu1SrsPqld2AhTWJnbmdf2QwZmeWT9v3VLv+OC9ZQ0dgu
bbEQPJOpVgdelJWkZDt6fR+WQCa7WYrVNRUYIfUuXi884NLTRQ6fXqnrRZfIH+osGDikw5/hGioY
TbvVQZpZ29m2+X/G6APbipXrGR+Jk6cFhD6hP9UkZWJQn4n6KbpnzvucA2B9jUoshqklpYbrANw4
aO7kjTBn1lOR+lx8vR+tm10pwv9gcErfU0rAC74wBhnI/iW1Zrys4k1xsJCY222gkjUETRp+r4GR
jGE0MVpeOLIjoDck46zFZx522wv+q2Tpv7ND+jOd1YIuEpzzXOw1YuvTu92/2liDMdm9H3BDodMM
BeLs7m64ZiPLUYSkgixCMBFUUObpbKsp9zZEUrsniW+1uPZXdTQQL2ihCdKDQS4hzI9vuBjHvfoe
6zaN8creZoztKkjb/vn5/b890oN09G5KEntpXipWsuKnl4C3kmaHmP5CP8rTFMREcUfmFJi2WYBw
9nrePAZxmWgADC3HOMfgSaSrfGXbGg0Qp/gLAG/vzf3WKPV/YiCNcsBMi63v7kPlMFyAKn31k4Xr
BkWwwvU8fsYemC5waZdUg3xc5OXQR5TKTwJ7UbkUbs9Za19pRiqgcilY+MhLuKcUGq7a3fwN9Ze+
N/X1tWZnoUhRB9ulSjstvwkuSCynRAsEkAYjctVu0k8cVbzsOtO3FqaOarkb9wxflQbizDymXIOK
QdCiYQmTzk0wJTs+QWjZjFxWkb5/KmfDSc0f6E7xUflCGNcAAYl2cMwRnMzk5Sq59ZXsBHMeXmPu
5EhAqcDeNLDDUBW1le7XON7jYOXg5OvmI/7duLC7W6cs1D7EJ85dBPbMQNrF6v693Eb+pVUyUKTz
hyJxpQHx4V9EG4fES396SJElpvATHReBPBMKOVlgWJH+SeaZYyhwg8BM5vXySyIM/q9LbH56uBoo
NPRSCA4bSMH1opc5QWyQaOH0Y0Ww/raCN7njgaX7BecU/xGxvYXHlsJFoNNCv5QVTY7VlI5K9JJd
WJWGh0+Nna9JdEhMTF/jSYpGFZy66WMi6zLhikE0jFOZNaVUFYuMp9vQQ1yrrHveRmgHrIJ/ntiG
o6viXMMAKRQ/43JSw98m+v1YiStcM3/EtU+cdLrqP7Nqe0P2pOY9bsgPEWy1l22/lsV52dnyxTHy
n1mZ4SoooMMjaxHu9UHz0tygX+/WvgU8TCE+7GHMqFbhYHm7MElTWLzKkDp5jQIXobc/7wX3DlIL
yOcrDX9wK7irk5tNQLFL1arZ+2ccQW1ObMjlQ33f01R7nx3G+FMAO2tVeYhMt7vf+bFj76uHYdV2
i1x9ts8hoBKScfFZqrXE6Zu4eUALlB0RUjBnpl2i4KuGdBeB8ToAxRrZn7eCT+PZfzs7lGCM/msn
jgQGnaHMrgepNrYZsA2YRG3uemDfWkX1lkUSIwJBOePROZOXhZ+dckORjAmXlmhRE5/LZJpsNvmR
vF3CHxxNHqPNucP6/JXmLUxbLHWzafwpLxQotdbTJU/LVrYp6wtO7/HaWl3hif1TjZ5W3KRjdWGD
Sx2UVpVKKouOURasUryXIt8mVJlMzB+HxGV/TtxPgsVXiPV48HpASBOVzlIJKyIgLa3izgxPi2Sj
cFRqh4jrN4sZWyqqc/puZH+EJfSW2t8vWwDXpOqWLlwdvt95LFuHbXIzQ7/WbjP1wggWyOQQotco
nzcR75CZ+UzS1kIp1TKubAIGGR8EJp2fHqXr3YBgY+E8ycFm95KNF1ZG5MZuzxqBPI7BnZgQVWos
1/UEZoeUvw1Z0T6mLFhj3Z4zopkjY8hclqOQ7VtM4xCwPdhWeMvV3y5wZfy4HBEqWiZFpwKaq3Lz
WGVdzw5CQc52hr+uHikwVdmNl6PGFTDr8Wthwal/sSpc4t2HjSRl4IAUBcsujgS4zbpsK9TQtmFY
a5i9W+pAMEpzIR4b62Dzf4/gmd+jSvO3vCf87Kxh6QGq4kirJ1lU5wb5ahqdS3TK9ErZNjj80HC1
PWxmkwOlT2Nc27KGp0r/hT0vftQHzXonFhWTMAY1gXzxxP84dl63pKZRmvkR4irCF54jZYltMxDk
x4pm1muiUc8/vN0GGeKNGrPJTBqyBHbJRwLy5fz/Su5PpohNjHh0EngaMHBtOAGXQAdtVaiDNsFs
AbcZR0IWCGOZmJcEuXjSBfsf9Zfffxv/RcO2MEnvKrdbPI/Gmezh0SVnHrtESsOvCsaXyJ33ZWZp
tD1OnjF+cKP6/g9M7cwlzyj7QVFSMou+FmsWCRzbrB6sWcqLxjjlYqetwuHms2AG0Cdgqkot0qCg
2Jsrhh79BgdKcj2QcaJtsKP6qXVu66TAQLclZhggb2ZOqRK8PWlq5zWuTknoABYUcFSLEkK4xkXM
M+EhKyn6RR5DlHBNtsfNuuXzJYCC0NGydfBOW6CqJIQM8cwmXOFTlMyQjHj1LY7fkHb+UXSsgPiP
/99ZIoe30N5Oxrkb1CrW+1QJruFjDmlp584YXhwSHrr9Lhinz1a1Iq7TBm8+nIw1KzR4spgedVAF
dLJFGj9vNLwlBJ7CugLZKVr3iDOEjskCQ9iBtqPydAJfp+fUbApZ47PLmhmBGnHFqhg+nrwTVkvI
2VE8AWOmFKb3tO1x+nq/Ny4YBTZqzxi3a+w4xYMco9HPuc0uyASU8ZHhKagOpCB9xkAGOuzpEhxX
G9RDFEdgrwHYARXeQLrrS4Gb5h8d3xMXwjZTs4ybqwJ8KqF70MSNFo/9oGlaBoGIvJQko6NIwVhq
APXuoMp1zflGf9AhaJcaLrjHYrAz0Pj2x5Fpc2TimvcT3vVl4zo5dSAZ/ypJ0UHOAmDM76uhYzPj
LSzSnU3GKB+udMD5FpP0TKUbR8oU1u9462FkWoOONUv1dRE3Ru3Pt3xDY2Y5x6fGHA3UPWDV0C7Z
YCNYgtvav00M3Exe7e0MLj4FwU0u1CyMqr8lodCiW9Ie4pcHLbp0GjJRtE8Y2x7BwLAdhKYvLz9P
9l03lqmq3PW+X4b6XyJBDDM95T+1FvhR0sVHUhtA/IXlTfCSBnKWcXTH5lO4xojvn6ZI4AzPHG9d
BfNBmmz3dsWcw/6H5SqWF4QmA6gNS3qtSgvVPD67l+DPKt5ZgoyXk9zH/s/R7GpFSdJLurRwghBL
E6Aio9L81neeVNHY8kqssmOxKlxsDBwZ/r7cBMRXoKONDymD0Fsplci4n+Z+RDXdn6MVynmiIU9Y
CwURTYYGoZGfgbfvgcjJWNUiasPncE6xIlQb9XFWJ+eJ7NbsP+g8vIyGjZhUH2cD/+dbzqOc+1c8
L7AX3GEDVoc5BWXxZGosxnDlFxs/FEhD9iIXbvBKx2crJYCAcRdvQvu4epuKJ3tUuwDLH1kYYyBQ
PpbVIAun2uR6rHGnZG/VEKznP5svma3+KVTyyCYJFWvEnvrM7OR2yh9BQkK9WUzlJJ2ysZK+s7gg
Mx2+40r/XLlaJfYtaO8ZG0fXGHYm1Dwfk3kzCXwXc4KqLlWOLZbMJNbfRkfRpCd4UIv7Avelziwh
Veec7SO3ZCSFdthYOflrHQX4nm9cG9ZN/vEDNuVfmUUDcH+F8lYBARHByUspaPRTcn2wOD5iwWeT
gz3QxZ8Q0jEmeRsF1OpnuDMNtq7Z5TeQvLPnTqNXKre4KJEMjP/x4eV8czwwBjsNh6A1VyrGV+MO
aR5UEnFkvvKdKeD4NLcEdm4xC1L3RBRKlHJ1HMybVF3xbhwnO3Oiws6Tqby15jH5J7KKH+wsCYLR
lL7dWRbYyxgqk9F4veNXihFk0eEpfLpxJqhNNHWqIGbOekb32L8zasrKpqs+TxV95oXDT+EaTj7I
O/nxBg3lEJiw06CtESwVOBr1sntlizKHwuI48b0tvKfGUEE/PBdgoRKPlPFI+lLDqAkuWciA1IK1
2SR7FhQAXif4Yg7HPFRuNyUcIuXRFDGq+GpCKze6GsacT2Uz6bOey7a/wm5eMQbVrctq+iyKHzI0
1Izm9qebpC9B3/Za6KwW7okl1aok4n8zy8QnYRLGBy0Et3n9NY5B9j/4v950jD/luCvCxAfrOiaY
br8ltV7dHcCRDIMCEUu/oFEYyowCk3CNRb5pQE86NFQTvE9XnxgaTJnDuBmxvkQRDrIjUSWttGqD
/QFxBXi4OUI8iedFFHGqhV8eglGA5Fo59FivVuM6yeHoQ+n/aDeOF+is4KRuWLe/zDC0WAJGN0f2
vAD4TC4ODh0XrFm6wt/AEHo0BYZ3TzE21TW+e2qsCzdvxtLjuMXvgLJz+7HkUqPY7Y8u8tf1pOK2
Qgg4iv+QXBJ4kXDJKxRWzeLCPk698qTXBxcD7VE76K1EGOEeUuec0LNP3IGknJ6weuBBoI/ox6/L
5LfTM4sk+tCgT7WA3AHdavABOoFLkePvlarJRPZjdswKdIMNoe+m39NEwDSx7rGUcDMmrmMAvgej
DmqD3ncwnn71+iGuGlZO5xzzhnhcmGVP5RjAoJ/Q4J8pH35DSjtaPdz5xZY1XWnhn1dSi3EyOjhI
o46V3nO5/7EI8liQ5ipr1txabDmsBkewRwjpJ9ynqVEmdHilKVneQzw4MHJlbf7sfcAseSQ4NZvs
kq6zXKZCVhknVYBhh/CzlMkCded/w0/nDNu0sKnhBeCIH/1x1V/LVLZuiCg8t7UdtjLXtsa3aeb0
BhMGsawr7uTkwpSEU3Z5EESUczYO6eEzAvx9B1TCnRfJe2mMj3wIG4GYtNF3H59uYZRrlXoqcOFo
6QhEMfXx4yLOhwaE0nUr5ksimygWwj2RE2qEhvNm7p8qml24JZ4L2SuJ6CMRKDGX5myAeqs739RB
Z11Q23JyBguSM/kunXL2FWOX3PW5tkn8GQVfE5N1slrs+uVrVh5h00L6Qf1AE1Y+sxwdDjrFlhzr
AbjaoLAtOyEqDzhEmRVnTiU1UHuwLVOrcuSTXdnW/9o1EUiGupfjwstRmU6DWgUDCFWRPYneU2QK
qGPFskfDVnA7cR3hq3A9MwmVPZDsPEaOFeFRh2IH07lGoCJN4eRlA0IrPM5SDxANDMcoNOsW7KTf
2x2d6ctnbzjbVC8arEQXyNj0bUX+yz/96D1EtZRYh6AMUXtY9g2AGnwVJEqvqoG7xqY+j2tluuqf
IqifNBx/n5VQmpLFgkbQSXBuVJxp3823YiopDQGjg/InEXJNcLpZ330RweQxOLCUnjFFll75mZXx
+VtHmIYb3XqcWTDP9hGYWC6Krx22A2UPA5EzD4jKyIcDSG0HEp5hBtLCGO5FJ8ihBQf9XAHavTo0
zLpTpbuDXparReC5o6TVe+IgPfLGX5y18A4HlaX+HOXQXyxx/GxaVs35Em/gi0zxcmJ7kwm8hPzR
q3kam/6ERMh9Ntnkq5hRLGEWkf7hgP6BK7HlvYgfr3wlsb2wa2ES4hmCrFVJDmsN8vVdVqJJw2Du
IGskDpry3QOR/+DgRCD2nUNBcWx0bBvzg5/kuEhcOz+ZSu4syN1QZs4ZIucWjRGqIxzQntnHNPp3
UwgaG6qXuZWR+lJobK6LyyYqM1SrPl/dUi/cbsqz14VmwgWH/4tkqZkzDCplwuah3BXfaZMD2pyC
+mPpbqOTuozUMfwQyvBL2ZKbLv9UjiYWpzKP1UgXMLb/CuLB6UCdbnAZJUpF0sMe952e8/8xBCfo
smxOGAYHPpF8Li6uvgx2q0/Jscqah9WA/MziwpjvoLNPFBwxbUNTd95M9A+x2fv0+w4P0NBfjnWC
N6Fqk4a2rQVy26sZjfZssG46NoUFTr7KGt9jR8jgWnXV0eAYj9FoGbrGmw4tsmtOFw5cg0dpfxBQ
3Ah6GtDYJpPSKkX4ss3QTCe4JMpOipMLlf7G/Lu6FczhnlSlG21Kv16gNho9I/iLCV1O1Wiip7Hb
IE57QDstUyvFfvK24zRbHUPGGu9gzaRgxw5/C/zSKtYf1oqRTOlebgNV4CHR9KULfubURNZvWOEL
rgNhndetTFtWeTyZlJObSKoNnE4eIDDTWXwQ3qWbII9xP3R8r0vFRhdKWvnVNikdQXaFN0npnbA/
dQbnjG7dVLMPRn4XU9nMIJJhz5Q6Apt4C3LXjc5QtjrnCci7v9xHJxUiJvUX7wx7wrSgZ7dsvJgo
bvKcrduk3BlVZhmeub805Mr/Ljz56ExLzIMXqAYlmOWP5N2/DZ4PVzMDlB+SftU1YbAW7lGfhewy
Bj8Ujxb5oMYgBW3TigbSojNb0nNN0VS/Y9VbvtqH1y2/J/+q6goN/58wE6+Vvl+fVZpTBS2SDWcc
Ma3q6kjnrGcmij7HRd1ikSFio9qSdUpbndidTvrSkHovkM0d0IHgdeeGxgAsmxiLI5q09iMeiiaw
PjfTVT/VvsyfHwnipbWRpXPB4z5T5ZfnUDpQY8pvU1SjQO+2Mthp3621DOiFmpt+W4FVOmdDVT5d
n5GeJLm9/p0AOitS1K2FG/eb8XsKVpBw6Y4QfysR+W7BjZMRw9m1Tzu8ORsWK7CgHgeEz735Ieim
YPkbqwv7iXYFiwGknfkagHsobbV1idDUl60/D4wHLaIWbu/vU+2q4UAtrkMbMl9gj10rek4m2x6/
dxvSznR4iTn03RT1L2WAAlQGlv1MAbgEVAFXn9QxXbG9B3GNL325sbQlbaDwHeVH1dP8Dm/mT/Ul
gxS8QaueS+4k/ZWKqOYF9nnghNFbq+jymjlUJdKXEwm8LaQY/bZZqYCQkbBuKWLktnUTAAqg8hml
Uddeqn03Hlo9NhmudHiiyF1YrmULRR3zZ2N7nzh9etco8rPEMXAgqr4cWSJojj0+XHo807b83Co6
b9LVeBrOliqEU4+6DuVGj2ezoILfSPp7B1SztVwzkSltGTJshzmgmyOGljZQUp76udoGzQ1+0XqK
gqOgLWXMOYFKMrtQKqXMOYeqJq/TY26BvsVwgQa9ybb00DA9Pskm8jFH7L68L1FeL3dOkYVDJssz
km2LEXS0K6woz9lUn0EVGFK8/FduJsE+sPMLbx7PcAU8mDcsDBrEIYVm92VweqKkabNn2/g0iBsL
9/ZYUOFRHhJdrrl1GzwocVp/6uwb9PqsEb3YrFEOW5QxKCKUehRGYXcbjDDQUHKyRUqW/3cGnrJ1
96xkTv/T9v7k6yWT2m3hbLxWCSIsruY2Vift5TB3f1rl29U8e26x1MO9TOHHOVJVpUF6/nxVNAZr
/zLaK6a0zPhXwpMb6oGh5VN7VH3ZQWh7vNN8E7oT5NDqnyfQed+t3ZEUgdHncbq7qx7uKrOyhmnp
R9mKbQpuqs0sv0kMG1aHOPTGs0bCCwvsYlrNrywkaL4MJn74xh2a1rczMzDrGLK3ofH6WbADEpsm
eOKe1v3T2MC8CrzAmtq2/Q9tFavlO4y+nGwgBFPqY2gI9Q02OCzWYvbDduwXtRpOx0VTy1Q02WSS
PgxvMglCtFk0VatHmn6xuD4ncie4minvla4aM57efGOaXGYh4A+BQ+nZr7JhPXFji+kD6NlC5Izr
2zVs3cVYQBczV9kuTfd1QsDq4R7SqCq2SRJ+gjWxNVtLjbOybRxV2cLY+PP01HdzeY3y28geEXdo
aaw6Bt4MoNdzUI9cv7NSu6YV/oYRZLdY+8Uu1D3hvAaMjKoexaQwpOYewEYhukwo0If+vWQpVkFX
h2A7oA9wNiryIWt/O1BMf4cHE7KMQbaAP26ky8d+ICf7m/UTmVnvQjE9FMPx/ZO8jW8v8toyKvN9
QO/7pdw3+Z5n15woloNnZn7GxaMgxGziU7SLIp3/UQtsep/wJZxBnR2OymgLdSvJEPaJd8m8bmu3
NgT0ZYWPeJ6XbZ8puu8H79fx7InAIua6XOvVttlCvPlJ6pLAQwRinWwRJNe6lX+RLt3mxOgVRZyz
SLzxPRiXeDzfKHWC97zOOhuCfY1X4/OfpLx0ddqwjmHzIaOlZ/Pbj7NlGYkQLnRqACDZ3Jw7TsSK
IrfOcclCucsqBRPD1cywyoLbNg0mRZU50EQVYrRTIwrlPxX0yXWdjQiopgYMtSgGIMgZFVMbWNs1
3+cdgm9X8urxVtWfabsmERqsLz8AE5kLsrrDBOsFVeHcvKFdKgtDSNHrQUOFjBbatTU5p1tGDLtI
4PZPozMYmNNXoir1nKhWByfA6QuAHyGVxZ0CiPVAKTLOGI2KPUPpvkphye4mhBb17GfltksDQdjq
nD8qF/jlxSRj7em1kMrMI8Bq85OZtvLKsraK5Lu4EKXwUTXbpkf5xdma9FvzL+iOEK684ypXbKXh
+jpigUjFHknKDaA6VViw7KDTNlZR/+KCvzW6SAyqp00x8JExpdICNKWytCNpn1p9xVjchr6aBM0t
p58KwLX9F2r7VBD48J4tjUn1aE4DDHJFAfh6LYyxqatwc2EZieUBL858KlYc6PWaiJfcGmOl575f
u+TYKSRt3DjxC0p97tLrcEw4kzP7FaUlPcW3NexbplyOkuODCFQkj6CsjQx+dL64u7DdgZFM6Jv2
S/CIMMnmbYKZEH0U3nVNXEeMiKCrF0p92VhpJdckiRx5LaYjUjX7VnPWeCVRGF9cdWoQLODJwN/x
1vca3z6jb9RnlUpRF9Gsyb0r9QbB9vlOcPOP9sZAkmMiD5ULnqYr4cXajxCI0j9mkRIl64xfSmrc
0Dcl+9fCvEolCea2Yft8RfBhE81Fgpv2PHJWRmpExEZmBEe96z8IAZDI3BMaKezM+v2LbovJha8C
ATSwLBD4xZLBCBO0+0foTvskrgWkKZLSusVZwPCdBeIz3y8NWJkinefXhXM316w/6MaoIY6imbno
+fcpkmvH1A9IYD+4DHvNMYlZoK6qvpCnZqrfs6gKhE8/A5AhMKdRZ0tbSennPCRcZn0xg0tW8iEW
shYY3HywQzUeSZ1NGDjeIA6A4l2TEn6AF1Tpm8sFioivvXOxFBS8y0BXx1Ixr/wg/mMFT4+gUvFc
KmeGnLS0TQrbhMi8ohzdxIJ5RHL3vfTslRysN1o5dEEVNDjrgdRTfzSjYs1Y6OWTNNZFUkCS99Lc
larRgkDyOf8G/q9jHu7vDUT8j1DIFl+K6I1BIdMySADoGSzXxBwcIo5CGrxeE6pf86/E3NcVXYPi
Qnau3ILqu7ZVgaL+JKw1vfohehybkcoCwbQtaYrmSU7TATU3g6xUn4qk47Ef0VJ6sKac1Gb1YoHs
uP2YkIANQ+I42BKVugJvD3Gy5wxwJQINdKqC4OyhRnT5lkwPh847lVa4ElwOYniE6SkUgcAFiwV1
RoU5kbY7741UclCuOt3d4q+1xb8KbKMCpRELrJehSF2EYae/CUoPDzBfszxP1xf2wDdAbA05MT1/
MJ0iBLqIyMjlK0N4wX6tNOCqnfTF55E1ZJpJBiiGx/Xi+shlIUZy+tQzez4q64KsVolBjJbtIG3R
tikERUsf1QLB/LURtgO0lrlILFq34uV/kd0zLsRs0Cf2nq8g1ZW28MLDDgRM0KynH2BrJExBxK9G
mFymDYsKAMyYWO/b2B2KARR7CeGW8r2oR2WP3fCrfKwARmHV1yoZ19ewhOtOqtpGMHQ+2SnQ8klh
1CG8O6XhojSaglJ+Pi9ioxln6AZqKVrkkkt81go1mSrk+n51jURq6zIhJKtIfsDnkLT9g8/+xYiP
PTAoyjOK1JB6vVdRsmEN2KGaW79pq/8NyxT4qCWuyXVLrPYDnJsd53jIhmKAj0MATo2Cvzg7+D01
tQRwdtggJ0ZDN1xGPKiiyEJmr49vgjUKTpk+8oe3jcQJSIOBAnVcqoShK0wbECPu//KBmnsjq/ry
B031UWA2LdeaEBo8kMVjYE4hZ4wL
`protect end_protected
