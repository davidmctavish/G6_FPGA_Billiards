`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bX/e7HKXt5fB+Vp/no5snmR+Y6bAR0gZ8eOu3RjMWMySuG4mXkvEOXNCMaex7kZCNF3SJFo1a3Pn
m6EtqQj4LA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DaE0+omCn38Cw3I3i1/jiq8uL3Rz0Ja5LKy7ybMjb6phupUzKGzs9M6KvlPul6XWm4YvTfNKO8hH
01RqtOPSZTDe0FOGXWx+m/M1d8qMh+sQ+EAZk9p8iVnSVRmIQmWA8Win9XtntLm+lo09sr5lJQ4p
edPOIeqHc69Pffm5EDc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fjfIFxZLcdJcOCBuls/T4XWS7/PfAntYBtrz/GHgqfPnkNFzLVEly8zNJIHziQtbMu/kDBU4zazB
guJzJaEEojtlEIVz2a5xOFkNgFJ81VcLYJ6+uayRClvCBYV9RGEl+YUi1nBLh0lz6xukVzaRcWg5
sUMoxEwKlepaiXCMKwA9ZmiGNb5DeCBhr4Idyohgt0U2/fiDxHyYwe5k0wXUaxdo/4rFCxdRLTWd
o26hpf9PZ//M/oOcUibfyS82tix6Ei/2cwcDvnCJ3MhAtaLaxCV6PKFXg327fKgN2Iz8XQN8OTIG
utfw1dqZ5ivk4HBbUQdnCqEY6qKPg/tCsOz+Pg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nf+0z41D75t3Bs2sakAG7W+75TxyRwm5e6r+E1esHRZLkYdy8dj47PYsT9hqZh8M88fBLOdcaelo
AfgrAlOtXG3xFneVLtwq/RkcYe/zAFu/ndKDdKp/Fd8h5ZIuM4KhSApgrPy0iuTlCPj26zVm03jR
zWUalXFDcZB3M7lxqDE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MbFcTBCjRb10u3WNKyLoegPmHGry4fS8H7G84zIIf+WnFRmQyQUZH/NOEhVZU3dCRYBA5aL0kpZJ
IoVJfFk+p12ly3tg0T+n/cvYABYhXeegKlYt0pphgqSskgypJdGASSMUKE2WTa12KDiJ+yQFDlSl
un8tlsKT+pISfuhXyfi+i1aCGNzOpCrDRYY7nxkXC8LMxjancXFCfwGi2lCHAFwhtguHu9NreL4M
LxpBpawTfBDaMUYrjv6JInU3rtMqyuYzyUueiLDdH9U3i5mRgVWqGye0SfM57dlMGKdrvXtRQFFt
T8RN30s2P+qQF2l4m/sBtli3DiQCGLphCz+/jg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 68608)
`protect data_block
joIEDx1hlsebdklPwUJQH/oGYbPXL8UT9L+CxMZRNaTHopI5lG2efbXXRrvopUMRxzhUguZ+CNJC
A+so8kxIvNm4sMI8CjAL5X0nsE2wHNerJUbn/V7fl1fZAdyTd/NYT3QmDJXkuh0fN6HySCa8RZRv
658o6Yjg0IQfl1mzvvVJf4G4WC+tspmoFD6qGSFW9kZupLVPUl+MeHjnqhDZzwFKDkYLdlhhp7ln
X6wRhwt54Iti8dpig6kk/ouHghXqd1LvJVeiLIdC4i3I79rvVebFWEF/sXl2vdm4Nie4RjRdnAe5
5Emd+STZduW5EdvbU7rkEqrl4Ctb76zCNoaL/2RzklQELw0SojXoa/me1hpIGarx33ZRZLUyEPRm
MBfbonq7yiKqc3e5MqbJfV1fnkDqpQmZQ7idKZaUOzPFzJlMj5+sm3RoD81fGIhibB5G36doIqJc
upicSGwcTa1LaXKsFF5nJFUadULgwLhuKxsWIS8tMloz2tE3eGhUhJ38ehIT5R/874pxFG6HuO6p
M281XEliOqtJPmKQWo/oOcClOw+6F2nkKEltVpssqVZMKy5MyaB68Jb980aFIJRxdXzThJ3lCAE8
uH2Aw9JJvA+v3FMGGR5lR9WxcMiEDZIhclf+wU6TiIcba6iKS1BmmBC4jtFv+ki2Z9XgAOtbj49f
X7Py+pW/xIjASQmE45i0YiyUHFbKUe030IBe4smCsq0yd72Yt40ilSw8CAFxpxTVbAlBGCCqoNx/
ZOy89zdO3ploQpWLEX0sf45gGQymYkTGA4EYIVFuPt6zKGhc1jOI55UmYu+iWIAwS2UOyLLa84v4
ykkUZAXSZaYjsKlZa3kc1mr03g6+U50MYqn++X/EKzEMMXKSsXSYm97+yvLt278OPqY/5wR8OXjv
sWkrrRlhlQnP3goZrVTFLD757gnbvDUHlv7FnETepvopT4bvjS0CdyVL6d29GKqcmLXKSpblKv9/
/2OKfYO1KkgeL+TMLvvYqd9u6886lSGhjV0BLiWesZMLY+32pCzfvZ7ojZWGXL6reA//R3OofzUB
Qf291Lxik5scnRDyv5uioWbV/NerujA4s3r8NR73AbXP5PDFD8nmVVkAj58t+4oBI+LSNn8KEQ4F
Wahdx87iTS6RmoS/kn0bW4R4mrHL4BhuP3GTy5jPXDFMC4mctt1qrrKEJEViZG0ZMHLXpCRy5Ip8
9bWtpOCIOvecfrLUai9oHmc1RGeVfkjgEemfdxZCmk9hI0cOBdabAc6pu4AKW1GuYUQxjHO5mcf+
Zp8Pb3gVRw3WxctB/VksTXhrmAuOV/CWZ9FJn2e/S5J5X/IxuLfgMEzoGcBMZ6XVp2UH6PdH9N4b
MoWRYh5qfXCeWwbmEf096NNmWRO7oGrlBxl5+hTwC6f0wCBW6gr7IXTS5fEFFVX7Yc/ca8PpBZlN
JZr5oaRpSTQunZpIZ3G9BXsnPHmvb5ZA1nuI/Liu/thDDGrRhVICzfySveqiCZG5huOlu67CjRnX
g5Ih+R0btxDX9IR2TveMclN2/Pz8H8FavjJ2mXfQAe2S0Gc+lrUjqJcdj/WNXHZLbtCA/XhynriZ
Z4ZUeRY9M/B9h6wMeKOzIe+FtoZJxZO8nOEqd6y2l2OiCSaOAxkYdJYDSMjPV0/5uVqNpy9H3KYB
zUKHEto3RcepapXUBm3Ns1EyBO+KylA90rMzO15/Bvwz077BU5bhlFCXhUSIvML9KWNkl3DMWcHE
uuuPwzlzhhELGgK4tqBihHxOT4GmLFl5tYLoKmM+HAcD0ZbzdDzpiUBJIUadzJhr+nbiQbScskrd
GHmgSOuwS8aEvIfWbgJBz3F52VOWHonDGyVp4blC0ttxsIuKHCMZbEUwUzbOMCkXBVykByf27NSR
tuyr5FEQSguBJ+At0ycT1bQaOPAw0cdplRiTg4PB1sW0pWPQu/WzmN8LgI00+l4ZneoyJbsj0Crr
XxoP/aHeS+7kqdU8/3cn91eQAcy7/dyKaotaqlUcGfYz5i2fyfm/9yftk+m0sz/l4zBn/56xK7rN
EH1A+yV436bXrVtdJjG1htBvf47+JgjBGQ+FzVhVRIVgXThaXSj4AFPaY04MqN/vQrY4elMpM5hZ
SaJAzAOrhHTARXHR9o96BNnD5If1aHAiDSm2wjN5xm5rsjsLhM1C6IO8wYkhJ8ruqp61XAFzWxuI
oYxfzs8RwYgX+hiT233Vm1gul2BFrXYe78kqgdbREOt0bMiQgKvqnL2daPaW1uAiqhSlpCYYwubY
BIzR4lIlnvHwPo1fBJ/LgT2Ns/egFLtKRkZqN3kos0qu8m8TRPb56S3b2EAKLZBz7Zhg3Xeaz0GX
tvq5uYt/Hl7bu5A6kI4kc7fsCO4fI9xec5oYUWXRcOB+5kAyW0/boDyEDN/FFqdBcq1LC24ITOz/
QiADVnGLJVT4iu15oYLzI8myIncMTqYxJm3o/wb2rdtSEKoMt90mnxMPluR1CHFwVTx7lr0r1HIL
Ko8IoFuvQ6RV4A8j+R/uCEdsLJdoWpE3GwIMfkIs4Oz99saGre6/fAsSRCUEvidkUwtDbJUdsWDK
alS3Q3RBvGPItRhOXRU2im/iWTVCnJvR90ZoYNkB7cpHRBW4ShhoF3a8Cbak7lb/HbsAFwB9mncu
tHQQUp3klE9z0gS1c6Q5txYKg3xrUzMyg8EOn5TrNtcAxc5Gqx1/QJosQCbFdvU1xah0KfQang09
EOPz6CLryadC++8fDtUpc/cPo4tWdfhrrCy5C/HsoWHPzvI9kQYQ9WPANZ6Xx/4G6mTXl92oUhhR
u55tclbfr3H2ay6jGX+X41Xn3pzb7MLxShqAv1hiuB9Jch09wmTOoLpKslPQM33Y5DBmkdfnb7tp
ZWmGzPGSZFcyTHFCUtW1qpFmM+djRn6XnjJdP24IXVHQ6kXdrr431b+ejddViellf7Pjq4Q6l5de
Ib2R6CaJ97wKfBDmOTpHPWFcveTLCrvvYzTPIb+HGs0Z0+d9SmAjWqtmjx4eYZiUSsyrNlTR5O1a
soc3zoTl9LpIpACgnaPJUelFP3xY6uJBAfyu++nNv7/j5GqmTeo6nCJEHK1fO85Gdj9oh4r772Mf
DX/PeCOMp4aUNxVUe9lnBuE+RvmOciL1jdpapCHuEagnrw4C+wtet0HZZOyRRv795Mc+N81emOSz
4v8BPjq8M648ulQJk9FeH+UB6XI2fFOOpQ4RYfH6YYwlQiQBzVi4pS3xZb80o9z8JlQ5PQ7yRHer
cWPEj/GLsyt2MzzBk6zjiIVGmEiGjIo8qBp9w5KasDuEB+D2nH+4bdWPwyJ7QQOu6E5aIOTPyebx
mRpwP344xjtMiEw6bFV+K6YLShQCDqXdu7OSNx9EApGIorFMaPKPbeMqCta67F5fcwln7yFDTkqo
bYng3MuA6sXVK3qjvURLuHQVCGi3NGZfkfePuY1HGhnEw0rFpFQ1N4aLa5Es7Yo39YxAZFheYlNy
5M9gexdTE2K8aBnoiHwV9VSyxJrxqmaMSW4oOXbYpQaSCmozcYC8ruNVQQUen2JROy864gmfazUU
rggPgbajEpdbm4pYdtX+DJeBc+LToAe4OXzltTdLzwv1Ab0mbXD4sbiSpNmZSNH4UuuHkEQcuHCd
7SlV+K//HGwnw1EIuYUA+AANun2e+VvMCjELb7Aj2CK8aAF5Q411oLHCIWIHZr5/dV4akkaqClI7
bWUeiV/PBs7PAVYa+e1J8O2aunIGNHTDzHXAQ1ghSlVPKjHIHZn+X23FISe7w381dgyUC1OeADY5
6ioRZ3f4hCxeBGCOINy4Q2XCxIxMhGyiOzG8RcZ4QZ/e5VEeOzWg2XU65osBqeQ60tKzbt+zI6/B
1qKZeQEo/ZdykCzWPIjY9uFecqclM77sSfLexkUG4eCBrd+eXH0l0a56qXItRnTeVJ6u6stc0LWG
4knVzCSoyA2nLofVFSArCccyJybSS7LJT4gqJp9m5bugB+F3WDefULJ4geYlUm22PzSJCdqoAFOz
V3FGUrpKA62SM0ZZzE/gOzLu8N4beFZsf6ZB543QT3dwH7cbXs0PzY2uBF4G9Z6cnqzBeOlXxdfU
/zTVzu6GbM22nIMJc43/S+Gu3E4bbG1wM1YXjTob4bnZ/KOnssDomlS2STkwpsBJ0qX8DWHILaME
FTe/hSemvktIicaxHd/qkNbqYtiYOSP2uKEyYmonziR6eLHqKK8IELQgeFGpacZX8iQINnpHU1Un
mDzh0JgYApk/1R6LJRanVcIsl6yUN1tw5HWoe99JVXTbFmTmGA5JOYTnIdVD8ZyOvcteb5mPgGmc
U0RsS2aoukND6kRRlCQLDjabRJ4woRLir49XKlRiwBwr7DvFA5HPwdo7g6n+FkoQObWsDbB8mJ0C
ltt1N0fH5roHaHnNxqfRvQM60m83BOruFn/7XUZDdII6UxQ7MDWcpBAaJNGFXy1bIHg1TrSAC/Wz
GoxjschgGyJU9MfMOgjlam8Y1t4kTloVQZ/HB1rTdlQgVUkHaoBWUvO3B11/yajHztzSilpMERli
/JnY8dRofNPnrnHCqU6NBzCM+ixqj43KNYQ5zAJ4qcmofAw9yHwWm7MOquiSTEovul3VaOmd+tck
L25gZN89ZKY4DCPzXvDSX4aQIUMPfzbr/XYFQ2Ly754AioE4A63jgZA+cU+dOt1TZ9rHVzVM3LhL
DMIWKG7Nsuo1cXs4IXS0R4AYU2npubkwXhvj6PywcHgxVkHGD5I84PfNOY509wRbVB2M+Zm4LvQ8
UuklaU9W/F5AZDGyb6zUwKKj5d+zI505+ausvdefm/bPBYVcRST+/UZ+MCa3V29ZZ9oy8XF07zWE
YolaKn8z2dcidMTS8REnt4o+UNjfwb5pgZaui0lX458CeMI3QXPtFsF7Kew1zeaUUcTi0kgkHEOA
w5w7etdwXWbd78CsXppY2LRB1gRZ7gM5YoKLzX1WT1UrKR6yqzEi4BGgRmqYA2Z/kBI/VCM1PsDb
5vIjp/FgBg7nrHq8d2lxj4DUijTgQGTet8JvA5Or9AaXZ9SQ3AZy1UvPdsMC44HXn4CHD+R3rJKa
bNw8qfwT4yWURR5p9OsQKgjw8Z5spgFLVSYc8rNNv6ynWL6UOa9m3k/rmvHDkLVcGQMygyq8S5QL
IILeEXGyuOZV/jfDeurvUeyRjbLvFVtoymF46Ttr6N+4+ufR8eWc+YZy1AO5ke3mEytdJTWP+9cC
gwefgUOEtC/fNr4KE+Tmu/lWPsyXqt+Jafd+qf1oMCfaBSuVZBpeh48YlG59rscWJtzgS+d5Jaf3
goy8/U2Ri5yTwdJDcsgc3BEArCRl/wKf2+lczi1uaNYH4MaEKjV1evKcVYp6cK6yTn4oR+BNCTAe
eymJNNWS9VxvlBAz4qyCYJV2pSYJRpQs9EPCWbQOiiwWbzAD5WwUoRcdX+1a6Fi9XClSzqLt4mCC
wkuZT7OPgUcP5Pjg6vILbqz+Hg/n9gPcp+gZoFCDIJKbQxHU6CM3nC3DAh4UN3EBSKnj1YKfDTpz
LGIHjyzsBc9xk3FyYrJun0b82vJyLe4Pu12P5qWA1CVwjL5aDlmw72pnCYXHU+cCXADhIjF0eReX
IDRK+2fbFvHQ8lwSURtDYaMLnJO6hMwPxdiVnAoWzKnpFfWLXU5ctwbYpshIYLn7ZrowwVoZLuF1
1t88hWFOySPVmukDwzwpDv/Kr6SkmIq993lHTh60gHGX47Nuv1DCvXqEoxfbISutbRgCxImaVsLW
QEfLgP35lRejZtbH/YTJWkl1s8oLMgl3TM/4B3IOLo5WIwWIfTmhKdzPJm2+oW6ZO7VlA7Z3zGw/
Mfdtg5ZtaeQBQdDNs1Mc9WiUa/qDA04HGgA0GAfu9pR/D/J4/JnfI8bA7hFwjxIhTJUS+pD73A9L
FmqM/l9KDR473/HU3y4/YuwXmhBHFIX7rT+pzCSl7Lvi3eAP5b4s7T1ThZ4csjNRrTI76zVPW9hG
6MbYhhLMKiiPmuvyLhKwUiGQPB7dKmVsTSjlCDdcVSHSXhWEqBeRWQscYNJISbeVvDwINJIthBkw
4y/b15sHQsAhKpLLBun23xiClIsLXMnIbIrVu/kNEb2A9ZaVEgL011uKVjfO3yxPtDWfIY7Jnhn1
zN3PGrHgiWah1bnh5KiK+oz/9DxrFjwuFHxH5q2+suS5I3J/oEZMAdyDeVUD53+cmPwNOtV7PvS/
9yCnUzN5+gw5p211tUg9ZurTmfzJzU9OWj5zx+Fasi4+RBnzur9UdJYEtMbzAGPUtKyXNppXFQca
6P5bcQ92RSV0kz1Y/dKQKiFASedaViFnXpAtqpqIJGn7z+6dg5EsORNWZ/z14M8Ar3Sn8fK0bu8K
pvH5ActeLFUMYboIVIWJ/R+N5jVfGhpBeq14P+3paawwS9TUYBGeA8gt6pcGM99+gCIFuzJQbuoQ
btmUhl0bPYM12ZQJjyEv08tZkqNeZFYz7f209zQT52xAsP8q+sz/vzy4laats0kRbKbxJ5kHIndJ
0KoYMz7JseY7h3fbokdxVX79fLRkYiInkqgCfFesxxuV+x7Ky+ElUYQnyNHesonM8C7fMlxclJ2s
NjH71W2IG9rAYZpNIUDdPjM5qK39XG0G/I3cN8dEtetgW/kP4hYnaAOUzbrI8Jm7fSpGSbHd8kaa
9SG4d23rhpw1ztC54nQKc3B8gueebBYTpMIK8J2UTET/xel4fA5MS7dPyGQ0zJmZSUSO0pE3+5Ae
tEXR2+0gn2WHMRBiuLrmVG1J8Z13JW5iQaVYSlMtSkybDd4BrlUIDZiXai0KbcMM1AhjMadS/spO
WrUfMSrl3dfHPeK2y8TGIlEGMJZp1uuq0qsncaqG/oYohmaYE5Q569UaUk6ra2dMvTGluvscAoZd
pVeOYRVo4Y7puLRDxrhcH2Og0QpFOga6RiDaroJoCtUAOlqMdoAfnL0Y6HEf0X9lCTWdyS7lshBA
XhBiJ23tfxBVERIrIme5b+gQuSS+cdKZXAz8N3MFZGfjJDHEEzDQTTZFtw8YYSb9IcwDv8c+Lg4M
2OwEw0UuV/NungYsQ7CBjEs/E8QCSl6RMZe579yLxt2ZfubsEYG4ky2rMEac1tYIKEJm76wN6VMl
ko/Qie76DpC+sviQvzbuO4Po1MvQSDh/WFFSaomadO3nQeMTooQWZ46b+W7Cn/+Ok+SVC8T6KM3k
5wEl5NUXHEBXmV5BP6mb2mV9tItNSKjIXQ+JMAfyET3RCSC5gLEekd1J9eaH0MZHlUdsX7flm+4P
opwxWyVQi7fj4yvYVSByM8ZfJfLbYiw1x5htJjcwonKsmx4PwaFTP6hOhmKjFiVVF7oxr/TVQkg+
gCQ/hcWpQT1TI5MsixN2yZMPEJfgLJHvtQhaKkWhGNyD8GGj5wy7FUeg+ZfKyhlhMhicOXOkRhIK
m0SdZAaWiQJ8Zrx8x/HC31/RpQYUT5+CGCbvHvwL1TdVf6pPeSXl4zkRRp3/QV+Zwi+YkRrZLPmd
6hN4DdQc313yd4TSHa3C0wGBERxSmyZp1Nb0+ZqoN25s/3l0bbW/moHp0XvOeI4pmwPSP+4A7V/W
ZjATFTa7Vrxdjr2pgpl8M9nJwvmpZG9agm16bXzLsUZ+m59jaIPSgML1iHdIbhkFHZxm/7WKIbn1
a1FKtONo4XE0A9MxIEU+vZrb2sSEpr/eD3Z5DrYSq/X+Q0flg6SIt2ZPo9kDhHjNA4h0sqpcT5fX
Z5+Ah2AuWkWAG81TrAGsN6NJQ/tRn0rhR4ArOLTk+QDyllvyJzhPQw/+Td48Z7DhUFwJ5q7/95cC
2VUvPsFGF3Rcec4JDEiBsWBQ6TJUcGfPkMp2K1IbI3mZ5+Vg1dT+eXUHvry8uVsXjLBgliSR6F8P
o1cLKLyrt4QN4PQVGY5t/FczKs4XaXx9Kl5uj/xJGnKP5lcbJTYJ8QH2DFFgsB60wKy4G7wH9S5f
OKL+ibVC6W2/C91c3EyGTbeymynlgYukUOBAU1yr7fjEvJwIUAYVe2zecCg7txZKJ3YQHnGPwCeo
kcH3g02pa/GYVlzfOvRo3/buwUgyt+tpb249DZhdK0PDfV9e30NbHvDFLoWDrLByqcVyTQ/5E+Fb
vndBz1iIgTx3jQv+sk3gdhgkGKQOLQN60Osg4u+Qq+rY4VASoLo3czvMwMY1RWuye3x7ZnLDWmn/
/54DPPxk/QGL/oow5DHlf1XrTd9oeo14IzdaaQGQlhi96yK3NXd3B1zJeQm8kxbZpTKhvjNn2+xf
RX71eoW4LbjX9vIkLZzXpI6LJg2VSIXaA38S+BEhyF+9LEDmjkadbPcjgbSyYdTCD/yABUVrdN9I
FVRW3Uoq59ZLUHXuxXx2Kz1pZ8v3p+C6y/9cBvHiEAVWcJWwIaGt8dXx9nk1l35Y4dJyvYaRUVBG
Qz1o33iYcePKYq6IFo0WFLqbOdm0u9zwT+l/jwiptK5GgxP/WtzrAmH4yzmgJQ9Mzi3zd7DLwNDU
uOpcezLYTsNebFYJ1339NvNxm7IUE7eYmgLCoG4bMPSYNMKB3pQ9UTMIhRci3y4flrkBjPBPn5xd
FizMdcjm3nH9seG+UstvcRDshji7REUmKH/p4KSFNkFy74IpqS+wqGKZCsFQrzKkb16jY1gtOiRy
WdxcXPG33i3tnCTE436F0uqLuiHUhZSlSDJ05Pf+QNR9LF/T39VKleaQ11VKcCxZagWqA7rtmC4j
q08eSGMt3d1tR1DLpxhiYIri/TWVvb46V88xsDcymm8+SB4DD58ifoJSXO78olBCBydSJn1ETQRT
lOWnAqldVYhOJOTS0X3QcKFlVKm0a1++Aq9IhBWmoPGPiThOC1Gn/k3Uffpb2unOEmlmiB4PrhjG
aNzF8eGs/OhwnKGTQv/S6pizhSkhhVVFsON+rbRfszenpcx1GNk7KuIpR6eLYvud3yEeuBXZcqmS
tjPYZ7cjYuOqHt8hNgekQpRCs4X3Wr6UWS8pjZIldpHdVxg4oXAm60SN2KgipCxlhjAysWQ4hMMH
Pl6lCJDakX+6mQSCZrzL2y+YDnJe95VKho9q/wgN71RhRqXzckzs0+G/8TQqNc0eoU0u1qpXFanO
tobsZJ0ALJslJTSDhXn4NeYQeU8l/ZqjXeMf6o33a6Gfi2UpOFwfcpz8ZehnfOLwW/AmFS4M+XBc
lvtvfGyktjJoexvcLZ23E9wTgE66WaSGmXUgaynhk24OMAGL824XclBXEEENUas8D5H7qaAZ+kR+
yrAefMectRa1wmZov0bEithCoVN1Yx7tJ5UzK5V/z0hSS0ZHh7rbt90MoagV0D448SZ04cQQyBQA
kpoAo74EI2EMiLAE8vVjRqFJOcmSYHlfsG7JqZndlweoWpE3qdm2utR3FyYsG6UylkyjaAZMRX3O
jaPM9/N0gGBZfeVhf+3ZVQlXsIgsTpD4r03zA+s4hTKyAU8tfltM9pRXTeERBO6uVbZT6oEzytFw
Yf/tBC+3VNvlbiH7Tbe0we/RtOf4LB5H2R3CP3b5MK/9o5KwMRXi2K/pSAsGoRo1RlHzSQL54Cnc
kxaMoY+KsdcQjHZ0hw3VXaqGMFyKFmfA87t/QLNJlC3zBpWrt/jM1ozHQWzz2v2PR00WtM7eouHb
7MZEyZ6zzDgCObMMUWcKqkt7e5oUHuC4YVSa4/TTcqywtiEZqAehiB+agFFhNVA5LL3Jmip6Erah
tv5Yl0VyUti5JtOfxG5nii96CH9a5x67L62kFEuFXvxdjRsneUxmTV0VyJp+fxFO5p6mmOyzCP78
bqydtkWQBKRvjETNDM+5P9NmqpHvKnnSPBIQ27ra/ehVCWUGS81axWKL63IKIofsjo7ftrzgO8kW
JDGRulj0jRWSoiW7EmcbA2Dtm3nSMtRyPUS/KMRgRLFRrRgD3wGzW35bjYSzX1c+C9mr8iYr0bjZ
WsPzzpPRD+TAY7zSPOAUzv1M3+zbQzpdppx7wZllOTSIC8490GmlGuxzGS5Ec1c/NtlsCcE3B3Dt
zTQWeIr37xBLc99kLm1TWhBlPfD1XNiHWBcXyCR+48j0KLyKLHB6I6/WtZ0zGfomhkb3HGfIJ5dr
xrGS3REDi3YcZzNoer47SEdIcjwbVyJt0+iSCsYmY/JhOU/7kcxv3Y6588UUjv/XJYnVWZ122m85
11Qgmf5VAzmbZcTCAzr4DJBDS/CCoUPNqTJGZy7MVxlE2WsGqBrsUCEhGRMkLoP8+rh2MMEoUP+5
M2bcudiVpBmsrgurN5s+d+A9LYteeIbx34gSq7WV5juSeWAe9m26RvfqtS/ArhvG6cAzgqQzxtTr
KK2y5APaFY1/Hd0AhAk7rNh9uzVTTLuq4hMBRCKvWsM/mtQwLfPwrR69FmBfY2uUPpH6AZg020pO
zQe2YwHs8NBe7DkPjAoHdobKr4LQHhBoeoAvSGv0BGMQr7UjHBgPFNb7tT4YsV70I/AUXhNgngKR
RuUFAFMc3hONTXSolMHO3SB3TDCSh2iJAOYMDiia8uiJGmIb05OeZy4OyNVNQ9FPonInzaXfJzxe
ybPo60M7mBBhxK9oKC66VH91zxkpWkRIChcR9Qd6+yE7ccJ6zf47kqiRlsidBmNJ01iSo/86+Eg/
Pj+MrFk59l1ksTGHJh2hArJMpynyTFycvjTHXGMzHw+oXgjPA+LmkEhgaOsfA4yMZdrUMfy/jINr
+Y0sBLHkeYiKy1+MYDN5VYBHXpc0i1en23m+DlT7f2LihdcdWigFwuw3jDnil2UADAa7/CpJL+Rz
THhuM/NJgx2VICx8K7I+s4aljiZ4yjrOzMrZBJIoxQxgv8U1gJ91fgNKtzXMicYkOegFP+s+ZjU0
qUQv4SvSCgnMWoRvyzztMek6x6Lgu7p/OngQ2IsJoBf5Uq2sJAwDFrDvQE5x4iPtXnOJopuMIE3B
fw5y8B68TfRkiz5o2wmYJZQOoDX/FwcZ4f9oSnj5REyNNQ7YUyYbLF7cXRfQ8Hwn5e8a0U9420Cu
RJjO2h6eZ0pkTMDtKUjC2rUFlJOJiil6/sHddaeZx3kvxF1l2lNWgyB9T0Bg17Y3z4Ge8nHznEuX
nr5Sh1PnDs7nop/u3TQ91kzks8EMjmLpP/NRsctBkAB9ZXeTpyZSG28fVY4ChtZ0u4HNyRjL2p4/
9QLmzkZxnGttkv30aS+M5N22RkMCKglzIR4mqPMmbW8ZyCjEwfivIKgQ8D32/jrjmqnIOjcJ9b4v
ZBetQ95K9LAbgGOFxeBqHxzyH33PGRuFep1TWTNSWspx6ZVzmBXyXF6lAAjUng0nJ3x1ZaZp/5ji
L37ixU0yiuM3KKTs0lcAUpBn53hkbAqLPE06GcJ8V8gZjJ8YWqV6yexPspp6X00otcpVz/c9j6Ff
MLsLQvFKhklx7aDTHY+Nus5CYeg54rW07M+sXeRkkH62QAb/gbCxiAwOpCjk6aBV0PVI1zA2Ry0Q
M1igOQ69tqUSxhxudL4yzF/lLpp/G1ZXXQpAM+nMD+fpzXGPvAi3+D0OqbydawXTrwP2dphTQTWV
MUsjbrINDG1Anbg8bxVRisMY2xw7TWMlokkbslXA6bbJo8QTZS8IOIpZjkArY4uH0eDoNPi61BLK
QvBh8LY6XqTpuO8GsEVAwuiP6sg6niqtXfPe+5asDxrSqot2eTS/oLMJKFIVm3qCJD3rXuK2jJxA
KvtC/X/qs8AnNcmbrAQSF0dxzAPBW0B2QqgxpFYqXBxI+HTnZ/edNYj9t3+zSvnTlzo9bduf7ctQ
ULiWP73pIqEpITSebJXJriLOpEFfsqoomDfjrnSBd2g6aJ1YAv7A7kkkLtYYqS/Q0vWvniRoKrqg
L5mJKS55fjjgsUvUcTDJQEWH6uwtImc5vF3urS0ogL1jeAHEwkEdSjF2JFH18LL4bco9Hn1VteNY
akGmFeeDO6ddglQJ5RHdYEfNBOowOC0OGhF6Plmzu6oa7yNILl6vFNo1WVWva9nrhthOPFBLrNWM
aFehSGbi463mjyG3t4NZrQqcbQ2h3CrTDOfXSe+icJKmc29iV8GCaRYCtk1xmJKPGXiEJSWllohx
xEbz4zZkRwdpHPEi4xW9pLDw6YAnnVQOQhCFwajQnWBhsh441MT7POa2nKbb7CeyqwpmMwpbOzxp
iPtcHRhkvfyDbuKNGflSGUinaeTH5wYhXTSrmV8A+9JdLwtYgX8TPta5QV05iAZ9jMug6neUAQ4N
EVACuKy4s0lP0bF82DJ05UCo/gRyjhFwOFFJx/xiHpyE7y8gmADVnRFZqCvyuPkT3tmLxo1u2YOP
ONjb3WRNbN59mJIXq7N+DvEw6SU0Y+d5ZkpxXBTCjAdGb/L1eML9q7e7QFzzW7jL449hCIFQLjTG
UYHht/RKDs/R4Uged4HPCHlOm0MToFwhYoZE047iIDlqbXyJWr8vrSnQ/nZTaaWYC/2ycX81QME8
AOArO+5yhOFQvPUgiOtxXZbJoYWKyQ6JptbI4TXjjoUHt/IlgoLyi6PuUw+REYKPAsA6okpXPghJ
eWxrWNBf2T0bttmAWdwoutc8OAR516fF8KIJ4yn73TFTCkDvGbwk3aXXKKB/TGlUACIGXCwevqgh
cpQ62PlQZpo6MUu1T8L4n39EpHHbuBB5CQS8577EdgSF7d1DXASN4VvRR4SNNlPhD7rSVmZLTshl
6MAd1caIoM1MpdKkXyOhOP0yoG4QKRs+NPJOB7tqNMVtX6a/5b1hXM8j/wqb7WTD1iqJvkyQNhKG
XHYcJQ58110ChC+lms0SV18Ii26twBVGAOwHX657HjVJmI+7YhjhPWJiDozSOQXgQ7PnOP0i939W
hscL7wPn5GjWoO5EsrE77QAjPUDqxpq/m41+pWuVevjs3eQcnckPFf/bwOez2B01pHVKQK7F8VpV
4xqOtwdcbBHs1Z8coRFItrErODl+/ODb0b/94+XqVgWDggeSpuOxeuVsRAXeIFxsZW7S5Pd02Up+
tyatvaX1lDx/7hT3DIbVsmMHm/QWVqIb8hkM4EHl685TLXHY1pKe5SueDmW/Iy78c8PN9xetsgC3
opkNo88df8wnTTiCFqZqTwEd0L/HQ4w0GSU37mZy+3rWE7xofWEOiqdMXAshm+zjSDmDKbZU/S3y
EVZtCU4HmdhnSVFXej/STZWikbq1q8SIPB3UdmhY4cuNs/7Ejw7sw8LcZfJpmPkqx/dx+YmvkhNL
im22xWnBOsqMRUb8tsFx0SYFQUIeD0vglgjLAikS5sOhErzx99IuXcUDKDZoJ+Mop3pJabuMe4UX
zHQc4Vk71tuaLsP+YXmZi7UNsL0weLhedtoeDc0mmhnT6d7UtFXErAlW+SMyym16w4M/EwLW9TGX
UBMYSe4tx9kMQfRtnIFcsNmAlScXvVYK0dD5siAjXDMDQC3g6qf6qkfUALAMLWiuzMtciu1GA3fi
A+d/3OuPooADPacZHTKaV/OA58PrJIcLPzSE6COod2ymcusWzEQdb5e3rnacK2k12RLwjpUGKwhu
2NnuQeDc2SvdmqWQ0TNlq5+rGQXPYcl8J9SPrO8aFxcSmwBx4AAOvCB5F8XGqA6agbA3eBvI2YBG
9a5LxrhTOecLx00uIIp6cz1fwqxqj5Pmk5G5FvPlvOOxkOJB+8XV8fKOwxMkL2xq1iMY+kBzQuYw
FXIf61T8l0cqN+Z9mMGS36Zs4+XAYQ0p2KLTAkW20Ba+/rg4UI0OPnnXaMdZ2uZRVH95yI+Xo0Ub
OJFT3wlRTXMbuc54xsgIGUjBZkasjocwod0sxTUqwACCQ09UcuMGR7hXaBnjeE/Oq7oX/zCQq9je
2yADVZokmclUzEp2nTBY8v9OPuo1pdbMXah5IpOlRhUIWXh/VpPSYBTWEDjA7TCGo+KY1QOgvK1R
nR8o+trcDTLG3a24sxzDG9iH5B5uxfpmnInyunLnpPPKqC9JdnmxfRHOM+HQPMGO/yHiPdRlmJ9y
RC0yNWD6Jsr6x4L7Wu3HuQY2b4vqUA/cf9n2/sCH2mXD+NUGexxjUDCt0rI2VhXDg77qDXlmtc2P
cTLIrkmx55Ojqwx98NWILBJCQhmSEBbXZ1sikFwiCALhspjimYlDcCdv8OYPO+U7NEPXTOCyE72K
9ELcd018PnFzoiHqcBagqOg8umaW5TRSZttAwqTC2Z436s+WgbM2HW8aQW2daAlKeDjL/u+ORYT0
2uW6exDYYhqgVETao5j3GXHkMcmEQ9g6xishato4dRf7I7GTBylgUjSCnG3WZ1YVLuH2B23JiB5F
zrA+L4UPnOfF/8S3hvnFV5lfsPE4gOgmsG/zd2SR86iciK5V73xYliKbbkmJEVLKMaL4Mg5h+BX1
yamjLCTds8y7HiExfrV3pmArx+5A2mntbrBtPLkWUqKcuawctjMn0Zt+uhIzmListWqF4ftqdx38
XlFEWBgU9SmdC1D9/4VGWEppy+S1Js1cpl7xxC74kYonFyt1O0BhnC1UzarS1Jl5RwZhI3UzFXL6
xM74yhB8M3nVHgWMhh37indwzdH+CEZLFWpz3u5HOlW7yXDmwmC7GN47Lt05SxDd1hmmvEhhhxzZ
aOZ93iePGXglCVBwlX2+bY0smk6YHnuzHjZAWxHrdzwspFifDLSir5URDDYFlaTZzKsza5mNrasa
ie7DZZcJkL58y62gYRLWwMD4e6S47QYSEUKcSNkh+JY+87sh8c7LFgRZee8GgH/bs7UDSTymB+La
a+2uvtp9m1tchxRsxzKLGH8r6zoGGrCtnr68ttYXmALITgV7/UTkZyVjAV/bSZ3lQy2fal57Hcz3
Ru8xZ1jHC5QSqu4AYvkuoQdFMntob2lweJIsLNh8FeNrkF3S1z2X50FeL/Kjq5dZf6cQc4w0mZnI
AreseVUPLiZX5S7L02q2fU8Bnsk2iTxmRJfFGcDnJ089RKi4atf6jk6ifJZIfzALC57DkR12HbAO
rHckQ/NMa0NCpb62ajm/WKPz0pETb9JiVreIMELT+97FAItnRFk/0P1bWRcyZwDjQIVvnPX1gH5c
KflHSQ/puBV2dPmSBhCso7oW7wQvu0jVym85EtZ9XauuoEYLECeTMWvt4wrC8tbzPi4g4nE+Gf8v
3CoMNunq+XolAvYdeORtSvPo/Lyu/6FF390KOg2QXWFz1UwjvqvEH7QcJ8FUuaF5stLuls7uLRFm
s513qQuv7G8Qn9PB3F76L08r8PdEOpGpgI+qIsVskKztUv/6V6DVkhshxMsaVYT4J1ojYFuGsrPR
JjHCsdw3J6JGvh4fbqSkl2K0MKkBDujo3R3CGbKVziD7bmvCH6X4qn/K2KAiytyenwJPtGcNQXCY
KO8mnPqa6HDH5ySL3Rzx1IOxUenfe53qQ7XiD0bgv8YWnSX3BBh18Qmg7rVun7cFtbSHJcsTlehr
QwnAYGz07ZPSTOvtF0tknSar308G9Bq4FIGCaS0dziGVZFqqvvgwX13NGKQoUsuGZx6Fn4TiaTV9
Y5TkZ5Ry9u998qrj62EE6qm+4/UdxNWcx9gjOfwSFj7duVieSIyzoM2POf/otilC+rOszebg+W5L
gs30FTjtyuxGv8R6YU25o1D+HcOkSFWCP/uxWBgz4juY3Js30IdInVKN7RhS0gQGYUWc9T4shoGk
nOy3+wtL8y5CvYvvVEzpHV2wFTzF0F+U34IjbwGwotCvScbAct/XUQUXq0ZNasLs10xLYMAlgMxF
+2k/50K1d3eNoHohdzPl5ua/GDgfVU7/nDM4yJB8RFHEcg1P9bkZ9IOWLXKs9yOoTiaMD5m7uqeJ
aTczvNVNESxNddy68tYRii2xzvYNM5xSGIZH5ZU6Ma7lWu9XKq0B3bed059wkRRgBhx8Aysy6/uC
05Z6BbnpneEh53mo+0o5PQ63YT5G2DtUBmdOF5SFrOVUa3Ri4Gfdj4sPmZa02ykkJ8OYS1xRZoQA
ZQv43hcCMC8uv682LWyYUxN5++qhfWyhAWsH8M9J10vz6jtxyfGhxRFjcmyaZioKdEbaHnEH25DU
vL0Hm1aJmHUngTySNURvIycuGq3kYyC/EAmbKdk9V20yanbt7tOz50FuBVVnUsCERn0nqqe6KJIM
lMWWRIOhgaq/eCC5bCC9UisgN38vUKDhrjP3KqF/NAAFuWByr+CPJLbST5aSAsDoGLJOW0wJeZV/
SzGZ3QdOmR5UCE+63eRgcTzI7Bz8akZw4drjcKtrkBzgeGAu9MoKO53ZbQ6Tg9N2H31Py1F2JpMp
uLZepQyHzgQWRFKxtKXk91guPHTgfIqCs2z+60WsTbjWSTCxkNBY8xKyyP2N5j580OHRne7qqOYQ
4hp0vupEjAxmPyQ38qf9Xejsb7IBmjjY7c1t3odcJ3n6DZaWxYj61IBE3hR8NMtfNMkca/wUTWpl
ZHTIVvGoaaU+VYqf+MYdQjZwIOF38s/EfGq8is5B9Ur/Hx8NIxJ9/5/7bZ5S6gDXbqh/5QIuTU4M
7D8gX1EDY+20RURcGogMGui1r0LzJb//pyT3DN3u99i2jnyf02KwDJ9YyygzlClfGaNY05QgXqhW
2wtlAAtchqiQVDARuz/io1xTRnjsRSQP80kWwYEv+6lsXkDt9o60fNtsp4PZ4O5eqKffSzgKsznV
vkKnm93moDaEt1vap/G8/UcTkATE5ai08YbOs2nvRiPxAF2EsjCAX1xF1+wR4tuB7iB7nvUclf3V
AU6CE1/a/+j85zjVrssLGX7hsZm9WELslwfkzd7oguHVJSo8KDfDsIzd6Pn0L5lCX8bfI4P4qpnV
RGDaJBowrU1bd5+VBSk90q4tUVihMwswuUPR3SU8vf5uI256D/JcE93URzqp4f7VZg4WpFPH89Wx
6RRD264+jtbhLTj3j1uZgt+fTfK5YVQ2jGDtXpVCR32OfMHP/Iu6tw7tKNwcBqxoOf1ANZVGcnej
cXP+iGId3ld8uU+dDh5KZ0G+RGdwSZylx6m0S0CpMUTBtiQNXCz1K3LNeiG6ChAWHwcPBeJh/8YO
JDc5RU1Pzyzc0InWkLcgr0jl0salbMAH9wSH1c+DquqQqwqiOCCzMwLrssllv+sBgXnK+Nok8X62
JWhndRdX0oBxF5M5XK4cn4VYpXkJdJHEs/eThnVe/lhLhcqph0UNiRiFH1Y5NeGUJZabQRP3X2sf
mCA6VOlTHFIwPRe/e8E1A1TZa1b5hiC2HhyyLTTVe4uA/2JMaPnDClO+byZ4Fnk3b7N/SOHwbEPD
HatNULGmJYY+lLF7am4NgvcN0qvTbLC98H8ZFwXnj3LU78KVqdFGC0C3TG5niINr7/YDmb9zVu0Q
c8TH0fRqGcvIdUxzxpWuL0o1cLaLN/tZLjhvBdeY3CICx8G51N5wnHxCN5dUkebENpqgiqu0EaOU
a+k2KOxQ2ET6IdZUknW63N1UGSsJmVj7n3LN1/mcJ0+tLwuBExOZgbIh+g7xBu5ZjsinHw1yONJh
j0zPJ2Oidb5JbZzUCe6xvU4oy1QlSX4AYJfyjv5YDczp51GzqNuzyvZ73JjJx5r4z+Dt5jHnQLAL
/D8jHMrk32uRhWrVmY+BZxx6JQKn6lYB2gTsn1bozTQX2n1hFLMoFIS/M3Kaql2f9yRo/aTU3OmB
nQLlVApIhsMfIFfczcv6IoJynYRFuoeP5pXM9Y2+tPr0mGHOs2DJm5m5bk48VZol/0xMZ7Ru4Ak6
lNwUVQ6Fsh/SXmQWnzVJFh1sffGrHfSbGYHq/Ngn3oFMCrpjSypDk/l7DOhFyuoTlF7BmBggnzJ2
FsaTcAUD3X4KURLVbnFfQcscy7sh2siyo5C1xlRFYbrSr0oAbA56bI3ARGzuP4+/43bPdXcL0Kvp
soMnSzjcHS0wWkJw/sUEOqtXwoQKs2mg8uJteimOMGDptIJ5+KgrUMXlSh7vgi911n8RHR6c3Tmj
dXz0Npcb3vW2mKfuh7n2Rwc55OXFysOYdF0MGFVJenLPPs5m1S6tT51tThzxpq6/QayzjKHe33xt
3SG74IEls5CJJpYXLbSi6zW7nt7mOmFHNmaEZYthw6PAArjbg0w0yXVjpRRi8ov7XqpeuGsajKPj
aFlK1CP1HFHbce2d2XtNKMhXNnEMd/+P/XaR8Th1YTXDTCI21CB04uQfUMpDNyNugBWM49yCa5NE
gTCz4gJqkohe74jTsZSXLUAOJ78Q0+SUTZf8rlDPL3SobQpIKnNmoDlFyxwPVU7uwo76IJ4eJ85k
/Rlxr+bzoSwCnrv28VYSy9fqjk84LdHAkW6Ur4tY1HgNixkxRgHIUNPOgwr2Y/Sv9OiApFagwysq
x03pf5xwz6umPrMSSkn843syCDVDlkSetal0I7S+yv+/Sf5jmJJiTPEzhhBvrV1u4wBmqjHVF/GZ
PgAC0smdCTUJBKO+g+OFEkhlVsrII8A7qRPKozNUT3swyNJzZb+vDN5SCWW420gboy3YDY6wFmzF
YIxY1w3fUOM80Z7KpdrZ59Dh4v+rZGHLmugN/sg8Jja5Rgm+GOsUkzUdG09hqx78aO7cR0pSCzvL
l4xw7RoYjXBANmNhu6oEWOMWHzVqft+gFB2u6U9dlwEhnqUXGtIT7wnWyo7dtgJHQvasYCfs6jd/
z9tLhu54merNtrwyNMyZkJmFbl2/FQX/t4awtfdmzlmbQU6uLqa/RHEt3vyU8hdTtGMSt1Sou0ox
Yd2imAjXI7onSp9jD/DSUk3C2DStBmRffG8kEMvNjpunmJXR9HJNDirEIeFIaql+PulaqGwUnzHd
qFSlj8sxFpsnGXzp/yrKhuS/Hh8nxeZty1buZroz4XiraOVTskHs5F9bGrMAMnVeKMRmpm+GXFZT
lORWJmq0HmsSs9maVcbC69usiXKuMdLOf2KzgfIvVFYnqfdqa42hGmBkA2gCE2NB547w7epkpCa+
yfRX7Ry7EJ4qh5rCc8DyorybMMqC4LXXbn4mSH6fLnpFWr4H0J6UcvnaNdT5xuQmag5DpTfNBp62
kL9W141NS1pL79+sGZ3yzVpjJRW3/VVtiXfmL+G8rw68M1Dl4aHaGjOfaumTdEbnvJN7I9ueyKNL
zaSgWfCzZNAs6yoc/uG5uhi5mkCxxvUxz+m8wlOovNYiPTIOLNzG/ojEhqy6ve1LH9/aLP92I+jD
skh/pTUCIGAd7++7j65UVOGmTHnqg4qlXvFZa8Fv6485I3LpR8yTY6U6MFii/LrBGk4GQnmzYAzY
NYcvb/UEKqRBm72GNnVAogyMZ70427CIDLoTPSHiFrPhaKcbj/hiGBpHKjDVVY090aIHO0xw+cf5
sTnlGA4cvcl74zlukb1er578qiFC7toOqy+2eJX06yZPZv60aRerukXz7BSkTVc71nkSekpLjvkv
i2xbS/F2lxm2aCQUsaBdkW4Fa5TBJXHUKNZyrQQbgH2Jz0o19ZCatXz/kLElyvgEpu00NG0LLhJi
/f6XgAcdCXdgkjm4VcWExm4wbyfMZ2xVg20YgwwvD+9JUMJiNgFPuUm31MIWkESKN+rG1Hy6og2Y
j42c0WnxwqnS/8JvJoxV3/1gDxdt74NpcY5zs4Dp+JrGaY1NkhB89m3aVJibDBVIXpJBX0BP9dUM
TP7iCHmJekvmiQR0glWBYK+bzzggm4kGj5IPLGVZv5S9ejYk/IWaHzRXWAbXGmw2TW6ml1NO6toU
8vjP2YNy8j/PVYGySiezR/9xqVP4vADJTkqBM+zF4s+7wHPwmK72mfYhtRUh2/eWPagHetfMA7r8
qdjEfeqm1bfqjMoRCsuMO9zVH3+wYpgCSAM2v0becnBC1hBvxHFXyHo/TGvF210/0lYV8lupBIYk
wbpN51OwMlzOFzG/i9MJ0rYepNKi5E0gTmoX3+FNF4PYlzNrnagnlGuRN2Ryjz3U75rrgSXKDNKq
LY+/6UrhGiNtDtPFIBquTnUkOWJNDFRnBOBmGeZL2KY/mG8SHyWgqKPZyzXnn9FwvEZaeflCiPXK
YwhtsOQhbLPfQHiGgffc2q3IvbELtZEnkafgF225ftztwVALFxwBjtmVz5YsuSakQyNsHx5d3r6Z
JTtC1ssRXxoqbw4cwoXRmcesgUId9APNdLAAkd4caBYvY4lT/I5QnO13b3WW7p4Go9GNIjOb75UN
lPQ0J7+EWcg6TgwpnkLC37oOKCbeRZzVxzSMMcoEgQGEk3HOK7ckekqzRD7f65nJyKBb1cNlIvFw
nvj+WM+e5mosg9qHPjIBhIGyL9qsB0YqzYOQVtvnuxC6IXaKupyIyOuTBe7NJxjcnp3rvhRG3GoE
ciA/mOWBEmb/f+5LtUmY2W6mNZa2Ctun8k3ckOU3wgfisG+DhnMFR1GFfmuGQ9BPsv3dhBz7DsF1
MQyAJfMWts57iC6oyVsMhUFQoDpkXBrzUvUt1ndgzLBM9DiVA52qzd5ICBIeG8YgIzIlpZ4JV6Mx
ub+AykIkgCxV5X5rrhHIRLXVt8PP84G0SCZQp8jg/m/lfo70P9A8rbYHIHINkJb7C/rh2gvqo9ve
1ZF2raAX8PROrClFdvgzdTy1RYXtI1mNUzceXSlvkA4XT+PtYJATed/gEueVskqmzmc8TpzaDmh8
v1ZON5P3q6d1eowufl6tJNntSk5xWM0o1mTA1b2QPfgEHOrOgYDxEslWTfhReiLHcr9tPGu4fwp8
fTd19njdaa0NJgJpXbxGweHLqBSHOIDOIobI12I0YkzuUqzrXoWoNltEBc/Rjik7370aRvItnCSn
KkXE1YaCqJT90MCB5B2LHfU2N3/fy7wnOKoS1yecnO7EK9ofWMvZSUPfyo3ERk3rxnRjsngE7Cmv
1ZE8XK5vlFVfFb+0IQd203t/ebTgQ5Gn/G2Xkx0Y/vRjka6yzNH6NTzpazxmDdO+Em6hyvnM1brY
QYTKA+UllXf/wpa9RT/buutCHGPzIu+0QLCXW/71/tS3Q0/tBKsiGbcQ6mwcmmM2OATQ4eWEXjjF
V8E2+4Ut2s+1Vy25noZY/PNjyAVXjVpOZ4K5TfJ13JxXIjHA/PMX/L3RE6eIyznlbfJ5lzIey1Qe
NAVFZ0IvzB1mcep4YB8hEaTDSb0gsSGfroQtFTuFcHub7Dq+PlY2BXF4x9aiSq4+Z7aOSPscSyDS
ksaZfPzreNM0NQevZxTUkTVCyTdBkf9Pjbu5pqybmUJ7H0OL6q4kmH0jbgAkbrAeavRWo729FZK3
644IRsaroPXf5n8KEi3H9ruGZZv8iJz8y3VlYXaXkvwFQr5vceFDmo9p4812fhpoOP8nob4qMuKn
ZmxJ15e3Ue9B2PXQ1U6c+XhG6tPkjj2b8lZGRUtTnccO1tpBXnZIY6WImlO2tZe9iXE4wxEiaEkp
+3zwFH8KHzrP7kG/P/GLHd178bfZzt8XeDMStutAybDj65iONivFrYfZo8LA1swVtzyhk6L3ufwT
MMjAwmQ72FuwH8RM85vRFQRC/ctHY9D7Q1XaqzEzePTCFzlVITtBXtkiDmg+AZ8uV8KcP7lVoRX5
dEiKm+U0hD/tozjQHNR/QXQj2bRnTWPt2WqH4XFeakHEO38v/1/3wIwkd6zzHG6n8vn7c6KsnDly
evI8p/0oOBrsut7m46vIU0mCtHfao237/QHsoekpBN3v4AVqnIrCiLbq/xManNu2p/efB9GdgrHx
en0aVxK8DjG5F1+qTa+lwKkbZdNLvMTDwsLmBihyz/EG9KPuuzoMKYGYnWgFunDTlb7XIIupxePf
hMcMxdsqLjLXCcvBu6YQW7XFJrW5H56eRipddmA4nY6De8HMT3L5PJHgmu4mN6VZYficnRvwsXmH
2Ue+n5bexcrF+ziedkRZ+GzzFj99sLjV2mPviFHmfcE/Si2ZDUJ+vAYm7dli4ewm3K6Z193AWJ8M
ihGs2EB5HBejgpDOjVglGTZTyZ8SJXWbqo1aZ2qVBB0vYaTlPJ3AIuVqcqPWsllqsuo5i9abYDDL
Bi3bxn8Q4AzKE5jy1wYnmq4QvvQjeAnomp+B0NCUoyarECwcAd1Gq1KrninwRdFkqiW2Pesn5bSu
JdEkLtmrbIPIUaG9O46UvcPEGgZck4ZcVIAoZrpldYtnQGXbOECSbsf8KUZiiIgUSI4Hlg4UafAr
bEhKI44RNYy7EykP3WXzjs9awFYFfcJS3KhxABLqHZZR47YKQcWIdRgk6tJVKRJM6ET63D0dtm49
1KYtH/oKGodEHk5kXQUfL1973U/jZtBLEDqgkUNahm+PkP19ruuvRSCQNRXw76DjBDc5JmIjcWRk
dyxY67IoUvz/vD88iNlmbL2PYPB6KV69VpUeRz8UjH10wA1oRLymYkxQy5sMjmHU3gziH3fxWnIZ
jyZNBvugVCaVju06GElMnVK1DfGc+C6OPjDXReVFg2NOo6/zJwmFbJhgD0QD1jnUNwuItw42+DSS
Kt6dU5Jy3Eo6hfg4jo1S220C7ETs2xUhNVnz0Qkq0NFMSNNmp2vAFgsFjv+3qf/WJ50W8fwlh7aX
FHTIn4eaosY6eDRhiCbtrOaMdM6mfCdkrjoIsMeAT5SEaF2I6j2JSeGGIb8snsbsebTcbdR+msg9
2lAM6JHS2KkWezURlDJ4zRVNA5UrLWhmQC4ATRjK80q6dEHKSO3RAXclwGb8iKMhsxbsQKI8pD9L
AVDc/tsBQCm6kIqbFQjqIfiMWmCO8IvAlhHDnuJFCUTR3LlXh4uigQl48xwX5PITSY3ppGLINWM0
QmqfkY4q6iUdUldvJuIgx+9z1ldLmIB2pqn0zdvJYox7nVHwYXzkl8XNjT+BiiWkewdkG+zzXD1J
P+Z9fQrdPCIoDYe3drdk3N69J1hb6mIwDDgZ9VYFZ6xkK5cKHU0+HOyIxgKpqjlfnZUHBBShlTnX
wGNHTZO9FNI7FnsBBpTIWJ/s8RsQxVU2U+BIh3PSWJLsHO+R8G8TM2rjKayxnRDG/agRGIq8IncO
JDNBduxI5VUhPYuhAePz5opFydVteKVp4g/np+fORzGIIOeGfI+gmHcESNqs9AAiiB3jbFgOnBsc
DI3IuKTZkG2UJ/wfJNIpKmA13JfIVEgG45z3pDENvvAkI3LBoMjzBP2ERFrD88uGZSrAu3Qpbzmv
lfD2yQ9koqZMtx9sNCpdN4jwZADeU34pO20TZLxXEiZBcrKaj0KS6eChDRZkW756Jh0LSvvAqrLU
QV3JVy9mgLbbMZyGHlO6FX0hNRKoq2KzEilAcuSuhRUgvsRy8aiCBiLaLY7K23K5mere2/OH9oPd
A9LOGuDkTQRXm3PJ60j7pKFkQABqEoi2HX2nPlSDNtruJLrIMs8XTnW6pp60NiW/oKapQShFn6cY
YO5xErbj4JtLOiYqOqYokFnlH9/xu4wHg8Vpz1fb0ASqPyzIr4kEIzgNjeTezVUGgPkPm+iISBR1
hnMJKO1rXP5lj2EQuxqgAhf2IBRLvl7XmJ09ZDpuXAxejHkvEVWSOSubmYYHxO7b2FddkNEwXah8
aUdq0VgTgQ6+f70AYfmPpcyad23xEuQ3df5OZw4AUmQZz1GJ9rx/NewXyHrhwwNTGkTApFKjW2eH
Hc4EXdY06CMDRWgfdsSFZ6NWJMdxNUMaNj6szX8GHGpwD8VXvebusMicSTYXqhUtiQILIIWuopJn
MXrxsQ5FbOqDRr3BeEl5nzflly1XIQTDdfe4DR/QPu3Lrzm2IEdnnD/+WZUrNDk8rNTQM6RuMYJ3
dmLKeI4erNEnYFZTa07sglFnMyRNZ0Hy3HYi2FAuBZSAEyaGxw5NtMMjOuFlLkpbfIB/HLtSN0OB
G0gJu0M0bgypMfGkHD5CszGm37eiRSkZhHDqp58dPjxIGc5cY5LO77Q+KSuAgWw3HVM+UJ9AVvcD
H0Okn/8ARHhHJY67MuV/iPDkz1+VZs5UEBfEo5ptgbQuYsmbdF4UzCwF3ZSvQehriZholFHUdysY
efyB6p5WUMSk7sYeuCyFtwzDfjJkLWYcb3P7lvNSqUpGXxsVgtZslk4wP0Vc8XWONqH94wnPL8WY
5iOU7PfqGPBQ5p79dXptDXlhRdZMgldq1hj0alK7FUmPcFqU0JQ/NkBN/RSv1iTQQ97yKH4rwRbd
9S5VgOs05wUPpUZTZjR3uw3iVOtKXzPtNjF/dzQuuIMJ82Kv02l5Abaq9KwbXdkmKzYPmb0onpjq
ab302+7dTUPwgr106hDRBq7P/UOW+9WrZUBL5CgxPVdPCsIEzcJr+BLAYXXD477iNnNSmrGOrIyo
UCxclrYigdbMNiNJdA3PqbTw5wvV9lqQa5D9KbS5zmJGk+sYyfSXYJKouV6GftsQsC5FBiWvJBCv
/cEvDBitvHllnmNAoSRy8pZEvbLw6CJYGBxCD6/n8ngQBqrSwUB5t1XZ8Sc6UVUUq+B8iAhgZBRT
4dwazIXnuYcaILKWzaj8wDbpf5Su2XuO1oXbs3ypz/29z4CUg1HPkPSqnAA3n6ApI3Rv5x9/gC9t
wsT8OpjlFjZgxxfj5jh53cCs4V/x3woK7k1Gm7afauQH2XgMprekENYv+Up33vKXLH2ScAvUTelu
iHQKh9eXEyJ3kNlk65tbiYY2mBaia4MxuRATUsdVvRbPaLHdLybZBJ9bd3nH39ddI884OpFRVQVE
fMilxuVwd2/rb6VIht60QV6A15y32j779qhWNB7lgFZPXw0onTemoTe7lJLK+R+V2/0gF3hzqMgj
zK6P9jq/bHqOMeyU9TAvzhFh7Fjwok+RZd0y8pOZrDOAG1M3AEzB2K5qqNqfxAv/lTsuHg/GzXxp
Fuu0pzlZTXGoVL0KPswt5XKf11Q+pXsozEMUvNrrt69Dw3FX2UlmVRG+meGYk5YqnxgH64P1+1Nz
DzfMiDwNdm4RyJd8t88zwEbUeQDhhrFZA6WCWFiJwoW5YIuy5Q13Uy4ZaTL6uiKej1+ECeuRd2mp
yaM4yJFXMp5YFLxP7lX+cct/GySaL9kKPoiho70VRyz8MN4/OqgK8iuFLbZVONWc7PhtvBqHzAOO
86P250Th9YQ5zDfZBfIGyE9x0JGtjp9j8PvTO5jzWVATK+5PPRaQhb9DMOPOwHcc77+H3kzcALEW
x3hCL4o4yfnZ/DhQezEjghBiTjBXaiGWl7igmlGilwQYqP7dLtDwxBj+b8jh2G68ETMZ5JeubPdb
qwesgkdZHpwPkpSwe0PsEbv7hTaYPCnqpUOqjr1foJgcXQ8m/l/08M30gmF+U1D/b3W3BcvpyRKn
+FiLFpZejuhkHDbqBvK+UkWvCYelGMPTIrSc/fSOYddX3TtZ5POUJCTlKUizt8CUvC+T1gDoP8mk
YZIlC+pFg6iyyfeXBBFPEUyj4M5yLiIJMpHke2VbS2Tv7n04d9oTeDK8INj1Q7P1AkgpkfxHZqFm
cD0XYcxj48SQxVDkmqBQJ5jjzlzfI0HRMIAmblJyiEF6v1AhY9/162rJTqfpLGisiT3h/U0X3L7M
xH4+wf8agWZk3RklS4SK28nXhBmMxaduHdmvKivpD2GsgIxgv0W9SiDUQE8/DprN0oLrRd4Kurid
kA3nqzXtv8n2iFgrkBSIezURVq4tMky3z8lwAz9A3kCTS/a4fHKU7y1G5Z3NeeAvc6NgeY3hp8kn
Pz34OEd3FG6spdJpP2JIsXyEMG/wSL4kO/hprTUCXllYLiZHNK5rl5N77j0X98139+G8BjjZX2Mv
ASwyXlCfnQ8RuceZAOPA3RwROn0gKenQcP/zhH0woxXPTRyt6Sto/ONXLLSRZEWc6wEzF1N1v2sk
4Yn2envSAAHsaIjSRtx3dyi+tjzfKmsR9F14BLmsNIr0F7uF4qhZniNaPR+I0zFvLPDFagGJedDt
FMDhUl9keKZaTdv/fe2hEjORQ/XHHSrWo1C/O3Crh7sXMxlxLEbskOorE0/yOG9dFCSaJ6w2sCQm
3AN2wbqkdvpzXj2oV93tj8X3/KYkGOMaxtxoaGpTfBJoEUaDsIpo3/MAmssSSLhzQ0kBXqWEfW0Q
M9IRo/hMJ5VkO9vSBIOcWYtPIrDS4KuBnzluiAOP8COTiSo47NCdiupz8SHXoBvV1C9vMqVTWbp6
t4CipEk3To2OH45JfFA3h8Kpgc6T8e7lVr3MiwHpwkLMdbKciRTrOSbeoWp21VqJlzahUx1BJ4Iz
SuuXhCGqa9glSYTPwpfyIBESQ0wQls5veCiLivFolSobs4j2+rwd+K/5L0Wyco+nLrhgN0RtU/cE
5+EKnvXRWrJhW8kcROHEw1G8C5DEWjn4JVEEf/LOZSSp+rm/0NwL4RNI+M/mzdnMFpS1nRuMDAIM
7gDORDjE2rpv9tJOaZ1tSxjnzAcRCCKISPu9quq5dtWcT7FIwR4p0Fva7RMkQuiKiImHndjPDXA4
mrqxGnl34TFIEtiiK8eqrfyqT+XaMmgm1eQEJxWPdbcqPp8jMLcLumdb0pddu+UPZ5eVbVbD1xAQ
3qSjmw5ROP42quwmC1DfBVmmaTkSXBpaTq8Gzl9r0zYMEBCSSB7ZgJXQoZfSwb8nMrfqX+QzPGhP
flE7LAwF+hTE/l9NVCGQAHQhx9huyZoLTxIsdmTHiYXwTQfjSRwvRuSVJ8o7pCnwlbUnYijXxzvI
iVzIvBpH25iAW73Ah85VEwSqJIgenY50PU9qgMuKkaWQcxaf1XR9GlXt8mJfNXypCjFgqClyt5oY
e03rpD/n975t/9Pw84iIZXujzBNZtwScYC4wMWWzJsZLKzHvH8bsrEHRefth2qQuAG4f48U5FQMB
l8YNgDDHJ5WLx/hkumQoZd4uwRVMLzT6AcBIOFL0pu9TePdGC5Cn2ztIHOTqkzc9AuEvRPllJIrE
EYxfrTvkJv/Nu1fDqq//dZRSLxcK7yr0yb/lfvbI1Vpx5uIxv/9loZrMs8u87HdFQFD5veGIFgjV
hQ0JZw/QSxQ3FqQXO7v9N3FbozK7dU01o2n0kQLoMylozUAXJqw4zI7HB3NHF0EWQrZRko4iQXEu
sSbbcjO8F0FSyxKgyZ7ur/PX4ngLEXVPAh7A7IgLpbG60zIkX2JePWkDuowA8xkAqq8l5MrFjNeQ
yv6ILh8v9ZAC6TaYaPnNKfnJK2V4DLXCnahgk02XYzPtJTbRNhWEgWF6OWHxPBBh0Ln23cpk7Cv/
GLC9D+SYaw/vEEzdF5DMhqCy0yIxznHw3tpIiBZSFWkLEZFyevvVEx2o9uhpy0glgvrQtanDUWvr
oSTa1/zf5whE0sUIuix8+mCrhm7oLAcNaoIziGKp9anNn3EOXfruS/JmX/d48gKCHgboAvwXwpU1
t/ziLABxVR435MeK1qy/ODy+gB5Xg+DcHFEubXEseDVRgW4qTWYFUbj8XxDWrNTgnqnUfiMJGG/E
CZIyTpzkM0oRmwMtc2MCqujWCzvyn3eTr17qv1EAq+gOYdt7hz3Pcg86kHvx/u6BCTuPp8C1ZLgR
uX7yDiFSXQjpnY7wPMckif3iLFgrJmScAW6fnS7hzVYqkqW+WAIXbp8+5XFuEbC6Wf4r+zfdWTbk
yYTE7ly0ydwwP4uHcgbOLLtSqYWvDX4xYQ0ZnpHjSTIAp7H673PfWwmpX3cC5epIvMLS2FYIyXry
8HfMvAE7IQwnrVy+CYz8RLEskj2NYP9ptj9WNkbh5w+izkXQeSktgpAMWHUefULN2W1yolv7snOu
YQmajQNWWCasGyggYgPnRs2U5bo7HMRnxF6qloow6sIg6/Yd1q45FXbyl8cfUzjk6vQDV1xmuUX6
73lDoNcgNMCp8t1xKcwwVbqNGuZLowhQzOzXaHkkXDkWhEHSR7bJIC7iixID83rhWro0ogfZ3g4l
Igqv3VQru8RX790iCWozNjOwsYWuquDkhe5JM9BmY+gfcf4CN1gn6R1aoAwhGg+LlI6gf34Topl1
qqVlgJovtG3VWUWYimEbhBIS0QdCAGQ8aKdieLXYftfe8aE829JKw4b76DBakmTj6rysaoB1JRYU
Wh1EVwArw7o2eXWuVw8dhP43CrLhwiM5S6KrnB9nJOUwKYGniIoZ9cJkGJtV/D8r85SbYXSGFxjP
PxP7q5JACijDvz93g3z/Q/WzatKm/qBRnhHVObJ3nbGq49QC8++fpU6/Hmm09FDS/JBGMC8W+SH7
zy6Z25Q7MonGSB/4/NAdf8Lw3K1M1/yewOhz1Q3o9FhrrH8t0O4GOIsrGHWEZP3ujPIsK/sPpLDC
pJ7iHR4AvFvrc+bW7HfrnLi2N7UBfZ2AQr+r5AqR+FfuPuq9L0OsYGuFJaiYH5npjNY1wELfDtNp
u6blb/X2df64n3P/Niehg6DPvRuQWh5pSlJz1DmB84rtjne9HzFbRKNjdVmGX3yA7XWPmxKYxU/7
at8qWMBzv0QmN+/+PHUBUgmy1DYQaaFXvWakwMt/BDqqv7TWC2SfjuIsOf2EOch7JzCGUzI7Pxy5
5wgMeVzDygLB4OCYoew/WP06JXcu4IvJ1mRC1gaC1LFeDjmaW2Ve0qblzGteDqo4ceZ9Xu2DduL5
vj3Nk2pQgIYOS+plAWZCHWXaulqmVAi4NCeuGlB/QjKVjJLhYGB/LxFBrHc1MHjvs+e81RN6maII
xXLDS3/Jd7SOLp4Ky4P1bzhMfxKtK6/75HgL67MHnG52p2S40IHaYqBu2WUgKC8d+MHj5R5iDw+L
/nQiVrqvy8ToCfNwZQhYVa2svRFuAJLcDUvTsgS/omR0Yg97SmydUj1ExE/Z8rIOuW6873UUaUw3
5jFj8l3DUXykNNlfF1BndOOWuEu00aLNDCNuTFSNtyfGeQc1P58Cj+IxjYStYMDKJWo0BuZRdEwR
7G9yzFmLrjGcM94TT2KuPaz4IEzY13ANbcHUXHgIQcJILrZWl2K7UhYZv5/GEJ7iO7VVQlphowgz
BXvteWfvoBdqpLtbrHsaWzESwQT8HZkWmMvSd7xcH2ngZf6JFvkHsqTM55QsXPlfXJy02l4O1uYr
pksjdZDivwylaJ2c8QLWENuFpSB6miCMBqAJtGZ+kIrOP8bzGwmcBXSdClTbzbebcYl5qOIdyTUJ
QCYHyB4ETgjMghC4sHl+cQtlGDLEFfuTpyFYq31QhNFLUecsqVH43SS8VibhK9E+hcOXyp7h7S+B
/awh+w9Tr4V7JuSy8ZNDYLnNLbkSYUELmJW7tdKoR2XOPoHoGx/qIUnU2XifJQ5VMZRaQsw4wiUx
DpCOXGTo4KhVOqsTRmMkCLyQbtiDVcStVkVZLm74VYZRhcte0KrJ2VG25vT4o6C49nIRs3j0PCWT
vU2cixUWl2hG8KghNhMVyvemlGFwoEdv2FFVvUv98jRhKkn1MNh0OMm80Y05o2ImTsJjJdYNKlMX
oBujBZ6ir19rh5vR8m/RozpmdYleIYHHMJF0if8bHlOVCSdImc0NfGsglvjDCKjjLBZZbE4URzyW
ABbxhaU0c3+o2c+BDhTkprzWJEE+1fzJkDqXUYD2JGxMV8z7307I8bVYQgghlEUi9hklDGBU7AI8
CfPC331sbrmzY0Fn6SXX5p0SZAbmpbP6JazXmR4R7RfbglxRba6bE6j0YTzDOQK5bVUNaTXfSXcP
8g5YDavOsBy3HCQ6wIKsdV5IuQ4uT7F5wG+uh2uPcuD2b2IcfqCeMYuj4oKmI5tYTvFHhcqsIHPg
6pyM86NpIRJ5Di+P8+LYk5oXWsrDmV1GwgzLmduDcyYzE5VrhioDVuJCuFyCcJCD1uAhOx/LV6Tp
mKHl45fCw8Qskwy90PAb5zwBx3XqVil92KN4Dg5pExrtujL/4ab16fxnAmPYuMTfM9h0q6jHVJql
EKbuzCLaDhwDzlYqJHr9emuFHlImUWglPYOTdZjOeAmsu5Co72BNfH7Vgafb4/5bgLcMS0dZ6ryl
jqqJ0svsntX0dpzbVXqBw4Z68cdiiHstnol+zn8CLr0yJDxHpAJxK56PU/BJnwCiCMjnjhESWNc0
MmxTnsuTCCOmyvbpzpRGsy3gM5RmyloZuGJW7Rig6pPTT5e+RYqyPN43yMbfVk5OZEcxueRl8fx5
T5GD7Pq0NuuwaKzC59k85h4KpKGbAyY4IqJjJKBQK56PvjGY5g803qgFk4+0BdCacClJ3EDY64mW
fAGXmPhpbOzV4W3uuU2V/rfDQmx75MfgDReZHKP5YWirVI2wsdCEm3/wGHTSCIUqCKwattJsLljv
1+bN7z8xfIVcKdTSQjndLic9nRu0qlmMb4VQ7KgXIqAcl9lvCZvdKA2EzkVUNol72/svA/hKC1sg
+Qriyj0lv4++Kl822g6Xy0NkbIT+MFKfKEkeC3ThGhEvwZsLxsaGqGjVH1TGlBBDcHMCVtQU2dAj
arhq0Czi1ldzzJpD2w7AFDTRW6xLjKjMaQaFDPBFMclzkW2y+MQ2NTzHKGMJTuzZU8OCvoaMSMFg
gR4CXo7Ku449afpyh6nYWMx8dStNvUqbrMLNiA1mXsgXNc5ozjtOAZu/Dem/Z4DkRw0IW/Gh/NQo
sLspD51uTYGj+qZYcbyQYOBQAka5wN7kXb30EXuWGI8/0K0yXQ/xMetHmKFAfAsjRgl+zrt/Vg9s
QGG5OpiIZ7CtWB2xuQCrFc0C4A0vyeARiUWRJptunM4eIIyp3chemj0ZLoQTtJND1ScJJRpp7Y3G
AuPURe7vK19NyLWgpmUfLFKLTnLEfTiUjG45tjqcN9xnSUrXhjo/AunOmJdxu4wdUSkF27YzWG+R
ipo9LtVtR9ScbbFwBkJJ2n+WtGluyj3XPo3lOgT0DkS6DKFJv6h23Po2eN0ZPHmnDPgz3EyUkWqB
EWMYkTCdx9W6fFd23B7mCVk4csfPsojAD2WxUK9dp02XJ5UPfKowVRWyw6hvJqNtGfWex2MhYxLX
hjC1h23Crcf8b2aa+ErO+yLkrDr2GzKqVjoNDzSD2kXEh5JECfEzjtN8ePlg1NFWOufxDiRkojjp
nn6Q6tonXMQqbsGXG4owu/s48F4Vpcjt5Sm9T4/frlAhsWj/9M2BBZ21GOjXQUZOr47TvniM68d9
qznFIBCf1NBWlACahvZddsSCl+MI57fq7xMxMl9xWgu4aW8eWPvjEO13mv0fRirEXLID3QspqLjg
rgMUQn5coT5KOyr9/wnW6A0dI6vcTQ2U7UIHgeCOcZ6ya9yNmvq4EmTus5MtTrylC0juz77XNdFA
/hM7pwDiGiAO2jVk1E/cfIXDGswRXLdoJ68wfYwDzPXU8oZ1Llo82nEpq4QBzd2Ps7Ygv3QYWin7
FZHwhW8NAQZObE1yIChUMT2HAXMT4sZVBvsGDameAE4TInOCRAcA1ae755+YNTStcmOvNna/VmEr
g5pE2UQn+vb0uLhcwmuVPzTOkJBUJaJR1QB+gU+tuOeOPnDBUTbOZDxbagn7XAVsIOvG6Phfcfbs
AI9xMQd1N0enL9rwwwtH4/v50wO6o6QYxPm+nidbklraKpRFhchzD3E1LFv84Cane1JSAr5jxxBJ
iiB8DiawJyKS/qaQkR1Nu3BEI0171BYnzSqMtt/Lld0BUmN7+fVkZ6QL061drmycCn8QwWHpeCep
/XuTG+uV+9HZZ4XyHpj2NrG1hnloxRf6ihctQTXuLop9obC8KHSHuycJ3Dgdbo7wzbKLUMM+i4u7
iAFqfPwC7fA36OL78O9Gu/5DjJmPdWVpOWnC3mtUzig/jCH5E2B7GooiStS0VtunJ77Qsa18t02s
nu7H2HbrDWANeQOZzsKbFg/jh+yufH4/La6S1IhQ1iBTOU0E7L59KnxtaoseHLlEScAMsXz17nmD
9HdjezzFcwrftNm3ulj52OtuAgSKmOz7VtrUKamWXNPAsTM49N2LhbInrkdHvBfgufGrLT+mExdg
602QbT67bRDIjQyWtZnj1AEUU9CzyCAr5Ul1bHQyPkqtWr3k/dFS4Gt34L8ldvM4ipYFQvEDCRj9
DaFzwlQBWN80o4tSLv4zzXaqwQElnBnG6RSOfntvZU+IW49Jpf4xpfEtw7nBHlCYqUOPEjpbSG5a
w3JZJDhZz0PAFYWX7M4L8eyql2jEobDkEz+SZNlkncOHQUBM8A24cgw+gosR7mKWES8bjf9U0d8S
73OyXILaSvonNrVyj8+7Je++GrblWpR/vBZiVpTh249bz0Krh4Dv5fnA699IxfiFB64/qlU4pK5i
Qoklysxh2vHM/WjlYrYrit4nCWdBcsYnxyr+q58vZFG/ln3Z7ZSxRjG5/w6+nCuAteWx4mLm0Rss
h7wTjxGfwuu8WSv0qFgwMGOc9flB114uxRU7ajD3CT0OPrhVZclgkxGPOCR2IsKltnxP4s8cOJjw
GTRvxo+kwm1+J0EBbg3Lex3tvJf3oXgcP1XlS2OccAoQJjN1/aPJjMV5OL+RnQj8OPGfT6gPTZ7g
nj+Vm/8pDtwd7CDc8PjC+giGPnJfxrEsPVg0513f2AdrBOAwqS7U9ZKcxL6x33+pVEJfqV9AnApc
KYbwN9ol8XFiMxWsqNgTNTNDev93/kS/UeCNKjPztFoSTqsaIormYlOTa646IAs1hZ8b6qgyAkqq
apvhNHlFsE/VzXF43iSLLSDqFGsawBVEsisX0pykNjNnIhMT41+daUljeWoNZHXYog8jeCx9fras
cEc8VsuVrkk4+uYaYAJhIB65GDHXHiWPNi/iiuQ+naKeVvunXjRpF5KFqc7GGynBvOZrZGyl7aEi
+4vR352QwQhozInSUajs8wbNsgTfGYf9HjtKgvUz/ux9Uvke4XWEdnjE9Y76WXzk8xHy6NLa+ZHX
c1ToghEqO3qVffNiBIuHE8IsRo7V6ShwreoOs9ui9qZ+1TkF7kE7XYThqlMO/M8L5Dsw28htHHfG
B1SsUjogqPpzo8EKREOvydBF+AZhbEN23XhK/ZQlGhutjIQoVn+5AJ8nqhEhn94pWaFvmyeo7lHC
2XmPmhhn18kzErF8rJcsUkfxYDlPGJXqDbOx2MI45i0BuAsvm+QdWdGnIDZV+MhqMJkioPTQC0NH
LhJY+VlOh8JtaIYKpPqvPKaNSbpA4bKwgpAOAbjNg3SImTVCVmOHTlbcxn5rHrGqMDT3VU2r8RWM
/XTdwTABgWMTSAzG/POTcxp9O7zbgMOoCv7W+gbau38B820a4VFyq7veRAPEfWkomYojUdO33Z1f
nrbO6BNGkLgnsGPualEfjUnpAoce/h7LUAM+6hCOFOXyozAHUPLbVjlIfw7Uq4Yb8MZxiGw/K7ts
hFgQAMi/3xNt7sL7nlJxhX1MioOnFQBgEiF/j/xpyUSSlDeUfw96vRCnWZyttVF1TnI3ZFyIMkj0
Dh3dI+m6171HRJxn7f0P5YMTGk85BJDCNiGoq9uiLSg3dBJeqVSipJyt9CEUpZrAR71kEv+64Bw3
4OjVhi+q9mglpbzaJr0GH/2CvnRBw4FT0DUqDb9g8DsvcHRi6Q/5idOrb0303gWsm9PzNUZ7tUw6
FQX55mWdgYslNVrR51yV+fGmCC53XL2/X4r2mVyahmJ4Mafb+Utgr5dTwN8YEKSLH0rJ5S2BOlY3
wUJcu2G0Zy3uGwSudzTn2vp059NnwNOkmgWc/snqIZgSPlzKOeeotjnRPZdKrTLpRQbiP/6M7kRW
qokCIpYjsBYy1SO1JBSqRKUasMU4DFd0iCifKXxw3WkRua+MfCnfFOIsazu+0R4Nv0VwW0HtY6sU
NDNfG0bzyxEtI/kKjsxyVmTLCNAAFhPchP2RJ4+4bhNSOaTump/MCh4/+bxAxhod4Z8JDWJ2l3Rv
fbUp52hPhWhRdXPAZNlo15e0/MD+m8c4UfQmeHJe2KE0597KqemraO8YTue/yJow1PmPdkTOrCeI
cmpAA6CEpCOYjbrJo+5QYNa1jZyAWXPzhNal6Vwamw9sPU0N1Eh9LH4mrEzs7DBz9/7/o5/mBePS
94B2DUfEF79zkuNRIineuB6YBE9/7GwIR3I6Sp4xXak7xb1tRkPQPJenXdjSV2HdijKD2G3S2wW7
fmt1W2gEaQGBSGgcaL3vvX3qpTn/0rwI2PBFut6Dmt/U2+KKZnhJeodSbPlzdCmwZwIQHWkca+cr
Vzhykavz0JShPp8pFo1Do61co4oDw5iPvd7QAVEv5O1CcTRz0cVTHjVRU+w/PrjulPOw5T8ZI4iE
MrWnc5T+XxTL4R3TVgSfmaFYwohLnLIssVGanBrcvXpvj/ZmqiQXXBjm+Q9tiH4u8iMQj4fEC0G5
Nxpap2b0pxbZnkGXoA8FhPZNl/xR4wu/o4RnZZaQa6zic1DSyugqTVxN1XW7sMiAY6aYlCnpqcYg
4F/BqFSX1r1oAWdv1cRRmqTZEbmTuzo3+7v/5gM1QwdpMtFueEzG8xgsl9nfaD/WxLrIKylJXj2J
EyT5bfTVczE4s2RkKruI9pkEQTI/XGSj57jMCUbfYtPPAKklSlTGDe3edjQanrnYmv/4W515zk2R
2Vktmo22YxwxskXGVCQMIwEPHZdr9MfQ+ANccAK8ZlrA9rEiu5IBd+6G2PaoO3bk8cUQ7p3tIdPu
Gp1XM7UxUQ+zH6WmngLuafR4Cl7IC2cjBWOdltivfWlDNPxaWGCmdsK1PQnFpOuwWzcF7NRWe9kO
6JgyDetqLRm3OVG8Z6aWvbdr/rLlNMXw93lNTe9n7lbFrUwTrOf4V87kyBsalI/XeP1q5VtdLxoy
tfiqc6/iyXkFWT48yxorLXA/a6qvJSlW6NWNzwIdBG6n9KBnBlgoHfwrHidcWLMrWWo4M1DK9jMC
Vav5s7TbW5UAlP4XwQlj5mH0cDNs6XrhzsDGhKDkEMKG7msVLHg+CnDp8eWtGV00+vAu76J7tEQK
H1iWLHotjJo9ENBrPf/bUAs3GBppZjb2EMNxq6NyMS8Lf2Fb6SL92tAbMYJYnfgc3L2fqeIARDqw
gcZoH1I9pQ1j/IbXpTDUmtVMJua5c5OQhemVTBlIl/nu+Uuvddh+PA3QGnOKGd29OIhQipGDnt5B
TGHLKIYkxzln8SwyWW9O9O7zPOBLUxTUEhxsBDd/WK5UQgAILgtmsAtKGMX9yfQn5G09+RbUQEBv
VhY0v21vdWM8sz31sM/d1vX9m+nacoSzY15FLxqX7BHpV+KYnddhuyx3ksD4DCiurfPjHwa3CV1b
0dNnnQE1ubnj7HOiRASjml0MasnJKSaPe6xF6xVUbysoLuI684owVLzCAaCNkN0iJ8BeNIblK1wV
VahXdc3NHS0sXSYLVpBh9rwcP2BYLgOlysbzpXue5uCXzqXWYYIVGdMcOGhCmCBKLmH5WVO+iuzA
WFjZdeWF42cL5TDJwAgt4S5zad/yZik+QWgvcjk6V3Fk1+xIs6Rx3WgvWfVXbrGDbuW+RddTGj88
EWWhupC5EeVtHMMOrDhkIyBigyjL2MVFl3D5DXogSpVB5Bx6Ojrihrwqek7IHzFBl70jsNZtsQ79
xFFRXMQvqrATq5Q3jCv/TNmzYOIQ1s9crOe2XjBewnD3vYOFT32zOa9yHj5tESWQldPkZq9OHnt6
uGGKs3U0wXr7ysqNoXl2djl8U/1jvQAqVDash7TQ7MlPrgHn4f8Z6QBV0ZMj2UCbZ5U4dXifaQFu
SST6qmDLiBI6zLK3Od77Q2fL46sJ6oXvUoEmltRgGxxUZKFsp0ZbQiMcEwsUUAF/DTq01f9j+g00
g2+m3qMwgXQcoTppOt5k8Y5Vy/z+LyCdFLrR3uUlWCvGNvA48/d8rb+ysG7d7R2zvfMe4Vteu9BN
Rdka3Lr2swQBMPahMDvVTwKu0yaAjJ7xRNOKSuLgxFK8MBdNdR2fdJhSvWQ8mtkFPeDKOQNxoG0R
DXWbqs4x64axubZyp1dx3c86lLYicSllt6ufeDQl22dUEoR8dG9KiBTxeCyZKM5uOJvwFFWD/Ci5
c6AlsZjwrypS8WNGM0bn46mR9HwLY1iJdQK6xx04DDT2u3uP/SXdIUP2aoB64hmU8rtYGpM4op61
vjAmbQzi9tGCHhtd/O82dsiqDVs70KWOnE6Tkk9H+fjkKfN5rfYEpqyscU0l6GV/6Qi+EYt7hn7y
S4K4i2BlfpAjzMRs5bv331d1hrhsm0CZV1hU3Jj/R5hEvbzo342a+kXjyY8J5U/KE19BS+A9howz
JkZGdaGs/oL0jl84OTSW+VbLi0WaGDIdP1OKNkoESQZLG1x32ktLsXX053sj5qK0+OGe1Ll0XDIq
aZjzar7kZ4FVgY6+yLZKcB2f7XKDyOIL3X8gc6+3gFB3hbgY+z2YEfoLvu5cfFZFuvFtSJAdo6+W
66GOr+Jx2kaJVXsd4ERBrHEuPD4/jf49iEeeZH68hZLjyH8JmN0lPLoLaKzg7pKZLv2/HkHTDYCg
nUShZs2fEvfH7NC07n8JL63M5tOhR5QChNBaT3XJauEyfM5oG13tfH6njQ0F7i7yMv7ODtwQNlF/
/WAGxuzjA25HVZPVV0kikbOcpgdAWNJ3wOQuWrXee25RLABLd0Eq2zTfizaT/wV/mBm17eHduNW3
aQsiKA5OytjBR7JE14P7P/q3zMb7ANK8qFSvlgBXVCUPDDtYOzQYNNgOT2QlGmmnqFD81t/H8gGV
m4qDb/3u6GTm5NBkah0AlfBUG4qlAWoTnWCGCAk/ovoUsVWJ7B4bpnXshzlipodVbLoyqiho4B4/
bKBsNhi4U1Op5OqYE+IBZZfTje3P6Ret0gJN962TqjFayoa/VCnlbC3TTDdZ0PMiixZa/Vw7WUEI
0pSGPqVHjTnUwJ7Rwkl+VmzvfHF0hMY3vRQSEr5LL/nO82fnekXT1p6kL38o8fqIAVkKi5jZgXW9
J0SigwmGai5GwUDB/Xmmn0aCGHWPvfuXaslHfRwowgYc/XpohJNnCE0DuVc6t8+lwg1W6chBNxXm
D66oh0uLnIns2Px9tTu9NkKADCHZWFpXrKIl199UyI+lx+uUi50Rr1u5anbkhfPdIyTckt3SzuB0
tZBdR4U2/dWkKgxG5B/JLVZRaYWeJC5Pskara00FFuqgZQMejg6DVpzw6lp6kLECW5EAjo/gpXW4
01ceqLB4m0TFjM62moEXj5aiqI6MKtfHT2OxmlSgRJftLfcGZUqYNYFPnYikuqARmgJD3eWG9f3A
wT+T8kkOXUS7HXq16m1r49r151aL4jFY5bodD/1jkb8ILA66QkqwLv9Cbmo1zmgnghdaFTRyoov1
nRWUWRb1f+C9FnxGwliTw0G94JiGHcmSMldx1VNeU1I3o9+f3jk0Uxo5MLMRFEIudCd2K69SH0jC
Z7/D90OwSBm3TFQg//DEGkRXk5UOtM/NzzDp2hTVqgrEviRvLzXotxY+nLLi7jLHjE7RVxNA6aVl
Hx2uDREd0TdWAD2hgIaqHA++tCnlxxBGJXQkUueM0XNDKFYV5IP1MyUuta6zH5pIe1BzrZwhmp8H
DCGoJqv3sYoxrEB5d4NDtCl09xlxkz8mKAdCTiKHlpleyLIYXFy++RBDl7IPAIwr39pvQei326Zw
OKuccb6daHl1oTFQYyQYKUPiqXvcQM7mUzUpV/qhKZnyrf0D/Qn1gtVXQ6J1t6XX0w3NGxYxQ349
BeuMV3GIaG/9pCTrA/wqYoujnFdNi+5Bx6RoAZegsmvzbE9jLpk97RviUeFjyR3EnZeRRUOTfdjo
oMvfIwX/+cmQlLrpsYPBMVbRSFdzmPaBeDaiz3cRFy2ywIQDVuYlOrTw+XvwMQ4eMyQv2SJoJ02o
g/y+pC39JixFv9Ur7aR2vB4kpinSEeFjQ77MAPEVWd3xReG37oDsYZn0mkEiyQdIZJXdwEAacj3C
6qR6pfqg+VvMREKKxax49v15BWaT6xML5pnjpUd/YI47/TctODNsDJsG5S2RSLY0ZAhTG+lcs2M5
gwa2+eO6q0tuyD5AlkQyK3S0A6PiD2Hr0r5nWbmGfUDtNzq6qV2x8snasERQ+g/t4CZ8ye6lIlP7
yGfUbNQ8RAUi41O/hgbux/fdSm4+1K1bydPDKs9ykV5ZBiJ1A58FYZCF9HVzOx0BvGvPJB1bkThb
EmHIA1n2uAf4SikF/pVGZm1R3XPJRegPHARhduTxg+GOCs8EZuhRCDH6CWNetYd/lx3mHpOGuLsD
EarO5FjTE93BSRIOZKAGlgPodJu52hLqqKfg5VlzMOtPK1LahVsptCAJAJSwiDFYUoG/4hJVSkDf
PJ2C0yR66cT9WnrrSVuYceK9bhQ7iznZz4ch3OvRHtPEVmyTgsHz5dlCKj6Kp2MpwcZvJLcBtU4D
6EBRpQJdS7lDKN7N85d/+ucBwxjnrMOzz7FiAhpXFcPoXgQvnk3/ZAgq0SHo4LwbanPTKbty2zsH
j71rxKHvfiVRa+Ew1aO7N4Z2bznhZvJRoj6Z6rs0CdPXkRoeIqbmS6lLijCn2ivwPFHMEeBx4Olf
h2ebEUwh2fXJSjTCSqLJY2n4pXvABiR8Jb5mhDDXU1vDlS0b+bO5GqYdVWUOf4zfFfdSQS0m/gto
9lgBf4RTw/aujYAwji/J2npPES2RJFxBlB9i4zkFaLx/0PtdmCGFJlMeVdeWx/ImbqKRY+Kj5jM3
TEoAsthvQV98qOJg2qcBs7AiKcR1XkdOYt1F/IEQjnoZVd1/YNz5o6fBsSO5ZfX5kORbZO74l1to
9iUV9bh7kkrMdJLaWXMNTcFhUxYtX+jQFoCJCgRmUMtPFw66spdQe91GG3iQhNwwM/O3XjOmwUX+
Qmbha3K/W0UtaaxxpQ0pNymDYO18iXaTvkkVHDGNdC3p+gFEodCZeTSKvJ0xAqC9KodkmwZv95Up
p6ezhAV3IPFnFcxJz9mszqztpviD1LdG0cnWR9XRRavc4cqiBmGn2TFh6U57evlahG4fn4KUGn6+
1CcF90rdTIl21w23iGYmkA6LIgweTHdZ1WzsJag0H9ExtO0u3RPJrCP3EceR44priTgnwiNkCJw+
Ho61wzkXwKedfHZaB+eKuRnEH38Mguengxl0JZNvYEbm0drX9tEHs3ZpbhO/zOlDPnHaaNREW+ct
VeFOqNPSJPVxSlMW9l6dcY4QfGvDF9mAsO4u3oaYwvn8L5t7XxHryMpnqKBS+9sIXbQqguwTvZxq
PlEdHECZ9OujvbDWqBMZEhjY4j59Gvko9pXJuimaNXaV77tvgO1JLdMF0iLaARPkLmB1wqwlHYLw
Lo0TIsK7G12cKGB6OOJzZMbfs8Ck28eHeh2NWxy5HuoucGSGN2xq241ePsYowFulsNYDcwiv3PqF
nbwEgWGKifiIH+iOeLUB32m18y/IlLLf7atSxlH4tKmboCNqX8gVgu0lGvNQUQnGsnFfjgjOX2Xu
DCZMyl2MEGQLruatO2XVoiSVedL3gX87bH4xN9bmgY3Z5X77j8hiNP22D655o6Ha2KP3qo8jSaTB
M/eb2wHUPJOM+l9e1Qsg+oKu493G1sMAiBorw5K6v5oApr9WtZ0ff0fR3fRI7TmZ9fWwwSfhgGqd
7l6wLJ+rK0n+eBKNSw+EhjOx1HD03qVSdouZ5jePyfIGelffpcwzGuT3Khdj1lNxEdgbRrZWnQ+W
tsYWc/xFQxXKBasARfr0cPnIDKQaibTqa4+/jr/6JSEwGiiPuMf9EDPNN7YOhR6XPIBG6OMmROVy
/ztEfJaky8WBquwHTIcwg9cwVhqaTlbey+eUWpwmvvpk4TYtbvBsMjXsEnMqasRyriZivasoyXp+
lnznAvluJ2Z5paPFPWmn1JPykaWsTN9E9GGVFCY41uypk6/+3FNjAjLYc6YncaUTFtnT2oPWYGXx
NZWrltuQLBPtcyxNdCFN2GoPLC2t6sjXairGX7kgRgsTbfdgBMLL1lCl61S+o79gbzX8FWbmdC0/
Pn1SlUVY3toa5M+k0r/WL7twrbdpe+QYfkVztVI7iWioznqFB/gFgZFN4RZwM5jYDxpWDkyINApy
+zNc7u6j5VXLntxwFgHpwevAM4L1T6iygnuUxHDIWeBDnwficGeFgd2eHhRqyymYL7Ons2HqCgAD
RQHQ1G/zuO/r+6KDZsAox5zhRoqiUhL2bs86ionweKU1MsliI5EPLhyHC1ES6XVBJp7+YNVvmrn+
k7HCxAL+vu2wGJtCsrIvTmrtAh9vB1v19KVhRujB0N1nnIz20Kw3Fe+F+en18+Q2kD6dLxnpp26g
2EjK/I4G3dU9owClfp0hXgJx1Rpfh5wfxXBEd46IT8Q/FcsINX3XKumKgEvDQP20SJEjFQ1GpPHI
pNGfvwD74WfjUPLum+oWyuPnyPLXplQzeNPJ/j1mV4I8TIe6vJiDuXYTQE/Vb63T0gKnsaM/WJma
hv9m0KGThdSJutzNX1G7l05jT54sPAYwtZhHV66/LmZF5mWZHjBsO71+1O5D0XjekKyqsTwhXQLP
6cDzcc0AgYZqqr2xLo5F5SaeFY2wrfDjZl2v4Zti8az1bAYIaEWnEm0VpYWhaR3sBDjYffXLIxRu
Pv/MZZuQ+dwRSIsX+m/q92W6e9DRbFmnj4qau/aoDNa5VPYH6fD/73httjSCtW4uh2RgSalrn18f
UROY58ZOjXhLJKxnpMQYWAk8CH0Q25tFQuJO+Ar/D+DGO8hkKNRYQRsKgUhv1GTHtzdfDGMVXHwj
5Flholj640uTWv8keN9qLUSmAwzO3GIGnl+UrdxmsGwumS+j6Q1zwQizXJc3DH2PpXtBxe8q1ci1
0P1c/1HBiIpd7cUpYnIe14Y07qZrBrWzYIDwjgi0XQkjcUmlzdTsYn1AXQQznVh3fL/FZI80U3DY
h3r387rNb6Zcs/QoonMsfz4/j3BuCaPuEN5biTFUw1sinuzLm030K5mkplySSIBSm0H75XQYa+91
77kxtr+hi9Dz6mXTtYaaXlJOfjTZG2rg3rKzSWvw+kyU8po0oH8gCBJVD6Cfe+L8SLRVkPmT7Pjo
DK3SGuoXx95qqAxdJ6TaFT/llP+4X/T2e6moOUQ6CavG01fyLBmVMzce9Ikz+TgE1Qb3AM9qG0sp
O0Bnxu3Dw1+GmF16S3LDy5St1YnDdu2CFLgvWEOUNnmjcMk/t9WhifX47m2XIoc54vdkC9qqP2g/
CX7MnM0xDBwuEjNP9eRBjB0GQFgfz6EV8I28FBPK4CX3iHLq0cznsH8rNgiv7zXNxSdlL6XotbQd
JEJpYwg2UE+19piuSyy8kHgPNqXeII6UwgRkY+FusTjp8ARi4GRjaqMzLjAoAeKZnAmw2KyJoaQM
qkAUSH5W4TQqDzvWqaDq9D63pibAClqbJMliLbVyrHDYYkQziucNm3jsWRZJQA6MnIbo6ZPvP7lc
a81xSvxPmqPF2soTAOWQ25tpy1J25Xl3BAlqaOB8iQcBW/KoGMHAl1M5dBVpCCc1sVbYehXLBUpa
0EXjDRaXVWr4rEqOeUHBRyRltWljuzjIE4Q7X4YPMKoxQUWc3hmX4dlDrLCSjdWkmBgqhkbRkSFM
LmD3ZWOfJzVCHtf9bj1hKw3L9wpwKQAJHn2ckh5lkCxE430hkc4YXJBY++SeRb8lpFtQKlbl59py
J4qL28ks2maPzkB/09i+k+VQYvdOxX2yHItYEhgmt01oxnEryjK+rdn4K0ZfSgtisjWJoSuFFoGy
AyHA+uA/Ib0iHq5n3TnPASrs9CJOTey2StRjAJyI+YqavV00ITX1lSmONMQ6ELvpWVGdDa9Bz9y/
eeokBOoGG9bL0b7C79P/kcV5BuUJPlrRd9abuiH9TvWmvK4w/XOvdFygsctndjQJv+QhL8BN8h6d
Y6/Nob2Y7WvevaFrgy7x6EC7ZLBf0KtZEt3/tzQr6mC5pFAnL+eKqZlLM85i5FpAxsayorgCnZuz
TpCm1bF/3rIwwZG35V27yBJ4d41Rpo7XcwnUaVQVorDZjV3wu1b4PamtYH4Clx7NDWHYR+lM8NQB
KvQutCilynv0wbLSBlGm+4mURODVT02tTQ9MNiLU+rBkAcF5e8CcseadxWZWef+LXp5w4W19gKMC
Gzhzgq0UZNXGWlwSFSd9v0TkkNqYptXudlyupP4We0IDWJWMZP8Wg8VG9/pxSJxPvl9BN7jg5fTQ
eDjrULtpzwEdA7WmfjWC8xNCGOR0iOx1Sn/xACA3rB6M5qXzjVMkNACYsXKBh1mPE/If6F18CO1I
3EYBIvOShKzuRhCcCDpjaNMMX3kff3/ZUjcJznZi3VPGAYXBneS6PU9iGGOcGjxdOWsKcXGAUfSO
AAD4B1UIF3AtgI7PADN9UgBN1wMn7V5OOOYSw9b0zqXuxgVAV+2p565UtRnoirY9Avx4Emy/DSQA
nbia1ltlUEtFDn4er7D8bJuQC5UjU7I2bzXuCRg9vKck5lg9WMJFF4cgnaoK2b+AVwiV7mZ2iK4Q
Gkjqh59/Adl2GkEW8zRlkfUkAEa/1SDcpqZV8qsGBWVpLSXO+Fv6zvbp0uR8XbaZVdKIoMuzyPtb
MOEHefgzldizRYKHId0hZVy2YVgvIJrMt/QUS9R6RqoXlsk3DJaKgwqx0KfgkRYl7Ol/+weuKeib
gOPloIAnsXzJegqjUcUDNPDPy1u7YjikqMlnGEztQq32O8nSFdIhkGy+c9dan5F23akTfVA5/WP9
mBD/6dsWKcIrnZWpPfjl/8wG23VCxAyhfPOL1JFgl0gVOX4kelT8R9Ke84YHhv9SxY6akJo579oB
2F3w/+ESnXmL5LFCQ9Jki0H0pf2iPYArTueHVW8ulJDzco9c7Qbo8tToXWCSGSSR/6z6kl97HSvT
vS/xAs09T6PT6F05Se6b3WAoKa1ktSNm+Fx/aFZvZqdhFhA7T9xuXCjD9u3f5UF0M7/f5PBemGOW
LxHJwTIzHg8B4mDvppRyRZYQCYdrF5zdiBLNhAgRNssGYtLCjmLd+3uf0y6fp0PgYGtTAHShKXUH
ehI7i2jULVuvihvIfmsu8UvBjwGRxGGFDa+4x46NxdyFGGZO7H4T1lSSsKJcYWCoZqtx8Gw4kJ5y
4L6SvMQ7DrzfYwfVQkQutHf5Kvi4+tAvhiuJMRAg8D35XejbeUyWNozHmzQL462wOh5PhV8MEWyi
46/esaczqTKavzDxaizxe5kN2ndD//c8TH17AEmDGuJIq1hJvlQ8MbsyCsHomcW3DFOHSahwr5zc
2opSXKSYUjiiF5nDCUtjyDzqV/c3YCiTLKb4Qof00AtsqZqXz9QayQwajwWVMuX3ejKv4Ymtfl/k
kLK1nUxbalWv2R1bifRSKe9Zh2rG7PXo1pTkEaFmhAU3pX6I0jbIkJoOhWXT+BagdiRKjcqs5XYe
x7t2s4bot0F1+MPqDcrchg3UBE7exs+fLOtm+jKGfZBLcKfQhGytgS9nvCS0SHx4wo0ei1FXmSyk
qany1Svfl+/8ZjQDsHktheD7Zsw4r7rbrerFwP3IMqFDB/rDGcyWQNOM3Y9CUuuY3uF8e7kkknhJ
TUFW0GRWSY5HQoQc/fumWaDz6IrmJHv/cQYC5IQDyfn0XS22Lt/UeYdTYCSTnCYDdM5RUhd/zsVn
E+NK2v4kwCKXo9VZz8mgSSsKxAlWGwWRURaVnuwh9o7bC6AlBgjFs5XjrhserAM2xDIIq69Iqr9R
PDQOfU+2v6aSP2278l8PASLjf+bDxwKiclhFy0PIlYHByTGZQlaH9UUkcQUsL1qtU9v7ZqxA2xLS
E7qWkqbkMwwZBQJksWhLaleO9GYKCJdVNU2hg1j6EVOWZm85wjturv4z16weSJOVMiwhE2AGHWqX
Tx1RzownsJ0PKFvGF/tJVQ7D9qSG6ztPfHBnQ5DHXuJNH0KbtjnUQs9zFO1n2toJmpfS0ub7sj09
FbygvbHUvO5K89312lWano+0I5fX8g2Sn86eqpRfpWhXSxElvR1kp90n9lRINWMoH6luRhH3kskp
vULS+D7ENng9RNUncHA3Eki7fJeFQz83EHgMor/P6UEVcYEbfpWa07ec0MA8ph2qdkPgnSSIdmQW
15aWJgBX8dvrP+1io/Aj/jwMFXL2gk9oreTEXTxB4YyhZkHK4e/fQBek9GLQwqcfTlAdAJISHyCN
Ng4joMBYdOxY6zDUbWrMSr89SbE+RDaMTWN8EqbIIsQybHZOT0W3ECJppstC0p53Zavpb7wzVICN
u5J5X9etO4KeI30zLMZ3qqcTr8eRy8fUU+55pJIz+wTAJn0hJPhWSms6+/qU0KbDyy5vLok2Huy8
XJpu/xx9s0SpuQ5eHxCarLBoz8BMqV+8cr1yr4ZM+kcjnXnl00XzBie37dOA/Ic8s1dox9sFuCNp
gwLbDWCeBuASpunGbkYIrs3TJ193yWXxOprLU/M64XqtPbCB6QyfbCioGibiD+WKw1qGZueYH5Qs
LJcWJRqOY4F2AH/hcBe2XBMsilcVTPPfxf5cVjLcEM8CsvUygo1hQob2IPI3an2lPSBtjb7pof1+
Coh9kb8SztxYgqW42HWAZCtAGNaONOfPKvAx//QxhCSNCil0IN8fVshc8kYH8WkHVTFQjOCAnbzk
lF7CWOT2o0wRWROeFlGusXrImgQLlAdKFZ1hhmluhXoZ45hYNgTQlEXFt8mVmq1eplpNYup8pOHL
S8bVpV9Zs05x8OgZXeeT20B1I0a0WLd0LAt5gW3DqmFMDAeeew6Fk7im3yI2AvHZrqm7d0Zqw4jW
WAyS7ESGbYwIx78f2s8wBqkq2MQuRL08p2CFHoYIHq/3G7zKg0X8WX4VL+fPa01XMQyF/6htGvot
EFNOvcmfXvB1jFJnR0TWgSYhp4SMemi8GHWEU39qfISa/w1guYq9GUgC14XJ5+omjuuZCdJbmDny
TqwvFucULbW/XDu8LaLwYPf9xu3d1vqwLvvaTJdAjbInFsMaoeEuxcjwZw4x2H8Yuqkj0cz85MkC
VARzl53gc39KIzwYarJgMFBOqsKOsmOUjNagj+DWl7jxhpNSOjfVGvKBvjQV4k8jO9Q528nUoglp
iemGJtIvGUHmWDs+9dKzh7ixZdXVElXWscBrWajIF6CyWA4G+N7dMVRSJbd9LyYz1nGBQANQoDMs
DEsoR9frtgNOeyECW1waf1bEPMEqHEkPZ/rrWx4oA7hNO5QVBSMza7WhjRIUkNaAi5Cg7pc7vuVv
Pzc058LDPZQFfSLpode36yhfybDj8p78Y7vGW2ECir3CA3gE+7WjBTVie1U2kmiZ1H7KNpl3yExO
BWXN3OEDZhINDnSe2ISCukAhoCI5g4wIMRrTdyd1bUN5odqFTuTM74b4qiLS8DEa1Phjmfqmj/ft
I43xsbfeZ88J93qB6lMpqPeAp+wPQ/++VS6glr4BHpw9N/T1kdBI0inbkODf9w3DjHFJEJuqvsBm
JHZiSGwyomKOwV74s9PxpW5q0CUVWLyOerbINz2TeNS/J3hgClUA0rd5oAet/gjJqDV6SANy96Di
Svr6n90yCjfzqm0iIMRr1SIZoUUgu8NiSmGPjNQwQNQBRtGEKPMlNlu/0fTD3T+mugRVdn+rfJx+
KBCLL3BK2MJanllfRkUooKi2LrNuhIJtEQ+amo8NAUzSgiKyHDTSePSFb30zX3+e4K0Fq3o5NFyT
/aGWi6VmwsfgpcCYz52QewE/QE8Ko/ms+fq4TvqOyRI9JYDTnLhbWyfBztytKcUHLezmktDTWAjn
qcja+xdPaUl40h9BtHmXKhXT+mI4kuExTaRKDNV0irqnDf0ax0VkQca4sqdz181nCdmiWDhCkwnE
JYhLAcl2/NsOkSNJftSeOSKOmUwqZgs4gmz2avvTWExtwZ5QMGr/ecyXXmKwOTRO1utWqmqUIUBu
QovmdFjN35FynLdxKROT7n3squZNosV3gSFBUh2vOlZcvlTKDyJaD0daRPVLrC5gyBBwUslz15nf
qgF92tsrb3dOf2VI4sLekUnmD4ve9cFK9gtp0076SN1+KA3DjbGkUYGUDfz/+ieOZG4lPy9aq6VG
HUKTBpsN//FGwp5LZJkeklcRevdsqOw8saBdFiXHJ8lC4ohuUUs44f3oJb4Hwz8GKZ+aiVySP7mn
TIUEtEoiPKC6vMuKGb16xld4/S+uVYqthrJoNDPs6S/m1QeiGbJq8KfLs+eahBw1v1wy97b0ItX+
Ysg8Fox8DnjpE0+LfrtSF5e4aA7iIqHH+5Qufh/bUkgitmCCGRvNo/MThTBGPIKrNxpRLCeR2ybD
WEiQLILzqXD3MdVd2C0hgF4M5YtOVnWmgvTWDvY0mQsgx2zuNOuvEqrlNePBqiH4l+boGzTlP8P9
ttrI9pycqa06NDP1LAzaeG4J52s1zyLMkEdzGhy5ZePxEx14Z+qy2B0ANAIsYPpq9T5IBckSohzF
Rn3PsiBPmFWtdnPfvIkI4Vmh7uLhPUSlxBNzX2/Dup4vM2Q1ezO//RsbFQfgWkBaxdkdtkAh8AK/
5vveTXbl4WZrSJBB5R9X+UxcKDMV105KJtyx7qfULjjkz2nRWJgmhBHZqNQ56LT+nhltcOCtOZdh
S+bhzRHWgYmN8mOm7x7q11QxkB8o26ldXlQnmRtdFAcBKa0S92n6peUEXbRXm4x+H583d8GIlIhr
xAcUX2mD9ChGa5DRmeK82rE9I/ElR/qjKE21UAFy3m1WeSRBDretJ5fElIJU/Jg+kHEVCEGB5jSO
C5Gn/UqB6Kec3I/ZDms7GqHLDapVwIfjz7o+5/m4Iu+oTqoka5+2C9pTvMZvamLOaDuMVW6UrK68
9EWovR6yF8lPQlFV4NV2DZJeiTFXV39ctCM1v/dSfenVnkKc24Ny73YFC/kbPmuBD235wJE+4nM1
xdL4eWQIENUfAPy1CgZLzxb0y1peF77tHLRywG2qRjM2jxfWrhNfhsMxIW3dNQmbc9veeOEm2kt1
mzOOrltFRWSIfVsEa/2lPx13JyVK2FtBVUV8iceJ3k41k4u/8GJl7TWDFKjCilB/nqVKU4Q7ga7o
/2kEDoNbA2bUA8hS1UumDro9rgvoc17WyQmKldzaoWYLnnpWjifGemj5LjXOFGQSC/ASZuRtpJml
ynMu5XCJoi+xViR3JxEuI5yPLvPbY48V+Jh6eAx0+buTuudcP2Cw8kk8cfHvefGY1zXmVfNPPiTX
lzZE5hx3EG60YRkfNzWhsjVdmLejtouMVhDpcgZUds60M4SWe2C/hpkhmKMAnGYgtPesLXMy4UJq
OsbpyiNcfRvmss03tf8EaJYAanPBvWdWN38/0svP3yfkwW5A7vlU5iW6c4uT20UnKX2AB1fOLLTn
CecocXPhX/5M9MCqqdJbS5lQwwxUWu+NIUTNCKlXTMxcm0J1+ckzTDzK1mGmHz/7bFmjpYzs+xH/
73ALcKKLglBFtszoReUG7Hn+SRNdxARVnUhfSQnNjzF5zJkOFyTGx/7uHaBIwX9+7PnKXjxbVxro
Px89tLhJM3B7wLaIt5HinWbG4N3Wa78gj6ZoIGr6jXYDCZux+VvJkn3yRuZUCiLNA+wA6i0dpd6t
zmt4PpLjxOayFkT/Rug/G5+7Mvo9hbCWesFmDecXO+3IeXiBR+x9Av650s6vcbIUfjXejCN47syY
kslpQXYyiI6SDhsjiq9u0eLe2HBc8kbwUqtENbPp+WWe1WMzljI+vEGT5RESQTEPETnnikKYMN6P
t0z/bsNIYTOVFR6B4myJjsh78dFGnwopuqPZ421HFg83OTcLP/s05OmmXjk0X4DcbwEVGalGWQ2m
pfRtPCTcDtMU9GpXpyWMwNwZR9l8S9OzeRJ1v5/2kFddweKK0+FrDY8JLxN9cSsMv6uGBDqUKF+6
7XAYTSE7unGcHHR8PMbn94iu61qUFjhvfmSsyy+FlTV9KVAhGjf+l+VPJSlzTQG+gnQaFYfFDSbH
BzWLvLqjapk/tjt36MnENWH61eHbfVeGyYBCs94NR8sjSWnoHLNl/u3S+tG8sThklrAgHLG091xs
RA/9FmY1HDXCKpLhhl23UJ5QmW3+tT0z5tH32YFrXJsT13ObtirqutWQcpvzdviBc+sqf0RU0dkA
AsrK46Ouobxo6VfRnnG26t5QgWPg6oqkPrXdL2P3Tjz2oOQEccmOQv8Zpa0UUHQ/tCUnknLklE1E
uT0nASjk8Yg3vXtktdLZgJVHLp7T7395+WANP99VER+uIPZ6wMQDqf/EqPGi6+9eon2BnB7+qpXd
LdxA3+nNR/r56TTF0YQcGPnfjf8g0wo1rgrruVQrAv33fmitmwnpF9paikaJWYuhhV7d2u3Q1Lc4
oAUAG8BQjmuMoOD5oStQcBrRV8/qpbIgjR5R/ksfSbnHDHrKebPmCMUHjGEvFMGhLmp0aChE7p23
aPS0H6nHvEB8Rz6jIRlnlRNT3dRyNcg5TD3+yhARcwEVmAq+pJIrDGYCCr21BjfMxwbtsqzkdrv4
qQ4FRXswYFkWpHlmeXXpiRZT8vMaVE0b+gbhJtcmTHLPdgUunCcd8ebTVhY2jgSsw5QsTA28zgkb
rzJfbDGIPatUpYcnta9eI2orClkFcb25C98Fbi1D7tfh+/m5bz8EbmymQRpIiLb7TYPcj91395NA
YWynCzglblARS/xeS7Pua8/l0MOojFoj8qHWs3RnlvYSAwru9MGQb/yE6YjwtB3YRqlcB+CP82Jj
rj16/cnxFAi0ab76cm6cD5QSl6UwzgyhwcGugfCZE9EA4SeCG30C1xgE/b7Xpr+O/IeojOXd3a7o
QVWKRg++8fwrFhkFFINioxYW1T3FjZeNdQTPBrNduOsFq6mY1S+xO14eb42pS5PE6GSXDRYT+3vV
ZjdGrbWCNmNPjoG4L2y+NpdFlqCkw+yUQPxZsICpagmp0EuVN5+FhHFMXb7pRIlqofSBru2/4lj6
X32y0Zf87jAMJEfxDvKot/BsxlhJVeykCwNT6k2CtcqQxPmM+tIBZ7X63qaILeEZq2nZQiHtbwxL
STbGi/eu5c0G5nJEc7kCmlYRLwTr7TdvTGdfiO0KdSSksGTmS1HqtTC1Ejdz9/3bRF9gboHitxnF
C8toTfz6b2zoU9GpQP7T1G4xCA+2lutMhwdqdviA7D4He5YiLCtW4DaafhrWG8R0BMxTTLxSihRW
+aoBnbncJAFl9paiqRy8y5+r7HeUjazrjIpfcqy3y9eyZxgwcQV+C/VbtgOBEdWUUW2ne2L1V4aq
VI7nKcEHZQL8w03fnz88S5bzf/fmbzSJOY4SzSdZQvY7Ov5NhMkFcoTiADxCQnfc4RHLv7jC4PhI
HbXwbc+hJPVvMOopS9P/pTancTJe4gLPxjuVAmN+fedy4jNCT+gwF04C4QFMCjDLMctshQbaqf4C
aX3gZaB7N1Jx7d44fsGQrBu43snaSfqHdS4owENxaWO0YzVKIO/CezSeS3qrnBc5kP3bMfEV04Nl
uJT6IF6B+UoDWw1tVgUH7VzVpSTiFbY9MEHiNLiSANzHNrsT+AOAIwvCzlmsuLJvAygLLCfro5ts
GXbZoUPe1NcMu/+wwVtS0sCrJqvCAiE3W7dU1mYoh8PZp0KY8T6w3jBYIylxtpA3bV/7E4tk9f4J
ajli70N9xxtk9cteabqPAxtV2R200/pUxVUBrdPDV1y0Ok+b7+Rou4W5fNzNuuRli+SLndfS68z4
Lc/+AdG3s1adXMG2ze2c2Sqs7+5az2bWVx0EYyR/x6RS1KCc537TNAFsX1rmnZ7PZvhfLsuqATQ1
fIBBb4maDyoYNFQdEPxj4Fi3EMhmkarKNWOeQgEm3PdCI1Hz1/2ar++HCX4PgZo8Qf8DwO4Seh4x
NTmlQIo6zsQ+Q16AB12vVnhV2BubjCKgiHEL8cAECXarBDeCv62iy8nv8Rbnj3lBdRD5iNuY75l3
QZE8SZX+g6zPRWxCtAO0ZPBZyeuN2cmUYNXOEKMYNzG05WK0e0TTeVIivzETGuvN6wy3DvmLVXo9
sClWCthQVTxzcjh21eBrdtlrkHGeQozIwc6o/M8e3Wivfz2gw1lOevXLHAUsgafrw7yUhN5s9+tf
pF4cVFp9FpEh2PLG9eiaAIwe/a7ftHQsfJugpDD/5/kkUsypV1OInZ7ke3t32GEXaDTQcL35Y6RC
/u/J6FULZ7Xq51bTJT4IG7U0GqRkGotj6PntPV3s5alcbpnwH1+guVxELMtJDQ0fSMOnUaCIyycq
nAAvaT1SH9HKBKWjG1vHFYQhR8+38KC1U9kXrnoBEwifl0qiMzr35Qr6mCuAOjsUkn3W7raEevMg
fLlwwOwnGT/5iLe6PXrRFshTIJVLbm44z2cDgvp0vLcWPm6RHTEM+R8WHKoCXGPy1zdQck7elSW4
7sRW4Zz94pzoi52eR7XS4R50on60fZE1MB8Kdl1wp3din/8FajG14LURSYqLvVWVVUCaWv6ss9WZ
iusDI1XqocwYNxeBxRw9n6rL3B/9YfNOP+jVkKBZk/IAR27EpLI2H2H0AiYjGrUkxWZEPrzLLzJf
oYEyppImMaNMlZ+a0x3Nesf541n57dtLSFG+EkK364MZ4l8TLlxE93ktP4A0OfA6NTOwXpRgUC4w
Kd3p5lMOcptMhLx6Rfh6OozeOkRqrgy+7CWQL347rAs8D14OUsRdS3jh1AcBDUWLCkYvfrBCzXrF
tjL+dPcRJS1+UeBbpM7bYgbkieIfNoBVbwLwz6e+VpFpq9/Q3K73g0GxncZp0O4aOgy7IJ6hRd8F
SpPOY9Tzf6VYvRjF6KWGn/HN9jwadg0YEdmjK/DXG8vDUcMO5ju0cyC74KVp89DUTP36pA3W+Gu+
CtS2ibtPJgTtWP0o3wsiFXr+YgGLBmnuiyYH9ycTtLmeDba5ds9/PSJrlqH4GeZZGeD5J3ClaB/O
ohaSP/7IOAsVGEW0f+yyDTfCTBhNB/JU8bf7nG92+fE78pPk6en15p3I1d9qLF1BOf0cr772/Smo
iv8tLKh3LoPUyZulJIGGt+/+M1gTl/J9LrxrmCOHtnzmelVVHGM8A/JLR6t/jmR2vpbhaPxZLHbO
BNZcF9gSKSNOr8+J3wXtBPuZQSxyQBWJmKkBsK+REHKxnBpPOJEYlMUioma/dGchX20Ic7a7bv8+
y+tV1zao+K6tn5cP8rgswR3qb0AzXShDh301cNu8Hm0iuXmrJqHeO9eH0cNXFmkFON1/NBVgJWQN
+QoOvypPqOx1ZBO7ECnULz74laqlV9IwY4pJNXu3hYhhFYR4ST4Dm72Yo6fD4vU+OIHqTUmnHdUP
Rl8GHgxltzyWVqEJSqinGcNDE5XDDPAVdvN+zAsUnXkg62ajBG9zUQNUxhJK/Av8lBhz3C5bfB2R
4dAWJ7N+PrzwuOawIIYYPLbmLVOw1ApNTnn9cm/BdT448M3Ba8fbCI3QY5DE5YOtPh07Hkl6jUbO
jUb55ZnKqg5INQ9TlSTEW+lTjuCfzkm2/zWokRziGjhNn06k2+ceJZf5LHsYcSvzzFhL/70oMqdB
eNPgOyBS2tCTcYL9BG7X1zMOTZeaqaA6LHbMJ/3X4kZyMyIHOsEyfxoEs7ZLRGgyzHeLyTI1DlZv
nurFwdIa/kQLhzx0IyaUwNkxF83QEMaekuXcSMHtBtmAmCyNX/ZLN3Yc380fQHK0pnNx+a53jZuY
BNiqvmcglYeuyfpSDi6i6hcdgsJXPROaO2AzYms6DSr6lGEHl7T1OA5nJPthu6w/uSxWcneB8j0k
J45LItp3iSqhV53ch+EJLTA25QbeIWUuNUN0VeqTWsHtG3/kj9KccTgwcR6suymk4NAqLH16/bTB
kZ3EBGsG1xCFDb2fyUJ6my8cdVJAo+7drfp1m0RhlTu+KjiKjSz0Mzro8YUOXKHGboLlC7vFDthK
31icStCm224aerLJuy1iNUlKaW/3hOiLhgOUmJzX+tCKz1zSR844Hl8OhqUSs8X8Uc/TK0kZ5vxN
duRC5aX+XudgjYHrHk2f4JZL2K/Rzo+8ryqhAM8WO5+KSIQS3WTs0XuYzu61nZXlqL0xT7TqUyDa
WaDkJsCY5ey1/KpI+0w02Vy13JflQVN+rZwiVVII4gES4/zHmv8uU8XXt6JNHsKXPYV8PzfJolU0
NVdxuABj5wg+q1xM0q/F3MTyRcrLhE47iC3cet3EmD6vABts14u+Ev9iBF24y+T6eetz/Gy+Fjy5
0W27ZOnx3u9AimhiBY5//FcYn5BBt1czGSPa4gir/OOtySAnnMsgReOwlmUpvtLGjkcbs9+h5uIm
Bkeol6NhjrS/XMNh/YPLxFLUZpVLJoUvhnAe1W3QZBZupM42IzYSTompKby1ZgdeA7kghxngyAJN
dvBakPtBYhNYJVNIN2iEaYdOlkxETbHCJMWv9pLmW4lZPS8f7d7a3lM99CxpZtRZVc3evrm0581E
XZ9oyDaeQ5vBINB+nnw78564rpTrqxxF9w3htvvbA3Uqrsk6bvL7JObmAnwxACfzS2tXktJumP5N
T73+VBfU8/xoOf/XStMiP3qSmLmnDKzAbO9Hxze4opfN8Kk9lr2/6DLiaRNhU/UYe26WFCvAKrUw
SNV+wY2iU1U8C1GGN1HJYATpnnlbsph5Ram3LiF1rCm3126A6DzyRotgi24KEUVKwr6k1zZCXPk3
yJ+Lqq+guor+u5LkKhdR3QFfk0NZmUrHXjN/Y9pB4o1WkThE+PZzp0tAnPRC23vaPZgBalGoAR4+
MiP6rgpXUtxB7GLh34Z2D8JOPyhFkW7cZAMYuemaRIODmcrupJfKsEb1xrklWd4UVUE3EUcXIr5c
1cOJbyEuziXAdB78Nw8AL9hFw/TOAe04S91stoEVnj1Zorm0s8PM5+cXeg9K0YvraGxBjq6FB31l
O9jj+SGfxo/6RpcEWAPMLnbYjshzGMbbahM68x5Mf6AfIrHqcZtKCWpbNKrlnYMAHY6/v0H0nucr
js3XXTh9E5ySwOonIQnee2BoJSqM7TK3IDYFsAZp/mT/aWSdIHmHSZfpGcvBtKw8LqqQBYv31R9O
eswt40Jdj6QVoquEoK+hfFlQ8aNxMMO0dSuchHNgVNTzFS7Nw1epf4Afyo22wP4xrY9DF4cNZikY
WcgC/FxT+92EvwWMhPOLED4+hCvPPTCF617zy+4mat9YGEpUh8Hx0wqbJF54WPfnHj0qjRDVGFix
5Pq10dOU/VrOEkTskHwnJHz0rFR5VPIV4u6t3x7k2KLKx80m1MiCuLndU+Nc/wDMnp+jg5OmgEyC
fp1e5T7lS+HNkEfqwJ84AlH0TBoXVqpx1L4sPUeOi/MfZNEb2uyqTQnBxM5aJnLxxzxZ/lZEL81N
fGXF2iFteNj5A1OpC73mrZIBL/cIMsvnBm12MP7d99EQMz5i3VL1YzpODdAalqaUy5E1C44qi7+o
F/ht03gQmBKXLSan2UtVQEErL0/CVpC3G1DfhXwtfG8g5DUOrgt2pBxaDu+Siiuh2EviNxufsYQ9
ug46lhdDesyGkOB2Lfqpl8IzSIKlUqNXs0J+1kKUBkJMHc+2xE1pKkmXX5O5iDDPhXVUq8Ot+QkC
HBJ4rdp5rx9T9OY4E25TG+C3XOxOZ4pXeMtEt/hsruk9rxzgGO/g85jX88U705xF2T9RhguEsuUu
Qwdvz9hRboWSLfY+BiwYfrV42jg4EyU11AajXv1oy9fgusJdeQmyYeGlqDcFaagjCMJuy3la++i4
CYpn2aeAFKVo5tAWye+BBuh4DzeuhJqjKVUuQ0cjP9nxF0SYDEq+6NdJYdp935DMIwO57yFXJ2aw
6bhG9Ko/VoN6Wu//FqEMDImZdvTE4jzvnC4s2x5Mgv2r+ccMNRXsA/Fm0MjXw5Sf2yqXZNmBgYse
O56NaQKlho2Ik3tZ6hqKmHf3yS2wLkGiehgttk0uoGhrHLPQi0DI+Srqi65zoj4y7NI90BYAzbTz
ca9OgUwmcXb5gylXtn1bSnI/Hx7sdk5qMjB8+iSOHoLT+ifYfsoaDOeac9nOqPVDZLeejfdSR7Mi
Cwt6Bjy+1vzgnb8+6LPb9V8V8CdX5e5iPeqcwRIsnsK4ZeOeAmTOLJKOfcGl8y4hpg68sguTVVZf
R+iawSi+dPcYp8EYIQEcXrAHm0oSNCZTbLAghI256TfWOYBTbokjW203Ambbh5StRDam2IdGoFxb
m4JxUWNQOGRZns3Z+T0uP791zNikYqjEiL35bvZiT1bJ1GPQU0Z338NmkXUOLAcziVulEZ5pXxB7
qUYY7UovT0bk8p1yfce/RLWs6qsqZ/ZlrUYOZKiZ5Tv4sBcDews1D2/l/cCmJ9i4D2XVfBtr/NHx
vYfT8bfZZLYv2tgLEqtieNyR+hgVNLe1rAmIRlYPzJSWm9GlyKXROQUEpEjGJkeSMNJvXGkzk2uG
Hj2k63syDWIl43sM7qE8AqUljOqP+eKkolu/iF/6T3mN27yMBAXFUvpLtJggM4vCrbYdf0fLJ/xJ
ACoYMkq8Re6nmzLl0e8DexRhzpaCSXSPnOmfzT0fPrUu9yQLTI5x1OIWEdowufVGaOMZDSww5OsA
DfYpLhWAnzCuk364AedqutmHj3FUStQekdKCMiIsDoluqjg4D7ohU1MGA2tfg3c0jZ1aRwLSjvRH
6Keq3Jx6I3b7bXerpXFPSmE4qi+FlJBXAnIkE6WVIx7z78DwYpDStOo9y91Z5DzcF0UVivTsLN06
J5CT5xPUrgFPTto3i3fANS2jfjCFKvnkPuegS9qpBFMH4QnfAhDfHjdMRwIqFsPTMcvqSU3Xo7LH
pesjWXu6p2UA5RH9ECb0sKX1V8P2Old2AslfcqEFmyZjIFBMc/kdLIn14KX+dpPTUr5jQ6k+mA5B
SBzJ0lN6zRyiuGnN2XVeejn5RttyEh4n1CtGpQHgxH2QqYNSTngPSAVYaazntcAYAEsYgQfY61Oa
B2vQ5TaEEeAq7Vha/YY4jSHzPby2KrXO0EslomwBWsEsYleE7P2PXeFQDyKdojewDQh2CD7X1THB
CCybt1f3WHX+qxVFIwhEmYDVMZ9QI30DQQMrVisUngRRy8TAfK4fTKVesVrheykooes3BW2jZsJw
qK4p6UoPnZRp5sLJKQJ+YQD78zQUkk4FPkHXlPlEIDJzt0vagTFLmGxuHGnjAnxvvCSt7xeZyXEr
TchmNcJiQvuBxmerFUqSgU+1NiXc0oFmM2FEhSWkdMQCCHK5Q00ZXbab/E2g2Jlsj0k/kTxBla5h
TILEXyP1ofLMfaTsrBgtrX50GMag5WcXH/+rNPKSI1T/Iba1PvHI1IwGMQ9WiPtvkoFhEBXcUy06
SxTgMn8z9rDB9OstWq6a+115ppVVATyWEYQTO0KvKopSbEmXwwsTOCWxb1vc8PAa2Q4iGF+xm0hQ
cD05Y7JbTwU6rNhwkQ9oAboXQkbJOr4UpXxT4adHG9ssjG5joV5hJxwSA493QvCnQS3JodeMP8po
l8f4VhMy0C4cbgINgHYPQ++avN7VB1vKFlK3g/ieSJm9wzsNClpx4Z7jsWpqaTOgk0/NOCKO51N6
rlITbwCRl8lBlE6CBYGFfNWmF7L6CezNg9VD9OTrCOaLqqcblP1ELJM/hMDEaOAi5pErU+owAEKR
yhSIYllebEK08ol6vYYEDxc3B62GerunQm2b1BtRmcIyjaEtFuByZlzvLjvF1L15vkvXN9TPBl1E
1qstvfQuVYyI+UpnNzLWRQ9mjFkZi0hqBNuJrhLQTHIV+cBH588nuOX1NvV1Jkt2F7dOhvVNBxNS
1ZG0IK2Nnqwu+uLzj2ljbKmIO6KJicjcNu3Tj5xkPQLtTnVtU395menapbOi5V2HJODUOgADd37M
imG0hNyHnSIbexwSFhNlCUQ3x0FkZiaY/Rp2NXFDK3YbgWpKzjlGYg20ITv6AI2VXQ5wmX673IS2
cj208PkVxRMWjGXlt2WYRlosVYl1PtdJT4G3Bxi5jso4tKBry63W0LkRq/M6c5Zw0U9WmkgM6jBW
xRxZ3pjEOfCiPXpkBz9X5XS1kn+ZC9eTKScgTGw3eC9kDb3Pu4vzNOai8yu7FxKrLAlnzFV9gI5N
i3tsfc/ncslK8JdkM7KstnWN7mQHb2f7hdZXykj09/MbuJM9OTm3KhegEJpIOwvYG/CL6RHfmHj1
JGs+misx8fQoY640WDnqx5eUTCswpUzyGnuIvGlx0MLvYMD+n0IX5gH7Z3kmAfSOYruhXHeiqQk5
oTqOxsgApsUJPqxojWLmEPXnjsal87ICpx3byijUudohcenhZQSUdmGMfqPrIPU23NG+Ov96dGCw
YWbMCUpKJm/8Mf+yPFEwgXv2PpOXFx9ON88bQk/yNMgjkVgbllw2Tbj75G5QDD+FHvbdrzfbRFKb
msJIBvLvHI+Aon+YUkWzSL6cwD3w4dDMUYsoTHeEuCWppo9f9MdDpOZuI5wtlFgG0/g4vYpDE+A7
6mAltQ0rkK9nKANr16bW6r9ha1/Aw2THWVXjUvSCb7OVK3zz5OUgNcriOCgIO3hGe5XrXsHXyqXk
+9FlOKJMjcs3MrtrpcVXFRbhosALh0PHUWOq5p8ysTqNXeYjoYqIT+7Wqd0GlOsGVkLJvuYmd4ED
Ktx1aQHr2RPR4TA2rjS/xaRsS8vhRFnzkkWtelPVKWagMx86+GFm52I97hkRzQeNgPx0pkjcyiRG
cV79af2bgrnUOF5QaeOEWTIBsNr+7+dsPzwYnWbhmikGA/Rnu//kbU05spCur6RxJTmDq4/6Ljko
qbTslW7d0hTMoCvxujWOhd97pAVOAFIPHsj11lyvs3qg4jorAU3VUFOsbn7mHX/qyrsrJD7BMYuI
kog46huhbKqWw1zHluRZNP+5IZAplINgdwJBKQX6GAa7xwalIWFM8GSZw3AEjzhQBV6s/tmAxSLH
84yeQ0d8UvSqm+tUELFUZantfFf2jwbb/NJ5oZZFAn7iKF931FspAOurXOWqdJtmeNzf4c9CEmSK
WxYA8kaIbQI5DAm5fWj4Dnne8wTYGniNV7x6QognNbNiiFDkOs5A9tTpvdlrj1nlQcY1BlrWlCZD
m9LaD3yU4DZX9gIxfoTEqH2i5CHc2v3UCh0AiiL69KkcLdLwXaDrEWEqiDhGtusAa/JlovjKN9uj
F4fxrnIeZGz3iJuMnyk9Q5fJFN8fbwTuV04O6gzgEoSxd6/QTaKcGTvSCpZ3B1kU/zZaYVRCHLve
bf7/BSBp2a9J2TSZE+LL+WA+u99qLX3LlSBoYGCjjP1AWmEt3aDBteRF/GD9vD+r3zPcwS6VTS1X
g48c/Er3nvKVWoHYjSPrSmJdZsQQpnbKD688W3QSG7zHU0X3eOLx36hyGUdYHfkA0s57maZceiR0
sIcj6BBWOZ97IhkhedeAmCcr/U4kX2XY01z5aT+YXDP990eULcT0+Ybi6ZA/PNOi/xvaKosqLYxJ
1sj0ZQd+6Vp2P3ypW9a+SSySW4cfG1BzntxgjR0PYioVomo1LHGKv17JEa5A/a3UDfuYYkkBn8DS
ic1WsOhXmD6SDnybTuYx6LmtUY3HxNaz0yFUuI8eOcFT0tbcX9NNUUDzgwiAXVNytIeDQCUs7gbT
OX1LSb9yo29Yr8TZQCV3KYYOCMxZrE5ajQ2vxTECVUxKflgD8GGa0HVHtQwl7McxSkHo3PFw3Ubq
qZNhgcPNl6CKEugdtc4Pbs8LGCsT4pa3UfH2Y/2D8gsR2Yj6+xdCXC8x1nEXtI4LllJVWsikkE7g
02ohMVZwkdn/P2MC4KPN6FZabdSUoTfML0TZAy+B0dCE+5hjiFsP3p8iwy4ij3MCjuuLg3Wqd/bf
pc8HjFUUlfs3NLgfGLQZpcEF/1bHnpVko0KXVcN8ncPN3hYZnpL8az4LmW+2mAkwdKBzC7XtFdov
GDG3kCrjhXvPpejsjhOwsmRiZNMLEUSmnIQlumT12JgGmnvWQdJeGmbJbe9NrXQadT8+qYs2lhgx
VNvTDKjOVJtUdJd+DtBxN0Ef/ilBjWL95JuysMYqm7XmO4qSxnfVTvWcVaUEMEWBUaz3FZuw2Cxv
3iZovNCqp8+BFPvuxQzkS4B+qr0VErPHO3khh5Hj3pjllrIuaR9y6gwi1+D5QcNNvz5B+61h22Jx
9Plu1Wvwb3wS8MwVBmPC8HlpLItwtxf7r3FKCR2dx3eDGQ2w5P+G1XyJ212OL9w81ziykoT/1Bel
8Uh5dDQeaOwJ9sfljF3TxSsO0o4Ng1BBDP3HUVM/PQ1SRf/r5l6Xgn/ccmt23HrxOxah+X08iYJU
A/zE3XiP9Iaa5fo/T32yl225+wq8PHnA1mppEO1qwFQmLuRIOT3YU7ufjReGXarsDD8CU6LgKE8N
NlmWb9RSLh82FtUsBjfmPNCWwdrkvlYd1QZfzPBpA67jCNlnnjs7hpJGTOotrtdFHUDXI1yUJuRn
xSvX8xzNgjR1KduR4mL8Jw35FIQPGXcFywX7TJLODACFkjIsSq3aNTJKWo6FAqIl4ZvMdiOy1pTd
Q9p7qgLkIxjudng4A8KCwDWRuQeItvfh6iYwyRbx4yK342/wJCGVZNROGhzO1bEduk3Hm6MTur65
Mip+uUBEbqR49Xf/TT3fErh9El3KdscovSLRfB5N9VeAOToMXbC9qiurq0p6ZMz2eMJFbGn2on9f
HbPOfThRRxSRv+ugt5I6owOP3+pDlEDtt8MXxdWPdIZ3Fj6mD9T7HFAtAlQL0NlYn0Et6Jk5XIVU
YWtCrjCMr7R7meoBUFuWQN4yp35VZ2Kd4VMdEoMUUpQTwlsBH2dYue6m4QGmujNCJGQEMHdtqetT
2i6nRguvA0D29zbjXqSKcfHD1QVGC2w/DUw8TwKaOjYrEHfniITeAzhNkfJd9KMvJ4k5JDVN+ONT
dM79YDoxkLLlqVZnpuzTlp722u61aFjySVHa8trYpg4wYpsI3kARSCusiBhgf0r9vjmdgvzxyKBt
ka2xEf+XAEBh4Cg08FY16naCe/5GSSlwaf+y5FxdGMnMhoJgGQtmhYAIgAnoVqjS0NirZ+gSF7CL
H/VKhdwYsDq4K95shIBpi7uHkzkqusbiWu5F8DE+hLpDpPvbGROEyu56iFQjN1rB9gG7Lmnme0PF
EtQDVr18dctf6NU7D+PNq6yJb7kaVnpBX1Mz+YyXxHZPMHTbqnBc7YMKsio3eW1AC1v9iX1sTwR9
UpzEu/OY+wbw5eziqBW+FrV6B8V3zDeleIAiRjqLob1KEyFE6Fnte06E501WoMRQViNnUViN7zpg
eyfD90S+ZONT+DI8l0keMLN8PCS2Jj7YxdO3ctUZ0UNm7m9atP7PRkbrXcTG/zVr3DFHpwzrV0Sn
W4Y3XNVU8eOvNQkHZpMSz0iNdqSptoN94prSr2QCF/tjQvIYOuFWZRYFXopKlOChtfvGuRam95yj
RWRvtKUmVWBDjWmvLvZvGiNF4esJCnpHkj1VC50urM+0WqO/3rPLZDABnZCLO7unV0pAx+JzCtti
6FTusjqUvqcM1ls0svmVYkL92g1ttxU28JTwT/IJIY3pLqL+Sf3FHw5/f8V37EN6EJaw48t1EIMs
z6mEdQnyWawZyDVPdTl8jHEm2saNbUYNhxNhnJ9uwSG7twldcbo4CsZtb49pwraEgEu+50OKZaZQ
gZEPKe5u8hh8oZDbwjlRLIB0M0IlebbX/OoFzhBiM89tW7wFkqLa+8li15RYFsj0VVL9+rrMDPDy
2BNkjQyUzzo3If6dJT3pARSpdCGIuYcSfX9eXGzcfd/9lQ1qqG+4BUxVWDHQbuGoKIn4StzNX2Jv
kGXg+AolyOz/nf0grqwfoQnHtzp166bsklnsfX1umG3myoX0KsPxlY3Sm1YUGe6cAHbZguIMeOKA
OW89F2aSCNeFLwesD4mai5heA9MckNjpAmohr79FrQwxH6ie8D0skCNdpg9EgibzhrJaVwBEjf3D
Yq8HarH+AwPNF834QUhW4sDQr0R30ES654cicboE3Ysc0JkIy5tbHRyHw4hKtS7d2BTNnPXfdjPk
k+vRyKq/TmyAhxUqoVvJPBQc+nwWDUTEqBD6R2aJzWnhipHa2K12TrIMS5P+4/Q4WZ64UxFIoqgU
KkKBaOOXz1TdoBvqaPZeKGxOagX3/GEFtsovgYAMPmzNLMlNgfQGi/ec7zlPAIXfRxEKf9tQj/IF
m6KHCKmHMkIYjBsIzpz9rQw5yGjWBF0Z+2a/r8mEP8EQV0PZqdf7u4LBiaSrDdkBMshPBr7E4qC7
+ym9kFtK6SMftZ40AHtmmcW9w+fBX2iUJNxX8pXm/iaq95zLScG9M6llC+V47VWL4vpP5qNvEMem
KG77tHm5CcO5jxIuQb1JU1Z9TaLZEGaKuPmheLsLMUEs2ZZ3IbmNhSpZCwV2XqCwk7yf8ocstfzx
sbMDxfYmdL1LHIKMq02pgeWt+4Y5uJMH1nbcFVvRHBLS2hBHBmwcz8iaaiDR8m1BJqCuSBPZyaSj
bxqjiL0llPW8KhxHB4wIXGUhT7sutVaDV8jvUARxB1beR2kDBXNaP5TJQPfIKxEHIdmYyxsp158O
YxriaN5ENUgHw1xkhjRo2CdksWeEFGM2EfR7xycXxnVEmrXgtC5rlS0Xn90ctDa/arnly2Q2TTo6
Cq+UWSOIIzqvMaSaQweasCHonOo3h6PzOhhnsN89wxM+/5yWPCN+d7rXVndyxMZ+pvjnm6vZuVH0
BGpSldbxSjCatXfOpWxFHQcIb3f4AToyPUvko5XzetPJta8eaIRvV5vBgzhay0nDl2qXk83KlM3Z
oA5MwBIMYrrIhRlYiJ6xf/kMSa63mFR6ePkfNjUowjw3F2/1GIwKxNliVHzqlEmU5RKsaEt3PtNi
rVsusut16LCLek4VyR6BlN2icsxn109CSh7WygQj0qfjI3n8n3YhkGsL7iMs3SS4lyniAX3McjjU
ZuLFSUGzIa3qlbo3TTyzXy45x3zdlC39t5/TR3aT/v2WVWyVDGmRazceIhRgduczJhLFajuGbRAA
OdIvkie4nQXBVqDXkYbOqMZZRrX8nKBjVtbufUnDQhdeJvc6K3CmN/ytY4ytqMDZMLiVK39aMQR0
vc+v/u0cyLub6cemuRf6B4sW4M1NDkEFN8Rj7KaXohFBPjyV9D/vbZnmO9Cgh4ZP12rMlHgCDZa9
kmp1X39Huu85e5rUfrTHSapToss3f3lz36wKhNIclRI8aGQO/FKY6O5H7fCElYsk/wfbAYeaDjud
u6xZbEenNA2Z8zciyDocnVRSl2krwlN5J7YhPRmH8prLXkJNDABb0P/ElxFziEJ+jDHIMjDaeNAt
/wDx2SgKbZWQ4o57E0Wd/SUHBZKJDL7YP2Cad/vYBKgWp2Fup87fYliJRDAlN7fbyC6ZGvp0Ey9K
FlbPNYvFbiaesesB3ImENGP3ovfxEdI2NMTSmoGrqHiaxi725XszUUzIY4PANW2mjkXCsvBFZ/nF
QUH/wBdyqHwev20ERpQjVHk4BNillr1Nn7IuAXuL5OEDaA8NVtccFY/Y3ggEhGj9espo4NwOHdNc
KIE+AQ/M2u2XSz66c1/oUhLPY6thh4HmkNSesN9m008ct0a2ykyeovcmaeI8BxuWUy6rxJSX/lfj
A4ve2irNlAf6AVJC+qhTxTK287+NrxSV0ixIdQ9Kkh2x7gzfLajyCjbau0u2yFpr921YU+TBSuxg
dlPnS8ziDbwwtHFLbP+itatRL9C6ms42px6IvCUrS30rgxfH1DmjXta+RTCnji46VObt0vrPCThF
JuYq5Rm5nxNYkMJTjTgVdBfViuZYa/OgfGOQF9jB9Vu21l2lR8/A4lZEn+uyRtt8Aok8/QpkEMO5
6OYnh4SNbEvmLsyV13xE/NckJ5CyoSST/wCIzDWXOn1qEY5rtWjKnb75wQOxie6IwGR9iB4xgCwf
0oG2oGSudnKerP5TIj79fnSGz565TAGjprlB40Xhv0YrK2H+E6LpeaT+eErqgJc+xh4ULKH99Jzw
4xSjComqizMonBaIqSfHxlBlKmKf7QEdW4daohAGNvmn4bB4ZouPZACNvtpc8cJ4qCjBumUuTfm3
e1ynNsNpC2gLO2nBf7fxCWDbwfp6t1oMtVeVt5gFA7pv8Yz1+3wNFGBTMfy6svpCyK3bJm5G02I/
IH9ayRD8Ou2QcQgGqcIlUo0Zd6n9sCXC9NiWkeVLxPWO8jVeX4VkDLS2myjOWmQcS//8iKKFBS7V
gtNFDxp/reulcY6O8yVWwFOmffpb+R0iT6swp9P6PHoKb9XfoCR3F3rbUQ8zO5Jt0Ezo3fLLdXl7
fV46x2b/Dw8GX7i5KFedKI8w2QZ+mhFhRHfXY8RaZvy42Bm4vEUIIWWAk8ftnb5LJNV43U+1imD2
HfH6YAQkBpqVPT7JEeikkejxoBWDdUmzaxmth3RnpSKAfZ/Imq8zI5b2f+5wiedLA4aL2WsV3dOP
5bW27StqUyEydBP/hOZ/HTPzf7CSDTsC3Cauij0Y0rfOJWZtaKRG3i/5sKljBidI3seeQMaJGzrF
Gkb0hGc4iq4PQ8Yfyu212uPGfS7smgXt1X4wQeFHXS8E/51ym/WiPbSmuGzo6p0k4co4A1mKmHjq
D0W7E5zqdu6Dvo1UMi3NSn/9Qhy055xHP6ZJNE9986OTof0zZzerIfSVE6ncldzcurxLy5bjULim
M+0XJ3bKCEZJ+NbdBTB9xm/csdCQ4dn6QGNDW/F8USBFr2SWvWFYef+ZDPwFHknPAkFSc8KfzpLX
NgRqLmKwgiG1/3lO02qywn0g9NmeIiceoDgPUq1zLy16iuL6jRw+oZmwiaI0lX94tS3+Zrd6QHs0
6ebicRODxzJzLmW2bOeSVuE9D49W4mkdtdsUmruxTNBeR3ktjz0bBNW3BkrbeLtRWiimsPy+p6gh
62ha3okI5atf87jeYPIW1B6pI5La7NcvAO1EkuvpR4bdKO2ycmUKEInOmH89HC8YEPIOR6yDNCNu
HALOCqE01DBLUya2O1NwDx8ep4tJaNbquIzYO28KAE4Kd/6R2c3avHsFwMFGNIJSR+LUaxZ2ZClY
tuAXOA0PpsFWdENNeso5LKhc63mxe6t1QjGqqE2lpieQHP2hkMj7aVITqt5ctd7EnWFuu15ouK5n
p9+sNaIqZPVUUtSQC2tDFUZDiEQTumkQKSnk5stgrwl1cW3LTI81yQ9O3FFnR75N5ICsTBDiddl9
PFAcKpD/7bHN4Vubg1h6wSgVKXYeOcYdfkrQSLqkJGXzS0Qsb+prfBhgLkJOYmysS3zCnHXWP5P1
YoUX7xfsPba0RdM03yDRWtuwX6lNa2Ea4S7QWXCoUX4IVPp2SMgDGwPpBOQfD9H1HbfUGHTQky8f
Ia2uqAUby9ikp1QE/ElDnMX7rCx9e17L65eklrgHPkDSXh29QV0H+yoHaDOfKbXlouWfJPOyQwXu
yu9TKFodNgCLshjYX1iqVeiooogWB9NHj7cjf5eQUVxO0wCPxOpvVHUbEWOmnHzoihriRBYeVPmx
ISN+l/1M4TVweyNdjGLUkg7yvbjbUizqw8WrQQFnjtRPwVSkDjVYpD9ZARoqLGpaKJY/V3M8qGw2
IHnJVN2OfHV/Li8RfDmc/79ywv5YdNkuD6BVzExJkMG6vnG7GH7yGaO3gq/HUIxjIXVPyFRf++8z
5HSCzEfDuw/E+QPT+VbZXL+k1ERg7w5ULkw+XVkYl3oVM/l7U/w03Mpba5/jtJqP+4k3t4iZBmc4
04v24ubV1FcDhsjiECvN/NFyC38UUIQz5L4dIrN1wtbSzsnVnZoIFi13E5pGGrAqWdUTZeclqpVy
R0iXYvldOYzVrboxYzsRlCAsEoxCvGxw1pyePrZdhdQaqmODKmL3b8QaWXLDWm73m77784qBdetF
5/i5H9A7aFMki9hGJ6+4akZQezo2Y8Xja6pdNjZFJqw4fKkuSVrnJiJbvnng9HXRuhIzmRmnQZET
khEb4mxt+T6n8e1uVDHQrhiFEu9IJF/u+SGFYx/lq+khiQzLf566vDUQO6/ObcS0cRyH4S4coSmk
VyKZg3S1f/r4eiBAGFxVy6xfxftBA0RCEuAqoqkjfZJSovpVa+6ac8ETt8LQWn/v/3UKARygRyiz
QjS68HAjch2REps5gMMhmhGUBew5JMu3PlYu9YhbgSQoY7EQBrE+hZvWIugHeQMVPmSTtvb59GSM
bEcXlPP2YMrIpGuHvEJO9QxZZlIMEoqFmRPvwIVhuYMgSv+Da5nSY8uCfdiZtG8kkdvr97nipuq2
RjfpZrwA+FhcwirfHuAaOQ7eYcj6xeHCZm7kYVf/AusxXVLumw6hIjA+4EuVBN7tObd3XUU2ZONI
jVq3gRuJvQ/XKXqqnkjNM6J97qLMNu02LP5pugd4EBSIyiNtWkq9eWO+p3ThaJDBTKV3a6dNx/ux
91NfwV6FSL0S9w0ZxpWPubLDSO59q27WcpnrrJ3R4t/NGGQCPhZqt70xE7untMYwxHBiF9W092lO
3VsauUfu6aWAzjIpKMB4V+HmaqYSoPXqD2x8G0Rd8UZLCtxDN2sToOv6c6hcQxp8n6PZ80fcZEn2
AKQTcWDGbUkWNFoGGZyg9vKZCtNpmJS9L1xe7y2BWiPp/tGdp1G17uux6+BcntPWJcF3yY94OU7D
e1dnTqehveQ/+JwBrOP9/kno9VOpgRDGoHKTGr4wW5aKXym2m4hp8XSPvySRsfcCA6iPjTZ8CNIR
wi0+LSpqodK+x9QvjCMkzUDpQNLACGf01Wu2ryJnc3+g3XbkGs9vmSUsJkWGj4gbSLEDfZfbO3G+
1qtTPYYrWFdggPOLLlDtP3+Pore4g3HHLz907g8WCNz7K02ADEKwMkFavY+1HcLCWmIDHxbjMmWM
53eX202d+2moMiMWDFlRZuhWTMeT8fel2SrIkwIAQgBKoHecEYdkTnVLdvIIyPrZN5tP0HgKMWAO
TUlrvHPfGSkev9ckKEYpJOEs0kf7UA4ieuwUSgcVVxueuQ1Olzk5MpDUoyUDKWBrj8zwThBljEWa
G59IgCKhgLjO9pSWz7t6yIz9sSfhAY1LLCcUtLnoNsTuAoKvIXxZ+jKzzzoyf/AfZd7boaFMmA7t
1KpNRPejijtA1q9lPvGy9fkuDEKInYZuYlynov+7HTJaJFKZ0EsiE95FLkgq9c4YzcbT5JnBh6s5
+zbOY8ruz7fnBrzZUsBANTFpz+19XTZk9SPo2jW4/xfYMt73al/E4m8qL7chGhaUb5zSoBJXyhTN
BALT/iALISyzyM9IluYUUyQcqidHlvjIEcCdsu73R8MdpPYyLxVdjxese4//PfWlpKHP+lpIv1nX
hoK4y18TlQ/ZR5RFnNQHIItSWd9v3ZZSZA3v12RINn/8lvoYM6br72YW/ExSnbM7GevJDqiiMJzv
RwqYU1/PiAhxSPbV/ZMVD2P8ZlpnTerplK989VBGeakZcAK6qLJvVqNy4UbpQ75w9jfAQ8GcrA0X
5XOSQWdF3lFEe30VGtVdW9naWfO4fw5psK0WAWfJVtE3/b0CcPuy3uLMQiMvGj9D1RZC7hYUf18I
4jm4n8dYb5tKtDv9HHgQPdzJkxvcP8KKKpYxHmr3xG1vRxcW6iWH1XC5HbyVKMtbJC+r7fYN6Xsa
S7tSBb2jWY/IsVDXeKa6cOnUlJpxokQOfLwCbauYSnF16R9vkq6RBOyRHbbtqSCFv7ew+6MyKI6R
JhpH2qDkVoZ8CkufOc513g0i4/S7CRWf3ub7n4wC0KuKAT09QqFxSTIHmLBhU6C5zWtSzAkU750Q
B6WWWtHGS0vnskQBUXYOWDYDdxTJvR+MOkhUE8ZDNd4YlSJeb2wftCAcYpzmxxKlPs01qakqZLOQ
kEoT4B0AJd76FPMbx6Sl1Lad4N7bti1xV9pKnPRUG1q2mRxYjtdVVDxbGPkx+7NRfOUHgh+qYrJf
d/Y2PYQWEA7V6UyrI1FI48kjKbCVaqU6RLN3z9/GxflYiFJ6QKeNKJTosLuNcZuHGi6ciirEcp25
gw1hPhYTOrKXX4xVpnd9AQHLbKTaZJdKUUeDi9S/1cGY/eCIfPh2mwSiEdazg79O4JQiilQEmKm8
ko+VJanrrczDSFZmkLQ/HPkMTqlJ8/3DLDFB2m3aBS0qozn6NRZOwrWF2G9jPY3NWeRq+fNmWdW9
/squ2OlJKMojEwyr9PZ3NL3q/2EnvhfHEmR58OdT6boEac42Di0+Ku08mTZ4XuNFRiz/cbVmPF6R
Hn+ggMYP9UVPV9LiDNAshUUJ4TGGvRdV0jB8kdgqshHEg2QdWwAQHO3DXDlwlNsdv1qO7lHTk4Ya
GmDAPAFBOZb6FXDiA7zPYh/eQBMvtD7RUS6nBrbOu8WECkpXJx9KBdswhAuWWa9IGY+H6Y35NY5+
tU4Vq0gyS3zjoLxac0giOaYDlNbqzq5opiKe/L7IeNbwpvfO24uT9Xpii4v2C2ZayJ6khyj4rlrM
s8KL4H6meQ4tokd9muRLqrfwcsG2eoyJO14blSVg+IYVEEkw4+T2fug4pNBNjjV20YfOQ6oRXDk2
wDox3IVhVm+BTTCCdpmNf0RN9QG7n/Hq4+P3ZNzAHiYw0pfKHgWVmrCS+ssK8owsZQ3aMN+EMjJA
SIRILirsWLix9HBsQrDbr5TT0l9DUnqoir1zEi8IoupNjG7HOc7+viA1sTZlnf99015KgGJ6sxws
Mhs70jWOFlMAzwyfW4lKBroYx9WYNBpouTcUxi2/jKRRsUt27F8enLWqX8RUaxO9EOheTft0rfz6
tjlzIj2tgokUrE/iNrKOP1oucC6/FMJNhFFs8uQ8qpBVKCdVGunbuMqwjKJ1AvvGWi8g/gxqNwpG
rW+ekqt1BsqlcPIhwu3xTr75LSq19jF4QQsyMXgUshNE1Nch5KhSQ+kLb1mFNLr5JSeEEcAGyGUd
sXpoLthk2Uw2mcR+6XnmZKNNoOFqvuq7fIywBUgs3L8R65RT5iw8BAg5vJqlv0HV56goMz4wK8gW
wUwA6GoC0KYOuBrDTdq6i2jxr8jWX/+HWXP+3BnI29eFWGzUDvUPKZM9OrApVlAudVLg/+5fjj1l
6hgb2gjXI6L2HtxwN4RRXxiSN7QYkp8Mpt7ZcguEI2aNliyIpojOudqJFxFJp77rRwRpioizaB02
wsY1OC8zMIiJeg2dr6z7X9UlRSPHe+Pu1QBI0ZdQtRj6o1cdRLTXs9kLojE3RlOdGBJHw+CqPXGD
OTPvFseH5HD3k0bQm5xUkh0lHj/Sdu7h+SwjeqB4/TWvW6ym6D4+9Y1CvKZpEYunPqlTN+73rdgt
MpgaegGgwi+EP9y6Kr5Xt9KB4bt+8QLr0ANuHj19qQ1XUPDNd+Zmzc70IUA9hO6csoG6PDxJnH1B
C7jY9XL8k571cu1monNukCCXjkY671uIX0FTOAZaF0Wwrp+w6cdIEUYrcewpqJaYX3MFvos3s5Ru
a5q61ApsH9WDEQLGuynFf2/qaFnDavnelavIe/9FhGWEsyDNxluddK0Igp5g12xUSV5cJotD/m/t
0a0Ir0n1otH1GHyaHzkuhQcMoXqoZTwcNtFS9KEqPpELSpUXfCkHv+PgNIOArRcxrNfeDdFEvt4O
I10OjHXmQ4ZelGPPvQF+RPbCWW3EA6dgUnb7IXgHIROhW87FP6xg4Szk72ej5a+sQ/euEAkib6XO
jc3uF7xFGnG+EoOnGFvdpEra4hxgig5bIi8HUY5nLt5FJUxGlsneqTWQFxAwEHPEYcDygyHJW3ia
EoR1PEmoXatS289jL67xXsK4xRhuVIZr12SsEnbh6JJL12Ueoa+/LiOaBNn13KdcKNkxklnnVRVM
ljBHZLyEuHqYpYoGkO7089w1nE5EkgFWNHcCpSV8K8iEvOSsv9WiYjHfDxIB91IeJHBpAgmfmOPf
yTgNQ6+voMiSczxUqJBe62a8innsajESmIX3Qpdgnb9/G5wmRfrWxFU0xHDdMDiNMyTc7Z8xTdiD
4o5uAcvycp8WFecSbQblu7lYaEaXhdx1AKoDmsCUrIi6KqLTnYf0CfXB0KVDPw/qiEB5kab9Sj69
V8itkcb/1zQR8AVj+uZSzK0mLPUicQYK2UEdU1BC1lIQ76jBj+Ovpn2fY9rLDms4/bnFjmJ3ZlJ2
IZq2vMAbgmoB4jqO+Q/v5mORDWIWZ9GYVjcJ7xAYEq/LWh5n0ePtgErPhmPx3D/zoSV6Y9w3zdzv
7yiEDzkmwmCzZwVOSUY8qGLOFxTMxB5lcwXmtax5qpUe4WA+cOtWfkktO/KDQOydhsIKN70IZ+jm
jZcLSGc9bBYUzAPv53JD6gTkkaHRRfBvdg1pRxYrT0aoKpk+X6yfFhj/MLJwT9K6HcrXGhZdve/q
PoHPXY2lirSt3iRgxeJZ6MGYGslLV0vsUZmeIn7pAIcEb/Nx3ardl5O0TO3THO0EyN6t+sA8rkUO
8wOpO43BnT4W3AXGjZpWvQjlO1TEE21nS/t2iMDbMEbxXcE6kl0i1yxTqBEhKereG3YDhb1FGRyV
8p4TIHeLsXp6FYOzxntWMnJwNOPdSD6Uy0AzaYy8/flEwyyOA2oYnl21xnukXoa+TvkZ1CLr/q/C
UXqWQhD52Hwqk5HlaNH9ax3Ehl7a3GGIjlM+T/OsqyG4wBGqLEx5HLuPf96EC1Bicp1ZcBaSCO/O
M4e3P/KntOgqjXe6XeYI7BeOAmXLmMph9VjUoCEdI5qW9wqxMeO3rMuncf/+WmnjmPHnAxa/+seD
HibmAwHnJj6YpQUEJAbo4+TyvmSb7ImGmn3rpbd7ocT6uxzfBsUFqPUIxUUd5aW9Fcgg9H9fRWE6
mXr7VroaO4KPFUz7wrkUNvmc7CHt4OVS0zzuxHBj1PFIKvZd/Fgig7hE9wZJRlkFFVVB1rG9h9sN
bQ7K9R+kDhEU2NEoyNsID2n3l7VJBWY+KyuMs6DRWhwaCoc7EUQHEr/rm6f/QxSvmdSxLMFwYk3L
Zb0wguChUyBLOJJ4lYFL7s+jlYasw2qTj0GwshX7bJ1e6kaYwuXyHo5UdBolWSHi1+yOpDXvHhmw
Ag3OmfdZOhmWm6GLPWaxO8pvdZT5MObXskyeOP5AEPSDPF/cgCVs3R4mXDe/mqdpVXyJ8Ahrj1ik
pA5jqAajg/eQyl+hqgovwl8fGKyxpBeXfjmFtxxqFcOxbR84/Z5MgLvyxgQWexG/UUISg15+AXV3
5C912Wr68QbOd0PAcWqNchL0PIhDAa7QrnHOwe7gxzAAYR+MCWELSdhDnr4ye2ze8lguYjDo1Lhr
ZugRESX1WVTdNgHeeWC2NH7wwF1OVOfFl4HQNKd+3W6SluSzB2vypq36AdcGw2/EJNyPpDCCtuGs
luprYL1xYppgxC07dBeVJCRzR+Sc+b9vO1u/nFCLQURfRWEY+y7XJycpVCvdQV+2C4sbKELv7Gjx
rzBtZzw/RdK+3VSt1vAnHjZJ2AOZb1QW9bGxam3tIkjvSlfDHsBqropOWzt3tp/2ZEiYe9OzBzde
zoV2kaRSXbjonWUmivdri+f3N0hZcnn8WOXuRP7q8AllRhUA7q8xu3O37+o/RlsOLCq9+9k36Nv6
WqitM3eRxVQD9Mj3rVBtIyM5f79sS3fDoxKi9IvTEnRBCCIIeNq70NaGibu4BRe4KpEZnDT5shSn
GMAsD2HtnIQtuAOKGkF1HxD62hiG5U81RzdJc/cvTw8MVmUmbkHgTBN1XYiQNdsCL1WTXpvnf+yb
81c6GDj39RR6OsnEEXe6t7NBrOK2c37CE4My4RqMjY3QCtt8WneANyt/qoljKxJG5PvvpusCQ6el
p7803C5u6WscVQP/w8VjgRaXULwgy6PJGhGqMlbEOMEVJQSwHII+90Cmvxfa3Z98FBUD4qgjttkR
kdbV8Pb3tDLskXU+UII6CYK9O3WoIMjEJ9mQjQ+SUK5Hnj2enToURbcsOOTOZhc39e9deVZQqPZx
yePf2vgODV4aE+6D4VnpPEwhgL3rL1IU2fIsrxSQehV9fJJDCoLSluGWvLbcI82V45SdbOIFdqeq
QdOjr7AmhYv1w0mljxgqlrRv+N9q+c/naS0Mj4y0LFr0WDRmdvXZVEmeL210btJ8AgvC8K+XDCme
VjWVIrIvyCw3963r8CMDutiKeidjvLb+zq2Z3juDifLHSHbuKectIh31gnt4SaJkMEssPj4VZkbL
/TzNdS4S42DSrWrzjiTrbpS04xzmQrXbEUxXBdpC9LogzmPWAUvdpMfiHa8zYzSiSM6s9DpuRasA
yW5kzVVI8+hyb2avPIHnd0GVv9BsTo1mcA+faRdkIyM4EDbCzIAaYsqj78Q6FdwYaWwUleuj0OI/
I1efX1oqLqqrxd3/+7Iwblxo14d76yTWVf0WWVNNaR4tq/9w4gVjimZ9aehyU2jjbetmDFFgl7xo
Raqylzh9DGqtflXZxq0iTxnF6H+C/V26MKE8ipQ2hqxZml8g8baYK8WZirEsVBxZE9fZZL3ZcMEo
I/Te2yW+VKVBANsutUP8k2hi6HL60P5Sd13q9XZr2KKpAbfHcl0xLNm5Mihs/By7YnDtXsxWEV81
kLG4WB07f4Zws+NbY6LMbXxxnEV/RdJ2SA6h1zmX5m+uE5MrtgkeHVVYn41+cYaJdOVOD2RTIcIb
nrFiMUo/khS/4N7uhhoa8x5f24upeBjK46eKUz7d2qzMYfdoXYu0Vy0gqJyAdKZslWy4aA6xZIsU
u/9CLuNHJ629bozdnrV03wXmD+wubFYi6hxONpVz29rqIPPkeEpn4qU6IB0KuUY8IsJbdfK2qo4b
tiPNbiRAsLuCylQpWTTlEHOfe/jb7KIhXTl40QGPm36htyYqty6bH1Je+myDVQlutHz5H0yNxZr1
EfitI7BTIguj3SXVIwmg1x+yso0y8i8xODbQOk4AVF7P/SZzSXWMz1z/jvDNzXTIsAcdLVJd+Bw9
26IlBAlNqke3djNC2NDFyALM4Sc3Q78KIHZA+I6RrcpIOccTpLj5LGLRjwTgIr7odm3UM8+syQ6O
Qn8vNdR2AdOH0Vk3FGDaxH5JpWLJJ9BV20eAuX4ACMS7ub3u86y/7vAB5ZAtKSdjJTjNqgab7VWW
O9t8sO0xFYhQMmPO8HzQgIkJDPzV9cuRghXogxdfZXf4LFyaF1FnJV+oLJDxHWOPyfQjJkLrEAra
FbQHaBBYyjq+PABFYVzo9liDgiq6I2VBBYfRLW2drzli3F/hFOwSiTufHDIifE2p639mswYxzPAr
n5ayfoxwknPCzVcroriz6wSuHol1Uqa92e/8a3BBNu35FV0zyAh8OGfPfojBGLYg6Gi1+04CoOAM
h3ct6yPwYAAGjyzgKVx3htCSNrhtUUlwDE+e21x/UhJt169BhnryNhPOQNMxQSgOX/flVXCz+Ee/
7xOkwOLyRDYHflzTXLNVZXfc8BvLxfYJbayHfMzXnOj/0qngRnTNDClUOC/nLoZ5KPzoqi3iF5s3
syTiwZZG2e7dRo2kiQ/Xci8pc+BA4sl6WIzduPXmW6PS7iS6dAMq4Rrw+v1sIPhcQ8rNQtprJ27l
h2E4IYgRJuaT/2xLM6ShZ8OxW0At8t0XM/txcQaMiAE76TqQ6NzskHhxyhVsgds4qnAr42j/Cfgm
Ztz5iAjSSy8lNVAU7jThr5NgIyKI84ZQgmhyAOW6hqQ1/qjZyJaHXRedpx8cS90On7QsxuxrJGTg
/nsFKJR79nNZWfKbHHeDu6C9vmJ0iNw+v/Vp3pjF5Oa2dOr4lpn+zYXUL8siwXipCn09Ns/IfJsA
ZDp+WUzUAJx5dmakty1ew8HxaPf3isDN7CCmusv2DJ2Hp5OnlzuTKkUN3lXDBfmG5HNc0KHMHgYn
Y2UiIPbtYIQ/vkh31JwAh5QP7Yfl2+jyeiLuXPJYcbHEPJ9Gym+0YtvvI4+C3EDG/RMkr5l4naAG
By2Zfnt62zXr8gxU67DEHVRjg1rcMfzMudOUU3lwwt3qZz7KLFgI1L0ijrIV7Er8VSM5VpzquG5l
Z9AFbKnp7dhl63ZxmHTPDcAvEEhLK2zLyZldy4WJLb+cIkSiUR0aVIKp8QRb0kJQ+6T9OGLU79E5
Y+X1zcr6W1S6NFJ7e2JwwvcpivCxHIPwNZS6emjKXZphZlzRA9YWwzEBbHWID0aIY852AelYKQvz
VHbfiwp+8iAU754hc+DkbNg69mCqDTZoXU2051n/BHAE6mWEJK13T2zs6ze1WXDqmp73VZwGtcHc
3GcNtc+tfawe1gXkI6xYmXjIo2Q7LSmec6DeUg6RnKWAqC6d4ycNFf/ap5yPxU5RzIAnZ4L0QQi7
gUIJNfHvdy+dZr6IgSVMtkN3QqHwTMiZuGQUsV6VEhNJMvq58zwG9m/874/ps9k5JwXIyNruZq0D
juAovndP3NhgLAcJxICtmXL1SosUOPhZmAEW6DT114jr8kOWZAie0TW0CHzKAttAVrR0vVznCV0u
KXJC41EftoqmdHn7mkdmWkUwkyyuSzCYuuNJbUCkrufP8R0Zlxc+FhCd49vk9VT8CLwVNc9bm1jP
MIHf8tFJugTcf9plJVosRr9hSV1YZi/hVGqXVZRZ3TKQljPf3Zpopy/utMVD9GLLIuzVDGa3X+qD
j1hozoj1yS6PRo9aHXywtaXImJaCk063gQvHuRe93GWysBbuOkDD/6R5/ufl7lOyrI2zCuYwcpuQ
aGtMYMM6V3oHi2IYkaTdViD5latjQJRqyAF9y6CAQyE59T9i9azEavc1IxHgt6SVz9TMCE/djK67
lzgnBLQjolwzKCxV4mfe9bBCn3ldtrG+dbKxglsnhN2P2OGRsgqWa8/Q/010f4F7sBHZJF8Hcfyq
A/Di1B0bKUdwTDgIILjDVmqGtKK+vXshahT19d5KS5JTyoVFg3txBclLGTFderHa6P4rSaxrmiri
v2SUE7QD1M0DWYtY5J8fKYTjCiAJDKH8zv+IOeJgO5OiuqIfqwKIOWZMnmkPnjF8UqpAjyV3aQ04
XYSIOlt1pToIJTxYDLofFRz7lA6TAXaWm3DLjqoEn4i2ReteBKIXRLj8+Fjb8lKDfInBdaT7jTbG
Wg7uMx+1VpkUfzGTyd7GqsWdod5RaVeBuHpAOtOO1Lau9E2UbX7tYlT9LjO8Y7kyn2t6aa+fMSrO
MnuWH+mq7+RGHaG5oMseQYHD6fhqO5cyLMWaf/PuZqXirCYKVqUtfZdakghl6tFQRdTygkp4ULLT
g3gHcTvGuzpFl4hY/el8aRsrQtODuCc+XXfx0kL6AsKd56dEfLJDtapd+OIEZW5AINEFzq+WtzLn
o8JiYDDHFWivZPONeKX7vX1bu250so/czS7YItEgA97JBiITABnbWWYZT96+3hYSKH1lEuZTHxBj
ynRSdTuU4qrYVOyKa66d5Jz5chljO1Ibl2GZ1kL4OEdiORzMAbz506iaL1Lwx3Uk6f+Ra+nB5Tk9
k8zojb+J1NTiuGEeXxPdZsafGshttqg/lI1xKE0AXQwi58zcxxJ7/s962fOcAFoWI407Ya5v065Y
wDkqKogGoqkNw61/EXwMgm3i7TSvJO4U1oswLADk/3wi+I/1tUvOawk2YQ4zxs8Zx2x4V8ElqWe6
3zDMMjKQMVy0a0hGkqSatbTtlArmZqr0GejnIvJl4YFB1seCKvwys/wjRhEEJ3IRLeb5j1NSn6O/
O5zQkH7la2RNl9g1EB/fzzVlZEY6A7QpjhamPCa8LqwBalf/92u77kMAA2pHORvMDvVuwHruqn7z
Khwzt5RebU6dzlXusonEu0oYpe2KSp7Tk2B2iS8WSzkHJhS1wZsuMUQAd9fTrk8ySysXUGj439tz
oTgu+Dq9UW3PFory73eAWtOU4/3Hwt/aQgz6CY3UVgNgOTGePc1sX69xvqeTv6eVSpz3DvdBK054
B4kQ9+ailBwjkEKrzx6DDKFVeMpS8Jsb1mhrDrW71e5LYGtTjJojnET+RgjWVT4If8vQb5f6eSXd
TKvKCOCtXeqpQM9nQLMbVCmWEujbjd69FUwJCNqV1X6KQge4Px7C+imiG3rTofkDevXIGWD3yxQd
l5VtBkbKm8oScpAHbKgUZUtf8SnfkUQ+QoUFO1UrZmfqYegaNlTVg0YFS4vuJ1KekGi6zoqNsqR1
YyVnTHeSsrSS6zdvJ10V4bGarE6+OFLWJG2/KqNA6ekgm7SIj9biKdvKXj1NFYLDbK1MyeCJ1HSi
Gj6ABXq5lXkSFFQhmdZqI4eWadDQm4KDorfAL813p7EyIO/PkYIJ7rE3fjme9MySWWAQgpfl/wuG
YNq67UGe9UYBkR6i46adG3RwULkJOMxKDQSFujP7tTA/zLX1QyJKLcFASH/KkauKCaUEYdUUHqkO
wGHr+SOiwf8J9WeDz8OaqcmuEkPSe9f4fuYXbNXQQVTlmF3onHpMh4DuzRKorp6bgILdNEW5lAjH
06BF7FjTk3j9Q5R4l4Rpm25hPgjxYAsmw2Hldg9hVZceJEQW6FfCkDXG7w4fTeHZRy0hfm/zGhSR
cRjgRBqnpEzAMUkWIE4NASJbOrpbPJHbuL9evMqteGDB+9g0pvroggUOdr53VAqqOZWqKTIbXuyl
Xbg9fGTG8yJLHygZ7AFf0yIXT7r0t42RGX/nQic6g1eiMbUtrzrTDHsvmYGHWtV8CGuhD5vZi0GP
a/b34D/PurD2EFpweUtGcCP8cj4fMQJaCpQYQ6lHybjUcrbrX6SXO8Ew6Du5bsoOiEJWoHwoeZr5
VpsqeB4q0CogRofzGu0jXDcd7vNoKD3l7S5z+TfKECkWPXRFt550N+/6ZBcWBqeK4hCATQ90Ht9r
hetDAi2odqQhlZO4qLr6+/joCpCI4b23r/AjATbQ1hapgkKSe505hAzvGETr5BAxl1qZBjVaZJSr
7kvge18ji4iTpttPzvgN9LTzuFsrhOxX15azihJ76elz4p6tOiaf09GZetHyWoWqbRqxtknAsTb5
JQe1PsnE7uKC+ceV3GdO+HZ3tpNnoL+kjZR4h3Qrx2OyvEeEIbHEwygnNRdYQQt1CyTNirLQqLnf
i/RwAH+zKvksDYCcjzOqa+cXcAHxW6VWcjUoOsOZEWSxuybxPa28dfgJfzn3a7D9amT0aHwEesF7
ns29pnONkyNJCvnVYOtLUr9gBsLVNmLUVWjbQWHHfL+TXJMB6IXD65phVxtOlOSDct1TgsZIVW2k
OkYU7T3Npb6HfxLWkC0NYEuO3EgFxUg+7kBzJJP357+/p/IYzrTPvzEKwnJ26pr64WtbW6O/Jp//
Mwa3IWXucF3oP0Wwwia0ffcNUDA4NEJKYt5652Nvkds20OybsNlkn4Q9sdrObRx9sN7BLYkxJSo8
bRjCPa+23L8cbFhM8GE6zWUZgKIcd5BHkiJhFnD+diWyU4Mzj8yam4sNHvsErfSBoH9isDan5JL3
PSuxKmJoqOIW7LQN6F2eoTXOzO4ZvTh4Oqe68kvgONdo17M3hdZmdsFOCkOP5i/MjBLkLzmJQ3D4
dXpFOEjG98EiEDo/nC9cxj52IKalaDqtUpIhPW2TNYGg8bKkG/rjnXvo+5MXx427HUzRKXRDWFwN
HqCoPYRx7aOacqrAzhaUO7UPJv1eEde3P7z7oGvPAVndC3grsTzFCGlFf4nIT/kNDSXn9t8IfIvl
Js3PHVOdpqrwZV7voM28CBf741AmxFj+tdWcnoQsG7Vxxb6LPJouhpooOHBDuoAEUS5wQdr+ET8q
7mDfPQVw9KxA0naTl00mvSnNdRdhoNGhVer4WgAnkrArn0Bwases1F3X1QjvTnYoOjbRgetUvQRO
r2SHyX0iYkN68MrS5B1bNLOgrHBiPipovabp+1G5JAoVMhfsDdNJi2lFPFHOeDRA1ZzOYQIQXq23
wTIItd6r0lInKYNM3Lxcdqi0RkpTuITuABva1whjrcoFYXOKbb1OVX8FNuuXUnkdHXgYtUT2FOKN
q/sHHjIPpiXlQVsOR5UrdZTnusLPI2+hW9ta5hO1MR507m8Sw4zGFAWp3kNqNiVsBp/Shz3Ypic1
bVgrclUzaaGzrVQsVKLW2FFHp1dJNCX5wUQNbsvxsSHcq0CTwx3riVYCLHC5J/YqFNl156n3Dcgi
ibJtG9DayEQsyCJ3sTBtpLKzR0VDC090iQPHvS5/86OF4TxqxUQaJ1em3RWaCBFo/vUNK2vhxPpy
oXvL6n4YafywdIpsMqehKVIE2AVwcpFZCwhnhlqc87l5SS14E6DF+1auOVHQ2pqWj06Vaw7NkNC+
0IFQUFJ8OIzkoznfI7a8SldYx3EYIyOJ8DDh0QBMwx5hP9tjUEC8/SRBVWuvnrY5i/CpWZXAMqIb
YAfeePNym/2ggqvSYgYxaCky8kM5yZDXXFNjK/Z7KfbGiuErWnrj4LN2M0M2VaOjIPnd1yQLwx/O
BM1Eq9bCGGHXs5EQZrTV2EJkX8ALr7pRMAgVp6MGfMP1OC0bJ6DxLRZ23AhDW15+Nlom/yfCDJrd
zjoVMxGbNib7GVczeXmjQBvoadBrUgTsA812Kf9lTWabXZiPy6/CqoAFwlwSIUuW0rH9mm0UXqAu
Iz3xadgQz6i3uawwHT6cC40hZiFqK3MpYJ0nscMwp+1SVtHzPdEFPgMcMKweIVy74bFLJWs8ud5W
0OufanJg6eiHBT09loCOnJHrcIZ791KboDwq+nakAEPK3t93lGjOysIczswkms2++mzG7wsmaLId
zlwq+yXwJTqb1JuYATJ0gVXqKtADvsqoRa+GdIamJkMQJ1cPW+NxM0Rt7QZp7aE/SiExG1eCw8yp
FnA7ucyIQc/HoRU9ogvx7npAlAeuGy27JgUFDxr7U1V9iJTYhVbkBzN5rdddv3B4NyTfxs9/yncf
TiH6Z7yD3v/T15XHmoOAzjy7/hZmyzDQpMA7s6UIsRfEE2eCAC6KPXEClyJu2t2688IPq5N9ZPW5
jRqbBKjF+M6pqMojrBNAryzEtdRHWBxxZvGlUMDP88QjAqO3DHc9v3ffB4BXVBSX700MIR0nV+gz
z9BLqAXgpke6HJY4x5xmufZNIVvESzd78ZV6eKFUkUJSN3LyFspsm/AVnGYp8YVVR9sy7DIcdWcF
T6bB06UY2/K4XVF/TnBJVH/8FyctlGKhq91Hfl/gz9kLkcwvuQLeWF9PmltR1hPaCqdQvfzVBGpR
BG8oYGdb7QXyd13TzRJmyWRCpF0IbusAI/bukqivVQ5iQew+YFRooNmuC22SVNnRkOjGmkqy1IXh
lIUmVnKLQMh1xhT1VVb9x4jdq7KMHZgZLhmQkQ7XJY1UMtggQHpPCsmPNmi9nUEIiE5tcvSkdD3h
G2/Q7mRguBtGwJyzGuTXWTsUPBOn9R3YRdlluRleFPB5ioQUaHKBFYvfUDPxM66fmr+u94x7QoyD
ZFrG8Gy6dbAccNsENEFY34vmLNwWo9zw5RpuVRin6zEEirGdzm7SHmX/y/P69zOe7np++xre4KQZ
NHjAaM+AO/v/cGGcpfLP5jBpt5/DcG7zsHfPgKcfHJ6tTAgbJaOySg8RQwR8nmfH4zCzuqlv3ycP
HwcWoVtyFNsP++JLwCHdD+W/XN1hFDVECK1XC3/9I7NjoSonX9bCR5sNGf0atTM4SuYqEdnO6Lli
Y9ShqobyzNQO2mwKKizOYEIyf+6DDDbAYmTAvVD20Litnt22VfvASv3tnABdYRMZEJeYjMMDerQf
iRky/If3a6Cs7aq/KlXs6A5pUe53j5mkNHgiWZes+o1+hxpQM/AciIOO7m34XTILMXYEo9Wgb/Gk
5Mjf2xzlH2eyOxLh5zaFgyGr2ULJKWEOC2QKfT/nqHwt8gtvNf4as8+2hu2gnXKxD38d/li6broX
rAcuO6aZjydGZBklQDxi+o4N1cJPBqwBXB/L3IsjqNlvdIdljFJPUkKVrf/940hFKKU+k2dt54LT
qxo7zg+SrpNSee7X0u0f9jtLxBC0tk0baPedWSBhuJVtRhwG34BrbakI4g1ldUcPuSdK89zK0hGS
qZm+se8PYweWUTiR6KBpXg7U3L+0RpIVCpq2/yqPwvMQ93GM7ZxdOw+wbM0ZLf5VJbYblCVNd2n1
J/pKejiGqMTOhNbOZaGsByOHttblVCIZcuac15703jFibSPU+/PwbGCp2ynpKNfD01VstMbbEslL
EtZlBZbtw/YFP1F/RepRjCuOzu8cGAmMKc+qLOioBG/4dFHqz5SCxsxWVpGRnuu509ZcQYATZAsH
zPnW5am7Rl/BgfgRDPXFZ4Lvq9OFckCNxVaFdsZRbQX/nZ08e6yzdHA6LH5AD6nhs8AJTNHOKZ/b
bOuddgHA7MYFQijW6CqgarZ0nr0dACs2K0MAU1VK8cwPZGBrirpH745Ryqw2c8RrmKvFrKNEPwH9
8nFNmrrCLcUuU4QuIoPvbFwyaIIfPLp4786lLS5wrkVVpQlAPOjfepB7mYhWMKRgeoF7lj+LIO6l
hD8Liuy5JepD7nD1rvfPrqg+OnG7Y5R4Nt3N1QiQ2UGen+jjJ3bZI1q9j4MQ5+W9crDXED+aseFY
KvDHzv7HzaVunuoHuHA85T43//xjB7Pa9Y6RBRj4zQUtT0jy3D2vpLqisYiQj8+O/I5Vc0KDyhj2
2iqDWvKnDBE/ylv04TKqCNZmwRzJ7Atc3HIP/2uBEw4+WcEcXAwldnVcZOvI4tbucK4HlTTBr9si
+UgX5j+yKhkLF7+5Ct3fZU57CgXIKldmIQCQq5C7JU4YtvoN44KVnW7lsON1otS81/XFYZTEGB7A
43Xlrt0hs8WDYV1/a53UPN01GZie6BD7/kx92kVPqZUyaIxXln2y0zbYVK7K7a71rsXHPFOS+T2C
clR0xa/15FD/TrLLriSednnTaWrwQ2B46bgNqBZZeW2CMZwrrxYvThdIsPYhQxhFAq7STnnTeFyX
YTuFuLGNSj3ShZv8U01gccXkVdmEtX83qAyApFzqEhu44sVzFOQNwKvabDi6jfeWAWMaCYBAss0z
soZYZ3V+vhPs96+LoprP4nOwQk6b7Q36aYBnY5QgpXRTzKZEAdApXo7+r4iDIj6UFdYWwX6VrblE
zwrwI56fR/RBHIGYUglkA5BrXZFaDXYJtjrJoijSt6yrVjHDk/tVtRPbWmEPr+hE1bbXeZOXiQMp
sr5c+hvHDiU+Za5QdMuioy3yYU4aYbsjQoN0+FtDtRuEx5jqgXkbaei2X42ZfGLZz+DEGV4mE4s6
leuTMAHMQsFRmjsVo/1KjB7Lfix+YZWOL39FKuuc9Kj6Q459m3dqnasIfhnpup4rlj8kEP7y232T
KLoL38pGfuM9Eyw+SaLLcu4pjn1l5bcjbZ7DWkzm8ry3znmarPo/TYoNSVreuPkjH8IjyG+pk+45
GCrYN1dEPO+cg2ST54UaXZOB4JJ5MF9UTYy2c+X7w4JEQkukZEWXWDZ+t5CXYiEP6D5MMtUcFRR8
SsLz1OxX4SCB7TZmZtzruT7INReEUoxlcv7EdlHKaxTwfU9KEt/+QIDe60QG8Qdug9PJpbqQbsix
7vKm59gXvtvJsk1cquetLSC/ThRAlbIn8NbTrlsvlCBCNIMq82jBZFA0sa9mvBMH1R+K1U9V+Vw1
uytcWD8OYMaWsXKbO0PUDXmcO8BckN/t9ZljC1yLu7kCe19RWjfguPAnjMYR3amOjq/5dFV/s5s2
S303m3/A3iw+R8lC36wtH1jhvj1EtzcjDEvkfPewlP0j1stxgORJB988AlDgbFrnC0L8OlcDNL+7
GZynnUv6nCKZKnEBC7rujB1ZWJoKvV4eQ/AlJk8PDzp8jBfUTSJqWXAsUQFk7mjY+iGRfn6yHjHf
9a2p9gakUpVc0vTZ2+tK+Qq4fSaAekejo24XJdldOeC830M6vVfKqXsMfSCmzuMNKLVb46POP6Q7
OsJpRTa3OMkdqdR6RJ61qXWnw9yVNgBkRgxnOFANl1wjEktcs/vYBr4hfwuOgwPUDoVi+Cki6xcS
R0V2J4N2bUJHXcJsbHdVJi14/B8Zmb+NFzNOsofl42JVHGGEoYk8aYR7KANzeduz2BcEaAck2hkS
tjfAh+eflxT+LVVz7Ge7BZlJVmmx94r4k6Y2Mzc9GETHWNUt/Z1fiV/7JTYdIEw2jI+x0Av9qyaA
HBA0FTNbL+0dmfPQ0PhiXdGttc0R8Qj8YFESjJ6bapAepylD10ArENrWxsrQmq/gBZmZXpsmfvje
KhmEdXRyqiUJKT6ckdD2oUo3/XEA/qblOf77Nn7DzJLhSa4DGzXw54ZIRMEYiA3jddEmKbiGyqEe
VdbtQsWn6t0FhSmRLxYRjhPhCbuwgtrkDZ8RZseuUy2TrOxesgXf/6R4kv6cPuccQyorAe7veVas
5o0cRKr7TFwoe5hf5F1ZuXfoyjiaO6o16Iqdih0Nva9/h1jV6+y1qLV00fbvbZ/v6YsvTqbqsz0e
ULACoTzKaBwy/Be63qg9We36nd3I5yZOitC1Ftpx1NyuoxmQOuVI1/RQRg5n+Cwi12N1f5XQLgnW
gB6li2K7/KbpEmcwSlEppDKihwzhAgLbFwdJsojXZRGgytq2tRgD0vbVOvfk7tK+v7KTF106F3DY
lxsjT8IbR3cW7i6iXHXnEXbrQClwErvumYE5Zb5hL7pOdsrTjoKUtgDwDReBBwJ6Fr/9ROyJBZMs
rzjnm9O4sSXL8jTK5aYyyAXp+zIoaoaGTtBztzhGl/T7cqJmjWuynHWv2DwR8w+3IQ797JRCrNKy
+79HzyGDbz8bKMDDP6GfYAOu9sb2gNvY2G/pGAylUW2hFVM6hG6g6zTORtTKDAImAAIooTZf7NmM
UXqjE3RhkCQhrOAl4aSxwGzYG9AAGDF/GSvR/rUVLrhN/+ya9W5FJPScUKoMHFUEijOBl0FgGgUd
hNMl+9CpVRqoD5DGp0LyDYl1+/tqPItzBWtcxUNDe1aoV5p5CJJCY1PdZrN3wi7IkWj81R7K9biF
6Uc+Uk0xsNR7RUeqzNGQy5zCi17WZJr89knSEwx7NG/F0npwVRtLoIF300DqpusmRGozwbtu5Rz/
jk1CiJhFT5qD8jGUSQHbY8CkpwmjkJpiO5388kC2ZZ097aq9Mb6G4wgu1uqVU4qLykjzlkwz5WM0
XWKRsB8d9+whxwcxO95KkrI/oru1gPO/cv2HnSQB4E30QRtHJm4Urpxqt9OWpxvGgr2UJIOGkxoN
2uqa2s34dRAPk3CWPAWFBRCpLI6uRhv6z58Dnawpv8s3agv330yEFNOivtjaL1lsPz37RnLniXR8
2oQkqeaRiHapnbWYO/LBg6+/bf83wr5tlyLvIHoxTnblGtXAMd8ORwnqAs8zfCDZDYr32Q08jrSi
28GPk9Y43GWkdm3KaodZ1rP82UUItU6YWjsqfAi9mRn2c/veL//0a/x9lZG1ff9057TO32Y1cBzP
SqR7G5VqJYM+/2ncW3afXfAQOUjPTfoo7UbiX2YHih9IrynNmgCa4Gupp71WNsuerBPY/JiSo4vd
HyuvZXZ71eIgpsUCjgt0BzQD0KA0i5pdmF6ML+MZKaIww1StJnXOrKjD3BkFs9fB2oWV++kdtR9P
yCgzHhjpRxCww+CDpv9YtPax5YzPAH1Hr+KusSlBNOD99a1iXbmknASpTlGs8TRjGQZClDiBDWX9
KH1SDpv0jiSs5aAZlGUXfS1nCyTzT+rWT3NdgQbuf8X0opb5u7c8nzP0ea/CymvFFSTzVYIyG2AT
8J8SeZ+RGrEl/iKwLoUnjL2SXkE1dVkLRlDRQuFH912xY1RIB0hqf3GQS+vPkVF3uX5r0um+ELcs
KRbFmdiHop7YGCxgXAnoii8cUmyxD6BKNo3f16jRmpcWJEETOOwBLYy3TWtWfjE2f9N3jWiNx4zw
y1WSVgiNUOfCzJX+wOxvT7jtdraINPRPjvaIZ2/kNki61eydUX49tpTC6TTiO3zxfxq5p2RtCR2q
hDdKfa0KwqTx/BpS8+vz6LaCWaBuWzXLV1iahmBscPnuztadOG/dizVYFJa1lEaSpBFq+J0aDof8
KQVhKZY+dzss95fdBZKeowDSO8WwoC8KCfNP/sz/HloSExMpoJ6mu8MvwImb93OPT/LLw1d6PVFW
X1yT0noDqrKx83a4fBSVjFovZSJa/wMDyDL36qjdCIoxMV/dTqqhjpysj7OHJrNYObGlmeBvgYxn
Brb6SqeiBokDPc43p04CJWFSblSheQ6iO3AbfNzQvKXBfmAv2K9hinsgkV2ZCVbGiivuEUSsoc6a
Z64Ce/ynZu0I70bRtT18hTIlxl+FhkrGS0DTkxJX9shhYJ1bE503V1pneMxrZ/v7zNiSehAGAWPd
RAaUURBe+uMc7T8A1sdl9xMQ5Sdc4XwqrmjKTHlUKEYw4vsSznQzKU9xj7s4VIS8LPD77RbvcZAV
pRkx0oxZGeDtUPq2oeSvHrISWpgE/pqfSIWMXuvzhXMUkgNmw4uyXF9srrij3i65d732WDExq3Si
KeeKI3Oa2EG7rpesxF56skdtEcfHkv2eNrXoNDONq8et1rF7G9fK/lwwtFnyaUwjESLJuPC/VakV
5k2+2TQELxu3ICPqtI3ry+V2W63mCQ5Y2bDeWgrNjbt3d67h7px8VnOqfb8zplf2iSkPWw8wNLEV
Onmruv7KF7pUg0tbUC80k78M1V1O+wEqQYUX/L6DhwAGQOH0G+Y7qetW+pwgu2Iug0n5OtVnCDLG
upX82hsN6cBh8m6902r2wNMbTXfSQjiBU74bcoUAq8arWZIfJw5DZX+VDXbX2CA6k36u3zoweb2W
N83K2tChfxe4woSs7LkO1dZYRZFc0DgyiUWICEoXXzovS6cHWussLp/4vJ3mAPxhEr9tniREL3Ps
3weMDLu4H2T1zTfyopsnkCAe/riEz0vvyOJt0bG9JVql0jl74zAX9Xzu3Ci91e+f9FAyAS4czzhk
2D6RXy+mMQiMF7qWIaBqMH0L37EgDcMrm95HUf5TBdEC7wAe/OhBHXCDXbpUcIx9r+o1Lw8otpqc
wa0e8o4WDBlL3m6POCaqbqi1+HW5qBlWJdKyDTWsZFziyiYcIp3BD6cNg6y/FdJJyskkLAh9LyyF
DKE7rwMQstbVwhb0L1I3DnREvkatvd2XsbzkU2DMErbFwH9KJhCcpEKxkSmdgGSCDPELlKG3B+If
fCLTOa+1/7s7hKTViHY4ya7HMhP1etVOo5iC+N37XsUm4qRfXpr3PozvMSzRKkl3JyJEKel5r+2S
R78VFv7aMknzITEqpB7Yc9Gcs85y7ywS+La0MRJn5QdKm8gnvisakErGd2gY/IVIIvnn1jyBwwij
fRX4OpUHRHCzBNXeR7MdeKCMfUx77DvE1dcYPsPKtOYc/1BbmnPJTEB1+P/JpMq4jIg0eoWFh6JV
yjMIRCFlC2/lgN1sD0GTgIDNfrHp66wh7l3B9g7njY5QKv795QZ7zqKfR+7VDdhuWbmhpV9KsEH7
VswHaRWqbsv9/esJGHo8nhuCh3YzWWtlbe4ib22rPRl2ERizczA5jAKc6Q3j/+N2+ZhIpddAIE3v
nMRSD5UjBm4sW9KZs3QWQK8R0OZEV5llcp6jkhnmWBuaczuY7FoFD5fe42C+49RO9MSw/mfYS9Cj
OKhg7S6dCpShTOrMOA/ZGnZoygpUQPdRJNIUdM9ozXNyc4IFIfQR+VmM+OXTdePXVvSuvlroumwK
sOqPMZCvDxlCsAvESNKoZAAd3UA4oly8+zeYLXCbaNdORN+Nbxuf9TrqHtjm3o9FGh0fSKBXxzr2
xN/VHkX/qXel3IqF5o+VhuTI++Dxgm7Y55xlxq9L+sber+5UzoWQGcrtoyxuFIjXc8uAhQeau3KV
4R830a6PEmBwvMb8IaW2NYsh75MxgV74bs0pqa570kNSX3m2RFKH1/orcEX/lZC9eEKUyi6qfbUc
vPjfNmsOUfxLT9TkwzXgDrUNMEfHN3GUa9tGr3VaXHeteuBrRLinuKdwzsji6UaAmB4LJDp0VTdV
MAER+UdJRII3zGVRtI8EFfNZcmrxJ/PM/pSSmikpAoU3ZuIu2kaGZA0MlitMPxpR1fsZIxltNiye
7n1p4k2KhmMqIu5Qn4ky1cfsmf8HBhYt+4pFw3HV8r3yEViZNCOqiggWYqOS3OlXlAVbYO9Yf9S5
S2Bfiv3saeV3rfl1MedCcY5IfdGIBIgOYgiBljOlKh9KYQaRfnj6vtql6lNzyFBiuh6iVA/iRQH4
sX7C6DKDMkU4hu8GWOnYx+nge0wX7dOHQ968EVGhQwtj83dH8LLTb978jB9vuOD718cffT9dr1AS
C0b3OjoWFlEY5WNtsII61MS3bBBf1k8jJpxaZ9JcWEwlmxBO03uhGkk+evaYVv6yqs4wdvCLh0+F
Fyiu7qOJihoqGWTLj0Wgi5dEtn3ttVn2QC/Owa3t1mGFixlN4kPTS++hy4VizNBIHCque9pZmydI
nVRxo2yg6davxD8j1DWyBBmuBV25zrCjYsviAFv9p8+ukyDkmlkxZ3JT8SMXoO/fzFFus40rT23v
NEWIUh0nx1hijz7M43xiCyHJXREY4IdBHPSBnYs5twdlX9NVAZD60tqOOAketPxldnk0YOVHsgVq
RJl4mOsEEJzOy/045XBL2w/C9/X9sT7Q3fNCrfxwoikziBkglriFvREZb2ZLwR7o24UnUad8BCM8
92/9jKVeNhG5AGY9r+ChOUsJ++Cn/QeCCaOhaCHUfqNdXhxpqraCdXEhdMordOg05w8rgRpLxPGl
PbA8QxWSJ9kiHMhiiFTvThBLMYYCJg4kmxSy2hdqjgangBD4QetfUZkMPf2wpop/TG2fRZizDdz1
waTQvfNImuYuSzkMyS1qD5MAtogl8wNEsfdr1TVley2go2zaxDIrx5Q5ctPz15sum9p8mxUrbMWm
7kZWtc0pGk4Yy6Y/d921G7aCyGRaz6XEZ7JYXqj7ISrieeKwbgj0JGr3WvNwjjuow82ny1sIqIdE
TVtjC5ZUg8Bb/pv3HZC48+OZ/dRx+xBir4HMY9a7A3rH0eajQ31Bc6ftFy7XiLlRRDxIAWKTptcU
Br5M2LKYRVMjF+MQ2qUjptiYllOOQyHHd9Td3Q4VFz6tPn2yXkkxNmaBKRQJOeNGitLVD8h/IyMJ
n/efkwcbObI0DMbqk3MbaeLvWMNAKzTUVvJFi2IBoETQmRJaV1Vogb5rwBGWWeE0WbDQE2Etb6qb
PMoJw1mUBl2Dxw+tKeNwgADnTWbOPclFfrb2zSBH7sMgvYx1JhckyWbFEEyEWHT36N6r65lTFvnp
VhMw1qk4qAHl9Ch0QbphrQzDQi3eNtKgMyLVoYHndBb59D9fCyhSNZnx6mg6yelC918K7MxolDnI
G1IXua59EcHSiaEx4bjyjqKk5wFVRwnC/T8+4crH301lrXegikODlNqAe9/s5zMnTaznJ5KhPfpg
ccKjWmp1e59O+iGMLcQLz1F+6w2hZH/RAgx9rzNVQMUxIc2U/JbRooEZ4YJQ7bI4OPDBKxJWUq8M
vrLeysHn3Dpu1EZ4/9az4+e9wTjOhym+7EjrftbsCMwwqHr0JeuHMWCwimJruCN7lKGsdAbOymOr
dAHZ9g8jlRNuzrehGpXX4lyhZOQ7gLorOFVAaaR7NebgyVpT+tXpZ1q7IKzS96HMBPfnUAAlpS5n
Nip03ql0zzfLQibw1mAoKDJTchjfNug78bTJI8A9q6/SzQbCoxl8HYH2sBFzr8iNqstSWz0Ie/mC
U+zc8uv0pr5d2CzuAzxAFo21NzqxfTKXWVAXQeUsyFGAsB6N9Nkex0TfdrguQfYjfcFbW9QnIh9W
I5dMq4knXvwzxqQC5pNWmwSl/iOgaQfoMZDA0h1AZs9axYhfBrRMWikpOL2ktbcxr6NeLlG1auZB
nj2FbW+lALqtbhC6MsuBIpRbYv2hXdxxPmng/ucwtwhrDau6j2T/+q+EyRjXJKn2NSK3nhaHSfMG
dBLR+eoYAfC20sRR4o4nRvhV0t3facPNHYaYYRKfIRZz2SwJ7/60Kx3HUjtROd49V9FvlAHfWmtd
qQFFpgkhf6V3nNzTHw1Jcr3G3/S5jaJ18b6xxjHnd3wtKSTb1i2ioLAs42uw55aSWnRLVdcZr3iX
kLVa5qgUARnPhgSAp6bwvNUbJU/bs7sIV358tx9qAf//qhKW5FOxYx+gWTYOw4q3BfransY0kc/V
01isLYWUnwqHtdnDVBwAF+z+kGiVCysqFMt6O29xgSxrJXreJHZ73rP6DCrYUA3iHzrH+s59Nigl
KF2ePuGRLfsLaUi2v22HNvVVSS2XuEclPBGtuH9p93gDkOKWmfPDSEc0ykM+xCQjPN45MpncRSMc
X2KT++O1OPBSx9tNWFva4MomTQKvzKNo22ypSEkcGQgGfD6UK3WFiv4uKg1woSDfXS2sNverAKr+
mFU/rZzAqX9q7F2Km4sfGzkuK+eQt86jeOKiCOqd3fO/MOyKBIhVZrE5JPb/1SG64gTnf9vNMT6Z
FRAR2jJaDF2KGPrXDDZIu1tnnhpO6Nl8T0igYWT03QbWh8G5tXkT0wmoRf6pbFcoE0bmg14fQcT7
C2uHvJaUeIRnvwrWQ/PvsJszLg5LIxxrauJZAuulAzZw8DaHP38Luj9tieCniv9d8/YeKGJgi8AC
8J1gYNjWySkR3fiDlEZTh3ZuYzGamNKsQMg2nEDsoREgyumVZRcY5MZtAH+aCkp30hSF/sDJGnQN
gHv1G7zBrm3cNmBk+hGXgXwOkX9EuFc82w9rk0uaCJgEAkCGkE6vAWD9KrrPD71OALjecR+yig7d
MokDwerMUe/ESC2x0XF0leaqruHny+7T3tqhzcnY/T1s9cb9pKgRB84jW4vVWlLAQOV3KzlvuHUT
BK4DVJX+hD2Rn0qBF5sNCgPm+Zej1Zw0H8iJ200qwR4FInJxwD/h9A5YK64b/dpW53lR+NnqEXBB
TkGH7z8yYM7l+JI+toDeZnazkJ0BfR0OY0h/XGBaVxdoz4wTvsAqvbpQ/VPKv4p1n9PHxcOlltt0
N60Q8Exv8BgL6jpj5P2Lp5wSls4h9W51IbavQzJ6KiGognk1cnaWtnetEAfJOz2H5O8wtvBzN4XN
jVfVb9C0PnO5nLyiTjRz+ySEyOxfVvAIyFaheDiw/RwSwYxrti7WufTOI8ISn5prXRtwXXdb9xRd
mOXtWbvDFMoU7S2/BOOgA+0g8eXWV7LeVhrW6kD6FM+eUyGzkFqm4vp2feSI4XtwGOJBdxs7tlex
WafzctJm0V02of3xIGy2F9MiLtuUAnJCgCw7YQneeFF/nwEQy72IeZQTicrN38fWv10hWic3IYiS
JpMdWWfzVw4SH2zlTJdKCTb/AR0CMhTrSFahG8IzjOT8vtirIwv7ReT8q2r0izSoBeNT5u8+4KI7
glAhmrKKQ5Sugm8I/6KkhllBlRCBFXBK/4pUM+RCqe2yml7ahfKzFgAnGeqi4lD1q7mzAJibjnO5
tXO778DkFkSPbN5fsY5MKOdTtXDEVfbxPFMucyseCInyDVEJFYGzLvtGsoC8sCyWkRlQi3y2rKc0
8GjMDu9YMF0vXzv3b/ubO8XjMZYlKgqnKaz6U0nCPU3jfYh/FfOmErVKufcKD8lGKnn/bxDPbBaO
1H//zTyiimULLlW88FjsZv3X3vCbSjQ1YX6x7UOUYbo4PO2xaReAT1Yzm0fBxo8zcb9sDabx9zAX
/FM+shMG6xEaS3NILhUgDT2YQh740qPcEbWLQ4e9C/bJ7F1csJLYS1X9hmyP7VBQ9UXKMf6vqFGH
eD3tNq7WQYzY5/zNBA18fV0is1Nv/iq/gRLxuI4yQIGP1hAcIv4+rjL903Hxbp4XN2A8cD/xG3OK
cW56NExiZIDOVrl7T9LnO98BFdnWOixiGrJPrOdS0SWoooYN3R3DuhZhsBBMgbaQdp4A/c8kRM+h
l78lF/zkmtzPQJ2PEXhB0YmAZmQaFLtKrxHH+aKahvih27enVDe5JXu4gYuktIUVyHsxdJ9wBc9T
fGqGufMnm07mvmbdB33iLbk009FQrgmgkP+AAHiByXtjpcXCWEqjDnf9ZbukIEnqryxpi5iNsvXd
INLeWTkmEtqjUKsixScll6GjUKBP3bzNYZuw7Xm3/vYV1GaZULhImqr46axl1rbAckxeGO6UnczB
aSjsCsvZvEzCw4K7KWyiA6JvixXo/NQQKzv395FyKU+kyQMo8Xfv3vWp1LJglmDDtLDHFzJfdbKl
O/xnypDmFeGJq/FOHsazUaS7Q9q2wzZXipE5Cjj4DEI8ro+FMA9kts6pPkT9+DwV3qMP5ePfPrHQ
yr5eSjjHODprpdjJz1ZjxWMo88NT5Y8gT0H6VgKK0B2z4/drIAlcEcXjawU+37FAZhnTSGJ/2m04
BIj7qne5ag8ORafjXjI6aNKirg5kgyk+XXgJxyltVuX6yM+NV/vL8nlK2O2+rLnDBinwSbH7o5UX
u5Zi7jaIg1un9jmFEarexOXxSmPvhSlA+g65zzBWtiHnv+jaU9UXycPM2ywi1DZ4H0HD3B/7Z3ER
zbSjXscxbQF/RxPgBxNLLiBeIKBVfTMzMcOlKXu0Xy4Em9cbJTWq8FvRe3+yHJYVQ2EOnblyfpoU
uyOS/oQkehqSWoRABJxEAEJ5H7HIMZsKcJJldDmi7kVb36oYYSgs6CwHsK+eq3zJOd+G9I0CxaAE
Mn0GCFmS06Yg+hDIHFriQjuG3Pxre+pBJPFZCVa0cHrgSaGkvmYyat7ZITWz5q0P0wOJOezO3btq
sUtHPprTMwM3h7DlRY8UOurgc2zr0/vK13ewuslYitadyyKA2pXXuXu3Bx0uhUiVyAnmOC+QjhnA
8LRm6xJe4xmc3Gof9aCv9M79zTC060bi27l1KfaGURlDtA36T5USvHf3mHGlPdNn31AI+CKQTsSx
LaTJyhxmWUC0uA76xNADSa6ojmbjmI0EMbKwdjcAJi4mNWFDj2ZdW9og5gEAWt36cYYrdRtNtnlN
Z5tT7I/NEf+N+jbMEcfsNkqfQ72U3EYP51mkklq4KvUYiS3GJQA/l4qbmTtT6kT/ONwVBz0tqoqK
gSQueY3rzpCGuaKBPNAQcYi0dgYIh4+vMlQOVfKzSZBgripkk7KzmnawJc56s7P7bV0hmrhTi24f
mWQ85RrqRMV+txbdMRUZMBP57wHoiy3ZdzvdtlM7xoscxUOL1RlwVci+7We7uzg4RH1PIWN1YRry
zB+VfO91gPZSHbmLXUMfQ6hQZ7Wi+IFNNs6PDJ1UMASgg3665J1iAiWBlHSZjYxIlEpweN0xOEtc
zmkfIJ8pAVqgaihPoLLZeBqloDUqofSfroeAwENqyO9ZiGXY0KW8emtEtqmTw2jY+UJPXLr8bBD8
n7AEYnj/Yu7q6ofIEFVUvKeYXoY9Gvp/djthOqqDZJAgLtvmOhb4pwnk7CDLbhJmCvGKkb62E6um
Mav6o+tVjc+qYllP/reQSrXA5IdyjBzdA248N9YTR7Zv68NTLSR2C4T+yLtawriOoPJRz+AH3HYf
QTu4DFJlIJvMSEv1fpQFN84SI7oAPRiMK7QigUPXpp8YlZCLbSHe83+2zShk4EgaiMho0PPR6eBy
SvsN5wvQJsSJIpV15WeOnoxGauixlc4qlztnq0dLRmvz5odhyC/9tII+LOQtzbCLu3kfwpKXdq7V
yPRAQtgz1fojW2lyp9b3WZIJGFjpOYaORrI5Wm0FPChZXDb1cOtClEZFvIuRSpjRh4+OeEKR+SFW
JkFepoVwG7l95Lc6rn7nfcQ8HCDsegzHu+QgAtlOvIcCpDYybNNDo+tmeAysnY8ylsGTGLyZX0Hj
ThwRliO2zxKFX/JG/1Zu6NsaJNfGsSF3PeD+5Mp+gsVY+OU2KbK1D14MbC3udXC0fv1IkQ4HkbcJ
J+wV0YgjuS8r7UPiNAOTPlr7PRX/utuidImQYpVzgSSNDsideVZUzt7hrZLX0msiIwRTW7xQJDGw
cazkvthI9HcpsQG679KNcxZucytTOpybuvyhD+75khSIOxScJtR1zsVWMpmo5w7qzxi5E07iE1n6
gIiabhh8F7rX7fSYDXteZVHdV94SNpNcLnpfS7iiB2K4Fgdf0nm2dlv/tZbA5eAdjPHCK6RzrsHB
JwqFmcDckzMPCFJcVRCKNDl0t0KD9TppRwyEtVjtL+kRxJUHex6f8BIRM7UEoWcHXyFWIsVGTMNu
m2VRxSy+jujFzTAVe+FXM9+5MBF71i7TM/1RbdWKgtO1TtIx+gtXLgP9QCYpDAyupeuHJalgdFc0
0F0da5p8ZqMy6w+VyIfMBC0YuKh3vmLK386dfkrN1h7VNz6Dmw62EL1BhYX/VnZuNslk/xxGN6t/
M0qScpmWHWClTMidvS9A+b0VMoaSsIYOa40dHvI5QucOUMKrPsfVf0NLl8ZnmaVBS9a2oEAPcPml
yaJXBFL8s6/S4krG4hDLnE7cE3Ogh3rTHo+DaNMLSWET4FR+3CKVNiU3Ypvpe9ha1Vg8RWHUmBf5
9Af9KDJGwS/Ob0xvp5vX+mTfAAmQx1bintKgTUdZm/oZicrVtqGOwon4MnQoUgOqdpzXVLysakbM
FkWvfzOWyBvtvJMxNdjvA1g+OI4sRNaEvp6lLcevMBaQPGhfJrWnIxoQT3nmI5rtwkNK0xsTEQm7
bxqyuQrmQBko9c1tCBknqn4HQtWjHZOe6vfi/P4FVXRqY5P27jdThazlW3Re1GMFANmeSd+jt+UW
HaHJtQg82BNVgJI6oPm42h92uAHqZzqhEPtM9vvoGK9waRg9NzN/5hJlk61Ev76zfR9vh2gzYXa3
Fv2utdcQneVaT6fXeTy2q5A1cSiY8ETKzOpYK/mvub2yxsGO1kWpkVxvziddfdlkaJcuQvj7wVWb
080ISqn5Istt4R2swCbk4dlvx2P9gIyfT33UWd516VwkLmmpV3HZO0m6CS6DGWZ1fflENfp6gWf5
Ovh2AHvzB8qL1apRKtFmSRNp2FpCRrYeVmRQ8T1VdJbldaoA2ynYjqjs+6aTXN/bXOIlksh2d0K/
AHXBC7QaSA5hfw7ko5FHlkAITvvXnagmi+BOoZguL1m+RibR0AkCzx70nPFW2UylIjLb97A8jzii
r+dJHTEuWeB12o3oHFzR0uhuBi8BYs7BkNdcCbqtMLLxI5cUOYiaAQsrhuxZSAdfZud9Oj3p8Cm/
iCjdKWA595fLPo1p82yeHyuuQef7C/LKkTI834eoEBxSAeoYrKBvTMvmCfdF7dOeCGUApyAEhyIJ
w8Dtd/Qy6lBr7dbmQvX/w7nsmwYoGJosmYoEsPNc6y5OOhwNRgHXFnOmmFWawYXbWuUKdaYKoqOm
pch++wr8vcLdjX5zxR8xgYod47xXDJSmpo9d5R0yxuflI9n0AfS+Pzv3Foe1ZGmisCLVBFD6VjSu
7DwV9Dsp3aYQD70ZKwxzZPkCnv7ahQ0OTVH/9+hNQ0eETxRIqOkSTZs/yZuGQihACzZAu+nrr6Ni
vuDzhxeHUcoA1IGOAOU+sbFVPR70Lnv7C+mjEL+ViByxaGUd/g==
`protect end_protected
