`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TCf5JGgj/7ugzS/sKy0pUT5UHsQVCij5kMFYoFTJ8tss1iq5w0ZsMUYUr3jpzKxBpD03WfXcwZSA
wetHjviYAQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UCJ06o+/kNN4HFRiq8296i5eutve9tCcrt5e2TfD/ql1IGfnmHwDww7XpwWxR95wLZ0hiU9nZmfj
Lw3s0XwfHU2NgrlFg0g32Kl0szP+Kdxx/k1o5CNONeIoyI9qzrNvwVUcai8HTb2d0mMFW5jqblFt
lCzqoWjM7rVPr35MTi4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LEotkU+GtjlZNF3pNiQmTk7PYmxXham/0WU4S36F1R9sCsEeEKVZXi743WQ0P0GmzMoUulsv8krk
WVdt+58hcEp8TU+GzmWp16zuY+PSFGDJNbFXHyxv4RdjvUreDjvBn9I6ZxMoZOsZolEJUph5KMDL
YwB3DDF4fxPWGN1ZQtxP6hBRKtJK2HMCeA2jW1l4EizvArXE3WTMI8FtiFNufmRZrXapSnnzzTWr
AsaXt/ydEUJMd94wTb/lpbwR8o5vY+RIvoZWTULJo8bednl2A82O/igcAv+YQpt92NCRiLzvTCc0
mEBDSjEY6WrQM2ePDm5q2EQ0v4khEuZvQ4XvEg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AlLH/YgHj6mCBY3xSgnGDnQthI+brmGsURwYmiEQOK2t2bIUGrPEGqF4YLjOuzqMxH9wtbTXkH0t
4FrZS8vRJyL84tvltEegmAM1YWNuU2HKMUcl/r1E67WcEhZULYJkTt17CDGMnNnafpjmJNIgfvsP
RSUpXAbqimD9ZS1O+QM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mPhPeZbc7L4U7Cq2HPffhm6Uvs7gz7fvzp6+KTcIjExMeR13Iqd8726U0Y9I9t/WGlzGcfti6G7N
KJv7iiK42A5gaFMX4M739rF6FQIKnzLWNkRfLGyazDmpufyaw28bK5sLrHYb0zkKcZgIpFCNXDB2
+YObeA6WZXZbkxcQiYPYb+YfoGi6XgdCGTU8qh4v6JiRF+mshmKjRc8hvpIKi75csaLsU+/z1q/d
LWI0wg05IFu5WHOCd4B2g5MY4eFjpPywXsPr4H1echWFvqSHM+XniLfD3pwQFljHXjOK2EnMYbux
5cn+wIrk1WZF76IlHNa6fUvO/qFzgsHHk9im1g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3744)
`protect data_block
AbABPLrTOfNcZjwEAXqGmU/5eXvcg/3WI1ly/7Uv3OCgGmKFt9UWiUdutQ8J97TqtSqQZn0od6jZ
Y/nKRqe+ku4t2biaui97LRlzeUs2UDahKB/KS4XbSFXKgJhptx9vBNtybs24dUa0BNvO1ddJhKSx
zXVvCJCe0fLXGrr/yq6SyJbxrXXX9XFvp+Iqy1V0I+Z9VMJDuW3Ikkxv+VObPVJmcyVYfZGiIp+r
623WIizHLs1PWlB2dc68a5HpmM7BZ2B1WGhlMOVCqnTiVQPrGCZZeRQ0grEPNULJaA3V77q/FP/s
BZI8HwYjoiBr9rTTdiDHXsqJ9unFBqiSp5WwkMmfXmLswzoXozcNy27XBQtCQ7nT6nY/JydKu30V
xAIV4+WfcCtOjptAxTitGYKXHcZQJz7AKiArf2Ha5QeOlqLjpD7XSVQF2JZ04yTTV54T/knCeydh
Op1UY+uFrAIu9xeVindX3gW2VgO2EuWE1F2UboXW/bhKP2BtjRTRF4xYcBEOZc7IOP7vPCGf0cqY
OMbCjJIABXiJ+UeZZpiEbxdjKmm++R/KfV6P1lo/GJQXkXC/MK6OG5TM84lngDjoceu7s/O0ma1w
TqVHLtCDk+cjcEl0KP11g8VpU+5BsVWZB9AIoD7RxzGvNxaqtwmKcoV/cCEoKMw+4YcUBvSjFhJK
Nb7DwgekNmgy59VDUzyksM8XD1V+a+rxux/FeioQrBsy7d9auXCM11TgX8cc2e7WlGj2UASYT2LX
RtRyENZGMcam7hoBiemM4POuhzdY18E3uEi0ASQTF52ZbefQ+YBW4Sz5NDUvyG5tGnc9Vn2Cmils
7eZuRDdGRjnO0VF5MfWuy9yP+jnkp1HL1nZjK2AY9cYl2xuxoG/Ow9DOg+9cgSQdF7LZ65pDNSEl
mPuwinD6tlLqcsjUTCmYKBLS/KWB6tLX1iw1Kwt8TRKViapqmK9ED3483rCTfEVsi6GfmFf+FkEb
DIDu4BJavWKtURZApzJt5sBblMWkW5it+tocnc/SSXzE0PFUjSf3XNfx826yQ3IMxtebIqwtKrc7
jTj6DY8dxENyCayITgy5DN1mvPbW3jrPASS4zY2uep3N+0SXeCxqqutlv3DCBEeSwcaMR/4VOKZN
Zr1qCEEHbF7brCF2umy0AY1Gd7pXN5Mwun5hE0DmrU0P66lNQjvdjSvmkkIttgpLBaVMIaoYkKLC
1I8bakO/tRV1939kBBfDNol6RJS80WcfbD51zQO4CbgvXUM7tjo+G7f74E+0LCmYePFI/lldAdmR
ERyYgzj/Vfyg31k234RgJ+fNZM6LyfDTu5ruKrzLeXjLgGB2P1kyuDRRoRTiTYlflWVcKBwgenv4
06ogHN9mBHoEqHitvSPgxhAi21GxSk5al2dkag6tlEp+Lf9IymCzzW7cRG+49SSjsvxm+E6jU7g8
/VThF8LyyjiXKGXsrwp/qUlhjrGK0+GMSeINaOUTmoSthR6GdRTxSpqRYZOpRIp3BEFBNoK3Cxc1
mqgf6+NbHdta15k9w1qLdZK1jfOGB5K6yGmiTv+yfa9EcyBaHBLyS1UXO2BUUZrQScKPKKmCoCzi
rbyhgtlLsDyNkZ1pKWisZ0E9hjr3CpthNRnG9YkDUfiN7jU+b8iLETt28TGHahB4wXQxOzATxSZl
vCh43NzK9wXwkL+rp+gQtF1lQ+v4tvVIbjheM7kea7mBgXmFLOy9FKOWO6WZeZa6QnPOteuIWX7E
n/IREfik3fN4rQqkc/To83eIpkghEaIlcQxjLU/HTj0JTeqykzDDyQcTiqxVLnT4eW3Jlis3HRTu
55wlVfyThdOALHWv7H3ffAnwfEIDZv75q+WCskrPSddnZqxzGJmfzBqEm82qGmDLoFE96PyXOCjc
f2F7RwFFT8YdO77CVsq28+fbJOp5S+w4vtUF1IuQMufqLajeI1nR9zX4bs4n3wY4/z9+Q8TzLLKS
amYXMUCi5Yd2nWq6o01tdwXXsIikd/JZVBS0xHp6669EszDifzpKSP1ixu7F8kyuu+VAppp1VV9B
vQFQ2qm+i0XBiqAQWkwNZfs+iKKG3yLO8nM9vrsLBV/Faq6fmQXZzV/NZdC0SBcFj3k3PtFe1bmR
uXq2mVW0/yscfmwilWQPjKboNQugf1zSCgXsYUdQBTR3857vsYuKIGS/NyPIP+3lCfdnkvNLX2q/
wGtLLivwiLf7qYTYNlOZyZGdcIOm282jt7z4P02hZj/+gvSsHaY/mvC4RqgJEpYi5r7QH2HJ3Qc8
eWc8ECpLHgugXF7fdf2IXeu58OFbCJHE0q/dCMz9ViNh0cweLIlvVzA0teu5pDpOR7a9jASFEuSh
wDk1S69DJUl3RAZZTQqb6p6K3/EISqq61Enc21mz9AfHyiz0HzTO+bhW9cJkJV4BIljQFs0kKr0G
5NyjJJ8EtDbH6UCVuf7ib6l92cicIqIN2CBJHgR0YvAQ1OlKadllIyMa9mnkBnJrUECMZ2UY8zF9
+wLo+5KWGxs4gTXcxIzK/m7Qulvm3HS+GvGM2ySxaVtBJVu/dbbUgNmfXxveTlb/XmfXI7DeRGY5
mNNsaU5XHh21G0MmB5a9eh2XBZI5t+3jb/5Epjgm5kz8uRpLZIZIVbMMS+EAMfei81q+jaE2cDMS
qGHD89qrHOm31m3nt8lSFKFLcWAhD8P9rztLsT0x4Zy9I3SsjdEVy1EfOo6dNjmHBgPhtO8AWran
nFE1adnf7XYN3oX3m4jD5W1nSH+ijAmmIc1GvgjWlKgd+OtrRdhJAXsRK4z/LCbUlEfM+7zqb353
Hju6f+iskQCAx0NAw0lj7i35zIRnWBb6KeapzSkHWFmTztEH+gwGnTZ4xUjWgiPO8+FQPNf34ASs
2YZpE20515GMUNR+UJqZDkVwcF2c016y5NQzYeei1WY/2VrVXSvUlkj0aYIYkYxZziyWTVBefYHw
t2fTmtGSyfQj/m3qOkMBbSRF0GtxHV4SfgHdRhZDtpAiw5GkdhA0L9Xmd1tOeaND1zQNf8Q549ty
zbNE5UgkJnUWrrO/ITmuL9gG1EoBjbDakJ98wzXltLu35xJ5Wx/X+zYWoaDoWGjhABdbLluQGq0A
zycXfi22qtdkxhd/schxDL8L/+0iWV16hzHSKScOeUhlSfTumvk7OW6afg5A2axzqoD1BRTUhWBU
SHDu21ysFJZA+qDkuUiVHWfkpXrc0j3on1EZUcDLHs15AGlsLNwdd6y2EHxMqiflR+Exnu16Lp42
wn3qthUL2iiK5Jz8O6N5nJPmyOfYA/qwmfjLx7u3/BbwqooVKnlO5pg2Blt1xFcykarP4IsCOpc7
FmTih9bGQ04Q0bEvRmz1XC1Qn3MepupRbnKGM7q6guAMKv8qAYho3eqtfoWiKOlh5y2eRSR0LJnQ
tZWrHxGPI+So/iqjNaEzF38XjpFssm2bI+vxS1owy3IP3iP0tp8rwJcVn3JvHR9+yBbh65sErAkH
WcnkE7vaBvEMjLzerGuMg1b1z+BDX+sVoq8w6PudfhuVwV/Oe+dYWQshufBTBe3df0FP/55afwy1
5B5ADjYVIOulzFzCplOkRY1x4FFxLFl9fHQN4iJMFHqneNOYmQKzl7jCchJtqqIMRKzNfLtATpFx
SJh21RTwLbArmSn0zHe13bFr/rYSszG8c19AQeOeIREgAxc8Ig3NNv9XvZYBZTkt0t7pZy3a/vSj
WZOczjs7zlYxMuxkJBcbgKzc9+nMuG+36NzUXxv+SOklLjv5lxS+jV/6Juy0paL5zfxUH4O/f4Ab
EKxLomKD/Z+8/6qBbPD/SDLFrLYWZaPvW9tyfm0Ai0FwZNCn/mM1mpnEjwJxJWbotxthcxaqvjgZ
Q+yd6SmfcaCyTWRj+Bn6QRKCDSaa5z2fnNgBVWc+8gYMXxdZzkdvkYS/Gm76E8V1nAny3L0kacLY
7iQTfDqS76wHAwO4RfFSSgFXKSyv/4tqBCpNDLUJDjCL5yMmK1CBnuRqEGXygWBQlnrQt+lCfcMK
QgDe2CXAYhlzBl1vK2XUbuY4QLrpk8czQy8p7Lglke/O7kpzR+RTy7zFo8d3bdnVMDSQ4MBP53JF
KrNBdivxEjohMpsKJtkOLtYg2gmESZ6InI/70AZ1+ixj9fOvCEDE7ZnrGm8mA/fuwQ9ycEKEMHu0
ROF9gCRVrZu3v6Ri46ktCi/R4vy3tacDtKADmH+JrRBIyctowTkANHpqVTHVvVp8HYcfKyv5Vm98
4ETlCYGU26UnLwiEn9aHLoERHtWHaiC/zB8fG/mk/RTuFKbOPd1p0RPAgJNk8OwlHOqXktImNjQJ
LgTgO1sdbmTgDtvqgnO+dw1Cy2sV8aoS5eQu8UYDEqaCReb6th0Fq36mH5HVhlMg2LvQleKDM2Cg
vEWCIfaNCgU6WePZUUAg0JIothprcIWilvPGJksmmy6XDMTcWJVcVzo6FCZVgTon1TjkCp2KCmGt
yVZipcPKSgy2ukxljBtbnZZD683Z+Hsb7wfiOdZvksuCqCftbYpDQyA268+dSrt0ZqWEybLPRddj
OMrZQ7tyL/IXst8rqSiNQfgG6rmEGKNbmNLRbXPNrKJZEDFhKx2upfnBTEWCZPlAFtCB+vVcBF8t
nR/0wNMycHRklaljNJ5hkAmPugM3P5LQx+xT1J6Bxds1oIyVMw+F1zRL2ukjpqM0QhbdDaYSix+m
I8OzsCmrKaG1UsP0QltXZPA0Xg3oDhEOED5UEpFfcEfaOlS+1MLc7JfIWfU2Wh4AsgXpSxSx4xdJ
5XRko8TIS7W/rXAOmqViyU0RTENWie29DtD2xtR8/MKGvkUQdjDcAj95BqReYwVcSjrCuLUHoEqE
pjaGUFjZVThVRaL8ZwO7IzYbENPgAzNt+iWhCEAgtPQvfiMDokZQyJSWqSmtrZXT030OUywuq34j
ek9+vwhbYCOshOntHAM3x8a9A3rIh2hyQflzzgsyEz5is2WsTG/3
`protect end_protected
