`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ijGsPeN2IsIR73K/pq7pNvIVfL+yGCBU9d2PYspGWocl4eglQ+ci1s2LKHxiK/khQcbf4FiA5kqc
aVvQMBHzVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j9jOQkhjSueqJxMr/PEFIfJ1lwfF7Y9tUSDeDkMS2PlN7uPiwmHvvTHM+GEqMzMdya7VIaAiCUq7
+t0EMUGllv682Ktjd6PjQVAnv9sX3WTHOL2DT6AMXFg0bNpQYhAkpk810eqyBTClrLcKov59URn7
EYWwi+9Rc6mFyHMHL+4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kPoG92c/oBOxgV/zdve01Jx7h5Eg7Iziljiy+f2Mr775K3XJFSArYaLzaIpJgnKSMHLAtIRqkD6N
69NYCR1DusSPZwdBjv9BpXBLkUCl3tnm/Lfsq8pkTsbqFb0oLr+4AfyGdFdPl7LzcAEAFSoFGiGz
7gaTG/dlkxVmmxllJEvUbjUS/EBdDLouJYG1TGYHBGcahRwC0gCz8TMnpSIIPcE/mbkEhWiYWh4o
aLtBKvg2c9+0XP/dHM4fzowL43OFN4gCLocFOV5aekhCY1LH4aDQF9tp8AE1ES8s+k+O8mDNRPW/
TxHBm31nat1dOhBGN9Chh5HOmcReW8Q3eYENpg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4Qy/RPGogfA2cO5eoM91ob4uay7VAZnCvwQYb3elAmUZoEP/a+KmpmspGgrShCSQOFSAamIqYsJa
GnmN3+toeenoDuNUzt39ZLrXu4sMEmS/5nemZGGeXzFFbiZS1wh+BdHTAFnFhoCVVkP4TEQ5b6Hf
w4WlXdspCjjsS/lMcg8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iThWEfjJcy2bl/WuwSnVnc13v6cua1tEs2BKKswvXSpocjn87BRf3HC4eJ9Qt16FX6RB0O8vjZnl
Q5eGo/YWfFj2nQILQPV7VDTZ+EwsHO4HNh9nmR5N5ibOIaiPCm0HxkAPkWcqg2Rbv/VsHcRNGaED
jbQ1dnBpg+R7NupqlgHDXZt5LLJ/RwftT8qZxUr6DW/Gk5bgg5cmI2Qg8BqVqssqykMgwZMQ0PsZ
HL1cVK12176nJxoZ3zACXuBfi6U2va9MyC71n6q/WDcHRSyEPzgU3QZsYUWhjGjY95B65ficQ94I
AmYkV6pMSJxClstFCHTtrwxoUro25R5VdQjbEA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7120)
`protect data_block
LLs8LriFBcBbqTuEBcCZ6+9ZawU41NQ4QLHKJUJC8b51j5g3/gzhJuwf8vwiqJ7hazjZe1h/Liqz
CC6U7C1EeQOxm9udNTPyRmeIpBeuYfgsuQEIoC6VieinzjZcfITk+rTnQh71OtY1XKPC7jEMnWpr
0NGIzxeaBNek5J5ozB0+QctTKkvvX5xZEainn7e0jQyd97yxv+UtF1GNQAobuMlyq8KGxhvYJ6Z/
uKE/CQbuf2rBnds/hbU5Xr31Momm8IXvYV267yPYr0wHkw2LKJuwzBkNmhquJrm7u5IPg7tqyj1c
sex7HVJfCEhpLmh53zXpP1HtfSYfIH4Wco1MAXggQgoA22FP3VUKNmL5lly3eVvObAAmCV8YUCiY
TfvEaC1ky0q1Z8n6YUneyLidPNFI00EAGOhVQWAklUx822Xl8isHGcYYwyKHWQwEzPLw5j3Oi/Lj
pi0MPfnDN5P4RtIFXVAu5y2LE/bZiYGMTLIqnp25nQvVsysE9o1mmkfgaujIB8FPpF72SaiQWdn7
o7+eDSXWYovG8G3aIXmNzwjYss54ayVfIDZaR4QSoUXKzpKS9CIAldJrVyucp95iOH2vxg+EfkuO
2Sai7KV+fdZshp7YN2kFSRUuyMllmE6eaVO7LzbPTU3px/gLENoDqDNK/rzKWWNJv3CskgXPqsrR
cRCyNbtpd+m5dhhDX7MpMWzEzk+TkLi4Vrps9684AOu4nfPr8yNdijuZaSuknagJX2BMsY+m6zd2
igwsKtrkmQUAQj19rAXMa+ATFfV8D9EoL4mCc2kz2OJvipK22wvIDGTCxvPHVHPWDVi22XImkuxk
Mn7C3cDlzQsTHyoS7JI2ci2GRX+pp8EGKazxbUo2ltd5y6WUQZOGvW+I8BLFMbICJBtVFDMS9Cw1
Bquy6mQ5L+MwVZupzyLEESYlJauFHXmjw4pcy5wALGpxECwI8ov3twCiBy9Jt/MPv1kliKvHdd6c
Ad3hkAoBURP7xtvdrTfAfJwd25sFbuow2/Sf2E3CPZhNoQ0Oe659/CEwd4HXBxXpub9t1yScZjJt
BwTz16rHhvQ9p6zHfGQAvwSW8/+9kk10WsNBDLV+g4HFBsTd0IesWuDzjieM54p6clHF009B9jBe
o07QTSiFekqcGTBIGkBWv2vywfkEWNpiGpOtdsDYGLdlQ63DEKi/GFzrVZD0vx8hjv6Y4lGwjMFm
5Kx4PyTODBfyZbjGEn6Sw3Uggvup5kta8ufACGbWVwFSxACencFwAMw2NB7Abmexh7tomSKqmFzY
12/kHM3pLTBwv221IKpMmhDJgVEnwMw5sQAbA2+RY68res9qCdhdC66PDN7IjfL3lG7zvgNt9xnV
/4Tj7GvVXsgqJdqlascVFRY00/o2T0NlxlcsoZVlXwkEFZKMCM6UknH0G/idjkCukP35CWTaJqOQ
MY02NsLQwL8kLgvPPVhoKVuhY74Fom4mFwMdx2sARooaQ5Z25l3jnLdwhSMOi+YHUJbPRWxDk784
+z6CQ0TE6+SPSJeAi1tOTVy1t44itoimMlu42BQ3QkyV3X06kd+G0sFZQiPp50P0U9egBx7MdOPv
qDF8B7ILeoCDGhfLW1qkKTMPs0icd0soBa5Ehr6vDEKtCJklV5j4VPTS7y9Mzp+T5bM50sAA+69t
FpdjBYfvH2zDzjQRvIChzyD8ceuE5uuQqqQTXgZOIOCbsBgWljxH/brSy/tbEW2K2+9n4ZmctE31
Q+LeKlBDOLVk5XnkBXiG6R67DmFAp9f2/0eRRLDGNZ8dCGxtU6vP5wvQmC3PxptjrWJbzWO2UJ5l
dcvLtmWXA4KtDdNHDzLH4C6F5ugdsltExuRUJ0docb55wumtEIaSPeC0Hch9K1N0wq7xqifNpM18
l+660B+pAitePsyZkLPhalTb6mFt9Glzvz69nnJbabdaUKG4LKhK3f/D0aKMEJxzKcL3arfBhDEf
flEXjU4wB/0bRWrAdlLAFPPnA+I7+/FUq2Yax/Y6dXSJumL90jnGSomAs1IlX5vDJp6GahEweV0j
D7/aWoOrnjmzv8YUnlDWL6PwccsPpXl4I6kIeU+SjD7kqBdaDHZMmKh//l6eemcteitTAh+VDmXX
GZCp3vHRBfVn1E6KVaL1mnpVehDLFQfeVkaiah4OiZfrckHv67BkbwErCL9Ciq/XmT0Hi3u88V9Z
kFagjL+LqNPm+xArKa8tmLgmUjrDVhavWEkfyoysAIg61oE1s4WGnTLWlc5mPTa4WfKQzPxc+sRd
fI333YBE59A9kGMa69QWaiM4hlXbEj9CMXcO74m83vFYtWyNwUbH7EEX+0SOMrbIS8fVbND2Vzvp
eKCSWND/on3HxpSWV9h77jSpNWS622GtzJTFWTECSicEogZ6ex4BsH7p+FXsdkPHORah+IeHewx7
13iPbbNxaJBLP1QplOBCXTCGL4MZ+ej30PuIosvsb7199tBLzrfMuFC2hYV4Ta5ln2twBwujedej
g8jFZZkpstrd4P4JNP2qDYmdu40ukiiZIuESEX3ezJ8KZ7g7sehqAi+nM9+bzpQob4VOwTM9Fc4h
G75ccIW9qO94HH8bSE5sDWvYRxiqAf+a0GIyPKLvQm6rR/CSMhP0ppeBc6Ii896fj4ouK8Ij+5I1
jl2E/O+SNgjbjSNcS0esrwJoLBl6E5X+Gjg8Pb0h7pQRb660Q0LgYJ9lDzN9TKkajrNh5fWFAUyz
WMUGF7WrW1O/fjGEhSTE03qMO+ioTCNsz0ySrGGtVPMCTetHrZ8Wv7QIQApssjoC2Jnr6u/9NRQG
PEM1qJCwkaXvLGvdbHPKpWVtjkJf+dhKpQZ0UEKKBcC/+oRFW83G8tJ0UXXwAbQMqdYVOCF/SQKb
KYUV+p6ixNPCeEYlVOeqZ1FJUaO9QjcBIYAcBcquTlS6/oa4eMj/n/+3CSt7WWRhU041tNX6YM8V
hRUOAbcVASCSF00thoceti2w2ymJl3ZGIgN0ppMP5/QQscLhI73u87G9Efi40puQueHKUr21OpDz
tMNfeYdrPktkQ7/UAcdDFF0jl6I4LWuyl7M1myVRalhOWO2Zqd//MyQ8/eVMdU+liokZ/WWj7V9M
izp3CwQdjaXuTWw0pUSoaFGBO7e1CJWGNjaGv3On9O1kchz1MaOVzrQci5JSCTpGoLTCLDqZj4B9
6rjBBfA8ad8nccpIURo0Xk7kwmwi68zhy9AUmFb7SGt5HLGPIeYkRNwGu1VmgGHSE1HpDSkVwyyf
juyX0lmcI/ftNh/nT+Fu5SJDT6M39DLhd8/pQfCfCuuvU7ZVAMazjKkLdG1cZEc+W4zD3gkQGyCn
y5iLfMro4f1fHbgPglNkRnYaf+FICZ4slVNJSt0zRlfq2qALzkPMZqxlEJnP2IUISVXtzEVQlXXy
viwh+NcxOyFLZuDs9BJQFhdcLLjWAyTaMngeN3Y/EFmt8ysh8t+r4plWnUglLwhhjYT2QXMq+wXn
oV7vSxPOc6jC5/yxkRSDAqJQOo+Vqum9mCccBslOJhV9aarnRBQ8wwllJduqDM7HX6iSyQv4VeR6
VpoPNkh5vv2ZWs5KUvpaZbeANyMRi1eVGeKEzaLyQIr5fcaxfROSGqTp/4JMSoNgMZUZo5lKf4RR
m63d9RYPq6kxeS/WqXaSmV40xSbfi3K5++MU7o4eAg3UmkRGLRoo2ysg/+NSVmZFEPc2RGJTUNKT
EE9ONiRxi7ZRg+OxWiWQ8HmsDQgCc52v+C6t2Qwl0E1zJj3/IHsWcltb42WwU84jLMPyAQwiIsg1
O7gWqs571he8TIW+4hbwD8CF4zbT5833qDDHAOBpGLh8RZD248J2BLn+AdXwQHBWClRr9t0GAPlb
wUONaLhFhIR9W3ryW6ZNG7SWVk7Yw/etjJDMvuC+XYtOXr6DqdJMYDiDYAkoQcLWqcra4G24GdzB
Q1dzxkykxtCb3vHNAoWLQJtza9t81wrB4ILM0lXlI4un1CH+UEZzxyGbOZph+VjmfLaZzuFh44VC
0O58iyq4p6wCpQ8gnjBB3bSvR2HlIZ5ODvNKcVffyWSe+bz/hViUPH48ZqLUR94THsJHT30ng593
KyUET9IlBJDHSwbhPp9RdVqhsS7EJUHmXAF7E5Q5W4z0TyBu27hPwUolBbScqq1PlrCM3yQoOyrq
jBO/xWQK4RgGcSFy0qbuKZc6LnElw2CyMx+VMJUOvJ64JFkqIRWHooapfVAVY+7H09I9IECbecND
NxJLXdw31T2yy7gU69tBisYVdcj/WG3t7VEsSPij8js/ptVzbi4FGl2k6vHUPTf25Kw3fx3XH9vi
k9yFM3ATdYUHqtge+gna5i/kFmM8KXqhtzThHe04ISAbgmfpZY/Qm00f+q+4N0ppTqguFwFIdp4d
SpRSRWdMQFYOTLd3tazbKoMuK987f1m3sFvD0G9JmjsL/t5lddwNMQ7oJT/42bB8B9eoMJAtOXfL
eTeImV7tD6NpkiDkOAHPqGdbjhGQ8sV1y36F6R+rwtf0Xbh3BBqHv+Y5rarucgMF1fR44YxtkcOn
EBNP5EMXXkGKUgI4t9qQ89Vfmrhe2kJDLsoQ350m19KNeCuInpVTIDQbO0BuH5K7mhz9ibE5cbP9
vnCUiJegA2DieKS5AiUtqfoWShxglDgeM04+KKpBELKwfqTb5uv5eaBh028yeIpm2KYqhBVOL9Oz
kt3uZsP1e9JzlJJ0cOFqfslf5/TlAOombhhX0edntBE4sXyLDlXy9xkFh/wZdSMuqwfOuUdH5cju
DSQ4BbxeQSdHSNOM04EKVSv31WpEuimRxmnvf1KXqVVhi68lavCzXdEQ2XIzRQ8tb91ErWgMVWoK
B5+fL3VjynEsjrkKKLADgbt3t+f9UBqER5lv9S2h8353X2N5NtYI6HKq6ZOyvugQ2MeiBASLLEAE
c+rsYlRygs4RwZBe3P0RRO87laQcCr5LFpvV8/xSgfTzOdhjZrorpIBk5V+R+i7gs3wxPETy61be
XhrJAL1oU8eB92of5JO/to+Z6h28NR+m+QVYZNwfnvwcL3moemYWSoQfVbht65rFswGxbv4t9VSF
ZWV1TeciTKWko4Pnho7q60gtNybibG/pzIEG/YlS1qm2kL9ed1WzndsaZICpTtMP4qHn18wBm8DT
NlJ1mz8IbEXBAbss5X0CHPL86ejlWRFmk0bIQ3CElVlG9Rc8SzdNvkYxkC1IBPZ6+Li44nI3HMFL
l0U66Bgw2RvQpfLKV6ehrygM4XGAfu5BgBhrIK7HTIJxzHAz40nO4J+bNYYashktx+o9GzMgPJh7
mA2dI1I0jVW1cwi41GNKIo0R688jzdikJ4RDNIzZLK/PLGVU3wJ/T/UoqfJjgDxUpVn28uljgu0p
J1UImOXVsFdn2a+vlRw/u195+ud4GnVDEZbuuik0Q5LmlMSku8zDLu8zV03xerqmt7DSlNRhUNoY
1ucGZfJIkaGdyCxVpPOpnnDA1frkjv/CsKvfUCvGYX2yzfpL0fzyjzHLEhkuMUAnS8RLuTuLi4ur
lj4HkYKYi+o0wwUqaQBudov1GABysKaDn5a7pxaqDys8fCwBLmI2+oY/Iu+pSkJEpMyc9ukvMZwF
79V1hJxkGm/fZHt42NJflm7XLdGKkiZ4mU2kNkFHzqH6aNIk1We/CYlTRafK5s/gij86mZjwXxOR
LtglWRN+LwUzkzAbJ1pAJLRSyYPH+/uZsTVfS2Q+37JPClKdnun4xaapIuDO+VqeZAR1KVvOecXI
1SDbQwSaLRU3JkZzgWuQ/xPLq0rck9JXX37sXMR3J14mGrQe1TbUGBUORHdIDwI1t3HPE+beTsaF
Cr0EjOqayTt5R+XDDUOXXIyTUJkFaIjnDK1yWhtRuPdo64fRfbFyvjTh7PTuA0vpsQ2AGxYigUR7
g6UhQ0XlxukCkuBYvx+KO84FODRWqH6K19y636BRv9OYX4Obv9XWqrtIVexo+7y+KCpKuQhgQwie
eJRbwwtPMTln1XL1xAIOLyYMcmzcvX/BawHMJMhaug1PVl+mg2s8KobDDDMpRBtJQgg17kn9NzYw
tvWJFESmCyPL+Np912fzCVa087i0hYT5aBt3jnk4ji0ZvARhMXldaaiy6w6/21ycM/QIBY7U4bZ9
E9MMblyd6+J9XB2io8+uI3PS5IHEr4Au5ZTunPvaFiRbNaXkAN0oq5VTW3oFEOWZzhY/syVI0H8q
d60xJ6YwXigiiWlk6kMsAolGS5zMoRTQ2W9MQz7jSSqys8jH/11ixDI9gDqnpZnla4prcd/H22YK
/SeddLLiq8BrbChV2X81RXR/lfXB4Ozb/63gjZzaduVHv0hZqyNy7r2FTJxCueS7K2vg+IBVr2/F
+bJdBnZVSCDA6Xdpgrek7CrC/F4t6wr3i2M2rmzv1RaC/qY9pWUUbjtGzk0ttccuCz8cP6GNJilo
Sg5NP8kGnJYR2/gPzqJcHnb9IwK4zf4Q9mvYRIu1LTgbx1/zeClT6dTMA4lbjp0NHEQW9TwVrRAh
by4vS0RZ3cidC39yVyg69vxAVXc1iexlPMsX90iCN8zzFBi/lphatdc2uZpW9ov5UqFaa6qKAU/N
lJj0x+AhLN8Z7HTI4K6Kva9+ksIkamXEhRVmkMV7KwCNyFFpnRodiGN6cRWT1P91c+tLK+ifIZLb
IXnD9FOT7vCb3ubnfMesXVBT8xkbzXDGxuVs6D6pXhnaITnRkyU2nZxDwBYuuyKNtBbuDM3CW9Vp
dfbChmTmuj4puiMuscwgCOMkWx74h3+mN+ajAGCFT1cJtvOqUTvBSCOELdIlpHjY8bodYDGgoxpU
YGBZXZNYwA2FBanaaRf9ptO/WLOYQiY9/uxB37AhCZf3kxE35dEeYQlDJweT2Kj95NBpWxpIngs7
Qo5nVWyLjyS2+4Kal4oiVa+19qdMFbaKjQsvU58BnS2kIHhPTEKdcjiyQWr7Bx1zuZD3uO14/J0z
vpumFUhaHxhZdCqlb802z0C35anBvBO/Qo2UA2DM4a7x7T683I7I+xxCBOLj/qHZ0drY4sSQRdNS
2L3QGAsFtUAfsqjTSJ0/ob1YarhMXf6B7WSKDS1WRBK2WMyWxJomGkrEoWLZ4rcICFGnXMYY4H/H
Azfekm2ykWbb/iQLl/CQe1A02SpfvcGBVH5Bt1ahMPLOSSLzrTsOBBB8Ka6T8BF5IPXmHnsvlyuV
UM1GFSf/VgjiABWSY8xP3/3B0QkrESo/KaAuHFKIXqCuk42dFCgC9q0aEIY+tax92twRQL4TXV0e
0sJ57/LnEqXUKD9DiXpfoDet0cqjRtm3ci0ZOTzboRTDdzBQFsZw0tbtBsg2uoj8vV95FnFq9K/4
LWQSO0XJ6Yq1Oe/F1piz0Otpqi+P3qcrHJlNugTj85CJzsvG+MApBpYTIHQPIqlr8wR+lUaqyLHH
lPvLVqkPmwEGEK0oqnbWmXtNMFeaiyTfMQpohmxjiq5Hlhaa5VbmYl9vG9nYZu+4fKCJtvw008wc
TbKkY0ZCei/jz64pRXWFNIn78rP4d2SNA0XMZ6MoV7DbXBWqtz52qArwU/LXzT5nat0/KNH+rgWj
fGgbd8fIN8Ha97NSduPx8vAPgaIdLmsqlT1DxuyGKAbGg+u+M2QuZc4evHOKcVi1fOLq3nQI6evy
7TxMlLXtHdAdyd54pI3gv9jmLc06NmUo2u39u/sGJxXv7PCv8molcZbAF+1AbLHucXPnJWxWf3KD
YW/zRIu9iA62jl5zN23K7NeRnN31p9KTSSFO13KHXoUtN0GwaR4kkTcmaDEQbeETAHMwuq2i7yTY
rxNG88hAvrZhgJoF0UnICT8GJU5xxckAiIWfJtsg+kbLfEnNTiVwgHPI2oqSLi8ofvWmh4UuV28J
Abjb7TJ2uqvpowe7oRIRsyjl1Da0Z+lvz88vOxiRw+/ZcOzNlHsuDZuLWRHIyn8HLiAnZTwUT03g
V++5wVRpQVrLLFeI6Eld/NOVXQ8a84HXAjAV5olFV2eS2bBGwj7dS6rmiVyjsi+qmdbM0hqe9R8O
p88/3DZpCn30FFvf3QV+a91F2QtrQoQxe6JAqZ2qIKqX1XtbTRqs0WqfpQmvHmct07uZA+iQpbq+
K/sldQRqunqXhXnVCe2ObMYVscCQyIiQBiiRXa0L54sJYjDDj6IY6JUoZKu3I7aIuOyG66tSHgLQ
S/n/X9LaagzkOCGowzc01vm9hNFvTKsHHaUYJ6r6+/KXYRct27uL26ZYXmbiK4ExIVAmGyuEDV1o
KVlt5ey1CVBdcvI6VrWwJtiRPKJSsj25fmWVZgFWNF9LoSMeFIiDHti93/eokw9OKnFPiNA/yvwi
t/5u7LwlHQTQ5HmwOu1Vow0Y7SVzyaWsijv5xGzN3uIs52VccdRbmVYlunSONQAE85EmB40pM9n4
P1iA1QknvqNmIE11NGD+R+IgYpd+PA1pzjLtizEFteEsehsdj2d1AQxt2IJf3k8XKpR9ue1Yas1g
GHREH4szpRpjsg9STvPPzuhRnbJ0t8vvfQYupa6sUsNcYGtMp6daR6EpN4Q0+v2jmMvK9iOtWeXS
y5qleujb3JQybH2GFiiK1icEqTQUG7JGxMA/u767tZB+SSEgzLXf+kPhIvEuMBOUEcxNLMMII3Tz
ED1XlOXB+7dUGGxhUvZp0OZNHyRN8qJZ3SyXnIZu06V8aeKGXxgGJ+fyFP0Ar0fqbYzusHYpaEvB
8QW2Tm+W1uxU5woUQR93a2WfDXGOps7bfQCMR7oXSRY1+t1Tkj5vA7NOfnlvKrDt0b+0lFK+JyMQ
qEizG13BTSUYxTYCbrro/oHdIu38jSqhDeLx3RunRnbNuj8uEQWaV39AiyICSgvi/5Srjr92mXMK
yyyKM3MLR5NIGZBbOJ7UOCX0fcelZHsBwMn8oFUQrJVPplxknK4koanL169WG/X5Ggm00cjaT4w5
9tT6xFl6ZhMFH2sajD7FhSangvlLAkHBz9MDUy4CpVEG7Ku6hiCouj1o831yt8QBKOcjPZliMOEw
PiH3prtGiyTcfu080OFdX6wsGkZ2MJJ+dV5wXuohg5JKwhyMuGOUx3KT3gaM4v3LJMrPQLEygFBP
FEesBkZWUqopqt5NS8Q1mex7GRCsqRIcoS6M9SQm5T2nxcINtxVr/XcxZ2IZArqjkTlD2YRtdX/s
NRCB5hubt0x4JGQg7aWcmgThfmzJeh7HY7kfm6NgeK8NRnPKgcyPtO71txytcC465XzS0Kc9LOOQ
YnRjhqnZiV3r/zQ9tC6NPo0Qaj+LUR/7aOSHvDIgffJ97l65ANTR8c7Rpl44hiDYdMO6gZ0cJklq
VxxpvM07qvYiwFPKvgZsqBSuROiSHGwIfEInlX1i2ajDS6pzvYIRNE2XfX6Ap9UjUDLS99T33i7A
eGZlgVPyEDgMKk7/40qDOU4esTKHdtX/ul7y4BTbNaNnxGANbplYveQodgf/K+78nHt/Gw==
`protect end_protected
