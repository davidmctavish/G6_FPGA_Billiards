`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L90xxmHL9tGTFacRTjHXLA7HVWFNIvRzRQ5sEFLRO9G/T+Jr5n2HdIYNX0/emi5093tkJZ0kx5ya
OS9QjVJ63g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VCEKZIcAbFBi1Z53jjCpJCZdKETuny/m6fF8/ixtiANtRvGyQxAIk3Ix2T4NAecnevAOHhi0Hqaf
V+xAyuT6/Z+WtYNs/E1d+0jAyNDz9pq0EG8YmOKqtVBhLMKFMPC27Wt2AhoL4YS/b0m0onWlr77S
hn0PGlkSKrwdeJyjKw8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MgAQQ1pUOsbrezhql1fhqigj+2CWtoo3nrumxAlzz5I0YJBB4hF8PvZoz8L/GXq5YD31F8BT/j2s
NX6jTlge7czjl6xuCNN6w8jCWhk2GKuFo/SxIPXV5PMRbJMZwNZgKcBf4CTwZV89i0dkAbZ3JJlV
5TC6uXM8jA3Jwj87SoL7bPwjlGVH8n0P4g1a6Su0B3i/dshMMbSWc0yzlAp/51vMXcVTfG91Vzs5
2Uq/PJvZH/DKnPl9PhFdopXOCriL4TeVPE1eP+LcJ/2QjMYCcfezmThZ5ZwC+7dU7OqlXsNDlkky
ahR3rploWPtxGUmRl1ErNorw2YGqzRwOI04OYA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
X6IrkFPPr+Gb6aUoGZIiog3d/LHRM8myTzKb5sa10bX486Cj8QaaRLr+l+3TFXZcDP6+C8igqK4J
NDHSOJv4B+SXMfkNcn0r4lgBM0patCM/oy0h6V/bDcer16r+Ok3ScGr7ilOfqouoB2kwbo0yfgc9
rwF27OBjdQPawPZ7tIk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S3qkO3zFykogStXF3+f7Xj5LjoTyp43LjfQDgJvB1tJ8iJulkD/A2ArzaT+r7z5s4RAh0b/9qqu+
N4CKlk9QpGqocztXJmjLwiNEJQrHuO2qPme/pbDVJGzZVX3ONZwuhb+5luW6Bwx54BhlP8dtpStW
NeFdm3W/tV3ZVS1Ys/z//OaIddSoZYXj9I6H1lLaz4h2RR9SVkThYj0zWRVfjeHPGGI3qioyiKkW
U4r7njSKmgORMjLW4hsRX8yoRcv/bZG3MGwdGoYWwlHIM1trx32IB0Hdwd+VBcUsUjRMhiu+mAPB
EwB6ALA5hJ2ta8f1HaL4s9eYri6/tx7ZuAxHfA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7328)
`protect data_block
U3S/A+zauYQxCOrnCyemJr3X1YqRDj/Pmm+BwxL2LY/IpSp9IgyZ67HmjWfujl372UC5zX6YQxsL
QecZ1qvp+9kSdQl7oBTjOO+g5sfh7MK4zlNve2jg+omUm0ifcnSkDn7ORS5VFKz2wu7/Zs6rRGSe
yGURQE5ibO87aF6lbQB1wfunAyY/iEQNLmEj6Nb7LE/i3CiMVWQV5qb3gLzWNPC6JdIH5IVZRArb
/Qke5w6nTMaE/0av9JlmeGUtiyLrRRo8xMW8ZAH1nSppCYkfOvVe9nvzMuyt+SNPIUlrj/UrDXWC
GcajO0jthdtIaWu/q8gYzPutukovG23LEdCQfQIIcRN4YaJaOOw2b0mmpO4I71ODiU9QBId7X4VR
b1BkOX5524wZNJLnU6wK7W6QPbvvtDtRHqeHUJ0NFSPDIcDoqeBpwNbR7oTbyMTE8YWSs2PEjorJ
49hjxO16tS0WyMioLv90U2t8OxfsKI9C/ak+Eh8oSE6DmF94nyXWXwSRDvouRRCqR4mKSl46WaQw
ovjVK2p/M7g62HwxSUXPHGeluI3ogn5MZh/keao8oQRD4rnjtzrEPS8oLmEnExHqEJvuq8eyobjv
UHiPyFN+YUokFE2UFjushK7ZpnK+AKpL0ME3ia0t/V3ntBft8scZ5APP+r8C6zzVVx6La7PiRz8V
vbdZV+8eADZqRwtnZ4r27PNS4M1B8u+eAYvx42gxCTZ92t1REtJgBjKmQB/0slLyswTBxfgIOgu3
6KRFqGNzg+6PgWPtlS62gKtVPqW/ovSx0j4bsk1KSpUxkvUdItGXEnxgvClwDdkLcsOQjLiJK+W0
7JHWJ4gaewRiMN6AQ+vPF110crOgiVStUIxHlb5oMFnzqxRAucJguZ1XNUeUG+6I9A4cD/8jlo/y
sc3ycEPgQG+ipKrNTa7626q+bBeMIpjdq2KNsE/mqzsyfCKhmwM0Ia+71GmVDvtgFBtG2oi0nF4i
F8RFWDQqCMpQrp9HfyceDU+MiTekjq0Qt4zMFwoz6pB9n+HghL43XEsOO8RN8vYnKDXjq+BtcDFw
kbjH1bpESbr5SUvb2np8Ag2NTminKh0mgbDuwmuMUlzU0KGBUVWe9ddiioYQi6HGfJQetBaud3eh
2Nnz2RBSVg2KWIHTmHe6pH4dv1BgNXxT/LcwpBtCJBaxgyo4R9OKwbmBtfpad5TWY6u2erVbYvGM
HLnq0DIwUhUjshPXjxteOYB0Z3gL1GUcdKYGV6XUSWC+UVgkzrqQlcl1j33o1kpe409NG9zGpCPs
JNasEs2I3HyPlpuOArGaJlE4aHjT0O/5QHxNj6d9M4YvRbZxOGvSIALuAlP2PXnX8trq/7tfvsou
FG5bfRK5GRb2d4KIftghLC3Vo+KOJsE7wHWJsMPujSgL3DwbMdwZEpiWlmsg087HKfx6LTjIC+iV
jSlpdR65C0CbqypEvRDLTx+IysT3gRKJ2CPc2gzNIs/HX38EIp+1lyqu1mkfH0QICRdhw66CK+6C
oqA2kdW7GDsNZG6FtVJBdVQOtB2G6VBqNKFz7xCh1iIEWGxNLKBAf+IA8qusaDt45qDseavk8VrA
U5zEDnqPnAjdT4aDRzDqnrqoO5RjC5q1UwpyZFIrIjRioQo1ZNS3WNox/7XQLVPpPDL+g9uAVk9Q
nF6wWVnCCrzbeqhjgYzP6uPVdRXK0oE9nzkFeeI26zYL7+AqAcg6hjYaPUq0QUovnwa1hK1jwCqG
aGhjiW+5ka60u+fOiChKepvtUxwGtkdl4bc9fxWW6gxBqpgNapgpJI2LS+BLKRZNKuBm0Kfk6fan
XsRwwA3YgcY4yqeZ4S+ZHkifLw9FKoJ880qR40+1P04FUvlsVQH0nhmcgTNAxAaMRUFwKT5C6nWq
zdPhsQO216EuEkrZnPxL5heABjWH3+FcHp7y1JpQpI/m9xp0Y4UMa/ksyWEfTaNj6N6rchNAodq9
SRrehaOk9TpupAugFuoz6RcpQsbtpmOI07Xo+C0f/i16jwddJP/MJy2ShO0uSmjdhj5oON6KssSp
qqMvKS6fx53Ch9i5GTXQbcvwvW3W/UX6KaApKItVMa/qy2KVYiTKYnWxqIqFvPivdaJ2JoZrNOLu
kl7WHKuFG2eHTAedgrO3s+EazMUjHJSeTm8nkkPr+ftLzpZd7H4WKZR/qwZnMSyqLGHnRxXnFFfv
iMWzYmtQZFIeHBLQOLEZp83PLXqyvovKpHNqe5giI9/DYTOBdwM+lV7Y/M6Fw3RacM7ULeipE/6r
a16sy33IlLtlHXg6o27ttv7BS8Y3xkUmFXi5f80A5naFMazsXJo6VCijoLW/4H6V6Tb1589VMHWp
GPPEZ1dHhsh0VfT0zJnFgJp9CG1rE+h3JkGaZdpHD3MzERpIzrv4KModKxReK0O4VqIJgvmFzJvt
v0qbOD+9YDXgRnOAaOy1+tHzZl5hAHZkt35mWro6xM+Q7Ptgbp2xBNbFXlrnRzFFJ1S6pqqwDHI8
MRwF2qrVfnYdHnO3Of8mNxtH85sKrI9n+WvXa2L8fHYTpVhPXpeQ7rDMWU6m3Jmxz8FOOA8Gj3HC
HMdwDK3p/MOBaXxjWfP+hL11teI7Pixv9FHm0UHUV28IRlqtDcVBksHoIIADhwZawoQcUmiM8Rtb
nzaXTiWtFnjUs/xcc7H5P6LwkP156HfOsyICI98nqg0PrXSiTPGBf8WxUdvX8DEEQk99Qp/Qnbv7
LQsX5huy8HcLpussFwir+63IeGqI9os6hACl9xvyNGm8VF2QBdeRlooTbxcxZER/Ifzb6DNDFfcu
GVTzTbByCQTDeClJwqDB+U85UjJuFjH3d8JsRveMxIGgeEV/m9B1Kns/8Zp9Xphby4yFd/8ulkgD
BcljVSB/UCQM0LdmI23ATZ/NMGnB3yzK2nCD6+tpnmR/bOJ/Z2jdXCe7ZTkJlSJqzGUsjVrzp5ty
7gMT+HHYIjZCbK/PhgrJ2B3WJqVBfD/GDcnlcjtFJsV7QS3T4gtum2p3xWHcPy07r4LgBtIg3AwH
a5nlY82xV0qCb0Cr4g841eRoa2/OJHwlCDs1RLxb6uNK3ZJMCeZO9YwDEQvSzEqwEz/bed58Z22h
IajMsKuOV3NCmYuaU4vby8vwfBIeFjFVgeEPoDL7M5qo473z54iT2rK4jvqiNeph0dph8D3oU3Qu
h7Ns51jKPvb2Zx88rHqatO3CX80QXtASwdMgYYZdcJonbxFqDYOFo3N3qWJgMMBJMEMgeXZK0YZG
Uz8xGFEWuD+cMc9N6mhNoxsJETZdin644ja/4WsgKrJzMpYl2RYW0e7y9Ra+jl+8lgtYsvHvtbA7
fCzIU9t9pVQC/9qPtvhCMVrhJTivSI5IPUw40ijIIMc/3eqx8wAPPRYGk9qk0jENlgK7rdm6rdDy
h+xk4tXd9DHHCx6gLzHML9wn1MzmUmWN36Rcbwp5+XjPsFPVxYy/eqr+s2kVqAWo5ZSLV57JdOPf
xKuBcasPgiWVp0dtxl1c31WSM2gHeRLUgbhWqUGb+jOpnqtz7RLv2PqbRMetJoHVXYXz8XByCt2a
sgsrnUKyEEDrb+s6qDIsUFfs9mo+wFnkreham4WvitZ9Add6rXt6GogDAPLwoRVAUBK0njeWjZO2
G4dOXWZk3UXUW0PkiCd5027m3WWTdVyn9//xBcSr9JvZ50DeRqPh4hu7vvr1sjDjUf5berNnrIzp
CG88FWKZG6rtluvsg0SIlNcfAjTqw74DjgBPRqwJhnkA6yE9OGUVq2sxpqr5/5qBPD4zi5TIxLAT
0kWEwgqx8Tl0FyOF3bcClG4YV+1Kz4H9D0gS0ZlauQJ8beq7uctxErTaOvP/b9p/eTiQZQaBOVMr
EQ31zNI6nofBzWCmjmMD8y9IzQ+Sc2umk5SFhDE3N8tjD7IGOw+KtPiOceBUnAOapSWDzPh1geFN
DrYmJVt+pZLD/DpBK+052SFJEVIaE1vrM4V3N366l4o8CgMy62H8G9EEoncXbcitV8WlzmmYENMu
kMuRjhSZOeBQhiShjT9iG8GasL0BghiZ5GGeWeP7qtI6elj6GIutUPAkRKIE8yUKRLlY06yfb6zG
ZjEBf0ut8+yCfWO5uTjP8xcp1dnnJqyaK+ENiPHdef2KkIHXOReTcD50S8zxPAqv+Q6MNJfiTu+p
nKMjZZOrRDg/GYJkNTAXlp4aSQYBIEna4ZUR8twAANkLwNdeZRuYDC7sShZG1Yv7rkpB536nfWte
VHTTmW0gyUi/Qujd2Hk6XTTMqWVLt4Xnm/vlVT/mmtXWx+AIMcBX39+dZrGOzOQ8oJrIgFaPryyL
+W89mhutAmgEtWpJdKscSODaWBglL0np4X/I4WKiDiRr/Pv1Uf7s1hq9J+wZaITs/lYPuuJL6y+X
eZq6me/ul6OF+/YFcudoo17zQ4J/N1sKyy4RCyUft0YlzP35OeKeb61Xy5XR2cze1okDZjZEs8iW
qYgahuX3pDPP4yVxxByYTifC1WkTkpswOZwagC3Pj6o0edSnnw6fJIZlULgO+O3eGOPEe4bKuPnl
kOsMd4T/jqjg4YBacBRsVn8bnywrqMyZ67UuiiMA0qQ8B7QroMIkoHhLwJ33BSqwdfOGBxMD3u6A
VDd2X5ZD7VmPDXtYI32NQ/COp+Ptf1+G86ipXDhMIhSi+sQYPkG1jxcHrC8Y23/JJr+cZVPh70XE
FMYN4T69MwTgD2RSpy/cSyliBOQ7oV27ctffjKzba8GIcEnaCcL5yV+0mU6Ithx4OAHhufCEo0sL
XRKaAN3VybMY63lCBeJLkEazuPvxg7YAijBjT9JTdhkRp99fqjlDoqoyVX8BOZld/tK3rE8LTv85
LHLvk4uwn+fJy2a6xTLwlmGm0GJhke2pWQ4NqwHGscySTEsA09LacFBvyjdvtR9hVAdnLBRDVR2+
LCa4+siO0Qe0rcwLbY+WiUz9QqiIqfMovVcfBh1sMm6S9OEvmnlR/R/CoEs8H7S+ckfuob5KE0B2
qqCzhwEsxap785B6n4U5YugvJnfedinI/PSW9bPaCoJASo3hIVMb1hfUIrdzPdDuBNnOIvAmFCfI
hpDWvgjFE/GJqyO8gMxliPn5HXJkxoxNtjGVn3hInojc9xngTWpbR8P+0ZDlX/SCn8bPjoTx/5Q0
rytX2SdI6YWLuVPXQh97z9ecyWJfqQF+GGro8MwhoxabMOguQy6Nbm1oOnQjBzcgY7O6DaJba7Rn
uRQb1p+PaP1ddIDIsS0kvOdFI6ZCMJMnlgP8ygyF/0huLEFowlbkPS1NONEKYGWALbnTQkZpii/M
Z0ytuoM+/kYZENtgRfdOlDwak9wJAjvqBpP2b4ID5dQiELrcgDD7ST3NTE/RlJeEjrV+CHmRLCLI
PVEp8MDgx/6nvxuShv80FeyA9tIwoy07DvQ3Q3dtFY4JyJ1tKzPtAbHhs7L7qGFaPJMKcVf0KL5i
Re0E4vmX1/NgUa0TCmqlflLmn6lyGgyc0JppTDT9d3F1GZ8R/cIx5HqyJoIf1CNIWDb0uP151Enc
BrNwGTKiWkeBoRlOHhwJwQ+n3MVGp4g2t3F+LnvGUw6D4vkzypRvM2xwzl5N5QJPT23H7LW59tD7
jCeS/+BUvrSk+lc7X1C1mmtY9eIhOhMUdRJkHai+FQ3Y6gN8WAYwylqvUMOW1hWdF4V/i2FY2/mx
2b1uto4eD534GqDTkQdQL8/ZGkCQcjrhhA3HSL2DuajNFc9a5WJeneJPB2MqlQLKrWuZRf6GNFTq
y0cJ4O04EVqZnz7+p6x0XSt7Jv3Kq96kDXsB89bPjp7LGBtp+S+H29tpocVVPtcfI869PM3mV/Wx
Wz+BisK+A8lbjWKdX3Rwn+DODGbu+Ypw/3s8ZY3wQQ8xdJeJ2VBMNKBBFdRvcRPw+ulgjho8aX5u
0kIchVR0zWmVbmvQ7OxqvbBFf8tv/UCcDSDevhypwRZK7NkHKy9AJ50HpF0PO6DUa0gR92yTyuJs
q9kGYS05wOnzW9DXtGGPQI3MNWos6iC74PUWqL96XWsdUp1+EQ/Oute3f8OQSihv164yhPQiIkw8
FGzLu96PayR1q8Tp8OGOf2LcrZLD1yaXjap5LIN3APdsyTs5CfTo63ckNSfk1Q8FqrVFJkeAPZQ7
2OCeRKp3kgPsIBMarqnI+Hbt0OAJROITwaJTAIqCcR1EPcsTLkKSyKW8cTNKXtFTI2UbElZL3u9d
bmiNhAhfiYiZYIloaXh7q/WFlvYQT9kUewTUSAYx8SYS7BvonvI1qAYbirxVy/Vv2huQafaDfiCR
/+5tJM5V9xeO1uNkOei/hNjPg0OkzZ83d2dZVswje6cfgAl54eNhFEI1VRyZUmUCx8yCwl1LD4DT
GGoNqJcvId6PSfk+UCocVqyl/2rTOIVlsPhjAx8SAlKHMFi8umGE5I/5qyOzjh3VfD7DMuKzWWJQ
hMs6kiSvWlNkoWv6QtwJLlE6qS5fFfvSWYUVaV7U9Glz39inCnbxF6CvoVQwlODmHIu4rxITwxsn
GhK8CAV+Hiqn7uE190YgtZGlQp3PreKsnuor5vGVHbjqn8T/tCfMESl0RbZWKf9B0PIke9zPsrer
TP45g6HTPiRNwR/xUS/QsFbLLiPRr+D6uxtURFqPi25UkMpArK3ueFjE5f6T8h3Y66bVD3ObZJlp
Ou4BlD/f1rnS/N+tiJO0fA9oZ5DIvlprgLFm7/n1jgjGC6VcBzNfACq7IfSiPYHZX8gNWMughi1s
xVjz+EdE/00kDPZwOy5Ezbb/lKq6FmKzc08790BTtztFmIhagu/ZN0WWen65WaRfSPqudyZo2K4K
1u8BADVo2QLT4slBv6Fj5oT5eTx7hJ2lnKkc0oBTpdJX6OiIsqaTrhMrr7zdK9McrNKW3GgkGC+Z
ha/NYDxMLVux7OjeJRpHqj1nYG/4cwRsCGihnXczcJU6ATUrQL4TDiZ0+2oPCUNEeD4UsEIcY/2g
NluAuBbH162jdNehbmVzU9SyuKEok4yJXncHFPUDbjPeRxp0s9MWJMFN1vNJIve3kZQCgbxDmJUh
IaFB/f4fpr454Lb2BU8+wu4Sduqs2rzK4CdeLuSlaazEmel13gLQckKA0sUyePE9QZGPiq4Y+Nju
NYobZIf6lpcXQ9T3N4ghSXDt89A19MA2d/iAkd/ESZT3ayjcyKGZWrV+XcD5hC4ElcYghH+L6wGL
p4SS08BIcMTMV0nytslVPvrkOVRITJY3n5BxlP/0rgKA3vKEh7+XVk3Vd+CU8fXZiwAQ/YhixX7H
3bvdbEDLWP6nR+UeXU/dOvZcC1+HAYnHAVHDYppzdD6uTPeW1Ud1kHh1xsFrtf23B9Qtp5Xl/3Ms
LO9hAQz8K65xn7rc7DQev5zPwitVH7XZnJ9nfasv4+HkYBX1JiOtNq38Ih8grsKNWV/KSQFsPFBj
J6E37/ZmW+CKLdKdSJytfkcyXgqBMV9ywTWYx1qYjuzGHZmKZ2H69t5zOBqWrE4vW7tbCfQ/nc2w
LSXkucVp7/4ATamTe3ysfVmJSayQqlOkMrH2mQ5qY96TvLHgZNNx1M/81b9OYlKnS7QzJwXj2m8E
kmibTVGfIgxriWLFswflyagymGNiEOuVJqOrPWNjYPQSNUxx35WpvK1uUfpdG5QeDZ7qtoHNxEpX
y0Ow10N9WRHmgJ8bVXHXoB/56vAdWG+BIsLcQ0R17z5ByMFwmAFrDGtg7V3Ir831yYU2htdV3x7q
/kpnZ/bUU2vSrdAivPV7o5sWR/WcAXJPiljABJunB6nSf6HbjOLnaRQEYnipj1qTDGzqpCAotfnR
9rVoX6qnbZxob4MoSd6vUu7fg4fTDwwYaWQgCqSeUCL5q2WBuLh6Msu+YjCV7fHhwNqam+Z5ZCSh
+dxMlLeV0FzN5Y1hSZXxBtM3sh21qmr/sdJU9s7eQuO1uiEbacnrfmSYk1ijOHnvdoSJQAuri7BX
V1EVLGckennanUIo+jnBULQIUHh9GUpmyb9CJ+6gKHbxADeSo1ePUyuU5Mjnb2U3EfSGAoGpo5qJ
VYSVBn+LWM7uhQRxo+a87Qkb7lNftdOWdDiVqxFSEXYsoQlPk29d/UpplbCNj5OTkOTbgeOOmR71
bVRNUN8mv7beFinHP0VQ7QKPPfzdLffoae4SZ0ir6WFIvq5TRVEfV0gCuvBgE2FNVbNYwuvQKcDG
oord/HKQkp1AFWx97ARBZPKvMjyKwuZggatqMzOvxTKPo+o/W+HfEUuE2HP1YRnPXATpxmZ5IX7g
bktzCZG8x/55jZvOOKrSDfqCGfsDOEiho+GkcXLRG5J4y4aqUUT/+SSDUAHniilkIo/G6CuudBad
L7e1TT3CFHThADBdnbMAS3qTkIa9y6RwGyp4ItUxqGKQIazqIpejLcbnoXQ+GCSP7DYgNeCZSvus
i1P1c9boii94xaszx0JVut5mj+cLkF1qjLuhbrqXGxF1rO7uJHvnTjbJyNUV8U2247ttCkBXNLb7
qRUGQ0WNksU5BPlNiYgksPFpI7ROErEZ6eJmSrTHock7L0xTSWRVsXiuGNPiUdWO8z0Ld5kwFaHg
UHFjfaZ8gSCOsVwcf6eQ9YZ9JAFprnHADBFa2WqanHClmO9JSqKo3GhpfRl2ZU2JO37Mec7sKf9n
11W9YBdmnziMysDrePGZ7N72UH1VGzw2tvtuRh58geaDBr9VELuJ2io2jISXMSqKQ/Q0TxCl6bA8
TAysB5cclSG1oygjnXjJLUlRwpm3AZ9/YI/Uodr8/2BjxxdTKrDVoVdhHV/9Em8c8bvrUvCJtU3P
j44gUbRdpTozHgjmjFxcP4bQTXUZNqMwCCBs4hU6PQy1r1ywqw1Iy+qS018bcFvbsNwH3frJKPAQ
IQ0e4q59o1BCZh3fh+0bcL6p3dVIqOe8W4s4aBuBVHR22OI0IK2SF+h6J3Cr+iFS2RD1nyGPFQCk
Ca9vib7agAJYhvVK7NhCpoMvr+FnrHwLTMBtMZu6VkT6+YrkeI1PnJJtvnh0CUxAo498GzXJE4tY
+TzGUZfUAO6gZrKmlnxoen2BAOODNykNEtJhUDflqmmEFn/Qpo1Sf/E0RF54JIfBXtpLr699Lk2j
Anq/ZkrIKJzqy4+tuPcwcZfz6j/V6vX7Z99Bp8aeiQflzdh0py0OauQG0j84nORr8XpUT5kqBoo3
uFdqmEpjRb6kYF8peYRcnDGOOygLtvnEAQ1jXS7E1CS9tkHw8BNOz9PurDn/L+rqbHdQwUh8VQXX
I3MUNhSBMYU3y0GJ4akKsy8b9L1K3bNSLGb9t5Yzfzz1fQold3pNIZAs7FeobjkSoXcy24NquGGb
Jl7ZgBjh7UkdYQPps3q2RCs8WeWOhMcu8e93VVL+HraThmxbIl7mOFGQbn2At9Zs1pgPsCeOXtdG
9MeG8gGprdn5xvbMQIjvqPjlxuQgNfF1K0hqAIpmC53kIZMgipo2kah50mFNUfEE6jwrd7cSay1K
jLlg7d1CSTcrtY5Kex3Mo3X1EhEkL4f9kWfOLKA8DJtu2YVvtXolfIaJ3B7XY3rQFesG9Z5H3wF1
RmrgQlI9LoGnzhjKZnhTgU1R9NWsWQ/yO59Vhz5NT/gSyWy5Kb3lbCpXB4sWlsCmxGSja99Hdb0N
q8affz6fmWX2b8654uN+OvQnaeam6Z5M7la5oVd5lOpCgeu8C2zUpmd4NBSzbPMLBl4PWnqZ0dlg
fPKW+rFAbDKaZ9rBNwp+FzKzZZ9QJ1Kk6XhwEfq9Cjo=
`protect end_protected
