`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F9J3PCfV1jQN5P4kkdsShJy78WSiwQ0/6K65myKq4FRT1xUOGzS9Kna0XVhOY4PEVKP2HRh9CO5k
U9fyexo3Fg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nbfO9eqCGRo3v06TEM7dw5/MGE4zsrG1QCDGH838IR9oLaLlmbrYd+zRMzN9RrHvqiN5wvQx6V3g
p6eoB6dPn6VwkZjH4Uup/aiAe5X2NZVqqRFimFscv0wbEM1UwCjajg6I+wE3HceJQm2hMe1kj30R
irqT0bBRkkZY8+nWxMs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iXEWlOaN71uLMcH8HFaB/6XOpE1RUye4Cc8FklPom69ZmLCi5RFTo3XkDm3NyffW52hx8lrYudI+
MxBMfw3fEjOn4NOFYAz0coofdmsWMEiqGmt5jZ0zOriTl3zPtIOGMz5x4zv2VFeB5PEU1dOrCZF+
+OokchWVh2Yo7GXZiyTbSmACovk2Xbk65vE1dSVnhI+52hrYaiFXCv0oWOZVLHW7IxC3JvXYfn2L
5AQuUDZl/fUUn7r9EbX3MR/7QUZdv05fiiF+Rh6aBqzwPZ4GxglqSWRSuBy4A0OQIWPCVGJjDgv6
NKAmgSzpJIWTXqCEB/5IEGe4lbVEGvaoHJM2tQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IstXNjQDY30yFhod3HqYVxBJOHNrRykE/oIQuAs6tzxrBq5mZmwdHXtN5xCZYQN62HRRqxPt07ly
VZo2nfKeQpFJDSkR7FwrwaOZDEFVnnmg61yIZCsCc1+wfJEVNIGR9Z50riHhscGOGem27PiZkSy9
FfqTJbGd4qsUrKvkz8k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OECHQHVOE4gfUhpCYJXfJsIgKZTnzVe1OQxSWG0ACuSvQL7FMmDDuGEPaoFnUZzev6b4jSDvtgaQ
51QndLcVmGl1+6fI8A0ymGuoem3TVJp5uh1l0+Jse0r9yYLNyqdalQPBALM7yPuVk6AszaOSi0lX
BQ39aJEC47rOdlruK0qbMM0gM9rmkuiJGFpnyrWO8IeIlW5KoT+9J8RcEAjeKgk3orLu/U6x2qW6
5SiMX0oSUGomUujV4QpNVqcSrJPc79sAfhwL5juJ5I7wrGlXaQ6jA2Co0D7sBgtz6tj/2gc+vxKP
5uxkQTcOJrEfvgODgfo9Cs059g42hMA4GdjdRw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 32304)
`protect data_block
O3dQr9SVg/B3EBPq6j1jpsReHCuZHTEgKP+UzB9oYXWvRjj4qYSTxid0jtEwPIFZSJI5alLe9gKG
Mp2uGicvk9kbZnqho4m46iD8XejInceomYoozgtruhswD0h5forYWgmBkT/TxbFMpFOFx7H0OJfo
HVbEh57mwh3t7t2AaNzDfIJgEF8NomV/r7b18M3VwT0MZJtQPC2q19irBKqDFsfq8BYFaxxAB7Ht
At9XQ3YC024c7lCBumBtM+JWpCd2bd948VHWUxrTS6sX9MF9x/MjJc+UcsV+Wdp/ryyTIIq3/v5v
6n2f+nxyCS7fit2JpEsnqeky8lpG2jCzm3msJIbWBrHwSKQnO94F94YTmsMoJ6XpV9A0ocbRYqnW
pKzp+GZ8A71Fn/C9I1o3mutgsDKabDczgCI5algugg6qRIs5izloCn3H71fqJB7DhDR5ikKYLTVc
N3c1pJXD6DLRZeUnLNYJW/RUGy3xXFif33MwNtjrmI22pKSL6Dh2uphZwEFE/9n8ROTp9fLRhLGS
zSfr2OHpJ/kLwWiYGVSplNA80IF/F/ggEVqgduWTVtXVaEIOG31HjEotee/SIYlpyqBpxPiYbFRr
xYLa2hHwVgrmHZ2tvL7UdywRhzK9/UljJX1tWQH+BBLaBsOloSEoOaoodU0EWZMltXvD1hOD2fu3
AtIB1k0RhgmsJP3mPq8XG4F0LTB+X587H5XwRMgkLJBp4ZejrJ8wCkpJKs9YoKMrj6to+NBAHBu4
J3nKZrOXGuSpzsS+7xW0A89RxKOOVxgvAhMgN7rMtSpWTPA5YvmHA3A7qh46KzbEjAUCBnaTBxdv
go/OEDKcbm937Zbx++Ui97JHzQxPxxz0y37jpoxAhacUytMlo6GlHLgL19sO24OyeA+mm1Fg6hCL
Izs1axPZ1ZFqyfcdPnlRaIFULJrL0o5ogZwkJZxxZH4j570Jqgk6YriQX3f67QkxZVx+dD67fUwz
xt7TdOqvJIOQxGQ3mq8XOJdH9MXcld4bGZzqAkUBktNW3cNCq/UXyu/tmEY0n358l3knLZsjG6f/
qD8ymBstyaTN1iNcL/dxHnxF52s1FaW70bNzpSvKUqJoW7TZK5Uk9oSRY7CkkbmP04KoM+mZMn9w
zK2oVfZBGNzDRo5WJFXlqe6NgdA64I1D/E/PigQ7vJtXIibjZqFZIUdm6j6ud3Ko2G04+rx/rnCq
OGjPTKGKgZ29P/aJMyJ89sZLGQ0NiIhQ9gUVNI1MIN8v38ACApKfZTpsgKQV2jiRsIuYx/1ZtKhk
XzUJ+DwXOY4CVP+ORM2faN/ZmG9dpLHVcdwSOOe4G4CuZ86eDZMRh7FcWzkbwnOsFbnqlOlxS1Bs
fhZp1nYmsRo3AT/gBtQ52F4Ks2kd+Vt7h9N+My4kpgRL/62XiIcFB0Vfb4uno+4KwnCTCCa957oW
NlCTuZjzY3q05/Tgwm6vr3CqsHMFlTIQjDzU/J7uzGpOpuRPqeWqo2nWAjI/COGnNUBFNk/HT2jb
BXvAw8ewDNeLeB6j5T7kSQ08dbf7i9xwJaeqyiXlu+ghD0veh/RdBEphRruH1W8oGUf9I7hCHZWX
99r/h/f9ffNIRCiK3LhJYoBrIwm36fNZESs0DNHrMXOQ1bhbHv2WZ2p2l9dPJ987RHU1lVV+czQ6
brrFZ79TlFpKA2flSVrkx7NYUPtEq1JHsdsaYbQ/hQgbAy0zk4Wr1xD0l3TE4Ms+loHgzTujlNDX
m7l2H0FQgmzZ2WufqrtqReuH9iwIftTV06loHxQbmSbQqRDi+qhxXS/LNj+hPpcS78GALmoD3U9s
pseJbi6ivuALuCcrP3N/R1XDxuh8r1pDRVY5yNKq1YeZ7/mi/Fw83dwpZf1DMTUvaNysuv4k7xhq
5X/1nE/JeQ5daNFqiVKSMynz8SlC+2WwHGOUxes+IxfUOClkH6b4m9/m+g4VGd2UYp4BMI6dQzcy
igKJm+KgGfipMBd6qO+VTtWKJde8PauOZkEfBgFlQpxOrrI6bT/jNI+j4sbwWpJP3CFciKdq65QU
qqTH9QRhYcZ8bS+2OFjOdg5Do4AqVQryFgLczxXLaIfcSfa7eeqY78ewZwVGhE4sX1rJe6/Yvc2U
WRR+7sCyA0Ut/gF6wQ1dS78iXUIU5wWKh/AWufCYV0TbNYbS1vhWf26YCHerKgbHgyjtrc7hRp8K
uKwXmpyUWfwXsdvF+lPZdbn//y+kWBOzIM+3IIcd9u6WvoaweeIDRf7YLq6sPVlgmC8G6DO3rBUr
Zr1Tvqa5Weljk/sXpHgWwFip1ljm/LYZd/IBojEHrR23NC0pa/v8cOdePFk8QrqQX5UVW6n2DY20
ZbvcSSwi+m8uJRszv5i4IZZhvcanfv482986BLM3TsZC8AgP6duoPRyTlR3E294RA1v5AnwevDkH
lafVu3ugdlm6ZpoxbaDsqTGfCJJ8xeK2r9XxKfEQfwHv6Xn9nN0e6BMxi8Idgn6NqyXdVwFZk8Cu
vhKKnCu+8kgdPgdCV9o0hsmNqsFnNIe3ZxD7WVvXKcHhgPLgRESu6dAUoDoXADS2o6QrYYkEHNzq
gAq/Jg7lhMxr8wl3g+s8K72gQyNOCOa+FTrkT3a3sLSesFzAo9qeesllIuZdqJNwS2ZzFHBOQ6XW
rXiKF/l2w6K+BoSb2JdoGAC1BzOLxblAHz5ignkYKO8nVvbJGY4uK21zr2fzJ5kASzNfSX7Yo5TQ
M6sCXcdbi+pC6iuiXTPg1wozROrLvhG5zcRZ67eHQ3Znm5rxw6WMNqXNjks1Toe2Lvuf9nTQerjQ
Y3BciO/yuo2JmkmfHsiIdfmY9d1iyObyHyjHtNzm3wtuffAQqWVPwAPwzOj5PpVAOUC/+jflzgWJ
qHNcdSrDZsHwEFxw9acIURWBT9rQWAI5Cf1ZC6Wi9vUZDX5bEP+esqy6mKSu5RpjahtlfGOSRKTP
KX+dUxIBJouCwnkxf17m07knnW9N0tennHrHBvxOP962MY5XEPpk+o0/cReKHnMkHBZwCP/4xh18
6xPoPYgIAIyz64/SAE91+QAhBKe3EeUcindtpDM84MdBX7n6IJ9gHl/3mq133L3uLrFmYM1vRzZC
w86uo/kg1ibjY82D1BFuKyWk9puIclSA7LzXo/zh0zSXfkM8t4b7qgaPVjKFIVGwbnocwO9rdguB
PVYyGmtKy7/KP3KoM1CO/yGmThPouVVQr/hN19P/BIakX+vEwUzbZW7powlk7dQ2zGZ3GUSH0YAm
7cVrrUYaqq/ZfwJqSDa+FeR0cFmODfXP5ftAhErF6stbtUkA9oVC5TgJVPGi6/AZKt+m84d0iAwc
NxMQitLyEfaDoL8x14n9PZWsy/8aPxedB20rnlhHYI8LyNFaKB4lGt86+vE0jMDYyd1WgSudorvb
wG6+Xoz24tYnoelO9mvDY5O55+D5BDAHLW7q8YqZCeiHHys+FyQN/3FPa9SkABadHZ91ON/OHt+o
trtUx9If82Wiyr07nltWqhPYcrLAroLwU5t8TtZZ+lICQ8L3RoZVhWRwR0uI6Um3qbz/zljyH6Ct
MkGWco84VVHCNaY43X7W0ggP2KbHbFck1X5oSgvjPzmVQDhb69I0WRMVyirVrn1MLaM2XArxNYdx
qNDXFEXqD54TOCAm5Bz78Q9duo+NhAKy5WlCfYbX0wBR5phatjMIk8+SEAW7vljUoJN8biN+aYOt
g7nfei2i95Kgp0w1juoY8nxvbGU6UkVTguBNGnxKas/FPDaAQVFdDAolBfTAahygX65RRVtI1FQa
I/sI9gwVAsBXozXcns7dOLBHGsBllvtDPGCSXDX++G+AYqy7h0QDme5T/WJhOitJiAcihDQWYCAR
0fa2FpYWdd540tvhUYnmwlqUXU9V4mtqhzaJ0MHNFYFbIV6UfBZFyo7v+U+zg5yn0dh7fKeroQpM
KkrEtCAe3RZ0NdH7znhvg0sY8wdDPcBNDAD5cC/J3qTa+L0iipPy71R+XCQ1fDbPOJ6Ua1FyXhAW
CWHgMYh/2utkkyiWC2r2Q3yyp8aylEUR7z34hYl2eBGreSBZ2NU67uOdRFVA1in9iWMNZFEfs0Hu
4DJSLlADc0l2nUWSSbYrH3GPVgZYhCknyPgEhgJXpCKzcY/BQV4QeCKorvuXHTgDeBeaY7naAnYl
RtJmiwH9q5OJLp5owCJlbtO809I7FdPhycIfvgh2PIxh9K/uCpvLi7hpVWVTcEFcfMiz+7P+btFV
b9T5tPOZ4TKfguD50tXiwI9Wv3HysaI+JKXaYmimo4Hhqzq4ewoQ7YIJOJ76RlDfkjDp0rv+PPEd
/+94BCdB5ffA2w7CmKfxcWNuwOaadbGGhtzbIocakvxtVAg1taRVd95bJ+DdlPJlRdE+KhnJ4b0U
L7e0WqSh2WfexWGym9UcYfdUm9exG+QnOi3G+qy5U4UrKrxO0fctePGVJXKU82k6JA1Q3ziGxvwH
sNvqbQqyv17eKVNas4QuRj6Oza05HWFWqM6OMdIXboG25ZwM8ay5O2/9rHealf+pTqPfabmHlTlr
zxyj9Ihc5zBR+yyT5A21AY2EDPxv6WlGI05dd07Bd79LZ1BsNWbtkwGBWvLE5RUflOZ9QJKfhXIT
mqfj2WiShtbGCrCIiCrMzlteNJYKAJla9o3Cu5o2LRWzA7rGAej0rSe4D9Q/5cmNRoW7Y2Weojw4
n7QxTfr3QkxDuMVQ0KijuBQlDY0TDx5P+oOwy3dH5cCNqur/KV2fwSrT6mDeXJslcQLgybcTwm6S
NkekQHeKr/2zSbArklsk9ZTpIDagy7L8U+qvTXCguG+x1YLcudpgzhLqpmyYyYbvodwpP71PwQJB
dSxj7cXHI8xipn901uQzIOR+UCbUAS22GgrBvHfAV6i2Qbr0sdg8mn4u0tKcW9LGsK7gOtRfDAjX
6yn3NYB7ITXuxQwWtPyBJQyhXlE+6GyM/JRCykphlkMZJY5ME4LbCevFLqMv6Aiyml8/n7JTDa4z
HezKgT+ro77v0XWizorST+OQf3lyq+Q3SjwRmVOJ6nCgcPk64Ond7P5n7bXU9c5m/fKChaa85DuD
LH230zcLSkgxcSDoPxPOcA//CDd3KpnQ+wvsBLlG49jMcIY6r86Binusm4fnw+wz2LlI9SU0TuHv
IUGdWBTHSuZcHMomb5aqzcfpW+4aiwEsdXmxgGJmcm46zKoMmd4sau64ObYZ13yzzuirgTRXHTPe
Fl1FoPwsS0gdJv2MmCW6FKqtga/tsFGYt2mmbZEt/0ZttvDdiLykkLTPS07SzqZVnlqc6BhgwIw3
qp7tOT7TiaVZCuSZTt7OuGuyxtiZdl4WXVqtvegUcgUNSbET1chwNCDKiHGQQV+zr76SbWWr9Zyt
LJ1llpuCFpMstfr5Mf7koJxLWal6sZwlPlKTc2SScL0YiN+clNd4Gu3LM9bI0cJANTRJ4ubevyK1
M/rvJ/PaDZ26ztz4aKA756Ffbn1FWTqxkDAhwz+drO5bsyxNwonYH4VrbclvkZjFJOU1/wOTw9/t
iDRdJpQVxKMZ+kuW15Qsj00DezGt6dQ7bb1f8KV5kyHJ/JIVg+JheEZrtFHek91jdHj/jKHnbOB/
qGhi2cfHtJQTPsH00RXT+670GV1UxVR8yJ2Pj3NPrjMoyjkILaoPi2y7uJ9UH4TvFJAm/vtu6wAO
6YKDQF7YtoXAaqTZ9dBWPRkJ5avblqqUm7xY759EKH9E0qTU3K/TAwU9J3t1qMzD92/JkD7+m8Jg
N8UlcWbQUBDPdxDF+hkHiMCSzZT3lDdtNogTQEqvH79F4NajdXQAmawMvvN7dATBc/71yZAatU2W
3ATJOZroVlXOkaQog54kU0K0WZDizGjZMSLEMutlkZkkD0jdyKEjvzR5HbesYsHlQpkKhcuye/86
dY/MDh3ZQkorRoGYk5tGNw0hh4HMRbD0IlKnHHUKYwTDjdBmbFKnf/eVMLauWasr9WRL+Fk6n7Pz
+hwx/9B1g4g1yNlabrAB763sP7aDeG518rf0xJuO56vffMV/xG3SfdNDrSlr9xeK9YAMhUROr/jc
yh+ayd7Cb6cG/Qj9LhEFz8XupKH1Mh0PLxClPQaTpqk0wjmhrHQtqmvK02qBEmKQdmHOQ0vyZe6A
AXonJFbooimDuUG6/0sCsf7m+BwcukxsMnDyeWciyS3YyjFIVccEzpvZRDBb+4Ez71zocOyXV6jj
RGhsG782dxf5dr4FzJAiBxFbqmcEIUX8bUqr/ySPsUmWpsziO1QfOlqfJRP+D/l3Xg1GDhKpmpXh
ojGdML5s8jG5TeudRYSiKu/b3YpUPPuRXVaEMhcWH7ngW+fmIq7OH4Tk4SweiYoR9Wdpu18fFyOP
2pHR8e8kc8e2OuhRFIHrdaybcyF3HQvrs1ZncpR5z0sur4/+z/XV2K8/xZyTgcyIB7shw6P+MAYF
Ai87kvWAy6qmfGEmPam/2Skd9sRyEh2KPZGPwRghhJ8+v07JaHkE2kq44fi/LN2FuT59UdL0qXDN
BlK0v/vwe2QmmHYZYBBrucmsfwUhY+3IBl1k8aP2R+WR80hHI7/42SHCdpDu/HGbUCwFpz+csdO5
lemXT+cbN6WczmXtyjNQuK8CfCKx+HdJKbqUuz9dA1Rigyz9rchK/tCa3b/QoDQnlKRoKDqqW0xF
yRiJ4tmqLZKx+HqtR+MV3/3NgaOK234JWFMQk+x11lOBAwhHl4n7OWiImbfugsZqrYnsPT6MO6gN
D/3hFA6NGMgwtpc+4q/O8579udFlba0b4I+04oJJGeVmNaDOP+Eqx6hLZKUkD7XUMx8oN/0CAnhZ
sRl8FLWZX0EpQne4hGOMC7IuaMMynmyNRzIFz2RM9unqp4nvHg8NPvg/F9n4EAqkR8gp1Lkr8Ntj
4O17wCLVoOqtgczi9W0obaE+zAsWIYCOFT9yIZbnyfvfRFzJ4oBOiTKyFCOJtOHcsIkcZqeNOJuA
cI51XGTbF+d0IfjcDY4nlS5yebIJG+Az/Axnj/um4KCGLHiORtJKCBqJbHx+udZUcSej45xTcnXb
VuUJOaXaLTtYKT4ocNqhBob1iZzjj73VZSDh9F4V5Dxm2uW+BSjfvYf2VRVaI2LW9JFm6RPHo+9m
1Cjcp71fIee+TK6cnEJ31Ff5Vs8m4w+ur8HhvNK0BcJZY11qPODTsouZxrM2WY6X80kTk8Yynuxw
FM7N7FBGbPN3zU+pOOHLbvBukxrRZ99gqRzbJPDeDCf/1xT0AeXy4GogoAhe3ndetZS7BfakFgDv
hvhVL7NtJEZjp0CAOpackXAzAF5CtRxo570W2ZX2W5J61LnX46hDFH0hivj6diFRalte316xPsgq
VCGPbLsB3I6ezON6/Eq5oyQ5Aq30uR5JZ7BLVRkF9KDdKmwE/vzitK9cNw1bSi8puDGIBNWhGDe8
G/2OCvuK8/jM35ka+S4mvmzmJZnqNvTUJrcaMK44Kp96UvQnydKqMenH4nmnJpFyVHyNADslD5mK
wKsBlpb55wfZ4lI5Bn9ct4VcGItvtwnY8HVqlykCwZqPCDQq9Dh1Z6BX8WN+iEW07HJVeucdIGra
BV0v4ljEZ5urg8XDGquVuEWR336ycUHm5xleW0Q+B/HHIY+VTdk3jdgxSZwn9yMPmEDdLX13i4xF
/ITEgTq6Z3Ui25VOOVzxJjZ4w6OX5yPhZoMyhKUCLG+0RfR8NOLkx4FwXdS2TjRc8OPoKU7yOkNK
EpTvH5tESKxDHWdEwpDwM7lpiKzK96l2lQlGawGKTpFrYZvZEZPDPdZmPj79mSokq+3b8RFOOKZk
xHMUNMaQIpWt/5PYgpplLpZ4fJpbnN0Tw7agfzaDz3ZawesuEUTIuiU0sIRhmuMvSaf1OKqf2JQw
U3makgORWAXSuKjtQs8WLn+DxSJSpIQ3ICJQ+ndtMqanzh43hz0OWNCSRkA07vVktDC3Z57q7UmO
QmjscTSBdCdmBs2ujiJyez7xx/JCPu25DRGQYdrw4bNwCIb0YpylmE6tzls/WcK7emoqTPaA2asP
KRMFmNy4AAXDUrf77I27awRdP1R4SLzRK01RyOrYy1SnefffG58KfjVuUe2XtJY6JSxh7pkUuZOA
Dz/LzPI2weGfHoUhQ4UzA0kl8eH14iwAUbyaS3i83dmYNXTJk7kGxMqyrUCgeY6KDqzt/6O61rwI
SqVFn4R6xbIlealpfw5vO+2l9x/xoMHhw/OkCS3k5/JQ2BMNsjA1leqeRZUyqoSO+5W/wpjcVKMb
nY2SteNS70xi7vhNVshmKIU+cJHOM6R+4etmfKc/2P+Gzjq4ukeqhT6uQ6EPxoyt50dbVQg9RcDV
vTsvj27NjkajSi6Fnrc7WYqG/ad5J8eFjwb+PvTVc6Vvqn4dASby/5rcs5mx5N6r6yNb2MNOKQVk
8h35WAvnyZDTLYIASNsYL7Wx0+4Re7TwuT9km7v3tMwl8amzqjTmrb1ghF5NtLsUuwHNTdgpESqy
EpRpvpKjkT/Q8jSkmkcE1hgUFkWU2lSgWIlZlzMb7oZMUFmdjc4CrWHeEvJ94oSBPQOXM9QO50jF
kLZFeGrskvqCwGTXEgHofueeQ2ER5P5u0sm+hKMgA7v8IBeqovjcVQS/VeH4ZbEcLYcbnQLuFFnP
g+qLpzoAa3ieCB7Ii7fxvkZxnpFlKANUA9HoUWLKeYY3jkqetga7t+ZevuBYH8EppiPYkrmpu/PD
O00BYEdiXJNS61/h8H3f/ZCHpXamE1sjAPIOzGTicigs3vzAw/iol9AA0TLiMMHNRm2YMzSeDFYf
km7ZlvnIGmbIwAQlgKbhEJK1XEESCqaRZLTufE0YqBHuS1XSDVElltyohDk2PHC4bnXJAO+2D2xi
P2UImyhwkVjAlZJGTWx6ZN/bMK7jx5CA1f/yGb6Aq2a4acBfP3VHV3j4rcGlyT7iJz60vbRO5EEo
jLyYB/N60nSWo57/emNCAzCczYgY/2g8n6lW8JDjtzZPoYpDAZSsprlWvI7tsCjLKyyGhytGenjM
U/Hw7bf51X/y6htj0dUxJ27Lq+s/vN1pLvtIAln0OXZOyBrdNFu6mE7p8y1lVKs1Udya9Jg72mSy
yI2PLio8wGJ+MdAAQv+sK+qm+45z4OTIE+hDAHj5kxRDKqfpSpJhfpjYE5Oz+6r4TnOPqgVa3KK9
tg6w8Dc+zzvz6cAqeD7fd0au+g+OwSPnC3cRd64P1V0iPioYPC+S3tr7vXZSeUU0r9fDHNaFMBgV
DZEgj78iWKn3yviP6PPCCHppjd2jtqiGrheg6bKnL5hRt996mACDwVg6PRVZFxLNU/NGFZbUB9RL
UZ6baNEoguwhrhdJjdGLeALh1qCSWXUUQOObjhlMQOkDoNpLqZR3L0FnXpG1VfqIkFCUgH86mSPc
pN1Y2tn4vo9FkHS33572bHbSxSHbio8vNeE7U+RM6a2JGiH5dodGIbrTC6nSv1I5EeKZCqSq51ky
FJlL/ly+5bS+VK5VUvhdHH0s3dl55gqBnOTDslRKbHzZdl1mOcyEin3yma7upO3ujx/RM2TtM56E
Xldp16jL0J0ImQ8EDD6xIGggSMdsuIMtL75NtMGu6+EfgiMesalsHfL7XlVArUF6zSLdK+07Sn/M
IjlJYHtkNuacWwjpR6XYxi71rM0oheP+Ytd0/6LI2W1tX9txP8/KgsXzIMxHdkP83ADSKfnvcOen
xfhxfoCY/ljDKj/DjonPSd9QgeZUHsztZH6IEVIKhC3vU9+33UR2zNC8qN6gxTQFm2c+Arnvt99P
uqbIKBVR9yRFKJbjrH/702Lfqjqv4nhJbR5Grjahe8TiwBcYft+bqvpBmH/O+/LsAwTuIQWXgFLu
OVHKrjDYA42L7e6uBAkETWHMfaHwbBYe/PzImrhAYB/qqOFhOYepa+9+2sSkqWGw6a3FIt9pVLik
R/80pMV64Yh6L+w4rjONrISd2UsoF5n+ZVzOKcH3blkRq1oV17BMTRNcFgQHB1GoHOEOe93Eyh/e
ZIq8BlNlEoVWoMCCZHRKW9f2RZ4YHspFTT4C+uUTrhqM2HelbUPpffYpavmCABxAPGiB12iDTM5T
WMTJdNPvJu2kGIkbRsVKmSt+e1gv4w6GW0OF+HMWmmeDzpP2C8KFsAxUpJiAW3zMk6IA6aNmuOeQ
ZcNryZ9PdF8zeSGFvicoZtUezduPAtRk97vRxsUKGSCqLgvd/CHejhNllEjIRxeGSZVecJTBvodl
l15xxNOUQlyzQVQoelkFZRYTD2MduYo0q0aSetw3KfWyH/FcVBkY2Dv6AhI6y9dpStN2IvY2Snvi
fDrX+cPDEQsfHAhlpwoQQ+jBVmVJy1BNuZZ29JE9jOdiPRwM1PVX+AmsJ0CVEwCm0+S7E+abeduZ
TqwFnrgRG9JldxqO2i0RfpK0EY2qZqcEfaPcSbD8D0glX5GkJrdunWTldAZRmrb9tw99Ti8rnAxv
Iob/cfcWmAicxBqWm4lAI3WwB/YhvcPlcdquE+7Z3Vqg+s/ROJfEFD9hzn6c4GuKOdNmiKAJL2X8
WHACbcfxUGSCwll8HFetKmg7jKkUNePYegSCkBoudZDR1iZ2EeQK4Qpgad/X137rWiCkwAjjXaAR
/vhm93QIKHNNd5tfZFRrQPIhqGW4h4BBYJyjerGNrAM8BPUS4VHQklr9cNvfMVGgdtby64rBZXNI
eGylDl1npGZ2Q1TKydkA/w71KchGLq8EdxB9VATxtMsg2chWlh2jnPjZcv+115ftj7KXCHkd/l9U
OvEvjd0oBRaSz3pztnGjKFjEtluwdFNONvvMD/L9kozL8shQ2POYnV+Fm2hAsZESiPcf0NzLrlIc
zYDTWU3iExWomUNY+mEUYERGtKImjZju0PgDwWT96N2rf6r2BFp/R+9hWzQ9T1c5eWDk1ehZZhgJ
ZxuLlIP5rppK7syzrLuZUaErOtpnqaSC+b5xkphaoD8FZcE418uVjYOZE8YDgCs4SsjVugR96sVw
DDshIkEVlqWbLER3rztTWSBZGtNVlRG9zreLaYYQo2kh76AJ48I+0Eabjf7GgNrFShxgF6ncgsuR
BhE/SvxmJGPAIapc9ge40dPtmnT+Ji3Wb8OP86HKTbqU5Uc8Jc67aeVoIYKkdp/8hOJ4h/KTdeCs
yxFm3xYad1bJaUVcEpYsUxfe/uz7BAl+IJIKoa9HOKoI0FJl0FSf/YwhZCMcAWdZ9n0uvGlBmYPs
12g29EEZG/R+fKW835tEocRcG7l2ybztwtJKjDOuR/6et9rFIVrGKvJ3yziQf5Q6GcPZ2vwjQuBR
cyn+mrk4bzAKCnL66MU4+Pf/1M9sEBsY/tnvZbRlanS8j38zmjJzSO7Jd0A6CHARnZYXrQ16l/s0
dlYGIlrV5trP9XJJKOOhjy0VwDhZAjgpWtSaiO5rYZycci++TitynIvrSd5S7H/Bu7LNrMFgPIQE
obMsvcpJUjCNCsvbUG1qTbAEUpKlvf/6ym981gXgls0lDYyBVtDbvPnlEcDvhHFnWHWzOJ8nrbyO
IFXpK9IUXYiGUD2Bds13H6KdrOHPlA8Qju+xyB+B20z1hkbqmS9ySa6Isw2UZEKRgrNLjF+R0tww
nZ8wt/QH8nExMwj2xplVcCGVb838MFGZdMgMB7mWqHPuRcWQTn3ySlbxKxSKO3XIUC+4Bx7NRlIr
JsSRHigGIQRYMmEQpacXzS69X0HQAkH6FXIcBVGF0fGR0yXoSx4T+6TRuzLD7wKi7H8xA32a7K+3
GePV3cf83vXPyXDJKbMfBaFrDUOjzZQDG2O1kAhdEQc9i8cIpDWcjhBQ2qNEC++UYQu6UZXb/EXE
Nw4xlDdBpc19WB8RGkPTSDne9DqJBTA3ZBkB29FtJwmb0Un/WEGCi8U5Bc2UQ0soFncKN5vpbIaS
KTu1duLGqOxk23FRvJ/SjzPPhjQatIGpv/MDtPxB49kj7/XNuu+veaISDV/dvkMzYZY/UwEceWBI
7kU9WeDpOJOmIvcY1Fva7/w0ReZ06F+zjzmPcYWgme9nzTL/4nOmIEWdynTitppGMl9FmYnFW+bi
VI3bzJw2T3LIaeIHEcUZdTEQjFE1oeAe7vACHj4eu259jXuYAkqzU4GJ3kYgkzI4GLha+JRkphBH
NpSWTX28O2BLS4FJ1kIjp3fLCtkynKAupcV8OAXwfv9xMGpT9mOtIzcFAXFn+/miZ5Gl4er+vJDt
Tm3eJxv9dSfZRTxMN/7/nY2PhT9DkoAPDZ7yIeYoEOrZaH4rLpss4K4xkWR5mnQw/tLTYlkfcI66
yQP4kMnqdsrOWOvqngCKa22dY14a50WZcwOb3+/3nHARpddyNGyl5IBIMVqS0aRIwYvWBCzCMa5n
Bs+f6Iz0+fbo2TBS9oeCAPNsDauPQWEMCRing8V2e29zabk0rDJSbFPqnsGrFrQh+s6yyAIyYwjf
gAbMUWvzeylfWeN8w0qqHtxfgIbV8J65h/LfOTG1F+V5Ir9gWJBaJKqH+wLKBd76bsgJOYpmaDbE
PE0YEYKLuoD7wlt30TSCHg9q8tueEspnSesYxWRmbjWbQzeHNvToTkN6ERYfsToLDhTYzvFRPwES
gj6X7ufV6BNShi82nl4pMaZfRmLE+VBhjzTkiyGEaKY+30mRtNN9Rov3DBzNs/eKm7kVXZfw6zCT
dfrjNH2mc81wXviqiBufvlsGX9DNOJRdYlqERyY+ZKKXEjRK/kNs9MFi1iB8SJltTf7nIrGMIlwN
sBMei8dK10fpwt9VORtsqWITZ3ZnbOH2skj0VCcSeDhdxj8t+2XsaMMnpwtYXUrPacjxU4SAiA7g
p/Pz1gCA/4dLYDlqJ4NsfVhRh/oX5w0ZXWwdMiCOp/OPNpF1rdxl5XHPm045qmyzB8hJJ6mboNE9
FcbH+gIfTnZJ2nI4GtT8vMIKancRjiYctM0juSTkmnxbgZagYY5ji5ovYHD/7wHLn6144mebutn0
8tgZkbDRqNbz1wfyIDO918CK5F9tp5mEqBYBodG7umuTRWVYElL17lJpkIIrpNpHUiD5uBtshxxx
mW+FCWmVix9OuujKbzE8ln1o7AtUwVWkoDRFFWoDnPza4MiyegaiRUVYRjbJsvXhsHT9Oypu82XT
tl8GnOVP/WDxxry4rAV0X3iOoaUsL/sX7xvTwFBWOBl6ZtLEY4jn1A/zsb16i18aGYvsL5sJJXcE
1DA2l5ObOBc1TtXN60n3cbSiVSXZcj3MdlhdcXXdEyMv6e52pXRwXwXE1xkK1hSAmwq0rjSu6HS/
pf6GwGjvA5crmSB8/+gqAYGYsvFchBAqIV6kyUvVaKgnxjBpSYk2NOpxZuZw8JU4Xlo2Y+whiFMF
3dM6nO9r83KHOaEiCD/93Azb0EX3fs//oGHz1Aqqc5/SnhrHGUVdHz2qEadSAnre4KHZlVbWsHLv
9jlNDbiBaeUixEAp6q9nI7IWacQhuAmK/EYwPzWGPDGK0DPfxFEHZo7xG6uEY8gtAeUGnJUBNptN
NuKJH0nedH6jWUhxFLRC3av3HhSm4fkyDTJWE+hV2i/nlmVnrEN0I50WVkwrh8Ep6fm1qeFLURKb
eRjk/3ZqcDadHwZJ8AydMi2zSjEny/ZOS7YPP8r7ht+pheoPTg4q4Tbeq9aF61BCAquYXWaTAi4k
6gZyWcUBakMRNJJFjFzI6ENQiMnDsj9T76+FFT+ETCEysCHCFUCH55yU4N/gntTu0ADC2AeH+1T1
mdz9qrByUrDMXzAIEd8oO7rgW6LUGG7Bl+xf4UQkKHvvoMoJ8zn6rajZS0gA0MYfouIzYJlUj0CM
OIfdwQCHr6VQpI8Njuq31fzRJycJq+RXlW1FxYY2XF6Ye4uF/tT1wM5AFo2+4Bx3+xEfK6mD3b9t
b5+/NVjDXN5Lm/UL/MtnhUlf97mWJQnIYIN6chLPm2fZZB8Q4vemj1nmYG43G1JP0Io+yxa2M1SX
62PMzwOPChN12Vf38Y4qVN/d/ymEhf/ZMpMXny6XD+SZHY5hGzr7PHFVmaJW+kSRxTcLr5DkAj6f
LGxxLdEktVI73rHMIZklvf+1Jst54WgK8PoiOATzta8plNlv+5Zt7KD9p5sLrLmbHboLKNYbbke2
qSqyx0C9QmA74fSgyX/1J4gLpKGW/dMBCJ0RyUt5dz4mjcpGS+6dCsnQ8JohLtF+brOzKTkbOlM9
9Sb/tShoj9Y0Vv/g+anSznpdIXSTnd5wP04KNO9WTr2DozDZ0Xu6lfU03Hy02Q9xczrj+WX3qyye
Bw0N3FjtBH+S4ptUrU3EcUtGypWNngyb3eVMzAanl/VgdnGReUTSpm1Y9JUN0JJwvEd7vSD2Axxl
Dt2fl14R2C3KcHclBJE0In4gdMBx+sPzoqzXCUGWC9V15/1AhEaLBTfMyWdf7gKKaDR2Tyk6iofY
6h5hUn8l6TF0c5LTF9REqZMUUOVmoxc6TA3RiR+0yNHbhpHIL0/V3P2CBcifrQ5fC0rlkiDtcDXV
mGH6ZcpUofLjoUfBQ+ErK1hM02NLZIN6ZLxLPE/rXX0/iu0pe8T2qzSqZXGtSx2Se8PaIRBZsPbm
sY43gWlj27xDigaL8W/DDhV6MuhoMssVIygs7I24h6yf082kVMEWnzfKKlIxkVu268cOrBHJb0P7
BC8AUgZOu0qgFYf/reDCholELbJsoan+SuGIsJ2nKzE/JlOL0teofLQYmOiER4OVIViu0LtiL7N1
9kDZosz9dMFfbmCept27Tm+/H2v4jPjkgnhBvCUE1jESexlX2mTwx9AmoIdB1fJDR1YDA+Cdw6Kl
Q05c/Ltbgn+gb+iKhTPQicjsKyvltW3ioC6suFMS1hftd3tEc/kggwAOlzrGJ0hkg/DssfjQ/AOE
WIKTtIj0cg9JoTTckp8tXViNRLUqxzcFL7frNAnYnmwNxWmHgieuCB4PFPcVajZ9NAD2VJ8b8rhf
8B1fz15TF6NB9iCRCrlDowQnt73SwsZSeVH5cG7l6UwpzFVxMLnpvJX4xJQzo+M9PfFM1kLh03rd
SXMIOUjaWgIJV56i+56H6LSekuD3Vb4OtXOKXTpCmVMlUpqUeGMBh2DhbmulCwJfzi2aDkJdEQZr
QWxnYQG9ItMrcmc6Nhjj2h74fGNU91DsFCtLHka9xlXMN9RvqkwR/DpxPKjnrQTYrx8/qkIdhK1D
3yyGx58GTIisAyKccbh4vx4f+Bu6OsvMYyREIYPQ+4iwpseeRfHBcZBHr8Yl74SYD0h0AIXLHdCl
P7EdvMxyDaMTvBtDUV+CPOEACmby5b4OkUZn8Jm8NYlXD7Vn0Bh1LrEHkC3wPIX0uOrhhRdBWL5h
HchYy/J6SapwOiI81fuE5Lzl+rlfuoyPSK5S5fu31ZHKlL1tTOrZgeOtQyjE0Plod/X1sdjGfrnb
5w7aMRxc032AKwGext0aBJDsOD08F2KQnga776iCbCrsqfX8VcILJyQdOoPLviE7D68lLxc7zlOh
ZGPPFMrW3talU6FlMAtGMPgyuiW39S/UEjD9c9xLPMsvoNLtIUUQXr3gev3xGn8P1lSPV8QwixsW
v4hMDyRcVbR02maAqny0AJKn2QgBaN8g7pIlJkVNRofRGwwM+Dpa8nrKqZ5IRyte9FSLzl/moJKp
XIlw1eDBEOGuZNn6natdc7dl3DjaOId2VvPVPYqK9j8gdoAJZWMeLHSxfcLcUPuQL7fVYehlFW2Y
yDpR3wEHoFYnMdKbybOvi7ReuimdsQF4DiI5ZFR7XEjz7SAnKfPaWkn5niPLJh6I64X2spd26n5m
dfNDz28swgJeAHAAQaMxDj8vJao4KIu1P8e5H0va9ZgqCPQmG0zTvSaRwDSZO+vJg+7HYRD02O5V
HESuW3VpTbMJ7Sf6Qa91+3PjXUTyWz1CXyvjejh9IH5H8ZsdhqVyYbRatKE6igmflz+LHKh00Z/6
VFsfmUCREtI02UMPRI/os3rzvSTu/aUzUJvJ/heWSWe5xgVnRsT2Fli5MIomP5LbUavnhMRfKtOS
V5iGZVs4Xxtb12YBQpT3UgC+QguW21s+twYpswHAIvbcjCcNC907CjXJHihDN9OToy+oFRq8pXt8
N9iLzYYaD5sgrOhQlJ7M2YFeX5mzsFNgoiWarjhSpAD7cSxKGsPw2XYJufnQolPj3LxvbZM7v1O0
BZ4WclQ3unRarMuGAoGqScGFS7+nhOLyEzdp9ZfK+oX65e0Glg6OXp9ThdkNV6M39JYQvov54dt7
k9iUd3Fflk9Lq8EHDTZ6afJy8HnU0KxY2l3uAsrC4Myng8h3tAX6pIxDlgCee5F9Mg5rkCvBdOc9
+nP2hyatvwwJNcbtl1WVMpYXZIlFGoBrNwu/gbUeFj/dsUc4EJ6XOpJL5246kdAn6a5DKbQx9FAA
9kexfF0PLLo1uREIds4TXEPFF7NcG0Z/bnErsuLvraN4SvgKxXKggseK2RkkyACjcEPA4VKqydzK
UJlvqHCaldPBrLV6Wxlfd8CBg7TYg86HlYTX3J2OLK4M8VhFkxMrA+6j2+/o3VBig6A9WVZXjX5G
KfMisMYQCjhDg5iZZLVA7hFcT9VZZGZk2RHU29C6cF4kwvyG1MFKe5ij1hlnko6qFEYj8YsIWu/D
o5Ple4iMYFI4HFUwXVHlyJjq8lKkHFaD0OgzzOs3hEcFPV8cBqfxGs9wm2OvyMhPQ5/3JWm7q2S5
oPYbHe2hHrMb3RUVBnn0U8q2f272h+EPbinlXqSeM2IPjyAEWNsP3OGwLeuLM55sBuVDnHsXW3AP
gzYWvKszsjM36xFZORXLhFA7mLkMSeeJRNLQ9PPLSqRgSMRj6kiSRfxR7aqovOnO0icS+FqL8Gv0
9MeCHZEMETO8u+5x/HtonC9MM7O9PakAlNYw+zcU3JxBxGglbiTVTEwonH1zc7EAyzThWVqav8U3
SMb2YHKGUfA6qWUFJVPbZiW8kVy0lfFppgWPU3wsOz/Gy+NtKe2JegabztJXkxHr0oRJzi5ZxD+4
T5yzkQUW8v498Kfq/B/I4MXL0ifhmuFlkO1/Y6u1yrruurhX/PEssXdS0hEB918dCOWaixQ/25JH
Wn7JofrDHW4mRV44xMjKMXWqUbjkfYkrTU2ruOQPka56B6LZIfqamaRkpD9bBQmCzmV0DweBwgP+
02qM1V6487W5l7gcmeCMosS6Uc8lJzXy09MeH7Lo8IOqlJeI9ai0+Eic/7/RmKqi8+B4vbEmko/k
SS59TynGFDHajQ+Bhjp9Amn/lkKhb64qPpxeYPzTbLUU0yHxkedo1XMK2nXRquaS1/wspcGwb0tp
Z32ZajuDzwRl1TMSmkC0hBtnkZm/OTMKHAkawRwl7aF4Zx67dv+D6y0Id70//bSnOsCT5fw+U8P9
85s9waYxSnJFm42+KZdUd2sj+4it7XOKaohbE+KgaGvR3evXF5L3FkCF8r4spf3343wGwfogLm77
cH5L5gVktlx4ehSNckytXgBX6JlRF9oycQpAE09RvqIZXU/zXSN0XGoLmVi6w8KNl9Y96NUHb3z7
Wud8tJj4Tgx//6U7w4GNlVWp9AYoQm9xaZW8rrHK2/AJVj9ydpH9dikLhxwy9albgQpboXI9M/We
IcaM2YyeGg7gpz798DYMOgxPSQ/oQWolEU0Z6ZokqVYuHl9RNf+5FiUyxTWdSvPHW61vQ+eI7+p/
wmFF3vpbB967SJIfOJQQNPnOkg9b4x6VM1CxPkYWGFQOddALqzQH3xRrILIkupQ51rLUiM6TK/Fn
DBe/6+r4H59fEPuUxW0qhS82zrynw0IiA+4ag3BaYHqYuubzJL21OUnURjfTrKmGzQJheBvilMVu
M2uwMpudJ5x8lN5ehjzDOei1jAsmK9ITU4jOe3p2BAEO+f2A50hybzgb34seiBkAqXytNNSW3X1i
8ZwedHycJUdx7LddkmtY09y1vIgjIEGtrTvN8AvvdJs7H07B93FKrckmftYotiUzXNYSuGvGcEAH
Zydsz+15ei50SvgMVxaN+BA2h/2SfO1qrfmfaU8tgsA2LT36yc2xJ5rQDcAyGXLi91R2K5Hy/ROH
IpR7SJ9Z7ZfEz8qUmfnIj7hf4fwcx5ggsXmDTI8geeMa/2HgZiffJwO2kEnjfBGD0zycsb8ma0xo
wFor0+KEIwYZkK3rq7TzEpfdt8JAVR9H3ixRMKJ3Zv/wpXIpewQ/TU86HgJxwp9gvX7w4zDrKNYx
upDVocuniPi8KXneJO0rm5IO06roimPgHhTRzCmJZAdrscVJmpMiz2NYWdK5xUAHImTi28D+ax50
j4RSU3M2cowLFhhIxPWLrftbrJjormbliLo9r+l9bwlMVkKQjx/ORrW2nWWOl2iK2D1dT/J9tF8q
XvZCfqYKjI4qYW0LIt+kT8c6gfdm4Br0J1Ed8QD5gjj+Ia4gEpEYyweq2fmyQtq9mGMEUPjO8HKR
1+jzEtNx3g7oFEVqibKSfIMJRK+E6QSLY+Oy3COc/6orNk5gDWwxXMcKmIou0JVUC6q/PRbgu6ir
CtMc8JQskkYzRIh8vav6yCHoqUhVajlEAeoq9G2VA50O0V7KJeI5S0gkwWkEym3CoqT7XDDjzihH
S60aYdLt+4AuNRoRJ58v01uuX7h4l+cmZ4op+fy7wRfPCoFSzyBkICBhW/pXA1DncGv6/RsNutaw
FJDiGw5RQvb7MPkLk2VHviLG3rP5qR+A741/mJ68KzLTFx9ccilEGIRkBEM77BXOPE5OvbOrRgF8
9ZM5h7x4zuQMcci4mA5UzL+nvkYq944JGHhyiHWCW0xL1JldSg1chAAUX2CR7abFzV+hGg7fsihs
cpcfelDWNQwmCI1BpIyJw2/NodBvgAeGa3EQ383SYWm8QiFkHU1h8G2ZlLss+eHnkEpm1nqdvxo2
lyj+TCESwCy27nW0pII6O79YYj2r1m9VXwXgkMGyiu4hmAk9qS3/cTZEf19ePxWn/0yk1tCpHnSm
Nv6qB9jeOvsnuWykXFrrhDI07zUTAwKBWLZEWPG7uqGpWzrnIYKTz2agevDnApcK8WqLYh4Glqan
g13dHo4sXunXLLzAP0PFWe1LqHv5GgDxSDmzRQa7LdXLy92l6RA4zoT4SbO0toU2tQvdT8A3hWfZ
vef/rzKaqJ9+PA37MEHcmgGyhiRs6Xgh3gUcQYWQAjksB4z9zd27677U5lRBwMecSX0KBvpj+Nxj
1OivfAwGO+2JWXDqW8Ixvyltj5kml17RwaGqx7nplCc8fCXBSLgxumO1tArEmRdNuz+7MwzrQ5rc
jd8GXeOAecALmo6IbNe+slbjIjutURCjbS3dLdfisY+COUjomP1G1/c/67qpNzIwvymyfj1WyZm3
kio1whsl5ISRQ0o2lhzklm0Xxpt2QBf9lwhwurbnAIYOuPzP6Xp7uRB3rw4EOeCIjSVztPKsmM6t
gRG7G6CUiSeMgtgzFSNc/eaErBJimmxsGFN6D0/Fz2RUZ0Xtc4vvYzwbPt8yLo3rnVZJZ1n+I/hz
0bthSqhT8EPJCD/0eeTi8FBZBIwqzfnPLn8FUMiSutygPK4PUFuN/0R+Wh1AL2sSGvkTxh1qLlCv
CELpeK7fe7tXfn0yk6WExuJmURoL2JnzC+I8qXpuUqGGGFNQ+mpnjoZtBu0TX9ohBZRKb8UmQgPS
6+zdGK4Z/pGvtkh6SNWASZu13UOzKermq/DRxdm3hwM5usF29rYV/1Qj0Sf35tfYGO5gdXkxP+uA
2ciLwpziAQe9Ft0YohIGgY3lFfLdfCrqXfpG+cNQCZf+m8mbweLFyu9ecFgrjNNUOJ5TzhayV65t
UpuE6jP1Ib+QvcO5d75Vv2U06fA8hnh95MOE1NkZZpQKKFlhhsJ1vp6w5zkXX5BUpHcc+r71t2ZY
C2+/ZCjo/5DifJEuG0E42W6//sy1oeF/8vmZ9rsWZdOuLy2eo8uPQSNTN03tB3hJhaJL+HVBfUff
UMxShfF640HP04j2V//9+OD/OvP0awPwDH5U+WIRRW1CuYV3JAf7zAa+aSrtf52aDhAaFU7TNlKd
4lAu+hCXcTONdvXLi+rG1rWtGKpw617puuaWR8BgpkIUCfL18wotzxYqfVW2XcFQ2bdrcIrzhHLr
BE58XDHUXkO0IHAroDejyyZid0F+3R3C59NfzEilMMw2sovuQ92/dLW2HEuxzikK6drjohRbAx5a
8waZ5LIQrpu9aWe/Uebqo/Zu9Cj0JvJnwFiR4b4zfp0sSTkHcBZVuX2JUd/U6VIkj78zikCHpi1K
/GYZS259OFV7CR+86JuYdCJR7i0x5Rm3//dUXluEDDE+15X1nOngdbo8BPeVgSCy7ELFC1G7GO2T
Syl/x0Ubzq2n1Dpj3u82W8gkxk3Ydg44301YFpCm0hKyb8ePEiMElmHWMZ9DtTrcdhzlLLBcydvp
hx7Mkc+poAt6So5qztqZgdkXwnWl7J74uHMa+JaSBm2+OiNEfS6dnUl3Z412jw+QPTVKgiHhun8f
Jn8tOQHoPEoIkTcUCtn27AQbfhQVCHTVbfSlEnOC4dcJrxl3FGeyo+9h5BxiiFbKqA0JoD3udQkn
nb9ySDgkuNRYB1BNiDRZ6jkjAbSabHNei71xdmr169alMzbiIuKw5VUYTNqy5SP4PJwtRW4tCyA+
W8L8+3+XKMzVz+V0LKZzIOYtMvnGu5YanBSVG1C0i8ICUmLgX2nCoFbevkv8DDAdwR82CjTd7HhZ
0D8z/3t8by6O4iOs3ZtPtY8Iw9Mg5uT0PgNhOGTa+tlQsZxyWn+TrF0yaJByWzhlpaTPX0K00C4W
fSixPFJP18a9kFonSxIt2Eb5YZTspESkR0rszCrk39EtbGayTrUEEkSqn5yDbwKXGu2ILZW4sl1o
a1PflqsHet3H/+HEzTHtLLEIrRX0RlNaOZGrYNp86xmlxdi0SuGN6QtrBWS18trFBXfj4Tk+hiZE
joUqZao+5gVkm8pida4Ua9Ms3oEofqNVwq6TCh85EoLXRjNXxZouPVRVz7JgUWwp+0daIPj1zMKi
BZAtGAEDyhc6xJz98VWt8gB4fqMDop+DX5j6aPggKsDDyo2Pw2opWPpyqQtRxvexUVMQOg43xacj
/WRjj1JU9TBZ4bFx4+5XKPaRo6uLuzOtNPOEyoDxBlhNYMSpl1fEb2zFipXr17H5IKGL5F4bZvww
RasA92J4wujGclfcQYTMZ4ts/Da7t54+QrscUrGYoyt5iXIMATcogffCMQKvVOw1YIubI7YVMvqx
w0cS8iY387yHftg9dWQK8mDdPQaYXx2sLVEozPQAhZMWLCybTyKuyoCvtwBd+xr6qHJOoCpsVQLf
AIAybKdTLEVu+dFVdGH1Hco+uUn7FJl1R2+aW3wde/+StSXvVmVDs/pgooD1nNvcVkCwqZtvvCfl
wERLfNNnWadrmvMSMoJDNVT6a0zqfkFCLWG7ElvK62GMtZUx+KAKANad9vgEk61iUx0uP1FzJH8z
vYCoTfGuyK8DFXMxbx3QCNoTBaO1R1oiGHXtmAxmdBqi5XzkS/V5DR2XwVmcTPRLDjyWUlmTLZxj
FTORDVypg4ctpQaWkrZEufJ1cHqV5y1ngF3l0MTRZdFXfievGS3VrC/ZMty9zHP29Fnpsys3mR1t
+VUPZqbSXaC1IPNvp3Qdk6LJB+6YWGsdbtBnjGVNonF+e5BecYetajBPWbHJzoJyRuAy8zo0zcbx
YZqWir2Cn0M37IwglW4Pbfw15qVZ8rEfPWIUOA2DXZBTvIz21zI8Hbn7SK2HN4IaaCyVMRzopGln
P8wwxCjXllpDoV2kQ5xWZFVsYQ9qAbK0VDoAPebkWM9XlsTnzzvP+75M216VUkUW79+Hp6vCN5Gg
OOd6Jhi0fiSCtn1TIcaTL/wcHCarpZwfPjMPvDT3oaWve2A282lSObNO0PfkbqfV1nojRjs5GIWE
owY9GusA7qi1t8ffH1q0+xTsHumYT5u6peLoNdXgOjfP74neLKT+VXhnGfgaCGHqXjkuA2XaqISk
jBt41JL+9SrryjaMdtFRx4qPedvyLeWYNjjzdqVZRcTTa3ToCnVxZ5NilYQJEx5MeGl8vTOjwr4V
Kkbw6h1ycqAv5pda9KgGKYoj2MUdS3+YF+1rzHZK4o41dHg3c7UWU5cE8xdC/vqVSb/kimAhwFIg
Lw+gM0N8eesaYX2ssMWdHdYY/7jk5jOyOxg9iNGQNsWS7ePqtHCHvoBX07ZgnNgj29/Wq66gatFO
sk4adu5RSDOxB+MdCox7cCUm6mAmD9yIbtKx+760/TQr+KJCUigDvvPi67XGJ0uiS/5kTyxgXhvw
+Mud7YSk2+3XuaQFywKdkSftTWW8d1Aeu8BRjKePEFk4LtGnCLowpiRBroyuLYRRSzQvCOrMnUtq
m4hCSHJ85KcOvof5/xYKXNJzU+ac7tdfKoZMfWRyiAJ+IVlTwn3cOaRuKKksuXPAYhV/obNXxLWK
WKxwLpRq8sLL5xBsb7rldCAjTx9extiabKhRPkDzQQB4mnqX+I+6D5WXh7N1WjhGgVbNjPnjlwev
3cB/n1wul3JuGOD3G3U/f2Ins3+LeRkXbeMn0G7tyIErBUXecM8udgnJSNBRgLk8aE2crQxba4S+
SJuZ/3cOEaXb1/8TzbtdjtTktkG7cyAp6I5rp+m68Nqt0xH/0Vigm5z6AyFEjmL+kJt5z7/hBRtU
KfHaaiGsGMLfPdLTj9gDrH2NELUFaucoMl3uGmdY7Ff/dii4L9lHUXuki39VcYA0+xpDO/wh5HeP
Sq2I7RLaYNgYciQZS6mNHgU0sV87Zoz8EPtrcdPv7BgO4ARxpcl15NcUC5eKBT9WnHEPYRYRMdjQ
YEI5hiZUFSaZaPgiLRHG222JrHCbhE7KhFckuLcWRzD8EYI7HHtZP2/ffkSk4KfY3x9KB2rHJWn3
DCpQMgpyzCuH+CepU6MOVAHHGoaXAkaBO7XQAVJzmCvDZtUdh6c27pUBLAqXWs0qUO2LQNW/MSFw
0kRVv6n0ew4G5CjxQ4ANSe6HvGwQ8piDl+Mia+pPYNfi4FxtFWM/83uV0WYvceqzh6f39gELr3lU
/stTbP1opcX0S+ymOUjNko7LK3EMP5LLD1tiqLZMJdJB/sb/TZ8E8ce4/SoMrxXZbb9g6SpPdq2y
mMuxftMM7RZdRbcG4wqIUwtxP7/D8zayX0ctIWrRHl9XgKfrXcdxAKS/jYdBYrXlNwPzHdbH8ApE
TYg4TITE4gaj8/o0YH+VETlc+N6x4us0wdlEAsyvt4FiApdw46mu4fEjV28Nk62ytqnGFn34YDGW
zIJnCe4o0Tf+OsIwRguxkYy4yM3uzGoySaY4XHXmwR+V16KolsgS0X7EAYGv4LjnSW6RHKxgXRpB
nOvgbJ+7hwXbS1jD2wYnQ4KPbKdJ0vMIRxQ//9RmXKUBhz8hX8COB2vtc+LI7PDhd3ax9GdIMmjJ
GgP3QJVtyiruUs0gMbIQ/N5HkZjiQ8vQxQr6HR1Z80jznDhq3faDbYmnkLiXycmuBBWSIiVVuqBh
/sXAVVNx2cq+6vrUXmmDpO8ao1HKo6xVXMmcnkguKzqwfAOErhUGCpmuWg3G9M3Tycn11absYO1Q
k6SMtHVIF1xfZBbBHnsZXu2RS8k34Yr0rUwaKiwf2tN/lio1me7DdIrCmQ/RlIIxxKRKowjuzL6N
/KsPx3klq+XZIefCfflrVDr4STMHRrss2bBP5wc6hAOew31frb40xircd7roGDMwoxl2jv5uWOtz
PCU4PfC0qO0XXqGe7TsUkDsUMXFZ7npz+h2sdaGKUS3GXQvPmqRsfjtxsDQRTA1RsCKP0/PhQE0T
gwLzfZXj8h5jCLb3ioT8SzgngulUBfSIV0jxcyb8ilbkjVk6ohW4GEPpB+jNX+UaqLXq1NE7DLoN
xxp/lXADIzLbQwEQeRFtvyH2vuRk7XH3nccM0o7xaCchOvveVzEUwmqm12ZIa95dX1YDE8rj8Oti
Is3NZVlv5wLGkmH6YtL6iXmKcqSOGl8yh41/PzMFIcjnBg+H+YQ9V27B/UgOYx+xZFjfRnUsYbt+
CLw+Nu3CEok9VHSVAVQPYFHKgI2yok/tfywD5+bSKw3czbyxeydlWleYDlS4bRJ+Btizv0XULu75
V7cJm4UHiDG59Wid2kkXa7csQwFXT4UEQrAr4IIXS8CGNxtG4b+whokf2EyF4+3/Aw3jhQPgEisg
bmQMiPn+DQUhpZ4xUn2Nxcs/w5AWTbuLkAevU3Ha0KhWY4w1nPviry1WKxfnyq4nR3zJkHBJ84Qp
d4BUuVvF67sD7OyKftJRcO80f4Jv0Jhi/eY8wgkjA1ju0+Uxp1m4WvoQHU7o7nGlHLKYNsCveO6g
TL8mCgzA7RNChf4wAcStVxhBKQ3tZ97XomtF6ObSUsuja3akTOk9vk2Dd9xFkLI6VTgIdeMj49h2
jnHAwpStVmkjdN+7XdjX31wRhW9M5eoq/FvnI8BtJ3Jdjlq9iBLYmigDNsTE7Fv/wC6Sxrcem74F
I+QrrjZYjnrxMsMXWrSJdjd+qG7XlIATdRYMF9QpCD9+p7nRwjyic5AXHuHcGmS8Jbawood9RF+m
TDVf3Ur8QR13BTthix7t3lxElWutlHahkzxMpru4dFE9atCFeYuFevCa0GErBz/iT74csy2h/os7
g/kBEC8mCAbE/AOib59Rfdgrr3lZelQ0UyzDU/qRVliSiVyfxp3ujrA8PVwDhQjXzHJhVCvoXaEY
3qSlWb5JhXR9mVTUks1UMDpV3vUH30d8hhZc/Y+PXeliOFXcsUcKa+b1gE3MpU/RVT7eeIpCKP2z
7HMQYleOoYDUq+hBslA/3S/Q78YFBwdrYWwp5l6VQ/jDB5BwzXohnIhpsrseV5tkbG4WcysldWqd
PCwOVvNUGfvAyTLKqw62QopFug/UM3/abHmDqPXKveZBS6nZIqVpX7RMVLcwGrz0VJDPLN8Lz7ei
A1yDfoFvOLSDlmGzuY2/L+Vq1/fHGxLZBsa8LMttWcNALRAqnWOM+GeCRXL+uqmI65O0yVKc1o7V
HOrQqVAFKiBRCsTvRupfGFA2kCf3kNWd5fU/2zViCAACkyEPWESIPaLUp0l3HD03fbnvGrGCVOxq
IeM3wQBArrVrEWGLpLoysPT9Y/jJknIqnemBfv9BDrSTc5LRMmifTCVX77GsVnR4nKR86mUh2kdz
PFRameI66UvwVdqW12kY0SwnNyX0qXSPK6ZR6LpzArXeUmOV2uzLvWGwpWCDqEZU4ryDkjVDqOXY
S9eEva3xiScOq5BbDdOHQaquY+G6GPucsdNMU9qSUbAE3lcWRaj2aRJDsSM0YDoRePN3EdXdW6DR
MAP7ltfmKd2Gvd82oUZenHw3QLw/itjUCmzDw+2H4iZmLtEwdnfqO7MhkfJ3xooRXAmso4WOz381
Zid4iUaabg879KR7Pcw8TZI5tkotH1U5zOdQSRV7r9D+6GCY9Gj1P7oawtxh6iYLOMNX7+AjvJaw
jmnzCTZwvzx776k5RlXuuUt5eQy8zFyJHKHTJZsGN2wtPbD5OSiBDTP7nY162turwQd6FurI/Mji
0TJEfpQ0UfYCyg0rVvlg2Dmv2Zv4Nz3oGfTzwizN4dPNknnDx1G51gBBSydwSGOIUl39is9px4e5
epF7BILIDikvqo/Vs+41nj3J+/43QkG84dRr0L6+z9bassPAh18i1TDKbtU/+Ju6/dgOkEfJG+l1
wB9LTCB4QuWgN4lLQCemHjHuUGzMCdlNVIEDfksNElEAD3KiUQUkXMES5lhEXNOnIYq3LK9bRTLr
EkObWV6/0g6eC9l9BLI41+UpgmEimSGmpl4UWkOrjZXmvMY90RW+kuOcOmBt6EMCw49hRutSvHIU
miIBfNhu9BHWP7eTZPnEkKidt6R8pF5sTs5dG4ODvvsEVvvKnjB0vuOxMPDJemIYm4AjeEjyjvLi
qzcjhp23pG/AjBu9HikHYRIWeSyPOP+vAdl30oBf758GVETIEjZ7FQlKG/5mMDHS1vL8bz/hdVI1
t+19G22JJ27t/rVlybLxKW+ZAgqdN5fpIwSX40LlAQHKsUeQCySoO2XPGQXO0bzXslJ05O9ZDhHk
qfs9CkjqsB4RRWBUiFLp227p8o+owIaB/xbRq8/icmPJBowVrNMAH1tXaqO8m5QBkAhmheUx93mj
oGRmCC8m0c7cVnzN4376jNyRnHOBvk/HPgoLwvyV9LnV6Y/chViUR8A8a8c5ohQyW1vo4DLHwP+k
0PqxdQ8QMq53VhPj4mI8wptydqY6gq4oBcgPygV5zIxtlJq+vZc4E3eRj/PTuu7LuFAxF8Vvmlbh
yP6sPKq2vGLycqPNe9idtIvaiTbNzmwMSxGh/ADmilak/y4jtBzfLU0Def2A87jdDDl5gzxV8DjF
22NyuXKYR7aIcLT5DJdOavN9TUX/35ZRbioQBlB6U3x7VIqK/F8eSuc6QLqp/1tsYOAXfyWxSaEG
aooddXpZuEl5wycuezmWOT4c6qNVhEXVwZk5aPXKYwpqxt8TLQUbim3WlgQ1eKcXSwGyzPjTkcLb
Z/65S/Mk/ZxVr5wSPvjgBYO+dCitBsr1QQMhHjupsRrjo5gNV/W5xllfcKpKrOX6nUxVKz16rkb4
46bIlCwKhRiO0E0CMdJA4HV7rY8exW+cn7CPDijAEsK94CRQVy3g3jCRcxOGNceHrvXGO8ORYRPj
+fVKX3flpQhaBuGzwwOWX3IUT5fNvxKX6gKd2S5N+ChGU7wUoT9yZOUCkH00mtuQnKNx/kLpru7e
wD0yGgQt2ZGCICoPP2qYO3v0EYj1zI1GdadgJ1+BWiY3IASmjgsmwtH+/pyiq/WRBqx//YSMmzAJ
5CTwMEvsiFtkJcnCG0Wn5/jYzgIHpt6yS0n3TUCSbVta21sW0Lict7MrsFf+a3sOiC2bEZGSkRyC
hA52+Tx4eoPcgo2OQipus4NskYvh0dLzEhOjtcNM/GDaxkM+9U4fthr82HJAa/QuEjhoTjP2mXkp
hsapgYNGOg8N/6Xujil8mGyPghO5L+Idibk6Rf2M3UIsTGf/SG8Z/Un5YGRfAVaJlHAgBLToiPld
KJeBrnxlDudvjuBSbim3aByxpH8XvWkUjsLwltRcl7g+cWkdzKwzqo20u8hi6hpVORch3vaLb7VZ
TUb3kLc23i+Yi9XU4dr+IfWfiM+iiQtOxnFmB/WFBVjHJD2Iqp2Lkd8+ujAfcxk3bo8/cLWpCdm1
3nbBK+JgE9lUp34deQMtXCmMK75cXTN2kidQIlV3D76HOSfi95aXnbemkBE5VUgK1swO+9FwajHV
JE5en8xSXV/Kr1xDlylBs0kePRj/9FOmH8HFztWgzrL7ogpP6zwVIPDaUFy7bUX7boTa4nYlTT8e
cEJwVzqln59ubpX4VzxHBRDSBpkKN7XXxKyeQpvBamszaoba59OODCUsoWfjnn/7w6Fe1wZgwUKc
RyvRwKYYzKcIfBEW3pc9JAqutNGNQrR4ODIL4gvCHrFOFM2uelU40dhjJJCkYfjuTBA/5cEjHG3V
I6w438k9GS6g6LICWHS/6bD3IBiqN5ASjh+Crze2/JAPLZNxgdGYfEiX15rIjCxgA1lfYdyEOx/O
3t60LrOclizV4v35ZD/Fxg+VDhLIjpc+oOgI1ryeFzRI7LDfJRS3nmenWPx0eC+o0/VFXnxg7KZc
oGc1Qb/C7aKCQ1GgpbUl7DHcHwy6Qp0sziGbrEhdloln7AMycn72ev9jbW9q792CJ5eUlBi1Ua4h
xgE5qyxft2Fcze6OYyeTHtXWexQyRtZ+NzVZp7quYfL0PlkrZUWFpJIW4GFZn3n+ej7AU99Syudu
1TvbvBbQUEuL943CbzqfxBXG72wPujL5fS76WiqCjnyLa+duWSEpJkeKKvPn833HEokocUyN+vb/
b/fpdtJAEreq0fLeju0TTHU5JlYd4UieGZMHsK0xQ5hBnFVTQx+dzt/P+UoYO3m+q7h9eioOOlWW
35zvcdXkq7LPyq4FxmaHyDg4XdtmhIFqQWx6gn/AP0rS6t6ZGX4hyo/VL8ga8VxFnTYhsI/xsWFn
3P7wlXU6dsm3HjU3aJh4qM3Ia4NOCKsY224K+GGMWtanDvp1td6iPznz39sJex88GAV5/0CQO+uz
B3/xP5O7/PW03cJ6xsQYB9Ty769UgtGJ6GRlfhf1UdqchrsYMUk/wpzMgikNX9my+mvBQYdnMdUN
2YwK7uoh9RxJTv9QkeLUgsi+QkgHhV6hQnVMtVW8wv3gL7ba3S04Sn6EnNVkK6Dys1TZRHBmuuJJ
2ojqPS6Qo6J4E09nDhOSw96l/H/5ZQhMBE0ZygtxQ+vgjHWPVKKKH2ZNAqHSOQNuZYaT85/yqXSm
i0MP7jRn4HYNOA9Zz4Yep4wzTWEXea+SIaUYcR+RvfeKuZqOKBzrtwIhBm7a8gMzsb4lI7If5q2G
UZ2u7Zytl6dNAaBDBzDt6fcAAMLAt7uWsfWAuzoOeEOPWLDcvZbkV4YQaPda3ww9KK5MK2qAleTh
pXHkW7n47+KIstAfeKPD1PavtcwDIvKTVpZcLuGMj8TuOTvQ1zmBE4QyPNP9jIkZL5pXi4lHgqwt
AlJrugqgQoyPEAGCT95CXnkXQLPXqTGTE1NNKfV6dQcTiDbPXPpx1bSkcW67MKa0vK+/4GxGSifG
WvOLEogEdGCUmFkQjg7OuWUVXpafPwTGqDOXBtvdNE3OxvXc/E6jQlAE5WVpIpLRgTiYy8kFE75D
lK8GPtz6zXJy6/lQQs98hro7Tb8337rDtm3QSQ6IuIKwmSNIjyJ2UQADk8ncF3y3onjlzpykJpip
Vqg++SZRXyf1UIoKW3RF3Vp+0L4+RCFJbTy3qvLWhdvAF7N7z4e0upRGO36HE13EOD2RBlxvex1k
1i2UVuVHdHfbY3o9WeYyE584o5pl+58mqzq++2lvaXqaetKlN1pnD7kS4HwDlpOK/wnqEy/Mk121
tNpZ3JxSaJoYZPu0A5KZEyXiRhf+3oBu835adN1sDf/oGStslJ/GVNUf76Dr0bgaop8ravSThtoP
aewnjwfkJGn7uVPrOOWcwyE7l0hIra36xvXBQtcOAf5IBZVs72X+BPjVtdENUaVdexhlzDiP61f9
c+u5D1Fa3jZ4MEACC5OxKILNPtiy0NwWIPecbz9qlSL9lldiqOZ1LNlG8CSRhifKx/+3tNon+5EJ
P9nNPwNqnKcrgTzjgEjNmn5ElmbD2UrZYGGFwWBVqNfAEXM8xyRtZGCSL47HmXkdLM8haYbVzKEH
YKs2iBZ+ZsihRGRoJvXef+tX2CAAYR3fGD6Or4F3ybyzEgGFCHpxkiSmRpkLAd/PqcePBIhTXzu7
m3G1d75UTn1FtPIRuHO4C0cEAdjsGr+xD+TV91U3e9+IPgnGh0PyfSB5ZsZY4u0ZDx7kGB3Ydo4/
tXalVXwhdbJIVHmcvogBajgCmc+t622oX4lBAJa6fNuedIgnmBvdE7FN6GL3UurevQ37iHH+R/fR
qYSr8+zx5nFRaio0qPr7MV8mY7VjsBTsJKX/30M296E+rDjK+s9cCsb3u4VMBRAsI+BM5v1iPCT7
hWeDKlbDU/jFgQSrh8bNCZQrO6lhYx3T+GNY/5Z4zsjJjQCpNvM4KDT/dAmri2hC+TyeUOucjzBO
iwyMofi0ezSHDLKOs721MytYUoRiq5m7Qtos4qSlw2qQETf9gz2cm4Vzl7bL/g5fpRItr5t4S16R
YibGTKJFzMcJx6QW9IStCnTEwI0GmHbQcrSWHAHGjw2pWmYqyromSQOuQ5sU9/njIG+BBcvVymj5
qbxOT1w/XLuy9kKjoQyD2Uqf5R8Ow92RdTPUgJR7X9S/qIH1TpENXmaF8s4Kbf1uI2mAMXzDtiCm
p9v6AXfuDBcrUiRCMjVA48J0I2IZx2HGZDhVf3bd2qFw47EdGFAIeREHV317JjNPCpDy4TdgQXVT
St5kAHrL/QVLSZcXYrd2cVfQApKyYp6P0o7nSH+TAQBADJgGvu/P3iw5iaadZBdCqc9ujsaN65Sy
iug1GUUHTz/VzmJtq+2sJq1kTeMTstYM07wUwymqlzwdFTZng3WezKdZeuLxFmEUHJNRDovFSo1J
hxdsXFzDZIM5wCQ1FXOrbS8FY5c1Nej8FlgxXkj8tVb+uoyf+IX7MBi1dGJapWkUkvRqzAqCYe/u
I2PHRY5krflgjrAy6KAwPkIRgiEbnYzajAzZsqdOjtwaOBDhTbtyUGFHQsw0Dd0dSBaYllsm+DnL
k3MJwoBYuyiTd3c2za5CimDzoce3BjOEJNOQQuYW510uwFne2cwOA1WFVjPGADyX4HyNajiUaKaW
H/7bhLON+kBONF1rBPSzJhphL0MEqOG5EWGDGQsclRyHY1gvM+v3rrkYA2HFqAxQlE3lS7699T8I
xot57xQP7guNKYOwE2VOJ/fLXVkwTTZPzGRDEIU1qP2cn6aZUjNhxE87zxWJMwlqCewl2OVsENyG
znedZeOCIeWVnzdMacDLBBtNghH/+s7iS9PRCs02RQjEH34wPI/fFRHWOfB0TDaSxWllD3cFb7CQ
hU1mu1z1F8Dt0jyufH4iC3uI448kZ9elPmMrbo8/3dvnTDwLvkRjLMYgEuNH5oxFpU5tbUR0z1tN
mVvUzSBYzbHQDotp5p2/vwddaI8Fwnl1PJoG0j5UoAAfPh8bAwHEu/yKimyE3mg32DH/4CP2teo4
FO5k6jGWY8TiM58o/4Awvmy0Qkinpgi3KfkXP8/82a8v8Jg/imnJAMLJC2m/1EJE8C0MAwe9FqOE
ZDxkcT+z5gWv3DltY3yEYoLXLr28vKz7PISqgRxtelvWbtX5Vwhvs1WbBv92ulKH0u9/Splv+uB6
A6FgrU5uclhULxusLO1HRliSzJNSAeVmi/gVrTTdYs1MSzQG6MTC9wCWg1ynfCeZkM/+LM7A+Gsw
EZJwG9xsx3gkZT3NnlIaYcQrVH/sKiv0iohEyK+sJTAv8HgEV6takLHtpUO0C8XYTuRBmyyZa4rU
ZghiLznzZTwC3TGLL7beJEBWelfOJ584Ub8Ze+X3n2Ueb4vVuAeKh5u73FJs+YN1UNynZzHqTzOn
2OdQOj9v4IlnrxoC6723JVnzAzYef5k9NSG2p4ROK/jy3g/SY5rpcMHkUIF1QJQW5XH++4qp8Ces
GtXY/89nvcFyFAcZXCiTm259sr98kYJRoYaoUd34yEY1CLT8c3X48IjS1wYbpuf4QDXdbkHNyq5e
HLJMO/LvTv/wwOF3RgGFgr8mcdole2sem2Utfxo3EI8S7N87kQT9VFT3i6b57+mYljg8Fg3YO/BT
pgoW+G2T9fmC1f4UCO9zPAZG9Aoe6Niooidi3WZ7fiO7uCnr4oTcwatXGfHBp1InRM6P3lT1+lWM
R65DizMPnbiwWMgFCS3tFkGmayfhvxJh00jbSWFyAYtnpXKioRs571JRIXf7C5+VjY+3wCzNilmg
gd5eGwm00jSTW5nDnyr5WzR5fZo1GWj76j03moJgMp1/Y0xB3vKHyyMOKij0yR3Ixvyu2D3IemkG
b46VdDH6w5Mrc0iYxoq4CujGK7AN9snWlrouOyhWKfDgQOJkCIXuzObKX7x+bKb/x5f/Fy23OXVB
r/6v5U7X8TmxaqnTe3k/QFPMMCqQxPdzUWS+b5nR1mwdC7dBYzaM4Urc9/NKZSCqAUHUrlK6Guy7
is8JZ4iJK91bDoaBrUV44tS/QLbe6r++8kBJM6RPFIBJlhJKTOmRKUe1hbQcONHiJN9ej1hv1GXt
6dYDQkR2wklv8I+4paO5+HZR1y8Cg7TQr0/94L48WaYur+mk0gyZEfjUy7E/I6MhLOX0veHhFVJe
lf9mNr2/HPD1NS95hpJPJf2Aaf9s/ytaBRp0LcAcbHeQ3GLrTTA0lygOpT2XYySwU6GfkYtxf+IC
eqJowHz/aXKVZP95Js01HgLs9YO8Sy5PeViEZCXG2CdMxkqAd4Oh1pcXUUVz2Ln/4ZqII7l8EIkb
m8QDkBJdsET3FN4rK5vPs59whpxU/hoaLwOLl7vh224lc8KNLcgZohkuoHfTX+9Y0YjVBJcHrbVi
dXyhxhM7gXBlW8MOQ6rx5SGB9LEEbufA1ggxkaJQ4xyCnXychPZ5KmYhKzDZ9lfKnPrYbMbJsjja
trm4X9Wn7x/OnfbKQQJFk5n6NJZ6bAfagfJVrVxxOew8TA7Wy9f4+MioV2AAgprsvE7DBLklc1aL
+gBe6UxyFB44G9usJKXv5ULoML8H4492oUUAE9iUpaTnv8daOfiSi/lhRO0Y4HKiQsYmKvjyK1ca
667N1Lck/Yv5/VdrM0dHQApoKqyFe4PII+xBo69JlhR4BbcvFPDh5+6lAemb9lymvx4ThmF84z5p
uV8FrIuLBSMPIMviHgXwc1vEjTgKkMB/JmuBHO0jtiu1XTjkh7awQTSBuwoRxJCyLUpRxXzlqazX
3y3SYx6I4t+d8CT4sqP+CjFfWxDfJMhhsTKroOM2JaZl+ijB6YfkuWvV+wD0QKqQT7u9zg9cz7dd
XcJdxbWkfWVfaqovwCtLbuU0XZZTAGxS9k7zbjNTB+G5KBk4zTe8Jak9CUwAvbtFBsNhqx+oiTki
sMxKB+dCi/Gn7UB6gcv8fBclf2Tr2aJa/oaex17T37jLY5o6DT0MEBiFHMwN/tiVMQdcuOy/CY17
gns7JQ5o7uwr40iCOdThRGFzVGMwY23sM7eDW+HZtceqqKhzotm5sd7fR0lujuj0GgR1xzoF4CtN
nlNMZsceMBtW0rM0+lAgC1A5uvnrd7yM2WTVPHHCsS7IN/unsIqfzYgHAecUl4GGTyevG6plTVxx
I8TRkyefteJLO4QhOPP02NVyJAvB4bOKQEF7zGC1+eCSzc6bAGnzZ/xUsKjbH9OG3iWYkhc75X7T
IFrO3pIj3vmXMTmoCLpqV68T7rY6ZiE2LYEV7BM7lJzgwvQ8C573RicKaLsZrEDmDw+0fozZ0+Xq
FgW1kuCc5XLlDQ1PqA0W8+h8EUY0VyDgxLsNfICh8hFdIuECqs9eW6kbKxuhRw4Fi+raTOlkhKdq
f59Q2rr1NVf0aau1gAkYQYUWp7FCA+CbXECi8VN6qFK3aUSsXKslxMMyu9HEiCNeA5oh3jP7B6YZ
ldqPNk8FA8cEgToywEQxcGdEORoGK8rIjgQ7iw6Rpbj6CgmdGJxyKnVVD22+1oePnHHxOBx12PWg
ZJ9n6qJ9F3xyhhTjr2b6+bx2U04zCfoYo5I4hPEoPtkYH3WXvhAaMXTt1GYrIyGsDvoCY/zDDMQl
kqawfagGGTRHaEzEFHh0NyzEAxHwsXOHZTwg4GkQxwOS1UF8QceBUdWtvTBOL1JXPTcS/Y4vh4rd
e+K13yhCCNP2LDsFPhr0/JhcqIeuz/ozmsweoxoedhpzyZ+6Dv3hyNRKJZkaofwB6ys3+nJE+pqW
L4HTqoGuWBtrVm0hhHQspiPNklvJZ27LxYcCmUuKdXnd+WVI68p28NKh0azqvnhB/j5sgSC3FVgn
jCUQruNyRwl5jCTPJAx3QCvduY9r7IYmk/0/C5H6p029ny3B1Od0+mi5M+vnyDRNyYicMudzgVIt
8kon2TegBTuhLmeuA48S+EHqMQIvyKrYK0O3Vc6s50tjlVzeHRNggm7yK43KIyY98kxB/IznusvD
8q58XpvxY9oLEzbaUWnDnrxpxElet735ppBnvzehgTjtbvyz//cJwtdO7Ao68iI9iFKS2Z7B43A1
WEUsCTDgxgGUbMe+HEaYM/apdeSTqM8z8+yConrwE4PBr0G+5acPigCgpcZz5RLhtGyGALCQ1nAz
wYWNDkfdAhfrX1jrpyWt/u0euurdKsbJBESXt6XYXFoebXfcpfN/oUSX9fDrMpO8/ZVgRsh1IoBu
AxkAbQMA4rk20aYRR2w3xuaZq2U9UnhafeyS2J3SQBNFn0bduQg4ZTQ64AyEArohmvQ77mFxB7Ix
1Z5Z64yY8Ds7ZEfD2ukNWBlNFCMdLNb3ULvvTqKZxfDprAQRBaAztVYErJr+t3G3kHxexsfQOGZu
3DoZCT7c7R18f0N9F2tnypEcMqbyBEJJ2bV/cnOirx7JQ4mGXHbxWTVib0pqbXVvIrBmDcv9Q5wh
qA8hdngCcUXT37mFEWQYQGG1psQH+hkP4EHsRYyqRh1azuYb8FYzzeKJmD2+1vVOHnm3LwyGegXQ
xLJrqJCEwduJtbd7c3WtnIebSWi1g+9i4clABxSq6NUNCBQtYQ9tWPx+Q93pjgyqL9YJJgY6rsP9
m9EzpUeMH3+z1N3HaqX+OBcBF4ZcHxppzxEm1N/JvkWzsf3618H7HS+yi57ytVYGmrA4E0/dI4YM
DeqXjy280PMZd/90DCwL7iFuF75XZgSUA2QVgxcjzQLtcl6SjSw58Q+YyPprHUte6CoSeNHWYz2L
TLcsoO2jWZ+St2HUxo84SQBTBXG+sM0r5IPH2wGgAHZ8qEz+94zzdAJN73B0l6h863RCtPhb/Zki
9sGgvvtmyKnrLtYF2ATTdJC3FqjyCN69CJi54TIOOp6bcYtPIjo4zYaqAxGXNUw2R18F27VW4kRU
nWcCKrFgomQdD59sSE/i1x8zNTG98+1xmAoyKaeJRzESMtRC9J2/yVlN48n3jdhun2dC+U/WQkhn
MV6iDYe7uWOt+kEFRQSGwnypkiQVfv6EqIiKuvRnR5LVB/B5EPkOMzHT6+9gOdPvY7oxFVVUTF6k
UrFf309bKncTfiIwdMacpiPhRp/aqbI/BbVd16qCQ/37XOY5xmqP5OBy/eq5loIatBqw9tP4sVb3
dmJLflwTqcF129Tr8VxGeQKBeqvfWP9XZFUCZkR+u+AqNKjOahp3KObpUEElUNzL9mhN8gWR5wSe
VDMSjfXwlVkUs6NTvFtS17rmodeunZBlXjqiahOlK/C4pqYhFnO8rNFDWa7iY/xNDnTtKDMllxxQ
mIPyWAvuiFwpEB/EV2ne4zlGHXuHIpVI7ADLU+OEBLYwQ/8iEWL5QxFvVGvsZ83WBfxlXRCBVkFG
d2e0a9/2QmOCwpHHkCXINMG9Vtixgnwbm8MViug0Vv8wdWZnfCcu0in4qAxKJZ7zBX5Fy4uX4Lf+
kmD/NIRGqgIAuIpOMlA1ASip8e4rKzJn+0E/mRQADycT9qMvhf795RZcQ0AAqopRK0wkTl0Go8O3
mADHXc8+xINi0sAHq/prapoQ4uNm/b+Yd330R4nnHHpHYb/5UzU6S74mjm+0i+9ddCH81T3T8jdt
y/kmbRRU98w8iI/HmjMIeRZSl0rH/Ny0TxSE1y13rMAJW+g7LimiNmOXFJorjxKJJgceUJYnMvyu
qNn2gWSBatLzLQ0YvbIltOhR4IgX0vEDpBif1kRvY591atNUzudA8O1BP/RPsVP0ep6qydFX7Fpz
rZk3D+0hL9xVBnKCIc7jRUGeLMk1QMj+6MVcRwAKMgi3dYKh/mHKZBzcfSYC5yyqGDK85104tqIy
dJJoQzINp6C+w75ldLk6BHuJ2hmaxRQh4tc7w4s+8u43Tk8iLFDDfiEwDQ9D+a/JJj/Qv086KQRg
aggD0Zfibjzhuei8sSPF5tUlhTX9A2cJBMjPfGWMMf/zIAPj+GtxL05xc0UEIHTZ4+A0Na4K0D9L
CLciI3xtj2wQvfF+zjYQ5sSk5yGs0Q1n+/iwOFwMLpL3TtwIsLgBbGDcJCA+Nxd2s3Zz+M69ceLX
nxnijgBz6V97RpJFoIiEM5E/3ywSGrU1rRS07fJ01hsj95u2PgVdCOxFKFMWe+zW02qVtCNHMDeh
87Qb/dkpVuoR+KJvZrbLQyGML4nijxywT4TM5ydO0phQcTzXFySnF3zk3vV8bOFRBGg7XDe6x+M9
tbHNEpxv8SKxIB6UrY3vhBK4ieXESn+fo4lGFPJNUH5kUsiJe/7KQN5dhcCVgOghrj+nrXhQ9UrO
XVnIGVUNJi9Jc4Ip79N2zDou3FyRyU2vyv+EGp9s9bPeUHH2uFxnmo/0RsFFykqMX96XPXSrwj4N
7v804Wka9BXD3+OxAjqWNyhTXAY97AkIE3jD+Ms5UkdHZm0vREme0jgWZXTbQ5D81g1suhaBl1C7
/VTyaKpu6dznHf0anpi9kMHxaI7Lb7w7hv1uqkDecihT8ilTBoNrGCkCNJrw2vn1IAIbFfNw7++N
ckCtWREBqcPNSUpAdo3Bu0G149Q/27Ud8thTlfFKDTurO4ctL74shaqLjHgYnLnhhXUlC9C5PflU
A9vVYWaqLVyedH/1TJR7CIw+I3MQ2ADZ/UlVHZfOE1XHAlQhR01ueFM+t99xlISPUM5eoiw941TU
D31ItFLfCfmnCv9cirRhb2XY0V/xTei8IzYg84iZt0z/kNJYwnw+LptXFfSEW/gfGaUhtmhIaAgo
W2Xlt/IycH2fQVZMVAMEfun21ZYNzuCJdT+xlJaJO1SF5LksBoL+6CM+m/tBKRXLhrS8ZbVVUxKx
CfBNiLSecwcaGlJNR+Tr/DcGzQ4DRGEEw/r/0dK7Frnv1IqlgM6X9eXF0z+OnFCqyZFLhKpYV3DZ
KpRjxrjiwi5HCF9J7D0AdcDCy1z8XaVQ1flbXEIi4FjnArZQITNstLJagScOXYKUhuPsy9anZrN9
JjdLf0jOCJn3jd6ibwXpibKVO/cFLbe5pG8q47b0CMW8npX8CacHCsPdN09z63UacvxZKnPxbwIF
8AmILG3DZpXNLyyp2uaOM39AVppJOlUbiSCZ0QiB0CjAI72nSSfvPvTnMLpH+Nj+zztm2X2sormf
bpUXmIqQ7wSerVF6ZE0zomiBtGj9krbKfi+R98Terp5M5gVVLGnSK2p8MwJBIiVnpBHan4O2txyd
mPC+/czXZTLV/MKRvV0D4VNKQlO9sR57hOxG/CwKsXZJKsb7T3rp6of58zBJ2280BhlZqASaYL5C
4riKRObyZKN2zQJPFWBc6PXfzeuFXNA3wR50gk5xj71pE/yhW4uNg036dm4EtrcY+VN8VxIY+FQi
iaN0kqszM9oD8F2dY1AiqqzzSB2GUUyM3Fk9OYqNUadx75vsCL1LhpBFVnOwelMQvkLZrFxkFZPN
GMrAs8Fdnv1FttvSFSs9WTaKVj7j2nZVH1jqnhD5DbgJAWNpW1UDa/Fp5caGdVIRnm3fKvReiy9x
otYtMWdCl8KJXEoQtzRrs7CDiw1j3KyE+h3lgJScn8at1vnw7QYWdFApZs834x2dVa12gIU5eomW
tgN9+YldwIulmvdgeZZmdLRsYHIkwLhq1ysjeW665a0D5fqbjdl1hD7NUhTSyFzU8J7ogke1Pwx6
8IDV2T1g4wowvxO8vqdwafoaQrAyIs5es4OR8lpCQa7ucilVRUzSLbBhdpLY/V0SCQ+M5ige2af8
DPLUWcLdto1Dw8mhmBYQLyRhDJ1ofjTdP4u6TGsH7EdlBfMDgj/um6fBT6Yc+XO3GSqfU0XrWZkB
31ipQAOz43cvfMelI1yBkqAXQvB7pvYv8jXOzNHERRI6+/sq/dNCqJ2htjBsRAVp9TnmC73lI6/C
HYNjtKlOJ8wjV9+ZiVMlHoEUHO45JghzA+TB7/psH283C1P3kd+az/JrtQLv2H6gTwP4/W8+dtx6
2KNiquInifoNIUS+jDFYWQ/Pwqonw/Ua1xyF52Dqb1NIx0a7aoDt+l+GmTIFIfATbZRG6iFrF+5d
4QlxzgKQTCMA7asubiwCkYTtuH2qxWF+oCStu57xUfXyOH7jsDlNgSYppwJ1hCDAjxIj4f2mo8AB
9xBEP6pOrFpTsEaFfm9IJZmMfKWUdTH5FnXr57RB7VOKFyevjlc+uuMbzJ7TQpM4stYdmqEIgzEE
5cGed4nf0Q/loO60tJmjqI8hEk2y9zNFB7DqIYYujFC8jwooTwq/SzjGd3hz+otW6nY/Ix0DQ/Ce
N8QThsE9ax1uvoHjjJDz0OnW/5kaiXesHywNW9cc5TXW37o2YQN+NZNIcRAUCkb2ekAv+227GTv5
/MeyIeXyXMPwnCJm17tCypsTDDbmT4JvFUV7eR9jCkwXdKpQr6YqbriCfUyXfJ2nTwN0tqFk7uKK
kiO3Jb1e+Wo7B9QvSa4xec1iS4FBfDaKYc2mIwL1qfVleDQSGbjOjoIysIO61EpbYefV05ZPPjuX
KOquPMUBZEIh1VQhwFJOKiLg2gO/slxS64hkYhWojZkI403ife/ZqwBKB3NQ0A3iR82Tm71d/gM5
p/dg1AK6rw89XbPTLDxxBO9qHBBHOqjX0irX47Xpd4RELZyRfQxFTaTrydGOM+/K25S1Vlws4SbJ
l2G2Hemnj0OHy4YO9KQvzS4ez21qGOBR5CcJl8CapMSviwgF19sQ40uD68VYC1MOd05GSdQS8Zg0
OYF6A8ZIB4MFgkd/At7dzGjhA8CczvEFpZQD1xc6uKgg7OntmsWpa8pns6tAsyG7DPUtPAMfqOcJ
/4ffU5iWw5JjjkH2h5J8RfWLP+1AWfjyJzd2hlXP5jtUTkJV20uqSd+ynLCXjK56gZnWpQ/9iKgz
xvofaMzeqGQwE4bqX4UqWFBTiz+iBT3uUD2++3a0UV0QvHp1gJ2FbtfNvB+HbLzSliPtz+mbBH8e
kxaV5oNgosNyelgOgX3FoF9toq4qMdCABRDCWQwgqSdeFfwCRVt7mKi+ItOPBD5jESQrwQNgWaXV
YB8mx4Cp6kUIPUdO1uD2ITOBqdJckS4x2vg5puvxE8KuIacLUO8x/yDHHWWhT+NF4Q19PVLYAAif
+70xPupXKLMW8arSlmO9HTOL2z6s/LEwXr3GszNeijwJQjNreiKnYQa4U438Gx9vQuD2XTL5HNM/
OHQC5S0gf3f64rmnENGhPIrw/BL3EYTvjtvJMCdnN7lIRAJfNYxKo2IehSjbTzQbpazk4EW5IHjb
pRUZDV+R3fISKoNcQmdTs7nH+Yzq0mUENLU8bEedsz82FCsj3J11tM5tGdo4Q0pVB3NDViVgtf4k
xLbwdzX67BdMaFDpXYw5tIcRwGUFZtTKj03IjYj5c0VEx+noYskJnrY4lzV5hphp0iPwUpPGkTAh
DYhPn+YpjcTz4gFgGF2j9WFQkL/Ly0bIxojC0pbgyZpn+b1FUd6v6mzuDq4kuYOyncmW02eOJKdx
azsqIZaMsPgtAz3vvjk/p/FD+TRaEkghdFhwwS4Zte0cXnmp07lx3lXBDFRk1nKqQrK38qlMDyxz
ISRGTTQZkmzPLcx5SbRLedSTWxs34UCLzCa77KL6ulsPRf3d1t5PWf2bv6wtSU7TLZaADxMMby7g
uPWA/xqo8cbupPiasbMNt0tUKYbJMx5VnSgKtmZNZLrgbVZVvaOO7rikCfP3ReWvLoju4HR066Kc
RCvx0O4kftVarO6MwTipyscSgZofY0tBqw8TifpJFo1wLWtVeQ1losCXMtsF6cRwkJsLi8c/Inl1
JUEf6WiIyg0DRzyuV0XMGPpQPdVeLYsf3gCKvwZESRlJ19cwt5ZWBiW3yiRcgWKIKT3BQUMAZpFV
6+vds9qdpTaPJiZvn/cpv6wtku8yD4lz3sbcJznDek5UjRxDl/QVjkJD7HR/anZYFte9Cv6lDsdS
zto6Z105N5ju+W8BzYfBjzLoaei6Obbtrx1i9UgCd0RnBJzJ5J0hXGLpXCWyxAEJe9/7K92ww6NQ
ief/WoVL+Z5niqx3XQXLEH4lbHaAP/PWNPtxQ8vfZaSvTfNIXguLxNalcO95pmvF8beSw1BzXZEN
9i+HeifKMx1EDQnBxZVG0OJt8xXwhIewz1SjKwwC3OwcCQgMttQ/qhECW4HLpvrtcYDCQOdIytQo
Hn/oz4xn+TwgPBzV8vQqe5gq3TsB/v402u6vq8ZbCCal64bRqpVP99IehCdJrjFWnS9ZBde9ot7p
op4QbnceNUUHGEzYc9akH9fC6BU5XkKFG2tRJDOMxiqe3n6vtWe0mHIxLkfC2q9tP8HXfGL8zPdh
PzqFUqHpIriq+K83oWeA8dhnoD80OP6A1hqh4SDjxqmL9x6+UT/2ilI8lMW7cNdvqMVTyjlXRzUB
4gi4FGFv2lukU7B43xve12Ld1XLAC6i6NYykh/3Eb23bFbCYVDTQAEwAbWXKlkVDlGmIfCrrHfhw
BI0jx9gpDa9EkDR986EPgbaPfLlPJB/qcuzNzac67xfkDJzHJArlIOG69wRit/upaSrjawKZ0MEO
YC6Nuz4jliO7kDizhfUAMaGd+Xl7AlNlBLjSwDrGvLQqPBLgmrpamG8hQx6hOyAQDhVdluPqpGWK
SFGhNvH6i0ch/6jfp48REbhe8MjI/mF2bApc9H+K4LmPLlZgI8JW8KgrzTlhTs464g0H6UEU4FRK
MPiT6Lifz9pOj6ZiAkZaM3PMeuGJ9yV1odrKgYYvB9FDRc6EObyuLT8zkA0njTDXGzy0cv/ddrPD
1STTGBbxOpWJAhv/G7xqSYHl8XgZCOZ5AZJ4li7NoOPEzWC/bYMbOFK87x6866h/YPDm+VhW3EJi
FKaNR7TMlBdOsuqiqiunpNXQNdZazyKqin9DRkNg70t8vRHqfmieNbw3iiUg1adp3fHFxKVBgOtO
+nbFXcbcdbmOssWra+s/iD2MCcsAn6ALRtGvEznIRHFLhPVtId1AI9BGy4Ab1HHHfdWUm/O93V7/
aV+ErY76eeIx5LRSwQhIqxmObNKkwmQEZrVAL+dfaFogTOn3SgiJx9KzhdmBZJkYYRWOjNjmV9J9
J0CRShwbfgrZGTfoKet089B/5aHY4Jg8JE0ayIG08Bvyg4b1/iJnZoBgtT17vzJWYPmTBMINg31M
coKuL92OKH+vnJd9CwVQXNza4jxc1FMW4t9/BtCP6/qqevTr4vAeFs29+zcZsMf9Rm/OPvFk3IOO
5xGYgSnYQZxt5SIBADke7YT6fjlpysRtXzxzJW4rk3jJpuOJ4vNRp7OvxGDim5EpRBMbDWCeU/yx
yQiPlKH/rRenWt5nasrn02O8/I6eRNBsxS9QbA+GrwWWfJw8Vp8VuO41O3zsEn7hHDvX7qngUFUH
uF6hV4VQf/jRcPnlGXwz4zDEMUG3tlUPVLFT+wbL942Npru1USgs1JlLZAvYzo2cJPCOsnGYtGQR
AZMHwg6KnkvQ50dFFhwIEqWjvzlmX3ucMrsvulImd1Je1ZncRrdWFIvsVMKwgpSBV5iMJdJbVAgG
MfyNgVv01Dx/kC9QM3V8BJxcXlRlQ5gFL2f1KLhUpwQ1dzRT8EMi3WtD/2vgS7CBnfqqY7JB9yl9
LQ+H+6Y8SWHzmWkn6qAqRtpgFlRPxrb9/Pauf90Ag0OkM+J9g37fnJv0BKIDYJC3Ub4JEunpYetU
lvyyI4C+/zDJnh6Tih/ZtjQ2WMDJztI3sV6kGOJpVp7jwDsoEmTRMmd9R/l/DzmGerCFdRMmY3NF
8TWSX7YHCe9j2bGQsAC3agCvdGMpDxLAJD6EHGH6GAxSrNxAvycwy9RmiF4lhilFPm2zXpEqdnFx
IPzb2pExK5onDZ5ioPSzYgbPOumQYh52hoL91sWjoY91I54OxeXxC9XCFXSTcgM/oODr/F0v8EIb
yGh9SQ2O/q2N0TJuuWqvsvFa16wudE+NNVkKUzmT8N7LTtseEKHMwhjNj1t8xyDlUiyAdsSlHJau
pKT0dr7Pmcd5+IeuBdA/Wh3WHIkocQdqMHDyS0a/i8t1VlpELOyYwgYTLVS81pUo/gcSzolXY2F5
0QdSkbRSlH+Afv+ypHfl9eRKXKpl4OFVu7idC8ee02wLeU1CGl21mNq4Q8oboVg3SxiK6xHbmIJI
FhKxbIATJxTSwP0vKP+0djOAv8ciinHMc5Z7dXntJDAixf/eRz1JC5Hx4NgQ/tVSD4UlsB3d6KzC
bSUJuixcu5HaveUpMS+q10qOgBYZzkgiJKy2zNHKG78H92HeaWIV11BEnLkChp/LQVczYvkNlnyC
3O4SxdUDq359RWlYLg5IDhMHqV9vO6VnVbGhLZdWnkP06ZquWbCYmgykBR3TY7T2cf2MOtu8+amM
mxAm8KjsmdUSxXFb1CK2DNThsX5e+bjRZcJUia9u+cIS0v5lDdv3bhinLRGPHrzXDHEvRkTldCz0
2Fk38dPFmkmmR9wbHeEdhg9Y/R2iMxWDn2J7AddtFgYQS8IPMi3y3NWl7++lQnHaqrd9tHpXOAnc
J/n1FqO1S06GacDh0x9XHJpdBBcnEyXUKQN2Q6InUUGCJ5Fd4GaljkjIdV2H3WwMkomsjnPiXzEA
U3oQ5b3C7xsrSttygAs/sLXK0lWvio3SDSPzwZF0LD2fYCgZxEJuSJZCsT5YpdkGI4Dta8MflBvt
GdPia/Urhn00344rXygNpOzdWKnf+jk8rfdqz3njEaaJUuy/Ua6dRO7gRmj47ERa9TYxhn9rB/SY
ehxZj6f5KWAMH5k1fdiy5BY7dypTtcjI3Q+89FPZmxFTvo9XghM4ZEeVYrVNfOCgLdbHUnL/ehYv
l4z50dGTDlts1GgCPvUiJWHp9gGEUuI1aYbeBQh9kST28mkiCT8E1b1V1SA4SkN3kiLmiSBFXkik
/5F5Gkrvj7hRYPUIMYJxbkESGLUyKCe4IWcZglXuTwMfMvW8O2NGLkLsI+DoAKGBG5KGHsADTGch
sxzLS0/BAPsMLbAQX+U4NpdDSSGQ0e2VWrR8HHXVHZCfC/rXX8bhxFj8jLrEIg3b11jlQ/yi5GB8
uQIvfRhGecb1gi4rJHHRfGEzARAEH0cdju0Ec6ene4g4j0ukNAo+239c0zy2DeAA1ORbxZLSBojc
por9WCfVOJIWED3f3P/gq4OQ88iuGSmpY/1bIDOuhLR0/8rDn5QkWIw00cWMuai7wMwTA4W9EwNY
J4nCHHzwL2hlC3n0fQfpn8Ru2DJyejpKc7XzLXj/cgaTGL459Kb/7AVYLv4pmKc93mqf83GX96VM
gsBAoVde+7mH8g6gaTKorKKZpKRzcFP6ngLtDLMNbU/7Cu/ooVePqjan
`protect end_protected
