`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hD9RhqnvqitEdDN7FgX82KADji1MkoL73koQKOL4NFsVV2JimIcr6uB6GTH4AvZpLET4F05P0+Qk
myQOdGGNwQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dgFeIUtjL2cEznbA0V+97wiMXTGu2oZ9BaEBxuccjK9FViVENVvHIXk159EkE1yXv2YxIMUnHJWz
c+FUwnvuSdPvtrZ1QVSsyIfoWMm0+dSW+pqejU3lFE4jx7aiaYXqPUYP8aimi1m3sa2IXiERKjyO
n2UZdQhk6jBQovssUIU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jXqhjQT0nRa8RP8/KztNYXITaLqHTwU3wng+RS8Lt/9rMujGxB4jjWv77KlqUZdxnsFIoJ50HRBT
KlXlkUBRagT7RImmnYzrJMYfV1cmQqXJtVcQo2FXE8nVjeNG/CVOxpbFnvSGDqOaJdBy3uQZeQ2T
NIzaMsKH0tBl6tMuwaph6NgdDw4ZivN6q1e/hPDxBmcGDs92adw74noi3pidOVslVGjVurzD3saw
saDKT41YgVtaTjegcsQK9GeKTF2WiCeybB5XTpxiKeIfxF3wnjtvpjidxY26smAoyH3zy/FmL6gP
OWBfDGt240GdZNo0W/RSg7sg4nghFR/OGTY2LA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iz/1qjNm78b8MGJ5dbtwai/0H72tbp6OnC5cXJhX2nvrFOBjUgpoS3Mfx192/3j9mpiv/pg3d81Z
wbk7D/tMtcIietQPFO3dcDCjkfPW1gkb2OxO2AqQBcBVPBWMyxltxLagEBIhkQXLnvkBPeA03utp
8abNdSF0nXa9sOZirlQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q/8I8+lMqEwBPFSaPhsnJQYTpLpuLE/ShKf2aQmOKIqqo9bA7WNycVqkrZiVmwRxppRDFpfUzeMD
TigEW8ofjMgiWMzud09x4DzHuE0wg9sbMaHQUoyLvpsbUassOYmbQ9vAZ/sEZhBbmap7FqaWSlQP
92ZXgUo3akzjQ/UeQuzvFfNE9ehb2vZs2JWo0MsA+/3WUI5ASptGaO9oh9TFsauWuS3CZH7Gyg4c
L8KzWqYdrT+iFWRcG8fS2Ewp0Cse0O9aAT5RTJdaSfmuzIEHO1y1U0uw/ZwSJ35zaX/Fq9Oqg8my
lOFFFIUZHXJEn2vPquO4RJ+bzBf9+qM6uA9i0w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17280)
`protect data_block
NaPkmvwcQllby6emUH4CQk9rM76Fr5uITZuP33ujW4n9Knm7zgDcijpzdRhvrrmzl0AactSpXKrj
il8lJZnlaK57TCvJ1pK0T9/Z9isNXo5EPjG6QG0YwWi/8L2GprFlBpmldPzo9/Voz3sEtto+zqSW
RpN+locEYyu0OSG5DFPfFhi11qJRiVKf+hM3EAag7q+FjapL0RuPDd0WwtEF6Xi+f2kme/nlvqlb
ITg4y4TvGEaaKLt0tG0rfeNelOJhKz0C5M+35C1OdgJnJdal+Kvo8QwbeXBUXZqsGP8d0P5jSNQU
Zaq/hIeYIk9uB5hH2u1fstHfakUy4aDBlXlL0u7TC9kzeWeNKGLgFOoZe6dpNciSce1hsRwV1nzP
W9F94bpbN0FwGZX4KwwlKWuHwSyxVyreZ8rhZcNcJrS04qktPh3C2N2lScIDIzTsDFnY8GprXMvV
45uu/QBXVTi2n3dZT/hpvni2Nph61MasqsGObRk8PKWAbrUAqQl3Xg7ilkGslEGSiXSh8oyunl86
FZxmWdziDDn2Tmz6p5PK/Q8YjGQReinkpnzYkToCZ3ZTpHhkD3CItAgLLQK7wMn4HSKAVlDX/QsN
RxS6Xa5GsqQwL/C9YMrlPeSuS4qqJZaONAG+q+8h0vItnUctutfxy6Iptedx4a+iulhebu5bp9NK
prTYXnJ707nr/iBnFnXgixMUpYOEmVsieYjIGzgFBlnXnsqEQ8L6mUFKKJc2CUDZH+6nzWGgLAap
i4NgtIU9bEWxJbGtrdVe4vBT5TRtC3+mruUvixTqxd7lY5j/LtR4yPztAQaKAlqoF0ISlctIDd7w
vJ9MieQeCR2ZlqBxIO4PtoOPRuXL0JnisSfuIcQpMEjdQX+P08trQwqEXrTrAjTgltmpkSwU04dX
XI2Lsn2PvgGl3uoWLGe1vlOjvBJysSErymotu6QxPOIfKAcA39QMS00566NBUipUOhENKX2QovrG
J57bN08LoJBB7+9Xasp49DWDObbFOdemeHkUSIkjcMj2iJfDP+K1QqC1PPDpwfyat7F79ib5Jo95
8W5fFLzJP9lfE5HOuqinRdQaUZDg7HCvR1a+0EGdDfvz9FSJCYdI0xI7x7hbwcbmrnSWyaKuqTxZ
Oew7W09/EKrvGGRpRiCvzjPySI+CMcKpHYwbTof4JEGxShVVItyx5903pEL2T3+idPTNNL+2QhDQ
F7ExfiN1KHtaE+8liEqOv9V7VKkn0bBXNaTMTHQUTRCH/sgEZWVAMyKUKBJPQgRgjtGprWWCmJQH
2wgePEZFi1CqmRpDKSo8qAnkjOpxQBCxhMbMALgFqskPYVTNzff6Z0AfihOKEizmNKu8TOASNFP2
+AJSHZKQHnkggHs9s08tTXkXSAhUlyG2XFDIl5qjhB2tgjZVG4W419YKwwUdM/x0vNh8mqQ1L5Yp
m6XMleBZeV8MWp/w1DwiLTgN/EmFPsGpGgLtidS2XTaoup4b69ySVnIJusE//uycYCOD2F3YeVx1
xK56qk2te66FEWZ/tyjLR4Sbvs/pY8oOU2F0jtQyaclfWdCpH2zjhPkcR+DZDmHHCc29AaMQny5I
Qbn8LRZxF2Mcu9/JmnZcG2upvicJ/8Or69Dnh6E4iobSTUPkPm/SHja38dedgtYUYLaeW5hNrZye
WOQqj9mCZqJXhqJN4qBJ4XUAQsJr/2H0KAm7poHEO+PEGLQLx6JUZg/BqnL1OI2tl6vvbZzgCPLN
gwGmSutC8kroAFXmbjSHMmnSdT88mnmiE5gdlt084R4Z8ePyXyTwVGWG1vbGNFT37Yd7ogv9MRYR
YbT2y7AgtmPXGZujr9wtWN8fKamp1Vb691SuugYx//UIlIPM3l255zEIjRj1QEhzWn0AMEonLtzR
yA8Kq422Fu6Vl7jEYRzS997NI2ZQmLo1TPbhJV1T+3CStJtU7/Soqw1U6RxuHvonX0u91trLyGJI
JLMufGlLiWUvDLVPUlkFAZ+8OaaH71NhJ+a2fPhGTe42VkI+XWml4MO/05cbYW2yKAhGqXSfnJ40
Y2Oa7Gvlic3yCIYZi6+X+fZINLelnWBCWwXUih/rLN4i4E/np4reMbu3RIqM9DhAq6TxQ6Ljz+Te
wPpt2PPsmC6DEsVJk6KTxwMu0ku9KyXAEPYM1K8JKwg5Dc4fg+Lv5XMNlMCSoq6/Let6DxfQ6P1d
ZmH+PbYrU8+jYf9fNz48fd1kP4yrKNAk9XVWQYAPTgcU1IAx6V+yOhD4d9nqtaWHFiCYUe+9vzuA
i9+m5oV7DK/hXSY2kJNWUscJUrUs32SI8pFE/fNit9r3KHFflutPzeCDBapiKsuG3TujX9VJjqHL
rxB+xOdTnhbMaml8Qe+wKGvOPhvWFc63ErBPF3NZS3AZRGX4IOEqWiJ5Xz88O5YbqvSdFJ5fI5Uf
MpKXd21iHkz0GpHqrGEJWHJJi5jLhr9ZK745OGd8hlnkfUcUiU4XbbzNApo/WB1gfKCvRTZl5N87
20tpGf9ziyYAOhiIttyRIOvJtsDNrgY261fyqs5q6582cXtja/2vIefPrySXPBrpl84uPnQUvsTk
66x59V180GoH0m2zm1zQO6qYtXfEdzRyk7KkCpqFJO4TIHT153eUMoEmUYXLtjP1j1NJjNXH8zAp
MsEAUWeSFYr/qcWNpUEGBzrz+MYKm3LfDGFjaDztGVJDmzcwyRS+jAY3aldHcOgvtUepfZJE3LC3
r91fBQk9augqBDxogrLdcCOTaq19H68X21EOFEP1cSXNESqtpdg0ehHjkrEG12LxxdcOvWpksM+T
b6vNi/psaIN+ow+SNuudF9DNwml5lvaSfyGhlrhOLlZ0/V140evV2Jetg2ldPTUzHVCXzGooAzYh
8uLvtM57BFaIqdH7uxSB698SxWm//xl/KBw2Un+Y5vAQ1IEAMls6GZdbcVuYDeXwxjNC0A05UqYc
e+MJny3htBCg2hKN9G+/qWgcFySVXzpfKjr3cAmvKriv0IpuQS/vI9H/OZMb9hTM+Os8USs8Cue/
GNL/3KiApQNVkGlbzz1yd8q/IjfBL7m2Se+/lNlVwEGydV+dsTSkIdauWrP9QUGSnAXBO/DaF0Xp
y9+pj7v/p15hxzW7Cv2Hg9KI5olZp50CL2aClCf9zrHjbBtxniTQcDueLrSgJg0MDo1uXOEZc7zw
+7HhR+wHdIYw+4Ow3P6tCPjwV1et0Imu0CcGaKZzX9yK4epnbJ3bWc20kWX2KdFPjSfr/AByt/Wp
THqdNmFVhP6+jMVIIX0Vbz+YHBuatpehlZStNR4H9r8hH8wxrx+xYRDcIdajAQEM5LB/Xvcy9K0N
IYx+WW1ws0iLO+k5N5onV2z/xXnlI7a3TUIaYOfsnnw2kpDzBb3b5J6OPHBKkuhbS/1Tm+IrYvyF
v+qDAy6D5MxyyKqI9SzrlmZ+Kot7CCsGIyYFMMsAzk1z0+FRQXwLX+JPjrO/b05eOOiIbUdYAM0u
9dxN+ge598YhLfN6EFNKl1Q6Q5IWthcRHJfY8jSoedMbBg/QJ6lIx2haYM/1K30M33fQMmFPe27r
3UE7KUGK2cj+AnO90WdkCTQ0DWEPfXBRtI56sf3StWp6Nnw5R/q9YmA0AhVwtPWKdOHw71l/rpIX
O1LpqUW0+YD9QRixjx4Eip3adKEgi3P3qf3IpazrJ2Pg264t6kvBB6i/yYgwqGuXUSx2gvNwU8ww
qCiJDFr1AFBTKxpeySYapN3xw1yFtHw3874/gsww3Oez3KEmwvMzTZpo3dPgR+J5EqbKmmGhTRpB
g0m0gdYKrEEN6U+SsitmraWTEl+pGbGfzemDqKBwY4SDihyQGx5X8tS5dMnIXzYrcJRx4nc5xk42
XiELxif7BRQ5BzYnfZlZZy33a4V6s+VErW+9SpUdGyDkDGxURTsACXqBG+U2nDLS9apgzdBbXW5U
q+P9TIZf3XegaonMel0HFrgTw5GIyBp5Xczlflyvs20QnBWHEZ11Akl6aefQE44+jbV9k2vhKd04
gjtedEcHbn/nigYo7UpE4r7FD5ZdhBKqGTMGzwkZ74EixqyLk+mjx4cCC1cLn38oOAwWac0LQGCq
a3Hv+gEy/kgdiSpX4927OhDitnF5RD29EilmaLbsIpBmlNFpMuj0F9j2HO5cL6o9QOVN8+4R6DZP
hlUQ0btU6QAdk7kS1mwEo6rW3+EflnI7PSKWPUfsAYhZekibVTWCOlDb1DU54od6x+u4PNXnoivH
gxjYBcOUPpQR1rIovjrQ0cCxFWa/16oYLqwvZYivZ5Ddl+zdQhaVXd3wCtuY9PNBaVQtrtKoOGYK
XMkyIRu8Q1cYCyWtuKKF5ubH81Pi1NtH0zw6d5UnHE7/gbU5jVqdMQwzWhxvaHztasw2GBP0fhVb
GLBCZ9Sa4NGtAOSbhnN6RYRmmGirHHUGGWbbyBSlSuCEaivDZksSHgntWw9U3JEpoGDHxv5XG/d5
7U/SNPns6NbXc2DfTdazGXEuVMbHb2xhS6M5zZOmBwISbancREcACNV1F3x8NbLefAiWZ9Zu/vIn
UxutGJ54XH75b4BAios8WqHeWkv2G+49Z6Xl5pcjfAacxvnOadXHvXrmks3Jj4sbpW/97q8Xcc4C
5sEI+VGvI8l86PA5BBrdPyeUtQ+fs4EeqHAVic4fqtgDATkNFd0Yj4WKyOGpUj1Xx66u+gaX55BI
w9fdPu+XAin8Cv0wyTU4jPUGHtOkz43V2Mlh5PYG7eTtT4yhOLeG3VTaZX6Qqqj81ZvktZ4DKYQ4
W2nskaATBY8LvVL+6Vh60ZqYF8y7MyEYi5jC8DY+DXI/p1r0SbLl+7ZonfyfO8su1CLDzIYYLbNo
6VWXY+qAq0PhcbbvC10JiDCyp/aO+V/folVU+eJ+fe0o211N+2w/d9b5u3NMC9DIkKNl23xZ2I6/
gV9KYYy1rXcby+Ae5E/w7n6K90f04MZtpjU/qgGHo2ky205YSq6TlxmxFWYPd1uRDws0UOA0UqWb
QzsIN18fEOMk8O6EPG71dOVeqfXiKEZDSo0/sR/z8fKlQl/Aljir2wEJejUIHotVUUU4qL74R828
TX8A65rjXZ4WOBa7Dq4JllmAVePZM3qCMPbYgVsGl9src9rE+j6rKWO+v0l0UaagTpeoJ59OQtQl
Z3+Beh7SOe6nom3+S56qQSeFugGd13eaI/L1XxTWBVV3vaUaMObD4g14nywg8wa/n9Au9eb4HUNL
GEQPSSNq3uLUWc4/tOOxtTmonOuyT+GRnvVy/vAyjJi03niB1EnbNEVp4b5pAf9xtkHPjmCe5hvm
YtYhGPmQvGmvFTiYooILXpaskj/nw3IOXHhFUWr5GVMRrD6Orl0PVhP3wIfcv0GMlLy8tyGRrRDa
DjmWgqgMfeunp77v6SqHzAi9CnwYbwERU8LmsSIPO0spHekHvOB0hnbO17ecwF3KqSbeAHYm1Pw0
z/pbxSGnmgwxZYCzGfQxuU5MTlpGaB21bTowX0hO7w+eCxq3nTkGpZ9oehJV/Qwh1Xbo/hzKYjsU
yGoGRwDbETRkPTpjbtpYSPqI29nchpIhlz4ew5zCejf719JZG0fsn2ZDlqvNN5hI5UPSKC30bht4
6WsF0/Omc9sv9dFliZ3fgEqzNjiuZ82FC74tA/ZL9iAAlIzgo0BIl2qQ2TiaSoCea0t+rHrUKtZt
eYB6xRUXClrTR2jacW8cPliix1/FcPNh3tUSs6TGE3TlaXGeDQf1fz5nfwuvusk17QjOtcOq0d1S
qDhmx9eP0dmXVHGLDPocRnJk9O/UeE0b5Fikuj3n8oksIrsxDVYi9HGM8Wv1ou6fnNqEirIc0l6K
diAp6fML+uUMnR0MoJ3eHlnMkJGqYLE+ViH9HT5GfZrNyGHVgUTVuAZoOFqx9bDmQh3guFNqs5xb
JsqxIZ+Uv42//7VEprdHQMEw90xXBxjtd1ORZW0Kv7DNlrB1G53BLdGUpuH/k5dPseZvLgfPua3T
nQ2VlUVXD7cw/F4ve4qaSupKf/eKXkoDIp5hXLz4GqkrkOhuhr/fGClVHHIHfifZyFVP96jybcUl
s5BR+HuJTkRs6jV++f8V37WLw3PasYt2098BnP08S6HwHkkeJ4DW/E4sl78RukzrA2PRcZ4/q8m3
1pZV/VLKZIqtOYvRGT09VbCqOdTqHwoSP52SdLmTYfLQbaTg1hQpelN9ef8cKCHRQZHqqrdPWe4T
t0Wm0mNHoqerS+uUO3S8Z8nt9kc2eXqM6QOFdJOrI1I+6+MzlLVXE0WvP9WgPy/fZ+YLdE87EOfr
0TZKMoF6qJlFK4ZuYF6duJwMPtU7yNYzrH+svUk8S3FqFb7skEUGSqtcPzDnSgJe2W3GQBlExntD
PFyrly7WUk5TL0xypFgOZUeaa2O316rxUKcv98GCV3e98H8t0vxksjHB53WZJThGeMcwKVYiM0Cj
iKNWLGaUicrn9gQLOF3Lqrt2iMEXCHnnaUb4OjV2J7LBL8aoEQm/xgtvSQpMtKkQb869ht/us5jh
xMMiJG4mjSM2Rbqvm+dQFa7DIdm6FvXbJGftcn7EDCeWMEhOKQqswY2iG9MKzmkJHvn/zFnUBSJ+
sDVGYPiLLFHXaTdkYO2nmBXJt0dUCnmARgEnVMnm9PLSy+5fvc7Y7tFfXZL7AhxlwvMsM6X6H9rI
r30VXyktjY/pcdBNDuCDb4BqYjnUUA8UpHFpfbqYpQ8OzOJBNkZTyLpB+24IXrcwriY9N4stq3Te
0F7VDa3N70eevWXl/drc04f/ELjIAOmt3dfJjuILrjXnjHhFNOnGbqKhAG1IfjK8/5VMbOkH9a2i
k9cXUj4FehePfVGBVI5UXENGVSqj0d2qWRAGp6/k0O7VGfCKzXzThz3CqmXN4MejcaVTCTAJ8ohH
1xX3iFKgT0tr6SFTB1CBg5sDgHbZJlQoKoP0q6yPV0GrCCxR5BEC2gqys55O+V5JTvcMJLoiggTI
8LHfwzSTyrl3wz/GUwZxne1CcDfaQ4YcUD/JtJBPMywekj4MW9CSzIm8OqcaTqPFj6kosXyQs8ll
rRBRvjHhdMe/fXVjk9WsuyWJkEFhu92E0NfP0mLLqeecHIc4GVqCHV1cs91Sf7a940GMcAkOUfg7
/bdWpQ9hS0kIJKhfD5wiYBPppkEmyAFHoEITR+9XtY/Pmwb2dQLXC2jIftM1Cq9RLkVVgmhXNoDz
LAof3PgZ8iTZ3cA/lWke4V+zQ1QUTFrqPXDfFF2W+ffcg5cwvQug3re8GCg/g+odDgeb0U6DdfPM
Lo/l6so0YajYdqGvv1bSAnBvM4O36Gk3y103N4hBDpv0zicOB5WV4hmy8N9W40GGdoufUPAsGkFL
kpBTOpch0Fu5EqYwfX5DqgZRZHhUNnEmoc5k9gBak+E5BssvclTSC+hdHRV6vQiHLUrxxHb/h0fl
pxdpSZqEhDDo80uH++aBPu14k5CralDwBWwTfc9Qz1mbAExvJkxEavh/wb4t5hMN27XlR20x2FGu
YUiRfkkUoqLit1VnRdQL/9yVEWZTezKv8sObc3rXj32NGRr9UpzyyVWDVLQe4plgvpRKbrvHFW65
iW9WMEeoKz7+g2SOj9kzrGEJno9q5OfV3RHR15GRywvgrSyrciQc6JX5u5RwpMnjKi58pNcLBeEk
o4V36McyeQCMJOSV0XL5uFogqPHf9VqSZB4TJEVD82lU2wrTE56AFosBh4mSzvpL/c+QfGbr1oN4
ytEsVq4rruQ2HdKzIvpOcSAjN+o3j1TRobkvvelj97pvtzZ3CLvC2knPM1k+0dL0t6MzZQVQb5Aj
x40Zt8a6VYIUikFJ128GtnMFfP2F3KVPJWXso3BV4lG5SDIBDBdYXQ7KxGH4oKqzZbpATaq21kft
aWkHqMGI54ZbDN9wTZGWxmyYKibsPZg8fDKMqja2w9VIFwD8ZUcvUPFU5rgAHXJAd1qpdW9WZfAO
6P6aeAsDVY29NHAWbAsT0HjjRhtf5FkaIO51UturJ/a/bPJ+1Es10gV8XaKjs5HBQ3LRrShdDah3
uVAXDh+JH1yTa1lwBjSz+/5Ihv+QD/hLWRvysOyMisnoDLd7hW/RWo6QUZnl3shQvKfTJeqffk5+
Mrmv9u6A+KYSA1ZKgk81yQdwFsIryOzqQ63kYkYq+l6zN9d28o9H40ecsqMBxdQaoPrbBJTThNCk
8NAOdkd+TeGHae5WFNKTHMmqBVX3rY/B0rsnb7cdrx28g8M8u0DcX1OL15s6WvgnoH5bVNpr9EqU
c04JQTAb/+LqzFUumw4g4057ROOfU3cNuWk4QvwZsusL1KhCdLKBz2B6zK13SqaMnLOz5dE49gyq
VulnjmYw5f6QiB3KGFQyMKjM4UA0Zdw+IMpDKlV8GIw2yx41rbaMs5kFCE/8ODRCNRPstk8Grf31
Ilc+9qc6bEGjTjTjwqCRCruZ6XWp2bY02a0H0zt8y2HCCuBPqkqw6JaInWqZaz2e20fvfFGKJVHA
mq8n6kVtdI97wAVD8+7dYqy09CzvVW5PualtUCUEudwWmVoVCL5CtR9DEYy7vVkYZLNU2fQ83lbj
cGTUpQh80DldIxBbVUZmzOwwkImrFQnUpRtF8T7rd7iZFaH6giV4xFfhSNGCtKCHXmFas9xF3rK0
ARO+rHvlTnWBtAtxDginIz/vpLkjTjQADBU7BG82zNcT87K6q2CfyR/7Wpyi+knO+OrJWc/UQghy
aDaH7bJRkMTZJNjYVZQtqqiyKPhi3s4jK21BuRUtsfe81PshOSNQz6gQ68enDwvxP/eyZ2YpA5Me
PxeMpTOeojaXKA9Uigu2YPRGUNB8agaC54pOLWqu7hSHuG51I8hAFJatTNn5i7gDON74AfNSmUaZ
s4QPGUksadr1Qu3w92lIgwnIn1sO351HAI8+hJb9JhBItpVHLM7zBNJVfOa54tmREEc990qgnspB
1tuhOe7RLgH4azGJJknVd42Zb5Mc5teBEDZn8m0c8VP56v44Wru/D8obWM1DHb6Xy/9a2eOH0H1l
TTIQZIPXgnTHiHDwwnxs+6K2+QnbfU8Ha0UXH6y0K4UAdurjLWLLfNbRkGEzMMaOxDyd4k8404g3
yAF9IhUYrEr45WXcy+lCIuvYSonJgZyT0hGT6kKbtnKG1hIwtd7h4BRInbYnh8ouVBEUeF5O9qIM
JCgW0chM9YheGCG3fz70ZBDi7uJczdjfqbv0FwrhPMUdkyBzcnnOJtJnRUmymYpouY+dVA82mjGn
UGWD8mRnOxWFTPr7dzUsACrRPJ63vkL4PewaBxVZERFOegRcDI/MB6GsL+KHZF7KYXl/cTfxAfS7
Csn/jcvM1K1lSMHsre8TFmWoSj4dmyA1VgLV3QqVP9u0jdfyplhb/2pyYp/IQ6JnXMpKVxlKWHBS
tYVU38St1MGQ2YwdPpzzPiWVs6Vsrf30l8zbw+5keUcSUE2Sx3xWWs0wiHSHVDowDel6a6ZgoihJ
eNSj53QeFeggM3ID+7CV4neaafgwFJl0YSzQ7AP8qSXrrIPC0nea55fxh2+mEOnZHk5ugWcMp4ra
imCrYrAddMahWN0UC29TJ6B/56xNOPnowjIPXOzZuzFw9HM523TdANkPaK2m7MpQQcvwNcxHhRPg
6+TNz5k9UxI6+R72pZHDuShKP4JlFrb2zxaeaBJW5gXfjJcaMj+YEZJ9iBb+PvQ1uOupThqPz5ds
JArYQlDjZtYZOiVvet3JloxDel7L92zfX//7H/7za+0y6mrTq/o/GcjJLe62x46OM+zPe5qSvs2Q
MEkcuuWjcgzgZN7X+lN/MasTafr0NnILB0YQ0M4CQWthoL/WhwJ+0dRo43f4lOsQDGXz2C0hgPj5
+6k9fnwetIPRLVHozTaHAn0CJywWhPS9WTPyyT9kB+5NqVoic+6lG1I6RxCdyLHd5c/VMMsstsuJ
rYHGFyISzL1UaP5F8Rjrd3jH36GAIb1cLbJtAjLVFzJJHKqkCZFC+ZDIMnCHag/re7TjiNcLOyzK
ZX49CRpQODdAExMP66qDhN4h9+vcEw+fRVLY8yXiSP3Xkj6kKEzPmHrKB4apIK1nF028cUD6+5y2
/Rs9efpH/hs3zi49NWeEAx8cTg7Ixl6yC+tKmK6PvLsY6K2rAoc07xLhgfnjQZsiR1na7qAl9loj
ZU713mZ8KWDZCeIRSHjMaTAUC5bPcR+X34vbBnoxioMSguwCiUF2mDAa7gyLdCpXN2ObFWxlmkiQ
6BFJCV4bN8m8ak3Scl/qceGqILk7PTFCH1FJSML9x8v9bvc8pFV2TLICqEq2yaEahFXU8dgu3qZ2
9DO/5erAmQHeh/p11SyxiYy5282PJfVkxko+zSH3dRC5c2QzkCQkCQuDw7PJrocbjSEmiBRESkeq
nq86wXZ2V5ZzxklEkA2+oYK7L7pMZXNCUXnAXHqg/upA1TFQkgnJfStBLEtHYyAALjH+63wyzaTu
74akm4eGiroRmgrWQBud5L8K/asQLYtFIWpZaBMbza1uVqucDHYUFVDNs1RPooxb50/dqfL6ME6a
GOujPU6nzLIlHEkOwXwJGx6JfekCPTrHCGC9LF2kTar8u7AqzbayHN30My8iyjMs8hkdsukeXas8
REMz+RXVlS7n8Uuu4X9quS6HQ7Krq+cGpxQB9/qqtMG0JeuO18l0cskIpX9b/q3TyNqunsXtNYK9
pzSsdW4GgJEVF7627iiN0DRiq3Z9rAFB9FgiBI1JUrCnIssYPIn1p8PuT/njBp8Bsr7iQWiZ9g6x
BbaMqPUZeG0jvnkUD5dGEysn1w6sM0vQYDmhniUqN39HRiOEIk4w7m0J8GUOePWRqC4DblBS4h3F
ZqR3bJcRZPxcHMpffKddtuPp1TChtbEMxBoz2PdukJWsQH2xdv4FIlRxjhcn6QmHJ/XMvd4Uu0Cp
pK3s0IsseLbMLJ55qhKpY3y00JcBFeofVEKG72RvxUFjQdW5diY7ebS3upfNA09wUFhqMMp2pYe0
M9BFXXrtHd1Mw5rXrOXUa2jM3neC/Jig/QMss31876vtwzSa7jJQm6GTNeGj4tduN17c/g4EQXuX
VBClY8rO/DEWXXR5KzE3hPPkG3SPCGDOEK5jBDeJG+6kA4igBMWDtlHqQ/MzVCGsF1HkphQw4IPd
TVvlPNi5TyvXaxTV7IyFUq9/1DQNK6QCtrW06HvCmtjCEfxzmurenRFFSOl386Uvp5mRXbrZd9KU
yXnnul59u7M/fUm5kSZwqHkwyCoEpKUsL2X0dGJXELw08prBQTaYy6Vl+Gh5Y1sum5gxT3eLEJ/v
/4C4/MX80HbT9wkxulHxKtQPNy/LpxipoBuXTivOPRuQDSvDmOPcF+YbreR1y88t4Ton6kPc+lh/
H1SseDU0Ye2RgOVB+HEyx262yA2bMzmyY8pmKCV1YLCWvLGKUyrMElBb2mPamOE2uMNOn45cfUpK
yXQOzye6c2tsTOh8ehOnm550ybzzFeeDgJ47UT2fsmmAMX913NxQhdfWiKZeoBn39S1ozD+Ao/6A
n9AhHFMakQo9kkYzjJti0FEHLGJxyW5T8DIvkw6+kaXMGojwa1NflCj3COqVQw8KdMEvKxhmZt1z
OJNYsXjt3yf6kniYKastUt/3et/JGmVJyNCv4m0ujTimi/cq5GJm8dlBGo6I8fYwpJeFvU59tYs8
GhMZMwy2AHcMLn9PNbE6XB1Glj4A+HuGyHlB3gZOfEa4k+htdZ6khR6WggTVFWZv9vsqYoqu2AyW
84wMlv16kxDU0iDM3Q1KgatNxpF9s4pQD7hr0objgBxVrjuwPQX8foSQD/Be5kqp2eAKdMHr38fF
8+dJZQUNUaYf418Q8oc/BoBT1E92jXI14PwDgHBbhpsIkoacaShRyOxqxdlKUAAGzqU9W1FMftzt
YSQrfuvrtszYNW1AT2KZr88+BAVqdWzkMzyd1TFrYIrn7HKhAnI2ClNFXwE8L8d5F1w3Acpq68uk
0xGN0/Pk8qDEZfYCsVzDQbkhBME8Ecdot4ARlA6vOhhJkIabtqdRlg2W9Hhunt2Yop9w7DF2ezPz
C6OL9/o70divy+G9UAfLqaPqXCv/6NOPsguKJh5DrCOhodyjgzUhlLt2Nh7HOq4TV+2L0PuYt6+E
plSt32ful5mu0Hq0i04CYtZBM6OK6D16Lscc3Zy3OSlU3sAe0AlwNEdZNDnQVjw3Y7XxC4O42NiL
jLg2IX39EgUvaSqP3zQknkiDPaf/XAayJu/xmiUKrc8cjKf1u30hkHOdXx2Fy5UcbpS+AJKCLuQ6
xQqrZFbbDicvwZsdki11Ae0aD5kyp9kkoSFXIjioh6tVdGncmTzxZtEsB6udpk1qvhkWWY+PRvgz
2cazfwmHOuk8kgWF2qYfWZz3RvgR27VH68883L2FQaUJT2GhGn1ja+QMwqFqSbuh915iyxycdfG5
UEvP/Iti7qjz28XbdXmo+RaPKslizVCaKitgXTMazTuIJL6LmPhq0BDTlH4TSqegWYpuweyg7V5J
63sy0fnWK55YK4Q8YYIMzM4Fn1a1jzkT8nmkqDVeaKCSga1vz05zHHoSOhCqQ2F0IluOcHFBhjY8
C9pr6a727WaQTH9Ok3WQVooKidRw1/WlR7rlB5CRj2z1DenBqNhBiKvA1b+PJPWkv6lb+Q02k2yH
ZIQ/mpfEkDWg1HgVx40K7+uumoTwZoBsqHf0n7Ne0RSzwrFvH7BJfA5HtlC1WnkhNXD8gljqfsFv
2WbYjGrpueLfSMj5xhSmWeV5Gip1Qyitn6BqQOvy8912PdbfUinaXJG5avOuEOFT3ReH3zQShjD4
mMUAEb+/7PuEkImzko7vJ/AFYNv67ma1Oc98cIeb1WEb0SgOY71i58SqZz7TINr4okM0CocmQFKg
lYsysTQv/qR373dVFDHA52hqkFLpqCI+AHARZ1JhQfelhsWvaRRuU+Q6KQoWDjnS/ZVq9GpFGsdT
Ipks0M2kR8cTcXO7+agf6Pyf+CrMG5xQIZhlCeYrsmPjmG6Jl64heSx3YGJMtSDVbPQf58mhukqO
12gd10k+X3FY3oTWrXRQgtCCT5IFeBJBRjXjqEkm33Es8jHkWv/tNRptBUoyA25p3jQJMSEhoSpr
u5Iy8JwKpZS1ECCRahph8TyW3TKDZAoTG5iCqYnJsjDP7uwEIqsZMSLH7gkHMGwOl8xSUsV3+FRX
0OBzgTuf0pCAFW9TCC4rx1URXbK6TevouaE7qsj/yd+2bCWzOCwLtL2rPXezql7yKCdJPbJFuJ5M
ZSAhyAcwKaKjzkYCfbfNpBAx3K2dVTS8LOVksFd7WwqviPaQVBO7b5lq76XK1TXGxKbxTkN0Bxcp
5rDkiFkgEcL9oAtwRCa2Sr4VccFAYXZL0oytoNbdX0uByLQlB8a2ZWHejXPgIcrmJB1fFPHNGgFk
u6O+CdmAPFqV+zbCCET1ssurrfzAQb1Rh+tuPO+ND9yj7m8Q/4a6sbTtlBsB5ZmY03C57eMBP6Ma
EsI1ITAVYkA2ieAi+iiuRYJ/cA9Yq1/4kuyjrTOnGgX06guBYlBUc92vgqrorPlmol5acfgmSikd
uK8x8etgdEq47JU7lCjFW0VnBXqhHufPEW0GeboGqoWnuKGTsNukxncosRn4VrpBciULRDa4F8QQ
ZV6HgWwKIem+p71N3cuySCgKvgHBxZFqdUFhSGbh3UgyfCq6t8o/1ITvOvPFT2lW6Awr0l9wAIMH
WFLJFaHW2/r6P/3qWfowSiGxNQRu5klXbwGGZ9B+4KIEv9LlAdsUzqkJkOjPQEeGDItUuAbCNV6F
xjNDGmdwpJfZtB4cEY4do+cnzQV+PA9cK8fwXhkGwOgL1Ml9Bbya+D7q+yQBiUqF+8bmHBiK8UTH
Wf+yvq5LOSED17memZoD4bTBHt0/NJN0s8vjfyAAAwB+J+IO21EDfOWdifCdwYBkXMhT3N2vtzRT
lIK75f77uFh7Zc51wAJDEweBb7hB0m+HiGlc3q1njgwvpLKJ4Izj9c6Jq+6Xk+UK6vyrcANFkZYh
xgrAaOvqKVpZKeLAhoQ9Wkv+2/JCcI2iQMTlYyCGD2+2or/Wzn22AcYlZ7KuJ+z7x/6ZylOf/5gc
I7l5+AWcF+rzOCOa6hpkQSWLipYNOHp6tE6HhP+aS86/BtUklsTOVatCpKEaqkDuBCzQDXwNqYMv
L8XU7wP3tGHKbH12KAtvKUMrpy/LWVljz0XURv8Cpxaf6wgaAcAAOLyuR2cm2dWZr4k5xVxo8pNa
errZBJGcj+Jfoc2TBBx/7+9T82rYl+4K+1fuytd0tlp/0uMx1A+5VY27ycgmJzFlTcta3sD7a/h3
pznFTB4JWloJCxJKI0u7YtNdNwXOESGI4v2bI6NLVUjrxp1c/QIQ9aDxWfqGXMyEdJXcKi5Hwkja
G9Ko3qE7BtEhfv07feQQ3K+D1tbHxJ7XuRVtSbV+CkEoQjPckSTscMnmhY1sbnNLZSrsGCODovht
o+9Cr1KbmIAwsWcLPh6/ovHmNPQPNFsx/hiVDtXhCuwJGrRysf8qgYTjh4hRH/ZEiXL1M18dXir/
Zp3aRBZ9kXb1WcZrMsU5gGFJ7jovhPye9Ve7c/aD+JSyvNXT7R//bN0438+J+sk9qJGk8l//oNCQ
l+kD31WiPw2b1IcAH8SVhVp5EfEg0GrLUgUANimjCGimbJemQQhb4lXZig0mh+0TJ4Nw+PFz/hAU
nR3FmJD9Sr855by3EARQ1Tj8Dm1kYSRTueQ8DrR1OMnfVhVvA63V4RD00vsFs+pQypow8EE+JA4+
PWdeIzhkCPRKFN0rkIC9gwx1O4iJ8j5QxdZO8hVrl0ob0c2beT45K4ziJ8j+JXofYPNj8Zr9RNt0
5F+IInAgDg5DtYNhpujj5eBuhFDoHAtSATuoi/JoSvkVmCW/5h6VegdURTTQzQ6xHFHM3nhEsW0B
6vmML3MlUK97hzchnPApjvOVwf6QIFH/M2U6GoZsLL72uB+l38yrHQeC8boGASy4vGfcDMTIfegX
uPXr7/5ANm+ElqZcf/kIPJpv4dcXfbPZdUoyo6vf4IoSmQ/sX4EQmD7+3rWQIDyupq8ocpOaAvA2
8YT8XPSJkeS0EDlDvPj7koyRUpnhE+CqtD8c+pBniak79MxmaNek8w2LWO9wRLcTlBNTJRNJRnWx
GznKgoCWogeEy1e1y4vZnbyl4utYETs75Pnea8gQOPISRt6YMATUMfwyjP9lB4f/aXBF5QXgltm9
RsOGOLK3DG4j/DMmOdcnYk45b1xHEv3bDR3t/d48DAON3fR2DOo4HscAG+xnZGcZ8Hq4c7Wl0Iye
x6BP+7Hqd9ACPk/Le6n8zC/zaQHtAoqfDoFvMSSgtk6fYKqLTIWQgjCnTpOPCqNstGYKN5CkyqAD
dE4YsKdjEW8L09V9e1MxYZZOwSc/lbv45dxGY5GSAepoPpHkiE/DkRyec9cfOUBnzAyG0+Etg+//
WErOHDxONwNw5VY4nRJMEd4SbmvUSZAsm/F8cOHIQyzYDQhzI5esTALB8IYR1BRN2yuQbj9USNZu
SqqGH19ouKt65gKIfpktzW9VFAQ7sWpKEDD+YIwAbXaLqkQvvNt0S42WBsZkEH7g9Qv9N3P2tShV
7JRZhtQU4Esft65dU+A0H4qMD7mMPNS15cywNiB9o39Sd08bNKI0yQzoupDxIMUx+8ilPQ1We15u
I7tbI3y40Ax3z7P3WIOGv0e9RQ0UNuxgF3NzYoVyjx/zFpPh+OrKWgZ/jDCOVozU1g4tG0VnewXx
A6gcZzzMSzGu8MdGhQqMvDMgWW+ztDYOvCrp0c3JxfbLq/koUmcLO4fSW2EoAMU5uqfRl0N90dQO
apNsiUn62x++RPoRAiuS8bgYiMjA3ax6oOOT7V29Svrxs9wDpO5keOOke8U2oilfaKpiOwNkX8gy
L+XCcPh4gviwJklaAdPFbB5NUvvDZVTl28duUx8emNsch9Y/rg4cYPhb6FdHRDCOpOy51sDJW7hz
hp/Zxmc/vb/Z9893DGqHSNRR+h478BBZgRNudzKkMUnEVzW4E3zmflAzG9c2FPefVoX6m2kWWyoS
8FlXBvpT688pPYs6q1fRl1RUTs55C2Lc9MlNP40Mk6HowyMo3OtddCteJJnFSjKZb2H9Vz1dQ++3
o/AdC+wvqe2qlp3IJ+fm/xqvbqdvNZuDPjufqHZVzqNIF8zn+Q+5p/DhcDAlFGVfuLOLOb65NEV6
Ew5HvTdat/vm3fLGvCM+X9vJCGD9MsO6HYd9kJOZKO2RghYIlqqA+5vuBjfeahqZc3QCFYJqQbWJ
+Pt59mUW0ViQdbTHCR/VS/BbSvoWoo3wyUKdE3c5Z8e6E0rOTHFIP8cmq0EIbDhiC2+bdfYdPbfn
7OGx1+Km45KV7DByNUybhswxYMbHIuyiP6XAtVN93NOSlTC39uMN2oonCr2HRgwuQYrkwd8DmrcI
2fVABdph0nARlqgwoYfQfr+eX3H3jeVYOxwG6esUAhqhlEVIJu24gDKGHm38OuetdSOg8e4mGUZw
HEk/gFYL/gG2F8O/4s7XJOkySTW/avoL30yYZBBUx+DMqHt76v3rgV6l9/eEU2L4xHwXaiIMR/ZY
UqS1ikusFSHTp5nLMwKfhuEIo5OzomkJjbDhFDKeqeitdOhVRFEqWzCF61TSwoJFkEnSq0/w1jB6
lMOq73y/qjAXC3atSh2vBi0ItgGnDaj6j01AiKxwzQW93ept33cjnMj7pRrIDZ96FGR34SvtZhPJ
ODuCAoPjj/4ZseyD03ypw/wV0JayW/xVbQZx6CfiB+z25Qnqlv9Muv+jkwA1c2AnvHznBVLioFgR
qjPo3Hh8D0uCAx77CuNmXjpwIAe4RX4KFeEalM5AfgOuhkJPXdHf6+/oPxHypXb539/srLPfBJE9
uHKD4q5GaQL1dACm23aG+cC/JDl/zwwm2UWXNAVkeODI5Szlw6+LiVZgCeSncwCjlKH46y7fc6A6
2UHx/Avxb3uxTLjhQAceWxthE7nSbfkplV4ZgDmLYfhk8UwbtR+6zI0mSMP+IOZQKgjFX8untjj8
vw3PuhNfbSPZ5loLHcpNWvQEAOsZYCPxHbMyfIaiAn77aSg8AyxAxlyzPnpBB3bwRYfHvcyNOae8
wFMzS+Cz2oBUI3AhFOuHnI2fTEFpV6z6q2nwVlmZIRFuctTXhxaMXSpshyfTWkPp6h6nPrLLuPW8
Igy4hYoZZzz0MaCP1MrCj2V9DhxAzExL52ybA5UBHWvql9vxgUNNxcs2ZQ7xSwJ5h5cJ015VQDNs
X8nLF1ff/cEixpxNxdryHOXpsP7QEeethrBlRab/8BJg9X0IhExKFcIdi+a5WCAj36gkI4cOqQVu
i7QHcRYZiWZvbrKT4HPk4hSaVY5zeDxwt7PHLeEFHwKo0An4Zdt3v8P8o1Q24GGcagPxJsYfM9Ac
NeshC9ivSuFcKbgBwnGTZ3C63t3VZbhc2+WG6wE5h7bGPrxLbkF4Jtq7DhhRigobtoA7UIYFghtN
6i8uoymzWk0eWmKHgHnni8dirfvNTFGI0uF/hWZzUPhOw3Dvengbhgi3yqlER1s922UoiTiLqR+c
1fHVCsVzr2iF04R3DTQfActqmxk/NQ0N17yZPXS25SOHSETymAIvJQW9hyaHgUlYfQC/1O4CXP90
C/xueYxeQpubPwQ7Oz3iqjeamxuBSqeq26S3/oKkEyU2/zG5Rgj80sPJk6oI2CaIqZ/KzTJ8I/gX
tf7HSkpVP4Lt6kuCTY/s3nK+FYkP9ZmZ31jsrJEjOQFuK1in1v/fthwS0xo/oaTPVPSxfmpJsqJg
5yds+9pJrJrUSZAgJ+mwh6xi/QRNz/ZIGM8mrcTAiiAtV4g18E1PqcTvFvfp96Co13UzwCBFl9t0
SWfio321+ds+6S3Ic9V412sNwcsA8xee3dqB7QLpQETCfqRmwnnVz6p0ox5VAXhhg1MUzSZxjlii
VUe9JXp8bzTFRQs3Pcbg1trYJRPrxwT2DPtCBcUMkqucvv03ajloAcTgk5BUjvFLHyM+VIieR9yX
/DS6N9cXmMZzIaaUY9b9ya7zzgTXExwmQvdxm/LkQsUblnixoXTuxY5M39MDnhTxpIrgmGiYB1eQ
dc10WGRxBbSywJS8movckgdHGTiaPHnpy257FWWoNFbCU/ulT7D+qVaYFYAl7rBtzwg2EwjyJ+1O
4zTxT6VwbJhzFnhFhj+G0IFwpoJVabsxIiSJx19MLwBi9u1Rq1jE31OuMKn4X5nzCThuk4R7LXil
dhBcS8VLC9Sw/Yq1mANRYhk0ucgWjxP8X7yE5NyvA5+CXJOnQ7drpKiF6lza2heFWVKS9GZFTyZX
3T9pWQtzaVVcact/+arBRB+2ZKWdo/2xU8YmyFUB/Jkkgn3LDqstrFaOKaHlkNWk+c12+FedTPe2
D1a+llg80EoxY+n7zM46IwetGnUiCSHVPUNWdkr88X8n/tj7rLMzOlEL3+FXpja4Y/eAD964foop
tItww2BHlIq9oO7DLDrb/JyVXaQ5pvCsMVMykTqyXY3em8Ln6xeVvsQp/Vp8VDpSO2OcdwT/+lUf
PkJ8AiEHwXrqgnsGBG0uInQR63NLMXmQWtY8XexbPHmr490m4E8J/P3n0S36EwAA8f/cN9PJzzIS
LU1Zu6jIxEL4qJtrGeunEARpTyPr6CU1qJBJh0YsHZUdlTQpdrU2SW9kElggHGB8GXxRz3JFl/AN
GdeNL5HhThe58Xv3UWoX5pJ+KnRaFcCfTBn3nDPHsnVcQ3SDP9GM6ZOgIBNdOQUt7KTKzlWKjeTJ
xbhjb4z8Y3FBT9b0uHSDzCxZJB9HpFJmKWFgingjofyzCF35wt1/nTn1thn7D2RdqO7QYJDmOiL6
yEQupD12dxqsCj/4uNV7/0AFJWlFpZ7VSsCAp/myvZPOKDbqxCHwTth1uDm7tQW8jWrvdoHKmvre
YWiXOu9JU0zqHpzATk5tJncTGFOiYo1Y991bgncpECkI0uDdxJuttxgz30hu99eBM+eYxtBmEGlv
S306+vBXdezAy+iP3NXyzK1orh0OjJFVd25K9xYnckQs/UhhFfASvhmBLsFJyrQY/rY8XMWR4NIA
+mXCKbeZOLBq+ajekX1y5b4UiTk4uPGmcd1ICaXKDhAmnDaGuxFXestb/PVxBzVYSgruW3YOObbr
o2UGxlkn7XP9yezio5SG1ASfHDMtOguXChLLSuy0OXr38ohvbRzA4/gX8sHBBgpisV/VKGkiv4WA
b6A+xGU4SL0i2h31n3Wz2JTLb/c+JYpTACBfKvAaCALUhM1WK896Edc/XS9CR6CfsGS5ozpTDnLn
3xT1/LjsS7nLR/5PPEyC+G7lhq8PrFPzN3RrIbVcQi6KY/l+bq3SYxStr8iDiEPNId4FLf6LKoJr
Cqsau2pR85sddGIKEBKaoD4yEZBtC+M2rnXXMEWzBVOCI+qJB0W0FQgXCTvZNfp1RmGkYVIDzhVX
GqjI7IwYiTmwmkBclg2PgdtmedrkoPiWt/BXqH3l69wbvW7NVXx5rKIXMXmCGKSC8pKz76I+pB/u
SthBHlMC3zxqJL3GHGA/yRHPTDbgZvtTfib1sAGL7ynUIJg8rb2tPYFYTimkXVeQ6a3/TzbuA8P/
BKBsLa5nAMiPyCMMXcJw1QMdsblPVIp4qzqfDAJVuJHiGAUwb7tfPDpSXDWSzsWhYeIQBczzhNe4
8tV2bU7uZ6Xy8y+XHA4Oy//LPFMtNZlGJirlLiePDSHL2D68owkFLW1AyvJ99ZjblHRlXnGNUa/T
VB+wK1+k1oKTYaQwTNMhGTYSKmwGgH3TaqR/Gh3attfT/7qoPRUt/EgDFFQR48Ugiax0NSLvgYQI
L9zVHTFOjyw/AT32NT48EYrZhTzq/t9CSvLHLVy+q9MEU9JkKoLXmx5pE03NfLpi+b5cTZrjFEWG
6cMUtxcU3m91vISsn8UOjAGeEDRhKxYTcGWM4MEn9lmdP4K3puza06yvhcXTIV9kdpNDy30IaNoA
YzmbMOEECvW06stJUTau6aVDILWS3d6bs2gihh/7jEVx6iOfiC/U6pvt9TIyCJhzaGHLSMxkzFIU
7KyvmVFyfPkiY2OECzKo1x9ipl+1IUbBv0UlMCPMAPPPN8e+uUqo8YxISR4uVCSZyPIoXecD7jIz
HJZ6Wp7OTzpzgs+RYBrvZtj68Q+wfjxjmgS6y/SzrWHdIXrxG+cptf2bl2/lgfBeZSDRGn/+s06S
l3L+X8XUnz7L84CDhjCkLAfTxIjT7Sti+t8aHae7s95P/Rjlmgs6WRe2li2y3cbNhodcGTt47rWC
NBid7OFdnw67Y36NndGMnJP4QM0vW/RxBK9LvvqH/5ijB9QQZqyGjWbMYGgbQKqANONhXzX3Utpj
BT1QYG9jXwyKFYw/Uy7+VZBG58g9UZMEOWnORdUApWz8991X7eXIzaTW3AuhMTXQiNzSNv7cMEA2
wo7hEb+pCgykWaAea9XdCEws5zvE1Ln1OyHiEdMFlviUeDefjD7UCHnpzaxcDXdNpgZl6ImpCKWH
yzcArgdWYUqiOGWW2yRRYEabzLF1GtQRuyZR43/iAz9z/p692mHgFylkrrQrcoQwyPSeitPt6NPh
TKIfQaYoer0xT/yNyDLWOrC2DGnFp75ItvhQ3+qNxcl62ESXdfq3+IvSFbLBaPEksu0wY13LSgj6
OOZ9pAAC5j74zVbaaOXUYL4u+g/5ngF3psanB+Vir7elYovHNGVJ4wE7q2/0vw3KI3mzjxZnAxok
fXoaqQ5ihcHBIFc+KtoKiADmE8M93xSVDCrxMR19VPCl6jY0BUYy26o1zjiITw1qH3HnNDZiETsL
sOGXhlS09onUgsjPvKZ5+Ojr8EiaSz3Tm0gB2iB+S7AT4RPyUl4Va3C7QwJYTtjCnKCPWjfpyOpE
YQBqeNLWEFZEjbVVpen1beScIOZvZIniTDQu5rbCgaxFjjJclcZ6wt1w6gDcIIw7cawPizaRTEgw
LViqBIWoz9jIw6krxmjG2QliUKLObxIn3GptqWIWBusBCIH2kNFiS64aLgO9MQDdv3eS5g0Da9Yp
L99iB3knSX91q+ktcRfM8qvJHa6NHRCiww8Wlf1lvppO3GfWOPpnnepRW8So4P7mXXXXZeKL8hyy
5escljjay0LMd9Fog8XkEiQVG3Obu4O0l8Hz1km3XV9ljJ66iFFNfiMCpf8ZW+k0NSDzdhdWuLCf
MyFiK2AwdEyagm1bNjm6xpLRJOxgx8ipwzXuZYWs+gY6Fn6KPOz1vl8aKVCF392bjKy8iyRi5nJK
c4t/8+QcCI5Oh9uM/ZrZDYQEQWnr1gA4NCgD+A38/xukbbvx58CPbU41X/3FdgHSTiJZ3rwVlilW
08JeCuG9gAfT9yne1SJCFIjr21uzvyZh3e2HNkB639+b/JoBrxnZR0tkOt+NlShH6kL64GlOIsGQ
+STVWOW5nC36LTScX+53jJgpEKPHItJZ2oKwKEkYAHk10j9oX0fRHSjJLRsVL2T5Qcl+zGYFwAv4
2TV5EA6BKJl5JikogyyEpuMbPyzyUQZmngaFLC1ciDc7oOBAXppuEYeP6Whl0ca4fdqvLGsjTTbZ
3tVqo2tMREPgnkm8N5lQCzBxLv2x6Gj2DLWANxQUdRZTk7LMnPJz+9pRuOmdtqr4FAA7WQAZjBWa
8oxYAJ/bM02t0ihU1fGcAZRbqBSJOoynuOwVfWzKw54Nbg5kOXa8KNfr1uPlH9Ils19y1B0jx+Jh
LXynYAXGCW7RqnQrdj3FqJW3NRrwL4XKalDoCvaK56O14nWHpwESOsol/r1qjKKJNNp6ACSh52SN
9J3vAiZrrsBZXHbaiu8+R8hl28QObmqFpursbnXH47co4o2hz3hYHxXRkDc0LO851xnz/wP5Ruqn
Yf5850ZemoNpR7D1BxQnngTLgbKbUOFhspU0ZNd9FRSoniy2H7UilVZwT2qZy85ZI1V/QkWUUjDP
O/MKOAeR+Tr+XQ4N8kYZEjYu7Qoa6KsGOQCJiItQvPsMmMD2toSof0YH3qLUUAaOlU5oKpEUGk7R
CiHOC8NsOp5iy3Cht89uOnlHF6LzE+qSpJzQdaMnnLeehxLAs/QRFT0t+zixHL5gnlXY4+udGfOS
l2yUX25iuxpnER9nOlEuN9AyPAAz0bc+rMq63Y9vKgQTOs5qRLmRS61VPA3M0A+tKyvHPr9UVVzg
xZKLk102gkse0fIA+Q2MSuuAs8Zlnm90nbwcYl3vWrlosHLrgIjTh5tWjm/1oyVH2xmA/UWpj4xN
6WkJ5LPbrp4JBfNBtN/PxbT+4PpIO0C1slFv1MSK44iz88SZB0HCRM6SiaKPyPHMzF6dyvtd4elw
KYlbtMSmu3z6FHiLpOV6F+m7lmag3mvL/O7I7Lh/vmjGP0wPirPhPbx7CGZ724+KmAbzUsRq2ioR
jSpI72+zrYmpSbSI9P00vUP2n+Bb5tZQIBEEXpj9co7ijXHZ5Foeuk0Dv54MBHVWjbMpahBUmp9e
idRZ3+WXMLe6oU+Z5ddj2MKFnDsxuMLEpaRcKzbr59ZCRmJM3f0VqdW+4gkSWX2s+O2zvzqL3goS
dok86tl3NhOfLilEPCer7KBb7Ac54O3j3js+zzFpmXVirQwUdOkgVl8IDb6WrVHUUX690sgYHHmx
GSP+VQZzxMRAzD9eGnWhgoSbiezpnLjPc760QFnP6aC3XNXvtW22ADw7+rjZzS3KoFjfEVto97AB
HGvmA8EkA/gw130KksXazrdW3SwBIHS9w6S1ciScTj2zZX165Mx3oY6iOpZIX37nQ4ACP0GWzeMM
T92KsuyotShx17/aZFKcCPWpw2d2xwMN4u2YyHK2RuhAkDy1HMmEiEORm2WXItilNwmG8p4BxDjQ
kZMIEEtHX0z1t+DdiRE/XVCW746oYiD5VdI/uhiuxRk86AKIxZWDEpPu9ZBPyxTdJ4D+sN0LoMPH
ycNxBWWEU2VC
`protect end_protected
