`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OrfJfJKbMEd8Pz3wlara/ZLrdZVMve16qt1GIFknOlfDZsETzc0jiPb2ZLN+bj/6/1lGo8p/uhPS
bugTtI5qAw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mODUmGnb8dY9RkGR7yX+wQMxn0ZVsP+CDypyDkIFtyFAd3tOU/9vvLtksCfoC28ulWlZ4lheBqTW
w/7PxZ5QQhWvMyl5mQ4N5P485hO442Rn4vKqEqIA6HILubWoFpxv4hHLTqu3nUnsxddaiNU79itX
pVElWXOSf1gMFNRT53U=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qh0ZvVh/hOQ3NVABeb+kjiIdTFOU4ClKHoxogmvzoyN4RBFavosirS7FUNU/atCx+Kj90jXXYIUH
MpnNrlU3xC+YRGKYN6CzD8DcVhRpvCTwk0wlG2hAZ8aGNn0IAM1C0psKsjz9yMuW1qilK9FUHcJ0
zIoDJmW9VThaC9wTWhjTSINYt6i5QKNyqlpxvL1H3TevmeFl/c1Y4AHrhnbFQahfp9WJWwEKnYf/
2cpAg24s8PdcyMVNvveBDj/MWBhJGpjdSqY06d4FS3guG20Oo3B21DN9lNLNR7t7j8b81ax4z7bv
XhjzxiiC7zYXtjJJ+/Xf/5ahn7lnSw3fyPP+TA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tqfcsGy21Lp855i+j0HO0i6g+NbhHVyptUTYghVHzQ6R5Auiy5R6+crkoXmSPLXlITNBy7ELLX52
vOhO/ci3acy9JVPvusljHrdjAv1M8ZoAWiOwY1aUrBZLNXwyw3HLtHZLEtbUlFNnvKFac+OyPpSP
Xq5FUyQsXsSVOw0kAHs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NvTo34x1/KFmah7dBwY1nJ20AmzBmvTK1RtNCB29pD30E+wWZ25Nktkp8A5SDpSaxwqw88Oo1qsL
aEL6xWopNVPPUR47PRwqSbj+jSoVaW+hdDZSqABxlcLnO2xazsrsNtZOZRfp7OSxUF/+XWecNbmR
d5R3h+20kGEML/ALMNFyPtWijPhCYQiLuGDlQFSuAIk4+ettG3bMc8cBHMHRU3QPTBPuUfKbLyBd
Bz00lvR2XP6aNVsl7d07Cw3iHhUgMKjuARwfTEyeU+BWjz9ojRB2LpqFcIM4fa9CFhjvWnRN//0t
JZuldPMn3VPxQxj1ZuOVpfDdQBcr+jSm/k8pgg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14816)
`protect data_block
Hr4np4Vv7JQro3a6CUkbXWAaEBIMWGJZVmvYztds8gkeKmxqrF+i/chgSilpZQmpMKC/T7rkRAhC
DOzejRpCMbSCPQ/COnK1EvnLpEidRk1rFgTrdKZzF18QTlzt7QjslUhpVXTQC9Ct17KASr7USWEN
dU882FjyGT/m8F66Xf501Ha4cGGiohYjLhweEnJtZ9X62XiHn3D2j/6+Qy9YNTFmT7vNIEOCX04L
T6UD4b7vbQIDVcr9q9jGXPAVmWhUEiHZZ/g+1c9u9Kl5Ei1YVEqDDfbiLlbhmBI2BYAYdbkeeD0J
CpM4oIeCEGC1un+1ao9uOWPOiQdQSzhj036rAX/x1OY14FzBlewzz0IRhYZYgZ9+OmA3x/3N+WkZ
2yqwrFRwM7/ZpVPBpO+iaduso+I1bzK1CrVdxotzEf/iq/pJqkhfFHSnSl+mdhoSVci+dIS2hopY
Sc38PvpMx5B1wLyQFpk1RATlQ0fXQSkrPWRR5sqHpR6YnNjG36nLT4a+D85g7uIIew32Z3xvAVeh
cAAdb+YqWQ7E3psOIda5Cx7pc3Nvzw4A2DMlewZwop5Xbzhh3Z5gLh/w3UvjUrMCK3sRNRbhnqUk
euNMpH4ZDrDehynK/yhnLm9tJkWnfFha0VNjoMurRK3MotjfMLjbtEREgs08abYb6OZkClnfUkve
uOEOHsDj28OOEvmrtKzvF7Ih0NxKNunZTH1m2T9i4JN5TwjzMRRpBWnZZKdvQQd2NbBiDdJCyFqQ
NSSqTfNSVRs2CoJYCXcway/ydMXRl+LW7uovuv5tdNI/qJiYO6q1Jb+cqmXK3ZifEPsBqSUm2h8e
/6lwMvsP7pU9aH7XZeA3eoVB9C/KrilB++wCZQz/bflDyCfXwtfFRUswULPzpScnf0nZOs5gddYf
+74Z9SQf/tXr+xpLACHl3N4g9N87lCYWvZiQtlLIpHCkt6bEuzTwst6Gy24DlPeqEzDn6wK7w5JT
4U7IZeRqc92wFjVwNFgFd34y7FEPVpX7dVD5S3YWoHi1BGgIIjz97XPWJfx5uaxlMwulwlPCPe90
Itix/YD20vOcRJmVfYSXZCnbxUH9msOD3rNaXTQsyoKObVFGIu5hbHg39vUBZXBALoNxVvgBRtZ2
Baz+ZiL+H/yR6UHyeVp6QmuYJPWYn+JBa3fdDJr8uLAOicHBo47DCZ/6IeI0aVuT0aDEEukoMH4n
HFopdgkiJSNwFgEoVKpoquehd+a0t+VlbeX+wGSmhAn7PbahzHoTBizQYg3XpbQYkoidkm6mvOvR
0mIG1wbtTke0w2xm5qh8P8w+UAxcDGZkuj7GqnMcmdWo0owOwGfjXYNojIQ2a6pINOPERif3x4Uw
mV/iCMu/CLFqzKZszpOx5x4rscYDrwryUMA7tq928j/gkW5dnwE7/nW0oorLWDOUhOhWYIq/oZLB
Xvih5bCQSD2MVRbd9rY4wS+/VZb3hghW/IH3SNyApl7kHQALfyerfSd6emgNcmVE1OVXpnuoE4c8
URueHe0Vx86QSwbeZ2bBBnIN+jMxYNKybTp2urYrNYwMRekzLeHI6qtAd4RDwaXZCYm/KdLeTPXN
V3C/MjrP+lL+ZHK95f2VcnGeg9l2u5sKiAwk8EJY0MKinE27rN04WDZScDauErIkrE+mqqr6rgLg
1Fr8fMMFaKZBFkNNUDGok7bOVl4Q3YtVXoX+17wyBdlaVyZdVKtNSPn+Weo4+uAjnCeYjpH5ZRIP
SnZO1raeVjgcNlkdnbJR/OvbklTceJPzJwRcl16nTPT12iJOQ703Kibq0Rs0OveFAtvUmdlbrUJh
yQjAovs1POxIOjgBlwj31pswJ1m7scLniFZTpE4UpVEk6GGQI1OPVyYx63IHRzlGiVw+PKblSszL
edt31Zx8JGWH6BdndUhxY2XMG47uNQgY1sv+nw2XNJllID1eBrm3A32oldyFCXFQeTvl069EgwmK
9CKyjVCDDmqq0mIz9uSDtz+XMtUS/aMr6CDERK3SK4xWxBqshM1d2Ew8wIhxzuOmTDrmETo+7PSf
Ncu3CfT0fhPOjAFhylYAO38rR6y8RIWYypOyHPcBCe+ZmhULKpzBnu99OO85iaphGPIqtsWBLlvJ
7R4+NK+PL5vc7pMG1/Q9kguH3BGxkh5izpAhBe4S4/jXkrCU7orSrvnnq+y/yIzMuoYOwLZ8vREk
rBC1BCTo3HlgBucsIrDV7v6xdtcJAEfNHas6gg36xFD+Kpb/M1MH1OXjzumWr2kaRDwFMPPvLSME
ZHcUMQtZloJw2PXyNZMuv/tf3CQJ5hHrhjR5Ob5TMkzFlZHJgY1BTL9mpE0tdV4VSQK4YwCv02ph
7Ru8Z4kBJ1av1Nv5S3IA3Xj0uekmK1aZjzNfSxYz5r/P5RhiljSdXfyEehSOYDjvSLfzj0QoFcup
BoFTNlBc8YhJC3aW4LTJ3TkGLo/V+l/paDHwCwjrLfGqxc+G2tzNSEqVFLZpaFMsUp8T91P/XhRg
vxusIy43+a0MYLM2n5wjt0I6Y97p9TAP4yBSlRFM2xJ+5IUfe2R4hckEq8emQowrmlMb7PY52aSj
4WgntWVtTw1+v+Rz4BjCEkec0/6cnpQeciGMDZ6Z0jFTQoLLJ+EyxBO169SUxA8Ypcqdotkqh1cR
oY4FopgjyMsri0dHZEjhFRIq1qybE1KuhW1WOhQ/ljQPljYpHduAFEHn5j41m+TcWtG5CbLzHBJ5
kGO/9fi5hXGvY8Wfb5K6dnDIWfZl/M+rE3a3EN+LHyayBx7Yx/ei693UMFX3LayTKb1NAsMD+71r
yZ4/lVeVtiUo3XgdrFh+/ctSrKds0JGcovUi8Yh8VNj55fT5O5PQl55TgVcJPbmBc8TNTlj3a6fN
UDpzfIrvlQQYpJKqGuQlM4rotJaJaZCGGtRwYEJkBotrUI3Fz8CcSPRyoVcYudrv5hFI0RwC4QBZ
evICCXPSgeRcUseT0VrAby+mimLBSTM9FaUSNrt4tsg0x8AA+EzzL53go4dQ4KQ2fYBcHh9aFtuB
vU3xQop2W9l8a3BfNws3xUdXXYehAr4uFxa35tf+HcGjNxPvre1GQi3wdXHYJNniPgKT5/AKY+d0
5FJXeKVwkoGt3Y7QZ1tWsF1rC6Pu+nH0uqoE1Bpo2XZQqq+ueOFQQIU91/JPIZBWk9ptCR0caZVF
oaWm+O2QIPnSA4/Xp6juHx42Rl0TjPiJa8xq+ZW/RWnIU0uK8VEyxlkHnUuven7BPRlXNaC2lMML
awe4rxoUUu5Nxd9KhuHxO5N+FkqZnpYK7toc9QAAdSjdOimObkZLrEQJyvISJMAK2noo5D4zuX48
g2YIHcP1z3gdxcGv75cDP8ukVdZI50FTmpr4qnEBArASOydOxewpk6JZysSAI50AimnWWXH8mkJx
Rp6BwDFSe+uhCIZm1w1u/0TRzWOUpcZGt/ZyNKt1vMcBn/Ycyt8mVIB3IRm0IpKcdcbLo7XW4+Vo
q0l+caLg1nk3OWzVUHNjECe53o6SsRSVzJxA1btBT0Lrc0ihy8Z8Htbu5myUSbBqjyIgkCnpUKz2
aGERnngdc3jUhxaSIPIGrijg8FrCAAi7xjNAmadO7vUmSuz/hs5VYZvtc9rFbr3WaZyOvQiPo0Im
xpcuOb00CwuZsWr0gfc43kifgaK/K1Zh+eO30F6OBGEdxDU3GN4dgLwdG5ZtXmmMVISULZS72rgY
4RBmfuU9CNFTY1KxW8OHcbWgpM3vOlDiDknaN+Mlb/alPhvkVuCG9C78V9rJm2IaH03DMMVLGP1t
WIrHv+XZiF/xCyaupnWkgvFzMm/nUtEk6aAXsuv2uxnKfJf+wFMIRAQQkkLV9pNQzK3ff+hxOoCt
ROi/lcwnZOE0RNMzvzxPernbXJNjbDWRwX/oK36/VtMVHj3VXRtLyk6v1dFynmDbRcj87iPmK1sB
B/Oo4eEG4C4FbUjq3vnJHrdLv7dbqlS7WLNZn1ZOYLcMTQMLY9mkugdxzswzJMYdBUNyDB4dPfmy
/hglgJ/ad3a264ogKK3CgMl5nQAA6LGZlBYOZX4SGa36NFM1oeqHS18r+IG9xWuiD2/8Tv9UVMJx
hDBzHtxOhvpLaIRa4FYj3YQib3r/s4OLEYx5YTKVNneK7h2LTReJ4YWD7A1X0WAFy/WHD9107YyW
m1qo0/SnRjg7NjN+J5tlZGar30vpqh3i+Bmiun7BaqopVEtwvIsGhDHwEt6rWpAos5ar4E8Q6r23
Y6PstV05lDirnBHDCxbVa5tmKZOLq0SvSbVnYKvn87EmGV3dGUKk0TuhXVHPQtwLMnGzLpvTwsRH
l3XJdfyI6qIH/0qnCKPnEIdbTBF2T8ZI1+ojcto2QX4paIo2H8A3y9IKda1Asse4qqiNVYaKNDXN
zaZhnsUyfEz1RsJYruOULFptfon7Nr8RwLGRUo0mf3EcLHUQApeCwzFN7uJQQDRe/Bm6oTkcL4fQ
B5cq0XonglBnrloHBMbn4XqJNa8jhU4Y2b3EpIvwajiqH3wheGH14/7tbrUyIA0Rjpebg//E0Ebp
X6cg+HAS9rL1v/Dr6Ths5fJsXnxxXV/sMUEFcPxlGQD4aj7NPt+27yxdubaJq06Pc3ZZeEedc8VQ
2qMu23qtYEgQVTriuF36r3HsY1/qktLugPUIHYts7+kewLbNbCR5Z7DKMhk42jc/CPEmyEt9WR9D
sXJTrYvNnsxHdRkNaBVtUvOn+zT70rxtXdfVYtSY/ctUNpLjyWarxclPx5++V6qqVGVD6Mevbt0E
vp4R3ZCU1hJyp6Z1IyfsJ8YbJa635sOl5oS4GErYbyjJmoCEcK6XdqdbuBGj6FhtwLr0GmLWKDzU
8jOTup7d9GJw53Zq65YVfd2iRgoN2SY3ZL+tRePHu6Xy8LY0qJA+4XWcTjhI9MJRxOHW+kTbVhsq
Yp3/B1LNhDN4wiflhWXkRabGtknNi291l3jBH2JuDE30wQyODwfSNfcl5FZ8zOSN8uqdYjwaicmR
Y4hgOXkB8Zdw3HZmD3GqbISEep48+lbspYrL69oMH3Vxj3dENsYLGeVpa28OBRIwCgdZIY9meegT
z79+5OhHiW2TZNg78cQk0N9ytPeZbI8uaenRZ/aMI4fZaHTp8KEeBT1tPNAGurODVWL2xdXGl2Fd
rbbPoJHoJl6C/6LO8BoEt0SMAkmSSAt+gihKbYz3gG1trJI6CbrXOJY9ZbDK/1o+MX+CmeWZot6p
CktNCP7CjeBqhZjkmCUXybdHXF2j50uc/GwUsXsg2x7L3Ll7fdIOo85N00Ok7geQy0/wySceknEj
gLEzT1C6eEtKx8MN5+jjDlltIeb5L8+mrCAH5XUcCwqDvLbPqdTkDRomxPKQBh05hrRxU1dmMPZR
73jfRktTI6yipi0Y/NFCM5Cyy3B+ZBmT2jsbzCWEXqDTl3YMlEbGgSZix+GBkb65SbtT5pogJ99a
xTboGmiPDa9KtcNnlWSnEwik9gIVrYH3K23GnB9DiMwg9mXOurmn7n3d9m+W/gWFWHHGFkYFqcfZ
MMk5CCvlj/B+JFi12qVJXFM2pIRpT/DU09ljBj41GW10hfNFXr7y27V9E//CSinstjr/dbsFxOKt
/6N3V671qXe7zfhO9lAhLywhDHF1KC3MDrkcWc98etFyMsqN4Sr+tJ7f8l3pkDJY3icprOHyfI40
xVk341FJt0TA+D/M00ylALaJuoJnAVY9IgP7aewLCbZ6Jx0b0YEGE0+ygxPcAIasvbtWgx7BJ+7w
poBZqNWtflQ2TYnR54VXGp1xy5mo1c7UbJp97Ceu0/WHcz90xWqGF49wgV3yW7qlBZcydKPVuQGJ
rQGRO5iq6kW24oHKCKCDqiYfZcZrDA2dHXcMBfZqmHVvDpEfQMLmQxp8EjsLy9dP9RnaWn9K+R0M
d6GW/EH/brvhwKu98424ah6PvjtXWukK6LZSq7d6U42+RVf97YpX9Kvi4kBpQYYZQugoijI96hZN
FECg1Bp8pHIzyH6dxmTflOsbeYAgqs4VUGxbMhyXDeg+yKGRoP/8w2arrAFHNyUsVe4V9JcFcrRC
st6fcWwof0EjG0dlUbyjb7M/51P/dd7fFWUzgOF+Jkwb8dCC8GpFupmbt/d+0bcDZoQP8EUb4eiM
SY07ILIKBGlHlbdnL87eEZJKDn9TAkiqt4PbunHtWrSZBynDpKDEI4HrM+SMuPV9+LOhVk4S/n43
PRT7ISCIyCeipI05OorSo/bbToAHDnkCL1XKzcDCNrwaxVUaXyzJFgf/MLhFXIg/Z/sf2u+QxBG7
CnHsjK2f9y/5bWU/nX9+vpJwvpCB+zN8II1hQL4qzComgCK8c8rrdxRAaxHa/oDsCqIExy/w995Q
2Lz6bHlDrvS4j0+Ak5Y+R9sTtvEU4hB98sKF+WPlEiRMMStZWSCqkAMWsPKfrtuHBHRX4SugRMXD
SHm9anxXz4AoHqOlrCsWz1i7aNbg6RQ/JSFQzPAHD+RkV0zQisacJGgLC7rqJUUqEiCTsA0CZ0TF
64tHcIXjwuH+nU6Q1po0UeRK4LTb3zERX0KhBoczcvlSltNk3lpdKMt3+5XLhMyr3ftP+V4G0XrR
92zoikK9cU3xXz/3YGSv6c0CegDSiGyw0EQLd1B2La3igbtSDs8kYniWxKL0GWercurwxPBD5Ea4
Pi5IRyYUnfdidkKlSfdRT2uvvMT000nw6etc89/jiTkv2fwcOVz65HrmrVVkpgIMETQjEILGEweB
a1SWHjBZ8mOgU2XhCWT7IqGHOBGh4zT7kYhxRqoQn059uQNEsQSsjnzzJAb1J37kK/qY/eCXjUSP
4nlw31eoL4o4rFhiGQLtB7HqT/KZ8fKBtyQnU6aMfqALVaxlBkadVrFvteuXpsSO4klZ6Hpz5Iai
foCQV9mYKL/8ekMTEc4VgPkyqqZuBqIQLUOfCJFHYdUCOmxIZ6G6sFmdVBoyvoMQpsIMtQDoAU+/
G22b9SMrYgaCTGLkLDH7hFm0tftL7HRq/e103MJeWl4x3TVyhqqbhP5nMNnaZy6N9M2547/skTl9
v5/7WeHI3zKwqKEJhvjGSM9IcjZUFUVm9/1N9IiRkKrRhRZdmupvzgEsoM5PLK9oSa1VcgXo4RqH
HZlJsv0IkSZkePnJF6HXmIMCpUcs3VvUefwc6NnOsZOHEpG2V11JBM1AkvEOPAyPPMiHhYCR6Lfz
KrwW+8U3vhknP8buhtvIidHftj1nrOdVv6+1S1bZwYmAvzLD3NR0KUKeAbH8P5cYQNsj1ikWNfm8
/eMSxxuVXRNOWdcX9xAL76YXKscEbM2MCkJG6BJrHP8Q2iGJqIMulvnbb+prBaxsoPVEnNdpWi/o
v+tKKfjIzZSfPX4IXdxl/JARP4ikgY1LrjqhcwsIUWic4C7IQGnQ+oy30cdBBDIe85fQecBHRP05
gVKNZdvdZTUt14MCfteH6810Ud2JPb9+Iv4VEheoangsLHhR/x5HJVvuu9t2WNw72TWDkNMYDxJi
8dSw5te8PdMOS2retsJ8UA9jST0BZijoR+VrphXUFQhEGMpNqGDdZTImvuYLniDUdS/9AJhknkFO
SIoRVE+5Dj8VPE2iEMerW2pgRm1JwDEwWJshWxCCUaBrhx03HrK3GEyIsEJBdgUrLNs9ZnbwLoud
BidIa/5pGlToE9jFVm8KztQEaNzVBdJwPUP2xXgxNebULEpZKM08DFtvNddoREWeI7/YGC+Lay2/
tO0fvadgSfTc6VlcfSA0LO1+Rc1AQyl2ufzQKA+hfqbjGM/p65x0MO4oO59qVNUaBlOa/k6fUIkY
0aV8X07Ggy6i5xD9xUSEGX5MxPKbGDXgKfzWx4XB4zwhAA1gtzpIH8X4d2ChjKGcFxVcn5K4ASwX
FddNrKsGOENv/I+Y7MD8mTEzidcWRO+0sJjHKh0G1uOKKfJGdWDZqVzOB7Hd7meRHjCj8hfCZeLA
YVkZj5iOa1qJiSQnGaetqmzZX8JmOOrjHTr1c+Tp/RyBYRBtDoqbD7NxA+iNU2K94WKlmiQozrJd
OeHiDBsqFty8SS0q+mWAA0GzFfU97PWsSZGe2A5RD9agGTiAHf4OqtKg9ZhAH3XBzsmqIzE5rQDo
RTmxeU2Q7lX7SaO8iFS9CfoAr9zB5+Qk6E76jAmiDXSTV+lqt6qjtphDp6SS7iD5dwjYC/+4/O0O
LtuRIyLYgU/4Y1OQdLrasRmihEhueE4YHu0ycRzx307JwKAW/QCuVEFHynVp/OF+hvZL1yyWHGQ4
i3WpYMZQvVL55QQFVMnO2yvLFNigtxZnoH9WoMdofXXRIbM3muUc9+JL56qRfoykndYuAnlK2/Qr
yS+4B0qlmXCnyO62VUlQ/20C2OVFabDgkG/uOjO9FyFKvxIAVDrvb146fezgm6UAMFPuh3PBQdWV
FS/LZyVMXTaTl8FIIT+TOQLO8/w7WqLVpCla8+GyDTcs6cunJZ9bBI+AptyYUvGnfk3rCc0b8HoD
i2DS/tnadAc49Ao3f5kIyeobRS5YuxyNF0u0iczXfyEDiDRyPhrVEhm1XhxKBAk+zF0V9KKoisF6
dbbiwOAnDGVc03RqmLELnHPtKojEDccd+VfHy9XPDY7060GLBt3cqwP2gYzVF5UxK8152/In621v
uMrHMSlrxXrN4aH9q5XavzMOGuGN5sYw7zAnYByf4Z4WxF7auYLrSk4cQPtjxhazD9HniYAsBL32
weCC3wyBHpLr5yf1XlvMzibbyZFTjk9Mopx5rdBwuMlApozvPb+OmA2UsnpySJCtNnNnBPJbrZeY
kurea4dP5vpUhvZw/wK20FIKZV8yle/jLpQ+iyOopjZfsE08JvifNehiUIDQdzjJxuiBQk0PkER2
vFwv23uyGm6fN+tr9Qgss31WuWeepvJhInfAPgkqakZkxknubxs0XWvtz9W2BjNfsV7yni9m6dDn
RhPxg2iTmmk4HoOrN8vw+rCgzkw0Vt5P17GC8XB4Xfnmd6M35f7MfIkr0K3OFitldVwemGy7s87R
NpNLRYgibEUgPlrf4cj9MbVlTZrAjSVpsACFLsECFV8bkjoN2PnMA99MJIItWP45pBHLl0fjEHnY
07Ghn8OVxTic07fMXeY8vzhSqqqDtQCOeNzKBEoL5doOEU44zrpKkPswEcufXFch4wrhQVoIYQ40
iQYW+RBvF2j0+qjTskk1e2op2c3u0P4FboiwCukjZ+2nJiAou765n93Ny96eqqV3HQYrXeWcBIyQ
yVAB3TR16n1uhSNIu8WzzyxJsOm6fEqBMeMUu4c89bX/GRQv7RejpIClfOa+PJQ2gcZDfXjoynCZ
ZTJ+48CTLqr1ueq8yTNtRtLWBo55lKSG9QM9W+XE9fCQcZH7ajCri8/WsllI0VQ0IFTXiMy+qkxi
phGLBwfvXC/U+2kOz66fCmRqLSrsvIPP1TnN0ISfXt+iRuu0F7uRQIbAgeM1iEhP2v7zYowBgBMr
EygYW9mWGI+fd8PnqUElBg4xCHJCxdUqfMCxj+TkD1Cslig7y67NHo4A3wi3vl9rqQe9sWJfebjR
lf1Bslgv8C8kpRVu5gZkK0Xp1ruKmwLS7rmfnTp1la+eEDzjK8Q4sOUHQ+A6UXe9zfCcPHCwMB+D
EckJi8cu5R2vyzFO+pMwEnmX3pIB9oDv74ysBFsycUtNzNNqATv4Wvn07cykKeKwykr1ywZoUSVx
vwny/ATC3UyR9d03qlMLRGXCRIJE36mkpe5Vwe/tLXqH8b+6fhNJnHm7J6NGRr5pZ5rc5wdb21M6
FVNq0pXgI+eqGoZpW6Jbe7ZJqd3FlN27extIkh8qMoFv8pak5M5bhjY0zfqjtiP1h9Ju6RbdxZAj
oWCKAS3/dRHFfTAVKMnE8WECDgLhh9yIJDjpcG8ynJ//HSzJhkh8FJxmRfVUhousrBVWuQIthBLe
Cige2YG3tlEM89JpB0SUaykcnb6F/6h56Q0f/uNzJP70s01RoRdkZ8rVYts7vfg1yUj6ftanishT
3K5qtWr79MHe7wt6ixbMYFMd6R8lR12jybvM7yjTjoIkPo67IDw/waAJ7zdaKn1ZuM7pG+YfzBnb
goMRqanbKQnZa3y1pUepRDi6CjCqbHE9XCYZUioCUFTXHWvkQdE8eGc4pvqCbjG69l1mGW7tVn+x
oM9BFdtCJArupHTcFFbwytedbMpNX/iT2Y550kedzhtOQbDUM0YuBpAEw+wotfp4nFZQApQliYNE
3bW13zvNaL593Dn3TV5/S7SH5ZPJYw7iuAzl3aS+FnargVqzfOv0EnU9VxTY4ByoSI54vq+h1qmw
qTUMyeDvInU4nIhU1v20t/+M/dchRDVa1m9r2e8f6XGS799nZH1YIC/rzvky/n6ufHGpHh4JmFUe
mC7re42KZhfk3fpTKiG65vGQxaMFo+9JLJyHCeAHLkHC08JdG9Mvxsg0+60m+n6lBdxjPYpeSVyj
lkSYjaR1ke432YMiY/74WTsTy3xpD9a6ambcadXlJk3lgUx6OLhhlJ5viOHHu3GQJrDgcVetumV/
1rdJb6PkWtr6J61pzQyZJbUbjWsVc+KR/dZ00CyTPB/JVRiJBO6QESr00b1KnsgFS4D4bGTFzNGP
Bk7Qpaxfdg/vUxKV8oUdi3RqI0I5aeL0XfQlrBycmTWGFy2chCeq9y7JBzQWRSQRfUHhoS/amx1e
tnsL3wCRiUj84pRgkYI5LRGB/mK3upLD+l6gtZeNxoYfvQG2Mt8eKhSPpgQcVYxgM6hRb2CUnAlx
1vSd/HJXvONQpKjcl0hCgiKA0S+oQpf4eB3+UmQvgdScPsw1k1dDTZBPvI3U8E85hCjuLCRPkHA5
hZowqzwNA1Cm+VrzWeoiksenvKTGpWXWXfTwW56jW7IMKgRSYhvHKBgO+EDvi8lujgXTalpo1qTo
CnVuOVh8QGGqc9GiWvnJejv1q2M+HhBglPYcm0k4IlyBT1CNwJnCUqg8cZqqLZ88ZeTYr5uIdGo0
pYC/1lO3vgBr6lvPlvMT8HQEEgdMb+6KIMlUjXJE49PVeTwuzwnDcG/kKz/c2qXn8yJVPVkCfLia
TcDu1a8Pu8K+Y3WAG0BnjPWmozjjYdiUgSZ4ZYFRGOswNYdVnw1JfVAPbhSKuw8DPRvgL1CQEur5
tZdIioWLySZie8QMitIlrIaIiR3g39C31q5mlXmNN9fiMWUjsHfddLboKh93gUIrXINdmyTcxdGy
ubLosVRcA9smmzocUqJvUx02J4a+Be1VCwnVIB1AuOncurnjeEtLHJMNv0r+A17bVsTOFISswmMz
ovYyi7ixJWILYXBgWVm4u6r7Od3FPt5zIEj8dD7pckT0CA+jBJpy8CdkBP32V5oOzGXL72Tepqan
Pl8nvuSBfkctOD2pZ12yIu4KmPZjTv9KtXPufOQ8twieXZ3T/jwEZLGDdjg0SIowpwIjAQEiEGOS
FPcVIEGNadR9eN+dmuB1Th2U2CZYIu6NIESTDtdWSSPOCV/tvEyLbjKaGas+KWmqRVE8f8nso8kg
mv5EYOvXuhWsBUDI7Ds0VpxcqPPx9BynBjpk+6aGWACPI/lGMfOeTo50D4jhAFXkH4mxD5PLhwYE
cnmI5zQx1O2LdVvjmUQbjHXPkp7zITVRJFUEpBYFiEuO8p5p9oxl4lfgHx8fjUiJFainIlU1dHae
hZij1EKTm65LG0QIHiYihrbRtLFpjMpQGX/PD+AdX+esaxsOGzuUti237VlDmWtu3oVohSL0qF5w
fPwoZVTIMUHUZIWk3QNwUMFbaPSWG1ZbdwX5DYo+lnvjmn6wCo4AwLJ4ZfurO91rmPTGSuwprDiN
Vuve4QEUzGJSE3xv9XAOSxpu+0wIahaZzzA7rBAKuvIk+oymfP4EPRD5w3sZ7oViUfAhn017B3fV
FoEjD4d8Q13cf3q6Irz+SHqLDiDvFxDKIO5KQFXOZTsrNdFwxWpukuP/G0WnA9SrmGGPr7sn1Ib7
qCNJO5iJGvxEWF7oDThl+H2JpM3egvcx9qHO4MucexdJayMiFXJTSf9MXQ/6sDyTaOGrb9VZuWLV
BBMmvuIt9ZXw8nNm4WpLVHyMgpnrV+Gu//D8ZW7ydyrYVe69TTZpjJBRyQo6e4B9uVSGFPX1MI+u
xw8r8/0mnQ1BYtI/ikx4FiCB8exrdIZjDkzb1yoLrTtCNtP2jAj9n3NVWKb9DtF2i+HtkwzTiuZQ
DOwDNukNyokdCa13pFzsP8frT7gx0+OTLmMkuDgMktxX/Q64LBkC23jc4hvMvSft01p8Chr9/G3/
Av5rnToHOWXRC7q8IEXiTvhYWnWwVQMGD2+Q1SWO4o2T3/hxvTmcNJ7NVCv5IwMtABv9ZHj+O6n6
IRA//nm3Tsi5dzDEugQi0YZCpfI2rOYvUco7xGSm6fgSl9BNmth24WLgvGE7hLlZWfrbnDOtPFSK
gUMdZOu0uHZkV/5AMvzEy3SCzL0A7C3G/1dr5NPseOkLjpzRli5AFXinlRc1mfKv7TZakYdlCC6E
AUOJG8WDYEtQKmshVoBGoI3tSNuJCqRiCBsy/r9bIXnXJHK1Aa7Ji7cW2kCVqxhmeUhzSwzN0sT3
esvMj/B844racusTffqZBD6G1h2VBeJX//h+ibAVsraSxyH3pcGwDTLMOKu2pSA6voxJ0wg32V+Z
4noICOl3dd3yTkRsK5acyqdwJABDRR6QsYM7G1HShDLBAr+Is1Od9xv9pddxahrKDWs/YngI+JsT
oAy8W0U6R1d/2IdGjbO9iqm2XDJCE4z7pARuDyQcrJO+dTPGJdbGN/oXGdyR5ppmmuf2mcDaL5oB
Q/JlmWuJf0kxqDFxfCiSrsi019XFzaoU27SeHq+sMtPzQwKxytM5kEv081+d4aRvyItc1R0YZwWI
Fr4x2540OnictpF8nggTDkkzBq/cLuNcs29yem0sq84o4FkFSJ7gR3KW29pBO4REMtpq3mTMYyp2
vTs+GBsX/IG21dNvVjQ0I+/I9M+1y19a0vbIju1y1qE0c/lkU0+bb5W1nsO+Ulwm8edbCfvYe2F6
T8qaOWtvEAxO37P63atfpcCuWWIgg0H/8pQgsPTToMIRkzdpRSGOjZQDbC0/WgD1WHTVuvQ/u2M9
B6AjSB1TPXlja8/Q58ek8wjzszwZsDmkesj2ZJp/KrZzScqwA+ZmFWQFrel5x1aCaYybp/Hr0Aok
k6LoWAOHiz9Qaoa9+MiW0aihSWli9yvKWzPj3J8iAffypiQ+n55JM8g+pEeo1Va/keu2CRKPA/1Q
/ByJV26OJw9T1OOocJo7SrqSaKWgp547H8BADfKdSWr2Z/m8vxfskeQusvs0JenLJRN7pPOyvcvG
RxONxrv3Uxo1kuCwSMitElD0q9LGqPzQmQs/lJhY2TRo5N0yASsVkXdX1QwpGwtLJ/N4iOaAidll
Xgkp69uE5eiA8HFnrgczUYPz12jfnjMAC5bUYvqtqb5VRt596SRPMI8FjkEB1m1poiW8aItKgmni
+t4O2FGxM3e+LRIAq4qcVkcqwvqPybcXe2cMjx6CRtbkwwFSWYfdY2fUHeDG7vIsKivy4GtontHR
iyUMp4+a97fFXULkjSBox2xX+P88VDtm0+SuGjf/DoYCZ/H9WRoTzGhGIP3uGWc6Jwyx+rWwEiAU
+3vvypAThuRGLqq0RNjNJ0sT0Ea4JryO+2L3hbZxiEGRUIT7XTC+l1Ld9SqxNVZXyuYgjz9a9jEA
iPxtSR51RMwW122OIRe+di0yH0B6usumFE2wVquVA3EUHiyVH0KUGLbkzCMCU4yBuPhc80r8uzgJ
WkEhlHZ8T4IGr7sWlz+UEkE+58FVDUmIVjkOmUuLWxIBJA4vV9i9M6+Ojv9kJLsfccWi4q0fodN5
syq2yRwlXFXvwvatQ9NDsMQq9t2ckg+fsnKPwzbA/W5swQKZSqNJzvpldP0Uaeardjt9o5cB9E2g
aiShHjqoPiK8FF/fQbLXTjgMfQHKvQLC/+2Tr566c0DgyD8d3ZL8vGubZEB2Cc/M9LY//02OpTlw
yV9GJ7jZ56ceTClG3zr59yFCe1BsCzIdA1Thl/RiuoN3rbW9JW26vosl7W0iXbX7uMPuEmrXoBmn
ps9MT8gZN1BLDXpHGIHQiCZQnquqU3GyiSz+C1pzM4dhOWBzunvXReW/SKn4icN4FPxfJ/27Ow0H
xmzMThXtHs1MTWjjCPj6zBZX884b9Pp96TsP/jfDF/jvoLsQpqCwdpYrvul1QAUUjbaGzsoAvO+H
eD/czY41GnSp5Mq1miJM8IkuPecO2hBGb/rivRxmtOt2pN/GBFeyMK4bABpSJijPD7umArl/tO1l
oXZ0oNfp94P5o7agOxAi0xRgz5RaEdDBo8dFoEvPEor53Kxa1NdWVbeLY6cysW6BAa92YKZZPRV7
bkZHSaopdsg31NwYmwCDTJopCwv9obvJzoAeQ5ALfHKi7ZcHoj/rnK54SSDh0DCuHHxgCZvnvGEP
tHrwVWzbAMdcOFCGk4Z2gt45xWFX6mCenwsU6Td4yW8+RoNOQDJUu1m9MkpWzHpDwOt+9mJ1c3Bs
ropQIHntmJu3zvTphCkT0zAk03xCKbUgP+EpBmH2q8YWvkBN2DuWb3osNhjvQhXM3GApt+w2VV82
W415aWdRHmTC2akjTmxaK7elPmqU45cjzBGtCFhAFE3PBCsnWquVSI2ltxLGrUidP7MkErR9fYFy
rwl3GjCTIIbpmE1I0UH5zJ2kgKbQ5lInge4NcUHFfJSgeQsfZyANRyqw0gqlwVNr2foKOmsn8YRv
4RKYQK69A+JF62M7iWszZjmhBU+qQMPlevw2fzbwYqW4WoRDYqAKDeRAZnmreE7Ap9DCcVsGwkjA
9XEjzbUUm4d+Tkbs+b9lWpNT7jK59Fj41ggy27jD1ESdTmGkjZXgUe9CkX9iSEK1qYyGz4JKtZXP
TIPtUxxCrGVMYF/iBAiXRkTY+WkDIGWoR1phRpgv1ahMg5WaV513l2CdtkShHfEJ06Z/9BwxijtB
ZVyG2j8IJMuJVz37fj4A8o550398pDGDeZfVBH9aWWiuf8fjHrtCQ6XY61Qm1qyU1Px0AGhv/bQB
RrT2I9pDpCcbbrF8Fbcu3P7cbKRWDQ2TRPRSE5A0D0r5TSPH5ycAPAAEnxN2Ib8aYAyLk+pi6xSH
5Gn8WnEhESY0awW9CjRwReZuJnajw3KXNRJER4G4KZMI+Z+E9KSuIqwt7g/Fuw7FAruC3zOOsYa1
zJeTzB+DJ1HBEua1mCe20kUWtCjxGRMXBx9GvFNzbptJDnVaOlZ3mVqhgCyfA7Q/hpVEuc54V8XU
TqCszAL98G2/XH5wi9EnT6e8UlNLqAuDBPtkLVNnqwhros9KMX+ABNd3x2wslT1zcgSLFeK2TRSv
Karsv2kN+duL8eMRqnt3NAbsxUD8+y05r4WzUiADdEfj1LaDDGLIpSBYw9P3yEmsZ3IAQ2aujA84
Ea1W2V/fcU2j4MYnmy0ED2H8PTlJUKy8lo5E8ANDgHEWTGjaJoooJT9CBdedy5e/AbK/lm5nJci6
l+Aylr1Zd+ECMmI3Un7OHWbD6yuv1hAr4UAaTOCJw3s3DfmxOv0QYZUWGqcH8fkpi8VhrqE2Ewo/
PtHSqIj5NEaSyy8UgOIHjXdVq+vty2go9LYQsnpMi7K/51s27Qb8PdKbrZ3b0UK4aCp3zHI7JtJ7
1/y1dpf2pv+EantBxniRzgo5vHsanh5yGG90Ezqw+9dz57gpAcBG3RYafBLPVZU3XYzDV0w/bjky
Mb86UKtB6QzC/fbYJaBKb9mvdfTw7lM7Hp/EtSwflP/nkh9jsaMzJo7/I3T4uBJdEsnGwq4o+1Lm
/bJxGLUoyQomwJSUYWjVusx9a7uG0K1keamlweYtwtORxlOFV0PWWa2WD+9vY8W0mDRwJ7cJTTBp
KHLTk0vZZ1CaKvK9X7DfJEkeKWYJbCulkLAaNu7ye7EVftorTmbQnm+QpUXst2SqDJ8323Z+3HW3
lNid9A/OYNqqdimehIwtL7sHccnnzcEOxz+CGiNlgOGAnKmxXvTV6byYQ+Ka67hOtyC8dEllvbgZ
1JiY/+ScNh+DI1dLi5F/MsLkQ2W0deHyr4KkNUCV514fbSrVHMGctCEw0O7F4N879SshAy+Imsfi
nxmioSKq+er0vSvk9Ym4OKiEfdyxMcd5Q0WFrYAnaNtFX8Y2lRJanxCdrN9WNSMslqvZGd/uSK8z
6Yv91GmxQY494QWo9xDrHSj+HQiHMzF6ZNHcbfOEmhTKGAXJPX5OChcGKyEus4YELBA9Ys3Eyzi9
j1wn4GrjnYULHGbTI4MXXNCPSCSpev25i4nub5W+4XEpGrDhJIQdfZ0y4LW4/Zoj+GnU1THAlfq4
P3ixKgbnqMo7jL31d1YGgac9Bd+bujnYSpuagW1uUyDpOn6fg11iAsVReciXbdN69PVjGmSWSE/f
+TYkKp8nw0QTrQy+TYUpQxFFxPdnJ4PbzHISAskhbMW8EvWXQqCGBOjdE5HxHbFCCGCzZGTx+A7E
YaKAtmpm6eXEZrNKFcZaw4ANJ9gkpCaKymMmtMBMXcyhfPlEPUk8cWE3l60oLOLiwfS7R4x6YUc6
YOjKWSEG4ISqrGyXDQ/pnC2QKL9AYQ4ZTI/SW3NyoIZnTNjaRxxvYUgwlhhWPyQCD6HyGQ+/MA5C
wAZlb7gEVE3ycoNhPpnLRqALmIOSk8XwRf7arFOVWxc46NbcC3m+pXMqxa6eL0tscg/yR+KlhjTx
uMErqAs+QwWa9h5X7XufJfwQktdsA+/f1S7XcYByYKngfv8Q954BNxZ+8m+Nj37ypAfJSm5oEdLC
1oojC/Be8BYUS28a0hiVi8Lxdn3PmtHJRkLJ2IIGCrlZGkfd7u2VlpPqtN0M3NTSqL2+nKQnTv4M
PdQ7gfVdKeWDPwcwzB3wQ5yhWQ3PCQcSJcr1mCpmyLHZsy3wHU+n2qK5lbf5f/EcDx8HCRKMkhLD
gdcNZ7JQZ083UZneOvzqX0ChSvRYlghRgNYQWwEFuX9m4XoiHCpBVtye6EtBrIeffMOHM+dT+Pti
CPy02+jUJt0B5q6vgjSeofkj2LOV6Ze06r8p27kax5D2+crvBBY7chL+OqAMOCmdIWUFNIcBtJjm
nvxbJ1I0Ptf1bW79ma8kKK6/UvEaQitd3F6gk6eJzrIuWtapA2CsWQHeu3AlZCMcc3zioVjQv9d1
fri5I6zv7Z3qldIr0onXUWjuPWHCnj1vQX4mBvQFLTFSTmRSfcdAp2O07lfpx4b5FnLRBTQlgmIN
NiEwiUorORAS+liwfB3zTbkReLDJV4zLdp9W65Ai1/Qk1RMFflPjqrE1HMGhVVeUWE+jOWrNJsDo
hjSxU6XlI1kPxQ1IUDLEvnO2+haSlY2kUCmRVe/1x+k9lmi2bUQ5I3+qA8+guJthgcLu74hDlBko
yl+2L3xElTy16gr9MiZ32+5X8EghZ1V+7TM8/8haPxa16/mDY0kobtLVTEeFVeeWS+WgH4KDJjTw
fqoUhn4Vrc+BasAi3T3XZjJWWK72nicLbrV4MdFuE9ec29Gb70Vdr6fwHozsF0iiA53i0Ukj9OY3
zheTxGA7FtnuSvkKbkkfU3ob+aoOrXHHioVCKoeR0B8/gPsnB70QoOxBmTqHHadXMpMXO7/Ik+J+
1On4opPc70v5aaqgJfc4fta35TBVy/V9zDSbOUgnffepLYWmV2Rcm2j2Mk3Hq9FBzc2Dj4QU2Zly
ysXVtCOE2EkaQMjWRyzY0FVFjgOjx1FEddwofKJ9qvqhucWozjK/zH/oN+8JY37cKofUe5iQ4tYL
yPaEZJJvHLvZm/SIULn0GVqD+hT5UnrKiNilz5vQQ3REkVUItjMhfz8A/j6ZAQlSABJitmvIzet+
n/5It04xvWRBKyIHy3LmHLnwGLRDUTH742s3MWNyh/lRkBxomFUuSVOWtpygNWuq/HeZ6vE+RT0r
nvMXqWE14C+gXzGHhSC4IwKHdnKk5MzJsMK0pgWgm8HMlDVHUTEEfryjWkEcRgLtXfxEfA4qfcda
SddiXBRW+P2FgzGnXKOoXhV9HzuJyHSS1frllQbGYA21lg9eiB+bAUWpzdtcbROp8UC8jQwSn8aS
OhrkOoiurt0Ct93cWU4/Z9PNUsf5qp9Nko95zPOXoyOdtHzClG3a38DiJkx9aIksv0CPw1GY5Oo7
nWM4AfQb7UoBK+KPZ/SreqZ0oKmg/6l4qpjc05+AhrZX5rmgvcjOAo56w2r3Rft3avEacmCGj3Lz
7oDSxgr5+rFuVkkWQmaXfl3FNA8m7zutXnCCm5QE2PNd4jiGqBP3s83dGUS87gBSJQT8KOl0Cx0G
P5POqyh/bVjc2+TPd/Y0BT7eaSsMhWFqUSlQ8NiJXfWrpswbZIyu1iyKkqr/xbOXJmcqSCYthYKF
B3fZVeth2pAbOWssW2+Xy6C6ulYZJb0rDkHC6XJ0ZHlWfYYPXMbzo/AS0sKNzojJ9hJU1/3fpVdF
Rdb/S9E5uD0+Y+tc6VUP3+7jBq42MvXTg6nOuSnkqQdU8aMGB7b/n5+Xm0MwUihgTGoTT1hQYfx0
ByPMqMdNyAkxZb0zCL4Pus4sJqwfue3JmFeOJzdBbwouTWSEg4kfSygBRJP2AA6mkbO8sT1ayCBw
QEy0WVnszcNG6mFB+Xm/GmE/2FqfPBI9FbOkciuShjkfM63h7Kc6F9O04OuM7FkfcCZMm+a3U5YJ
QRuIDOy5R9BlgH+Bbwq0/KOTJOLT5ukxlRSVyh6W3bcsxkoBv3SdNeo/QNrp3MApGDSaF3bzQYO5
u9BNULCKmS1QOmBSq24JlnsdYPoNcIcQnXZ2r01c+WZGbn3XNdOAd7RStq9VXZZtAjUQLG8HdLsr
Yf84b0gl8zNifan/lVvyqUq7QSgUiuXH++8lfy3mJHs0w6YJi6OdLGV0TPgJOU0GaOGm1WlTlEe7
+2l1kUAdnAX6iYY28rZ6SiRHesODhL2Wi8klfP5S64FutLE7Zp1SykGkbzcor5JYKt0Hj4VXxjDT
Q//2aEIdx0gqZ6DN4pS/iKEsurPQflZLNyWP0NmV0vpaYY5Xmu1dM/NTHAcMGXf80HpnDi2pzHq6
bjpCHARcIZAdYlHsOVm00e7M7DXhQWzECsw8HOt6bDiQrSds0ourccqESUcYAt9p9C7JbczrY7bB
qun56x2ol7G52TFeHC5gpIex6VzlaNcqnnvVf/P/J6ZBsP1Y2RO/uYTGWD1UI1q5w9I9uskNMi7t
279oblJM+Heoa2hZkjrKa1CA+pItTlymRRn9ChXONTVZNclznSCwSfNz8REqxwk3rvqRX6XlF+pa
ohLlUpaOBCQZn+YXdaafFmdmVh0nqAh+GpzAOa5JqF2y37avVQXDr0yF0FT/UAnAsR9zUam5BGk0
3GmSAiDSFHQVosdE+kBmzkx/Wdc2uzHpSALWaAsZ/ElRnlKSv1A97+ao4E/PB2DvmwGJYPxgvY+x
0QYUt5eIatkb+N06dRZM7jXXIM4NHoTz84i430NYCqCNf3Gm8uOxiUokxVTzasNJawt1/oK7zIjZ
QzbP2Q7M4L8lsymQMw1dnY08h6SLpEGl3D5sdQDgcrj1yRiz4lvlj5ciEI0iXvToKRQJiBmox36q
PsiMR4c1k0eKmzrZLKDtmlYrZucFwiIUkJnT0M7mjWY/nEJoKdLpEnAB5sbmKo92/jvsPBs=
`protect end_protected
