`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Qz2BKiRnThARufOnA7iQEyAIDPSTg3sSshbI2Dcevp4Jr/watwsRuFiUdvFYOdQWG8pCHuobZCB2
K4Ztcug5WQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YHJ4i+8Na6h2LAt0HqovVcy43Gr34FRHgfGkDmHpO7Fggtql8beNbe5+yIgWpSdlo1CREzKM6mEk
Ne6bqdrsZ0mgGyhoUfDDM7R8zBsuh5k10JdZzrlfDMv1WOsAoh/TyowLuYz1pdi3QiNV+9mdOAsl
seY65Z2NhmAaEYhgTBI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iU73N/RoQgq52F+RcqswoLYgQKN3F+3qA71Z+nQs1NNjCTQA6DjPN78bjtNlNxW/T81lHFJcIYEs
wwY2/PI2SWYj9t5GABmDTzN+2xqMsQsYOGcu98Guqa9WZY3L0D9lHq9TXqiT+oujmOU31dROj70M
Trjy2qAwlpPTX73GK2hxqckP8Lj+c+9lRv8/Ve3SxH6Ih+5RnqcecwuEHOrnTTBMSs2mEBQp9owe
oSDgPyRlzw9ZzZO3v6x/ZQWbnNCGPXq1YidEU/7uKEaQszPwOoaw+PST6qJs5p7+X6s6i9wc1/IB
L3tgtYEXbF19zAHo033QrEPy/YbUSGKNJkAXYw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
s/hEs0uGCOr5TpwwqVd2jUmOmATlDoq/ePtVKAr1hmdM3P9nWY5XEQ9OsWCgPNk8JSJZJRsuv9qw
EbrjJJoakEBxCkce0f18nKBw4twpyPVN5j5soeOO5SIbfbFpA9NaB55RZPW53djmK2EQkSFYzn9E
x63eQ5Hyu/DEmyB+gjY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h7rP0M/4j7FKc/sEkLUdF2UqxZdnKEJBfjXD7hDca9KtwgF8duY38C5smV9V5XsU7Mvivsqf9Kw0
hb+E28IuMDVu3X0mc2t0ieQClEgzsNuHxjTNIzW0kJ5qQjryKhxGzuar3w2BZ0Jj/7vpJnmB+IeZ
Y240eAtpcN/D+2uo0OHWLEdiwGPUHPj35FU5yYQsLuKuqf46fVhohRpw0EYje5L+w+FfkuyxpcV4
emnP60vd9BE4a0oNl63lj8NMu/xBvUvCBNmbnRtzK0hi/hsUDsYE1H6jLTr9U/I6CSr9yJ0u9aJR
GvlX9qbyb+sLmK8Ep8kHk1N3uDp7hdOFpA9YyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5200)
`protect data_block
L6w2NClT2nYjESss6HZEd61vfW4DuCQ2NtvDwCwuvFwIqLppz/4mI6rpQHuca4YNVxTbrsYNiH+4
ZFI8LlW8BjZ9YHsgti0olWEXCyIeFilaCUW91PNy+e9zYVOtt3ZcDICpqL1r0kY+dnDxjqlYlW7A
MQCnrJRTsdSXCI3sAhxvwH99c5DiB+5TrFIv/PTK/Ty+Bo5wx9dNXbwhc8VmMJRnyLVR6mXDIwOv
VK6gxi2JHvDQez0lxNL5BjDCoKKM7fz4/R+t1vr8uT1unuL6CrnG6J8EY5X2mXjOMwT3wOOY7YMO
hPhAJ7t2Vsuh2w5W/DoHxaFQENLk96bx9Ty211li/SRRa588G/C8qz+7G8gQmhKadrdwJE77KmvK
D4Rfto1Aw3GKKEsX1rFGPQPRvx9B/tfrj9lyDRC/O9xEn/KBZz+M8FhVmT1ycjD6gLHXcFPD0wn3
4ivLMaH62HcVrf2HV2XufMFA4ItI/x0vKsW+HCFk7s2meIMkGTrPnPmxjxCwsqFDHAsgM4bMKNES
6jZT+Fl0wt8YZBaqnDggQ3OIYMXwrFRoz3XFtJfAOUAKNRMGcyeFjWYLG0UcRYZ7FMsXViP+kmJa
Ku1ltMBpJTEgMQvJpayKd2xVjZQZEwuJtkyd9B29neXcPSdwJwtBWbKwOykScHkYBkW1p+ApxCmG
UWPOarRVYOi6J/buKaeGS1CIEcM3NusATBrTT8HE4VqumNMIJRWX8Cb2QFynae2LIc2xq8ziIQ1C
jG9KJsdULIypwKWw0s7ibhdRsVVv4riHZyP8pWgSV79ZR6fmAcU3Xpu3QjztYkiYF1yGr5xLo//T
P/uaX+kyurplRifhMzWe4a4ILSKSkvbDbgK3ul42RsZjJKn8/BavVgI6ZyfUptiG6v0vJH8bUcu3
sWuKbdIPn96TkZrmY9Q53SnmXmFFhDGo7lHwOl7OObtMKJTlkVwvl5gR1XfzZcKJNBfa8h91LR2F
mAtH5P6PlOxWAGzE+IA/0th8Uu2P6DM7On+0MXI1QY99inAGZ+x0ytiZzVZyAu2fGXW3HiMvKXDe
i0G+ZLzzSfYLx2xQqA2wvHhu8iuek++3eQK99ecgePRYcf0ZqUNYqxunRboLRtVEhWn9QVYgbEqa
n7GVmbS6nZhE05Ea3FDuVw/817l0Z7TNJ/kwxOvZy7DFFReahNUXDpHd9ltVp72G+w2NIL0Ot8HW
33+u9MpexUfEf/Ctv4DIFXGrLBvfzUiJ3jR87tsxnfEviEOcYs5vKy7/NsJRfLLl9SChQ+wcT32C
VSJlP86BdTZMrH7chaHsoXeGNZiolUW5xOm0tGGiBmsMBRt4G5i0vmtQn5qH8ji/VUwNobBaE+XM
PHbRHc2e0K0ZmwkPZ2kQcKfjQ7IOTCJOMVCEEsxoOt6+UIJ0cKSpRkTYOE9w85TJpw8ehtv2pxrY
eZ9K5+J3UseJF43J1PfuFTZyXAR50AQxmufcN6zD2gT+/JGO9yGWnR13ewExNo8CtcVOqHEYpX0n
vzm9YkVEXskAB0lJ3mqRX1ZumpfYPQ4z5n1Px4slWiMWhl80Q+puWwUdWL34WAMBxH4mBZIN3+Br
Z14XC05PG6X8an5vrpYMKSa1rDtQQIE4ZbfGgHpwSOPxYihY2H+9wAmK3uBWhLSCJ1bi2I4ZsHwb
up2Fw2YBa7j27WqyDnLgGw8KZ5Pd6PVW+FhqjOaL25LCrlvgTNrD0t0w+WbbauERp9gW/w+KANTF
kAcDCsmmDG3xBH0bP8tQx9wYEvCEpXLiAVC0kvZwFTHpzSfHkhV14MPgvdcaFOAdmtY9uctpvll2
hb41vLTtKjqUnHrmUB4qlGAZCsg1B+Rpi44SxECb9QlMq45foc9Pt0SBWzKa7ksqxn2Vlfj8PCDY
p6fAUvM9XZ9vXU9Fp8i3h3La5CjRJ80c49R/oxPDSXXY/NY4Anxfib/MIKSu4lCsSsIpFNbJB1uH
uOISh1j2rIeVd/Gafl5fEwAs2VLj59NjbpM5gVhe4axeK5oTWtmTelEj+gvraQaMUbHi06ZvVD1F
A/lTtr6gcZ6NJjmvDbh8wyiD7G4yyHF2ASsP4vQyNRxqqv+JpH3OI+rItPDEizdw7AncTtcQ+n2O
J+QxanU24IsIi1one3OfI1URPUExZjQsleRqnPfw3SNqdJQQuf4NMe4f+5bXwJcYNxGQHElj0l9o
2dNT8F8iNg50FIF+F0dz+WLzItVk+d1r/JqHCPv/pGjI7Pq48UP7YYbaOdA+IOkpZr1jeEbnT5R4
LySJp+ONeX60ZvGdNnl4LduzKo+xijGxEqTdNdIFEQtuYvISi9+/RXM2+FP1N1oC+PXTF5IE1IA6
QkvrXQu1nNfEebMRtv4FyVFyPJEaQrlWrIPybhfNrk9yDZAePciwoxl8PyhnxDixoh5fUl+uUD9j
qoDI/W8ww/rkj3pdGbPiW9QeJB2KTdloTg1gHK7HtCxcckQ8HRxITCPb/q6TzEZbtROePJqDUWeE
yBpVH7ymaUSxNNPfeNVKU2EzhHvy9h7Y/MMJ87ZPYbkp9r8E4s/rlKau+91j6c+JvILTeKY7a39/
5lsMCZB63HK3ysNN+34OHRe8E4C3IRGxyR+SMZd/Fir3tXtFNuJs6EQfph1GHq+tXVXxjTIsIQ3c
4mj2B7hcg25aN8GTGYB2eqrbgdrhM/ELRqgz4kEQZ6duKa0s3W5Sje6vkUtSVwQdODjrLKCTzLlN
6Qdg/Fna9FXdBkxA8P+cBmuT6nPj6dY7A7EGAkPvh7LBg39K11Mt45bEUay4qhUpLFyqB+9DEbBY
+axA1a+xsuEhB7lTXQMkWOKLLnuQCEt0yTxjAkqD+L9Nbf9hpjl2x+WBW2DHV+8ZT1ll5Sm7P/0a
No8r9SzD8Za/pkhwNF15oONjE/v6+fuSlW8ftX2nGPRgFpUSeo+NJumGSa9yEK3PcRqe/4sRwnQ9
ptu9g5UV1HCM2I4DKUnpuOgiDWr/0pBDvoO4q2dMam4LVaAOcjEg5+tW62gJhrkkjdUiuf1jwYAZ
wHPfX4cV47hdniOAupTHKMdcmsyxlTqIdHd0rgLMM/xUdVtj5Xx+XYWY+1QA4GDzjk8FG37E1SZf
IC/9xP4PKtXaa7UsREKCVr9qTImaUuznr18V3eQBBMiqjjf648F3Tmjtq/pUlqeGCL5xTslUZKBZ
zaPq+9R4tReO3WG7qzb0oi+jCjDsoXs5Koo9PKzEvYAaPIEA9W9tqkrzFkegmaG1gqx4out4nCL5
XrZcA+Pn2asMLh/0TWh5VIf4p9gWGY2mYrSHINgluitqvo0fXRSNxW76Semdmx1rRMGhl5dUQNP5
D8tHD2eW+RI0vlubDZ8kLvQSz4Qlir42ptHwJM1DapDkw4vyDcm0X0aLGsmd51dTbZzcXQRFnP+d
WjmGwcSMrjigbt9+aHtL4IFy3lCW/sus4AtS8FiKpKqoGWhlRgRr9GKcvfQxbbnnzGTC74cklMXl
xnFg97qlxPiWOQz6+ph/iF3M3OoTCiFMTwcHo1N4SVO8Asdnb7OZIe48kX5yGw9zDdYGdjgcdz00
1ESg4110fBIomU8Fmd9Je/oM3SEupaZCHVAzbgZYvrqyPUyeH/m1dXQhjomll9w29hxIo93WEGwA
ONyBmGBWF8LcaJMel/JfzexMu9RGi2Y7GfG0zedJGsBHmf8e8g20aEbHYAbejPBmBnCaA8FrrZq7
eA1yXpwVLBXazBEQaOBbz/W95kDPcc6CoxwotHPUkSKbrKbSY0cvLJVCbHdV55g3xin8mKyp0406
ic3iSdRaIxh0tnXWosi2Sr4CC3boVRO9qY/4p/Gh5Oscvidce+kvgCS2Uw0+arbvxdHfh2J0koNr
L6l9vvq0pC+uxrtdvpYb2qYzZatLdVn8hxzaAo60dxw4DR3p+Ivq2cE8bSVz/azDCbi6HTw9P0UF
98Lmpb76VwDEfdIjtEIBjl1gFkyM/HW9YcOiQNQTxZcOTo7Rye91QHdyfG7Nfxq5+vBNn8jI6+Zx
Rs9ocOaBK+ZcLt+Fm62rMWksEi/X0BqrHlCf/v4gtX3lGVVTPmU5mD0ZjseVTaSRjN1SJTVsO+iF
yYc7tGXmFPB5sNjpihshO1vBMGyN+Ppn8+sMuu4Hslvncb9kYoY24tPx7adJLmlBijwh5hcrexUc
sC7yzFd2nvjO9MRYbW+c0444vzz/S5OZmRpefPnnTdWkVPazE0QDRdnzKEyMEkzL4gi0p9yS9Rxl
2PJ6Ks6SqP/WnVLKnVmp0Sz86VF6GnFQ6xmtfoeB6bl0OLPjvD2BxLLk4/v1XziGaHyNPDs8lWFs
/1s1bpQG8NeBQ61NeqAnmDDXeyoS6iXLMN9JvVNnyh1pMuT24VrHrnm/F4KNXwrtsxr4TmWhgSsF
EmQRzHs2OhfnRocGlPotGXm08Vk4QhDiB7Wk4109M0wCzC58e1xnqeKrjCT90cPKf2Lnt3aG3m0K
/nCFxlQgGaBPNSVngkdXcGlEw6vmMdzhO4oanxHblJNesORv6AQW+Sb5sBHJQaRuMDDsd1rnK7n5
ZE9ZpIp3K2is1JzRYwX82XA2NP+1LbzhDiLsgCaiDVFTDsd86HUvjMbLyxpUDEhsujily5vwFQ7U
eGkUmBXiKRsL91j8MfQcgc+9O+gjC8Tf1xj+1zBH+SFtZKdoFphQCEgIUQw/ufZCI4X/MCSsnh3Y
iLMbvT84Tedvk45rSnaVCcXId28TAAw70gerlt3ycGvOyDOFOjyOGT57CTI+LwZyaFJ1lFNpobpQ
V6zvJvceRniumhikRz8Ry7rd+UnFoozrzKhRukqvjK7Ec2xDRHh2pf8BaXNRbw06y8b2aWPN+RY5
4IvilbrAJjKZnfzU39mRqUZwtKlm+9vkT2oWFHbaeyscy+OkjPDmsRStE/h3W5NTGnuh8NYh/7Rn
2jJbeet3YRa/+gXoPpYq9gab/bNODOANpo12Fk6qAq1BzIxnMzxwqvJ6sMUJEiiDOMdrqZzdgIy8
Bi64cHicu1T3bgqcG3icN1lmEXGSqsUqiWsqh0OMc4KEWj4YDPJrRAu/UVGsC6FFtJS5zwIDE3Q3
cQ23hUcA1CJ+ofrvKM+WX4u1LsvXSvZZ0PWskLUvdobbYaCxOU8EWB2Hv9ysbk6gMzBRLtBlcnFd
e2DW1ernRybD9p/eMUANwXElykwQXZGqKnw/vGv/jiL+SdXIUcfWwhpicUmbijMvUl2GSqCK9Ui6
Jf8DHS1HpnrBPHga54pQvPK7gsLyAcZVXcA5yKl6Zzd2Rxb78LovMUlRfjn0ure7KGj4pdAZFcd8
w8tCnYFTuVr4JuYzJNj9a0GXnwXY9Mz5RroVl9lBuTD/3l8EEHpjtnuNplCqSmP7n6x7XUHDw5N+
/9mt5bnSRMpDONm5NUCzVi8hky5u3mV5jvmOqWTnbJLCsMu/zwcc5IZvxjqvUTyZ2I38aWa7TpB4
wiCRyb81fcDgnfSl88KNTbbWuvzrn3dX5mtS6cXPsoqBK02KtOcKuyHn15JtJrSoyBgLOfMeDw6z
WI/ww4rATsNsI4471lWmg4yHitwMMdJkQRNPFzXuUEsrfAt1Z1lhpk8lVDxD9pY3B9OoMhspwop7
MJFxhHAqUzmAseg61RFnxC+yRV2HChY1EHRhaAil+MLmCmG0W2p9l3kMim9mcOBtoxZjBfEYUeTO
WqtqQf4INs8nlbj/+uIYBdGlx+mDtx6yALDkCSdLzGCUHmGpqLFOftFf7uEha14U1ybrTnJnDlsR
8gSEcef0Ygv2Kk7k1RIdpKPfo5x4mYs9S8nb3wt9Czi9O9OOwtY9hpsjNAYhKowcri9cHzqliTLf
mOaEmd6K+AG+tCdFO/e0cPtAL74ER/k3YBCaWXffYsISRD+mWf1hn3hwtuLXZqvjQNVXb81dFTeI
UWNN4TRuoemxOUqgxqjKhd7townwT8ov99maFhq/INd//+bW3BU+HuYwaCxlEwl6RN+vJ78NCQzS
PzEfROGhpxEJwsU2AIH4JDGdESAoKAo8d5IM7OL2AoGH6WxpB6W5KvPT1dwnXeHxVSLX8r175DAC
GD0qsDXq9khfKLipGjVSLSD4cDVUAt6YzVpmqfkcz9n+2Wg7j3wHGhyHSAFlALTA4U4gEC3oNYT3
uK3xTCwzTr1s2MrErVMQTc57jI8/QLemtvL3RchTPjGJD967ZKc1TQyKgOFOzkmFZBBvvWua31o0
L7n8dLz2tyYgwSDJ6+gf7cD6RiYEytD4TMmmoXulSUlCBuVIl5ZR8gAturT4K9hChW89uD3al0vn
/khxdFqfpHKM09OG/cTZM1B6EWJeulxOECf2WqvRSzYtGNODXXJ7dpWbhEZHUXaG0/j1001YlRfG
YaT4av/eqQ0LFnwdwk9S4mjRmWy4cULeiHUXsmgNWGDmDKYN8I+RaVugPhbwTsV/SnqHi1R/1Kl5
KzQLs4O2HHITC6ZL6ekwkKen8kZfQkgxV6344RYH2C4MFSN9p7Z4+iYROkbbb7KR1MGGCf6M+jii
c8vvCCYT60zWb0TS2vwoPYWpeC35QJj7s7i7xLOnIqHLtEyoReu4G0hxbAXDe0/WDgUGzhUWzjHG
aEgxHAoUURCSS6lMY7HvyBUfK22A2OOI34r/1oj+VZ4LC2a3uIHSnKMsdizBoSeyrk1uO0qozZVM
6m0sl4Hg3DABa2VsNRFKf1UI5MQm1vkvqEqJMF5g5A5bZX98tlYuOQ/d1Xh4JDDeVBJCMzW/TM0S
bF25nw0NsgwiwhPryZVkvXiv1dzhhn9iyQvMFqGNGEuYFu87l8q/O9TPq82u1o6BB7+p3EQwWYbq
uWY6wyxAdmhzf3gl5dUit/yC8HVL+n4EkBYahmTC/s6b1jJT9LXghJ04Z0wUWGDMwKdeIMQyfF8S
9T+Nssetg8OFjmqB9Q==
`protect end_protected
