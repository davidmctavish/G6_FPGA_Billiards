`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gxJVQBcSQzsbwH1GLrg1ZESzDvrkikrA6vdLpp95ue41M0lmLElFgzzCnPkJPvxfP02JEfCkzu1s
pXyOx1+/ZQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6UL1EJsW9MY/SAJjdc4y/0ZbchfPWRZ1fO8sgcSvmzT8PhDxHiE2Qv094M2Mf5UxTO1pmguf74
HRrcuhkl5xTcz3SUgEh1WqTgvNR8v3I22HLFetAdFeAfwtFZ8WvCSLor3Yg5WhjacxKzsx/R+B3A
Ic1e9ERorPLK+2OWDXk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VKtFT/ad0mndSTNYku9P/p8pTsvri9shyNk13WEjbKiIq+gQoaEMBYqKlUj1txesDW5BSN/vb2L8
WcR0ho1RI1AGo8y9tYmqORrdmk40Vs1+gqMQCfIiZwlKBZmVSoyHFg/uvBbeY40omXist3OrVmLk
ek7TtttpRm83fmMK7OGVEehvqtEULYY3DOqBcu2re7sG7LxKpszndoH7kfBnWA+R4Uc33vWeadnd
g6Oz3503o4HZjTYzqaI83vGJuKxDWF5lpNA6grtaK6MLeulhLJkFI34NJnCbFwlIH0j/a6X/NOK9
kE/9xzaRMrt2DXPz06r1p9zWXUaXULkLZNJGCQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSxesrZXgYAQp6z3s+Mn8TPb3bLkqza8nC5XgxzWq/mXl1dMa5Ml2g5M80mUOlkXRmUOZymc+Bc4
WM2y1HxgX5+JsAIjs1wpPrFSHzjHRcHcvowsTXhTMQ12m5t3+UzDaDcRPweSUjf18fqi6cqE3nVU
Sfah17SHXQ+D8FjN0Ig=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pw16GfE5lmct+1yHq5aabqWplAJ9NyQFSmc7ZK86jiJfkiQiewcVOFWOaoYaAbWH8NvRlUTWxPDY
IJZow2AxlsHQYg/BVCCfi6Nou6nItiOvPTdaycyuC2yVki71gI8y/Hb3VqhrwCJyz+gO8RezkRKT
K7icG5iNkHF95Ybco1baJF1EsxTsjmFbbCqBjLdWPS+4hZQmoZ3Ifbb7SnBR+mh541FCQTCGTC2j
d/LaIIFECqkijQ+ZFSd6r4keOeZDRlAd90xaWc9YbUz8EcXsrFGvk0cfiELaenio+xWCzcCA4xZj
1RA4VErN6S6k0GdYguQHKTjRx2AHdBSjKkPAZg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8720)
`protect data_block
eZQbj7BZE/w2yRRmCqT/kugimM8hoNG05eTOM1dCqRFVkd0+dUXdup0xmX03/Oh3IaFgKMXxrnuC
fCULAdqNGWbZgQGu1DYuGb89q/ujzsC1mYtQ5rdtv132hQg5JtMyJIMo4OL+QxrEJ7waOFgxqH99
hVDstYdU+VsVHk9MLMt3Sn+DQia1fXhn3bfMhtf9Wyi+IeTd21Og9b2EAVrlEcTkEbKc6epc0E9h
ixNqUm2SWsAes7ifxrGwJa4ZGYw2RFtCP9T2UvKEWrIIz9ozGyALBB5KWcxjpfUAZonDqUAjAbuq
33Z+V4qzYdHYiqHgreNylqi/HwkpohnRh2KldTvPfKGM8sU8Bhtl4diW4w3Jawjt8IHIMMAbmEtX
ve1dLlEZq7rLginu53TBXA3RmULCCf3ajZzt/heRR8EfnYu8KAW2voRHFoQz5XoUBf6/BqN+OP3C
uPA20tfs3ovIFSS6hL9N8hziYULaTdk4tIzYxTqy5lPyoAT3k/nqpFcXgPqGimFSDSvQ9mBgEzrJ
a8TBPImEKLxcns0vJ+JnO0LL2zF5/+OhJYevHfsZ+2CL7aPqBDUYUV++q/8JdhJiIl6GMfsPEwch
YaBTxUFWVhHQTNA81gPILITyaIxDtwRrI96ikxZV68IUIZM/3/5WQzMF7g7AePXWBAAGCf2eabx6
v/ldoXk3iyWZsSsq0eIe+PoHpz9DPgHht0CECzvMerEnh/kBpnnqdcB658/fgc3jAWz3DUfw51/l
IMZfkcmFmvzg/1VROkJhln82SOCN9mavxfB7COH9IhhVow3Eou+JDNGyGvvJVIfgUIzFIGVrRLj6
AvDpTgxXPmLb3Yo5tRvybgTxK+YilDTg+xy7weQYdAkPnyuiy33twOxUpAr2qd80udTouq418ZS8
Qq+bkaRSsa/1QzUjMDWE52Mp7ugpbhExxkjXmPXshmqBwkDqP2Ir5IPZiryTFVFcFgokZk9qonYa
s958TIdYa6ucuBPNgR/GZGI3TLjrhM22yQjWG45NYPrDEstRDwzyc6J3ajC2du0xmXQE6fFsjHwp
LN5lEczqSzSDnyZAaVDt2Gene0jMYhUwrRalD5YVIL4ZaIV+elT4GsPSwPvSIR6tOEDNtn2UzLkj
npeV26Cq2ShrwEUpsuhYL2nPo7LCvMzsD9biFkqXvKYV1Ej3aLKj/713jmRk9T6KhzeCn39uSn9Y
69cO9N6tOSczzK5vk2+ucpy7/dJmp/hR6zfBIBJFqEpqkLrSWUl2WjpTg5zAwn9pI+OmyMCoUTQA
HL7gcDMa6NFxP1USsgKcruqyDUxmXmlcU0s5wW5lWchxDOaNgSYD/y2zo0sHNAsRGY5N9KcfiFJQ
ojoSkyAQzgdoOP4Ha9Vzun/g9YLZp9KuDO9EP/KHybnUV03OMMn2aZG57GhUUX+mdbeMaXQ7LaAR
zcyfpxRbcN+fw7RWWDMbIpZSjVEclizmQTKWkT7Zgy5HVkxy9ZRQis0/39VTHU2BIQHlkVBGE42X
xOlb9GnJ/dIlCWH8eXzQxx+4dlWTevibg9rnwF4vueuQlbZ0WDlvzVl0TdslLayQ0X2ch8Sqf9uq
kxdcS8uWlMDeP99O+O6QIMtOAZmaU10K9uZYtvCh5NWhYetzu7MTes1xUT6ue9V/5j0ToCNHlbeQ
SxmjW52SU6zKlfn9k7Eu29xscsoUPzPwCi6uK7hZUGFcBv3CQQB0IJ40OS9uDnBnw5Vg9PXh0GO8
pflTev/62bU3NPKxdWu4CX4GH93Kl5dXF16PBOkBtpMvcdmV68/hUyvWsx43LzneXMrTDZ9CVQi+
X60wNgYF1CZqF6/b2knAC3XbvbjWCzGpyoEp+J+NN27RRSVwy11MuU0+5zmqNIpM+sCutF0T2s1D
01imHCpYI5kLmS1BZsO2T84hzhpXQdOkFPGA7r9jkb/Jz6nqJ4M4pNe9RambCLU55yPz6lRJ1XCY
9ICJU3ZniaoUXF7QM1oZnJcnx7dObYNCDuPrDX/pLusTAwwbQ3Z4QEaIAJ3K8v/fNTLqneNxwYkf
7nW0YUjLMTtfliIdzjbk0xzz0JIf26RDawPaYHbr7u7tqwMa3Nf7QqFy9JLfGwaIed8FJF+E7bwv
JWyLtcymOxydgD6LCgMSO6LMNLWtfisXpsCW4dcGImJHZ2B5MjEY/JKPdnGbcamucHMG/q+6x/xO
/MtywSkQnT2wfJavTAwpZyC98lQH5jn4DVvfYWHz/DeDsgoMMnd1FafahCkmUE2gsVvbBcsLAeP3
RhGqrXjMdi9uTfn6d+U3AEvtxpL7rZYRmx0hMUqpZVZOUGwF4kIUdYuag4KxyLR2/Q6U2xxfdn2P
Q2j3Yhb41z9Ow60JALE0nqVj25X38VtUaAxeoSIyJXhFCTu/Wpj/P9dh/Iq9Nspyw8gAVu1UBsVw
1gBQ4u9g23ymhS6zLlA+k6UIE/tWvtVBPDgAz0lGZXN6rL3WtvB3GusLE/CAHlyDWNwZpUJb7YBe
BWHbfZX16vwtBFIWUYbUiV5D8IXX8QxA/gIp2iIg2X8kujzI7+1yb955MOEosrpZeQouKlC0pLZU
+ud55YB3EcXP8Qu4wO3SzRqZnVTcQGs4Lzj5Om/IIkzaxMQNr84iB8t3ZR66y0m7o7Ozz0U+3e4P
vP7ShqOkkY9g/3X/oGln0L7G9jtt63Uo5rrpp0MPiVdS3wEHpvcE65BgbIavng+AThX5/7s1Uff5
1flupMnBJ8//2LnRikQIFfmxvuiiqL0WgeHvZYtu+TCVhmfQayPRU5kFczxgNgkM6JlRAgbqGtyf
UJvHOOh5KubhFZ7VKA9GsthH5bwznRgCl7ItwpyIvLY51qWhKH0y3D+LH/dIl02qlWKZTV7tKEu2
K42ZSWcNJVX3L4GRs94TahYcbKGxpVTK62aJO5Omqz5YfviYAJS2t2MgN6VbPiDy9mzCpS3GFeGG
q2xjkbtfUREsKGIYWgi0jmN3SME1HgA4j2wylQp8ER64TjTE+ty8B64X9eV3kVJVgynf6ggGNXqx
FQmiPFVhCHSdRSxo1HLEcLvaWvCJnFNcf8fWSR5nrclnkBQy34heoMG+wd0qfYt1HOkGw4nffcFE
+QKC7NYMCzvKT5agzmZGybsbUeMp2uWTS6RiVVJdWvXVyYk5qfYj9mzKZEU5bdV/4fZYPnVxkaqm
Kf5+P0jw0T2exAJu2ldIK264ACN2s5z0O+WDtpbAxbh/jc/ZO8TRGuAbFSf0vwRkNDzcUAsS9CPA
4Cca5nh3DBXvpJc/fjW5SlfScRBJJfWoA2A3bXAjoLSFjcJt9DcbjE4FwaLqRqIWPMDJuw0uR4Sm
8HBcBpkX0ynDeqykkdm++P6biS5izQ40DRbwjzsOtlQREMLMGwLJumVCpdRefG7CfJ4ROTDe72M1
weD/Z19GBgV1pAkHD8tiIB6X6xyXO1fDa9bLbmGzpSi9QiagutnyJojGJyW+wxDib53wg0jpw4T0
JCs7w6fmwAd0zQJ2Z7LXJdEgCrxx4VpBJs4a2gcZICnFD3Bk9cZO+T2FRJc4E2W2Xe6WVu93HqPS
hHU4CZUqom3t/MgsljOVrasTKdZEgpRGH8ydo3AjPgrQD2cUgD2I/7wxrL94FfhwisdqXevtQdcr
miAlY5VtMWNQcKsjSl9uR05NxFhQ8VuTHNvJ/dnYGzuI+fLkO7qyN83O+wHuYP29I6H6r9DlgEWE
wYkqYAehNSMZPinl/Mtwc4PjAYDoZIx8R66zHuNqfVE8stBIYj8C1HmPK4tfDmdOKoh/YCgho9/I
6BqWPzM4A+8r+3gi79R1m4NO2hOUB1NbNprWgjRsACoXKSJfcQQzMwX2D9oMcBl46JmhXtS0RAVC
yZIfuiU/mdc3MI6qTyccuR2H4yVapkyWfrz9BuLRy6PEkv8u6uTuID9pQleCu5MSYT0YjAavBTr5
M5ah5wNrkDAmgF72RucffaY6Prt5UjxMABJU4BfTzSp8O2bC3uTAVzx3K6vuADOOMMOeYI4VLltX
DPdPcxIH3FauIPNavhYPXs0fZsMsxmiwpHia2RiRKbl6JP1Pkfn3txUFik0U3BkjWNrNWet/o72t
Na6kZoIK1gqucJwryjH5WpTTgdwxNZleV/FALkSj948J8/sSj4GzoQi0L2QJ/4xYYZuhnVciNzo2
Al6jOu3WGE0H0iPphpWokpzFHW+mLD8MtVCLGaH0rG4v0QOjojnHlkfwyz3c0QFJ/bx79Fip3JGO
i42dKnWPNsVJxieMVdU2X10dxF5j4L9on2IUEVjONvSSjxOdk7+df60vzQY7Khyc6P4y9y364MoN
Vt/PLASM/USx80w3ohjumD5xi/Yyd+ruC0cblDUjlywHvUHsd2Z87w+/xOkzk6XFYz9xpICjIaaG
T7sG5CQc8yl5S4+bjnoKPHQXRi0Ln1npMQvQ/vI0X3I2maFlACKOeG7dcaVtAj5/BnTBHSM09LIL
nc0jF8hMe64FpOW66zYyuQ9o9XN/ukOM5wB6+ATIaagl6S/Vt/exR6ALRPEd9aFnZjfp65aWBBb1
Dh9MQ6EjAAIMdwgfBHf7XctNmvlCHgjdqoBL7II4gC5irhkMFfkyIIDRLRDnAg02XSYiE0eRFR1T
4wU3Dj57POUX7U26r7feArSYt+4jVNXfJazvJyx7bbH6ARsieSW90dWtu1XGO/RdwytqP5FCBmuk
me3ALF+xTihC3jBUShsTol8xQZ5M89m6800q7bjVLcXFXSR/1tTPxQ9GTilBqQT1cOcZY2e6Yp7k
ySPZYjLwL5vMtVfKq0WbcTQkDFjgozSPiaj/eFjibDkVHgVgmxz+AjHsLMM1sc8//JAMKEtOEQkv
uNY9zsAZefTFY76S5h+/Gpngvs8SAidSSjd0UiZhXV/asi6gygw+3ft6NwsdsimFtnMM1vCVib46
i/r9OkHjq3LEA7w3ZZSZAd+8QL50dhT8aAVux+Y3IF3iFNIE7P1dbK5BBWJfh0tCg99DKxjC7f7z
MQrq0ooLH9EcJ50A/4drydp3CMDWSFnCQ4ancullgSheoKcxoFxw2+OZsFvLFwtKrGQn/yWzmngY
fceKaM8SQjVdxLdbPgLc1d5a25grH+DdzUvmDIX3CoBpXjclN6dbL7Rm7Dq5UW7TFiZQi2Gq7K21
6Js/mnJsj9diHyEULBnYCXpH36JhmnxyE/bweufM8IEFlTHMcY5RXxQ3V/Ic0dyyhzQYgz22s9f7
LZiLJFtGJS4KFoAX1KrKL3Wd8Ix7Y7Ui11YrMC4jljglHMNYTFlBLWB0Qc0nV2UjuURme5p8Qd0c
39aQkPi5gfbO1FCKBm1itnaQDYFT8fpesw9c2+enBmt2QUoNnAtHOPX6let006WBsaEGeXMXL4gG
iJYXhk+JyWgARxRQDvqAHDWY3tfhJloXqEAd8J2rT/kgfDrGXUhaXaB43fo4gFlcP3Qoe2WNmzxt
KvTvofkRZqwtbR6MHWVdSvV0+3ZTVSx5guyQ3M9kBrrbJjgQF/guOJaThUF+ACdzrFK2RkiCkULh
4p7OumxQgvWR9VKsCd4UvxlhgEU9X/ReuPVs66Z75WxgGRvRWmVU+5TJfQPilPytMawWTRk660DX
+k31inIZG1o3BHcEXdgK7oU4SF+1YSBu6TgOVRCKAD0g2mTfKMqv6AN7odtgo9j/idQJWCFV0K2D
kmD8a9EFv7HpZyQ3vy0woGbGOeIylNhGGTcYUQPd5wQg4A381GJDMCRTLm6LHOV6zPhPgnRfXjub
xeSbd3N9BJkFjf5uMLsKuqr9cOBxJkFQDPzyaRVDMXtgkMxOUJtyB306Ohg3jC5u5nZv7mQM5VW1
iyvDIHvXgu5Dte4rZXxdwQk1aGgXrEN31JI2g02QwzDmseMlvgBxQlb/aO/46zQ+OpQerEIgUakV
EeKVMAMcCMkC9fTx/TWN2toma20KicUK2MAIq2wcFAvzYZx+2KaAlAKFhzds4YvRbf6HSKrsRt5i
MIPBg2aIzq1W7xHFOhCcG6xopuvSPcmm3PkbD6Zhx8FzcbsHe3nffA4qIWz6V6880bHFw2r089zH
02G+PBmYE8efsUwdv/bu2J5PNojuzckMd0fMTWgCFSCLWyGA+qVf5JXHO8TDZ6cU5//J0ic7GhvL
4kU7IWE9IqaBby5NGs8x1EltyIEgvfpHQh0zAu8ksJH6sRmGvOdridDO3SquwzjSWIhzbGg2J/7c
pmWyewK3QL711faRSh3859qa6APiJOFHKXJ/VFD5Q95/74X080x1CqLdsccQ7zx11S2JbFFlFpoA
9LFAdDN04pxS6ru9yY4Euz7akmcXGG7aFbSWMatThoziLzW9dmT2lN0wCP/gf5QAyqN7MplRgIKJ
5Bht4nnnEtrjzEXH53StoiTOTk8rqMPFR3rPHI44pN+AXknQQQxVCofO1J3+b6I2kadNu3/toss6
bXSswvjr/4CG+7EWc9iHn+5WlTTxTkYMLMb/pmXOyhUqs+7AFoU4FJbpNu/Ro7ZRtu+/cu9/wmkC
wQ9qhvJeud6pa8IqW1k3BNjBzxOsvaOCgj2OiobEeC7/0uV5SJ0Ap369oKGaHXtf9A7L6NQ10sHX
jpyBD+HlGa37Uh/3DvG+YiC00ukyeyAFDp3gIC3JDk6E8LDXVTQ5ogWJZOX2JKfqeSnRgFvAIUY1
vEwqjJsowsoIeE02Wg9gAjzko0YueFDHVroAPKJu9jN8j3CEAc0dRDn1pN8AYyd1XF54AA4XS/49
kRE9oTINXz5WdNU1d0iOcXhUBl92rtjnCGKSNuQ6aVXVqVNtvIxvnfE6AK8mVivbxYKpHHpkCaqT
9gWoE1jwrz25idKx2+/M9nWnYRx22Gb2ofl0BPYWcKr0JNB6uDlTwzRBjE/f8soaP7Vrke3sqHOd
r6AbYce50h1ugxQVJ3IQI6tms+j4KWfNFJrl46tYbu+QTd2JKgYddf718lClGEY3hzuzT/cCcXgh
tpfvlF1HL2t5OxqhS2WbQct2cCZKzAJ5mbenOFm1z2ajQlFqnhcgEagbx7B+oHjXodHjGcBJPW/k
isAGWV45RKI2yAsNdJNpBDfbVJ5qS1vlnf08llOx/L0gHvq0rnkquWnpZDKNgdShJygnoF/mItmA
6pE4bH2Oxs9OQXq1d8C2CUJD44yj5L7oEhee5fCrp6rlR4rr9rTkXkGN4303aiSmCQcxgFABRAd+
pwtVVxZ22cCz/0+H45VXW089bjU3FSCqZWi+hMYvVLHtuGSV/ilgmnqcbQnglsLuImvID9w26ezG
ebHAfuxIiwhG2VTUya3DATiKORwJZZmtwRymw/3wWrAmelkXwqQLs0Md7URGSfMfa1YhjLf+Eb7a
gBgBnMvPCxr2l5GtmS3o6DNGNuEi2kUZIXfpZkNuaENtamIzfuTO5sVM7i5KFE4bdjYJcZGsGTn0
eXjHpjPm3awf/P/3JuUR0uISUEFqc5rEtOk1l68h07KKiRj4P86plDpj8pplJ5S0ZJmA8CB7A1x0
aJd/ZdF5h6Rz2VJ4DKAvtzQ5Ihj8JGH6iLoYNTG/eoVau+n0A6KopyhQurdmQwvyVCPcj2h1ovPW
+WU6Mxq+3czS6967VkrXfG1kOyARl706npzYFYHokJtzDF+5N7sgFd50I3j4KHKQ6oyj+GalCEus
b1vzzdLaI96BGX0CRwjxPilbsevVO7QLGrG7XJzIiVkvBsDgoY0gSnffPl4YW3Ex/5ggqM0okpzV
8PDNZQbUo2YmW6U5b272Zimrx4L3c+s+qYTUsV3sMVvy0Q/NA349iQVIjAazuUfW/8WxLXEONvZs
clLNSfZStTYCIWQWlzC26A39LDc0mYjzxB+p17+0WECImmiNHL7xfzVVpLJYssy2lALcj+iu0MF2
zOkveQibPKc+xawN6ed8aoHOb0ktzrqkNR5p8Tr2yEst9Uxxa+3EyjLlgqP7L2zAEFYcDCR7S4Aa
HwDTZR218ZQiu33u3gTq+Dr0pujZP0u3uu/bz7FUoFOqVGhrCyXk/9sRlU6d8SxY2n+UUZxo6WFz
RsITZBGr8yTyct91ECuVNJ/A2+pe2JAdi02QlMj8RO8+vMJo2HUtzAHcUfdO7QJZIlMNyKiDd4QT
j8G+8RBstF0uj8dXkqd1nFR1RA4CJi/rLOsga5kkpwlPPSOSSLMsq7nPMc7pa3TMKIYPVhj+rM8P
Vf/EFCy0J/bneFhWuCp8jh/GVpBYu3VsPqfakhnJqq1FcFhB0JP4PdsQGN4YUczLLxKbhSBLD9E9
OpOjO1s69qBSTaQqTHAB24rECJbwScX9mFZLQ2m4GNLnXbpZf4QCIZR3XK4x86xSZJvVOp/rkTD9
zEDRfUnwEUNZWF2HcFk2IeeArGVPQKvGqWyovTfhYVZNaQH1H6F9O6in3KFQSXYKeeHh5BKsP9xj
Jiug3jc9D2wwAhoNda5IfcXmSWLgvJ9t65vj3u5chhF+u1f9W2X+2kZ6/XXAuRxOwtc3YrkUXzHU
/OnUxw1iIFtiYiHEhP1COSB+BmPCwEqIYuo7gZbhJIMb3XNo743dve3onUzo8pXut1S1dRZp41ec
kGt2/nPCB0PbGK3UyVa97JkvVBJtHW+wP5eStpNhLynq4Bce/fR/ndRuHXxldseCYo37QS9efmKb
S8CNRn1krTtaDhsw60agGu81FAp9e3pw6qmCdchWH2B6fF9TlIwB0ktlAwKZBtVRC6qHpgvGuRkd
vypBvm/vzqo55/aiX/6U1GSJt/Vj97RjH4Wq+0DfhGTzbKwcj98KbEKg5cEg4Q3J6cvWORuW4W+8
hogtjET50LVBVHqQBqnCTDaILi0nRNrbwT66qglJeORSj5165ecCbLI/RjhEF/elfYf7Ffr3Vdw7
w5fzTnJ6E+29AP8YESXktaBtFghUuGJFSowTTRvh/gxCNx5x92/wJQcBQpUXDpgGojysbcIKcxqD
O6RXucGqGsEl5WA+pdsgVFFysZ6uKkf7cLZBeWYzZfdYBj/Q2qyi24U3Q0SNfiuU97UAZ9jPVLJh
95aMpci4iXAj3W4qshSMNP23C1kQsLCw0wSBKEGVRftMrju8a0D4R7f9QyAEgGbFdy9Dzv14vNhi
2RxqbNAzPC80+TvTJpAILqFH/NRF5gJSY/fN7/x0Xoin9UJlZtmfp/Hc0ShLZHQl+HdI1hHdMK+R
pWgLND0cbMIxM5DkjoXfWO7X5FVRNX9E1c+WearO9MSZ7kW302o37NapscwVelOTaaX9Wg2FkLmz
4Z37/7ATxreuPtlC3ev9UBhKV2AO9CBA7KKkObBKrhsY1bAPDb3UowBK2HanXPaKPBY+7yGdL6HN
9xEf+Bj5bm/k3LA+/QUsG20JMoTy8m/zju85V5jdwHIf88WLUKEXIUFjtwri0RCHUmkkVGDKw8fI
IZwi3OsQizbwGIh7aIOJGyi3zg9O9lld8ak6L1AOJ8ooKzz6P9fQ+f8jrIf4eKgymeFW5VPPvAKm
p2p/8in110udC1B1qU+TWqd/AFtwgxZ0H1PopdVkpUYcO3dy0GS4bRwfVHkGATYCkox8u1TeSJL8
eYSEHmVn+Uuz2FY+S2racrN7eD0Sg9pDLpDrEEliIUaG78waewSet4zZugzuaWDsFn+OxNNRbMz4
c3PQK48Yq2kWlfF4A6knhnRspQ2Q0NfXi4UIpnJsqoAGI4PtxW/zoZBxaFdUVeu7/7gRQ1eMVZzO
pCq6hneXM0qSjwpQBueiB9vVEoOZxv7zz3GHS2Wz5oi+a4BrW1qBPrRGwTfkOtsmhJOWpHmsJfEh
wB9Z1QYNGcnaUF6uzIEMqWSJyRf2f3+Y278klBUjXLWhXjeXm0p/8vZLqgpYWPnvqwtXTE18iO86
Whoea13fUs/D0wh+p+BRSPxe4t3jGW2Wz09lIVW3kUcccciwvLwtHfSFiO7sOrphyJZt3nOw7LRe
oi6ebUvbp7A8SzWM7+AqdSVwHuYZlGMryvz6qWv3LzleBysYt+DEf5/JZMWcc3/bd2x/wjJiGOCC
oGbM202/i2G+m9Cxp2xhBC85y1Pebcv3/J7ZExsD/qCZUO+6tp4TDKJsPrK/qqrOSDgBghZpnFgx
s58HgbDCpJRxsC7UaqvG2PoYznmnLLIfbZgLGTAIcfO3958uELOIIMco3fFlT3oMh4pQS1/sqQrL
1GNpATcasYHIaFDokE6vOglVCyxlpZRoQpYpSzpRvlx4TuSwCPL95wmoUjaJDntj7fQnEhoI5MOr
okNbH6OdJVTNNTAcE5CgpNy9yxmuIGQKdEQphUPLS6ZYP47XjVPC0/oXsa3FPjp/r7frkcWgx/KR
4InyTd7CKY0b/qx+7nnmKHZeQAOqf2J8aAAAgtX7uqqDW1YVbsIeQ1LGPLZRQZif2FXdvzmJOj1m
ecHKpBClq4j71phP8erbYZgvzIuvhnbDwxIxaO9IvqHIBpoCFhs8/RWqV4qkSjRfCxC791XhVbKN
Xzgb0Kzx4VY/qSE/JztpyPLJqg4hgZkkUHBuslnJzDEiJ0K2pkk5TzZBBaqZPFH0vhkGRohBg60v
VpD2faghHOkbpbU0dncMlpMaJw62mKfIuIvrYyl9eXwmlx3nyafjZGUxRX0kf0n/pi6je9ZlWhZl
yf89lyqhOBlBU7dGkFxZzdWKPH5wt5WQg2wj8WAlDKm6RoSadwpWP3RvtepA2w9IaEte8sjUOHSE
O7BeJR8kXjQZDwajZn0rkAr05rxVnX0O97ms2vtNZOjq3oSnH06lo5dME1o022Y7tz968lmae+zI
NaMrX2f/GMbZzj8qzyXoNnD1kUAuTjDgcYf4oNS4AzyRpgqzPH73Qv1eMlJ4vrhAIWnha8MPrvsS
c2cgAfcFMmJ9WzUooq7h5MetzHGlJdPY4pmTcoRtf+jI26Qm3wlYEvYVJmy8eiBiw57ZpQ1uRd8y
iUezBe2qwyigL9wMPAjyKhKROEC35iXrQUW+vPCO1PrFejyvCoQyWrKt5fbt9fKxPVWZc4eKMG9N
rfz9RITKKceHQUJg053mKTk64xsPNU2dyXYbsb7fwzNO905vOvzJGMaGLRCR9gsj0spdfyONPhGo
QzJZGpHAd++jIsio2XTfiUKhUchGU4gn1Zdpzy0aXGPqseTBCKH4fUWvvAIFCC91RAZVtdZli7Na
AXb7XABg4JpR58Y1BIh7TnIymlZbBiR3pTDdobNQoPLlHOWqKz21YLTwnyxxbB7RY9AiDzekXHAV
JmDGXYhOTI3Vb7f9h/U8S08la97/Z2p4lZPcEplcduGA+7fqA8KbbLjlxkxTPXgA/lOuOC1SR+b2
ayr4BR7U1j9q8CCvGDFNfzlhT8mgGOBiZr9TBWfLLn8etF2dtzJiAPPZ/8cJbz6gueMD8EwzV4bJ
Dp1DoF29nh/7iNME/3ruCfCDcn7PP57vWwzR1xxdO+GeWOT/28HYrkMn82QJMGI9+YwNUP+4mEst
7Y7gw/zHfcl7w3WJedWjJ0WJfFw4hQ6Fux6OJieEpmv3Mlhix4JUDE8iXurL5xDkB2FnF4ezeUV2
P+mqVCYNBYKRI426uVoDAec2sObD/vS5TRHuaH2ANg49OKJDSheyYhwek+C1dxQezX8FhxQbIu4=
`protect end_protected
