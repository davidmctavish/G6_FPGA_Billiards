`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nvOgv7ZCjWXhLig0DqIYarjRIYNMgvBL4t+RjnW9dPwbE+2Dmh32daQC+cRejtTj4d/pTHalxJ1U
DXmEK3skRQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e0ToDGmlBj6NVat0a3pVKyDwHKrzEA+UGHgXhK7OQgn7UuBvEGNAv8O1095qSG6Z7Ap4nUxIQGWO
HN8W9LyttSuXrYZwxN94RSwh8LTpJbvnyIYi7UKCvxXR5Oy5cXr7TEPpgeaKovipUGiYLgfC2CNR
3uJz/3+qMM7torm2K8Y=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fv7qg58PT8m+ynJ9+MpU/vfVq9t6OiKELULZ8eRfbgNQi0mKRfhO0U6zpHfAktl8i6biNbgdxqUE
lewPF3GZGKzH2NZ5CAy46Ey6BU2Uu1o6ZRPZPAz5O1c4YAafngpK9GxjijwiWyDRgJqYlLhfos+1
TthFnUdpgqsAoQ9NtD2kMZTv4trJ39rcXB5r8eqdA3/HjWFo55/0e1t7me6QYGbO9o4j02WCJ/2Y
CqdYVsXDTWfDKKuct8YE/4EnDinZv5ViFX2jT2xSj6HRofzKZ8wBHZo1qFMDOMZPAHxGBF4o16OB
G6fknQ749sUZkcDpaNI6KqkBUxthfVzLwlR7JQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vFoT66pkN2So8U11U09GK3GCMg3zGvtB6aww0ejFwkp+kCApkz1FUtfoW+7OurvLGha1nuizzFy6
JHqpRCC//bR/aAL59rW5bZvtLumUP/OfHLcpog4o2Jkknfgi/m4keolMa5f8rve6bl1KHM+P7zCq
lswSgclYJiDaxrvBzjQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmbUOreOtpRj/pbzJmDDVseOMTkM2iF7LTkKx4RCEXFMloMUOexcSsWaJjsuaCTUV4RlVxayjIKC
1Eu+tpQLZ3yTZLmqyMw3/94wD5Zc3P/Wung6Wut7iaMBcAD30CTI2i9yGrWoZvfm50+oD0lVDIey
yaJ7Rys9XXn3JxgaPWzVNJcXcFQajItPukj+WhvVOIdv39b3EBSWI9tNjZPLBLn8ije+c8Wgd8cu
KSmWLEix0GbbgKyTg3tTJ/hLjsymY8YrqsGzog9pkhMkWi5q+ZzJ0CzxzWzOn+s4HOFte+NKmRdv
yRVnpdnX0oQ28bUB6dG/ePjWYdVfyAokL+Hm1w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62128)
`protect data_block
TpWOUvIS01QcBtrl1Df5IIHoJK5PclsDcJ/CTJTC/6Fwp0CE/yDy1/lBl2k2QSeUM3deDGc5XAL6
78SISf6lHYdjiUXsjQcTu+D6tQ0HgeNcCX9jNN0SiMDG9Zy7RPDUhKq5j/badURsitf0c3QFxAgP
V1yyqEEjt267s0RqjJARG13VCcp7wsS40FsmvJE3gUSG4ds/KW/J0qPDdT3tYfkIrfEA+ysNP6Tn
qwxVE+K3Iyb4DCWTqrIz/6eDSmjYZ5AD/2EJ36yxuytmcEgLHBbG06hObTl5xHi5hHGM/wQtGxqg
EPDrY3jKdWgWC8XsNwk4kxWpeIOuxnxe4z/gt2KMovE54MvVl4gDb4TPsfd4ih/4gO3S7dhBqrIK
oTeE1mMUdX5H2sw97Mhxo+2hR4jIu3GgvbFagk/6u096b5f2OP5SEKDT4Z8w/HgV7YU22u6rMmhg
XsfhsmNCa7QJtVakeXBso1pto4wvi5B8wmbHdR97XNeeMumybiFOMyaONBxw3YeB+z2TIMSpCMee
YT1jKj2cS10fsURnSPEjp/+UvWzFTrPV0fl6VrL4VsXu0cto+m9RRqxFyZEBpKVbpCV32wxsm6ni
kGfMrYKUC3YsrUn0WXj0Vwc1VVFtFkm60tHiUU298jZr+IaYeZJbwp5CiYS8Be/A03jiqUz8KI+9
MCjI9nfrSec1Ji7gAgFABgQjXFQz2rT2AvqJgvFL4356ysAGKsoss0iwAY7I9SDVpj1K5Au/JWDw
NUVm/4Iruhie8qbgXivFa6UXkjdcd4BNy6YNITm/84BNyKYF64kE0wOjyCqv6NjAWB+YJzkNkKaX
dMoDKOmlwJFmzmriR7NHvjJ3APidzXGyF5eDz2RapsJexNyB3G1jsrLPkpjkUdNfIRSpyGVcW3cL
oY0hqQvTfctLGcap3hchumq5jEb/5Qvy8Z3feHkBJbjFyZ1B6uW5cz67ryzLbSQZmc3lJbOqTAmb
/3y8fzg/4zOSKzrHKj2pjVkVvZ9L+FX8bX5GHNKUtLW/n3extDrEmAyHNCZbNdUJzF3xdaMi7HFX
N3L3uQeaKkGaTKj+yofhdBPTZWZv7gGGHWktOKGCtZgwaY+xEfp131KJkrSavHOkaIDwyjINrrjF
uB3AafoFm/R0pFJ2uUdY0gosSE6nXejbf/ZdyBDwKnLCMqY3UeW1fzD6EBdl1jEbb1rUICt/ExUj
0KW2u91A8Cftqm5s4D1/yxwcrMSwHmSetNuK6QuJlC9kcpEnnZAZ8bVjj0HCtrREWGLEH1ZwA6f1
XaTAbfLtzwhzeCyVHNPafjE+eHsAyhc9CaFEo331U9NNCmN92kps+67MCBewkLQbUsE4Nqbi4rOP
z+dMWxVRIONldZ9NLUJqa1ndKfu/RiIXP53RwSLaxznFlKd7enUoosyP/D68J79JCxLqCvt2l1u9
VAlMZ36/Jnw7jCFzWl2EUNOI3DaqmCUP7dt/a+Ct4Lu3sPKytuDJxX815TJ+nPdN/ZE7x73teGvZ
ltgsRWFre+A1bWMxqmsOOw7PUX+Hg1rZldSrptzxzOA05q9yFSso7IIGAuRbg+6YT1JG5kXfJq8s
Nm1D3Q0zqsR0tItdTnh7i+kKhkQ7lu7P6A6xLNeKUH9C9vZmyrjqA7/5hQ7Vvgy3AO5UD3r94Lw4
YQrL2MrSvqfRxMKxuCYeCWi1uXPwkTlB8ry3apAGZxdVkxslmJa+4rNlgHf/sx1O/6ynWS/PEemQ
nu3IiI/+PQtXkfSGBEWBB9AV5SbwC5kbviBhOVqP4j3F92FmgOf9h0lJ/m4j/Xl8qnr2SgLcdhKj
X9gqbwcYBGMiIK6a4wnU/rBgH97gzfj4w2DWsHhdnbl/nq95OA5AYLo3pOkufIytskLDitAlOTbc
8QwcfrqqQ/RpfxzMDO/Pz+yyJV89n5p1wwRMxN/fIELAXyeVivpaEfdAnzirCQqUNmGl79/rN6l0
F2FYqJNTYsxdRpEZsjU7drDduiwhMF+lx028XlghOcP7iQj3EnWNKBR26bq942E74vCxt+AfNaLi
KiPQW8myUz/lSzqJ2/aIkgsW90p4+W6PO1kbb0EjP12ooqDnwaMUnCjCsR6Zx9ZJLuPxYoUuNvRb
JCmU6U/NGvK8X+GCtDnzt0nxe9BFwsFT7cLQ7Q3aso0omCbn9yEJzFm1PSZ58iq8+o3J02faJOyx
mI3Ll/ox6PDXxqXSGf2m1LVr0VKhlR8tKoOxZd6EeGcpN3UlfPZe/rGsI32B5TD8/rJqMRbhAJXE
e681aU5V3VjZlqvLTqUbYcd9gEsxrK50ssr+SzfNDcjaBHLWdAcmHjKzDd9QILNvfbvWWOFGQfDz
GE/ywCaAM+KuOb8LqLviTP91u18svTv4/TLQQNugBTjDkpPIBCwVYoInoTukgv09FgZnIj+D4viy
L7VUpvcUNL2TrzrA4S/OErsvU6tsLOhkQ07+s99k1Rm4pZEIldGFxq5qWQjKLXcHrncTPz0sWJEZ
GtJL6evE3WbzbURuhZOhq+fLP8SwEw32vaBEO2GqJVSkUNBF/k/x8sIbYHeDoZTZcfDVs+AkdR30
/aIZOeNQ5JJcqf3qTQULI54EEqIsX8yvUvC17mukj3YYd+HK+9UDsWu2krKvjwB94+iFUCujfyTF
cPAzvO5Qi4nOSTCvsoJKVNjD+3g5LlAVIMNji1Y7eSQCKFs4RBZX8q8gYNJWj/F7BBCXNEESaSbC
42ASvPvxOxxvkcCtNaxa3XyeaP0ZH3nQ7HstTmbB89SG62G5qm3KNxkCBCLXmk2E8kmiOHLVbIuU
ipQFZ8pq9UofgA0zhR9XqcNTuLFvYochud2aFhrKQtogKm1pUuS+7STsHcpsy2Cu0qiuHOifs6Ug
5JyWo8HD8O7Z72Azou6QQzMkIvDBYFa4NLmWKfj7R6H5tkgTDU+dHgVeScLDYFCXaHO+Yc9+S5oV
sZUPdIuzIeoOcxqcRaZs8udt4AEzAiQKuwRr3D1Hze01KFAFQh7VVKT4x+l14HiPS6MAPH6WBwSI
tU7HcYKOQ1iIFQ5pC+pxST/03sOuLLRh1ZfSQhsLoGRMg7OB72rW72EKs4F1V2WRiWFtp+vhDpO/
n46401ukVL2n2myEWT1KXotEuwMZ66m6UQN/mFjHKDDNvQDUmW8FdENobvailStoi2/4IDPgwnT9
hQnHcvvSurOWeAf/f0A6wVy+0ARhkLuwJdnkQshkhsxEaNfssNEp3rxswJGSf5MNxfq/Lu/mLt1X
m72MuljlmEMW9uKpKW+XQurFWdIXgGfeS/BszBuYJXJM3UQNz5Ex8q0FE9uBbt+XouLL8pIUwSHh
MYXhc26tdvnsvyOYAmMzxF+MLKGGVNiTgy3BtmNu5PZHS7yfI40tY8wOzSRr38NCBrt0EGPa16qe
D16oS5guhDcyf4A12s+pWlN2po5Tfo/vKdeahcN65Dwfe+T+qH2QyEPl9E16u29NMEZ/psOPc9fL
LX+OLgFQ6gQhXhmPGrcju2iA6X6X4972VnJkMssMQnY8oL9ng7PTfDaVNB6inORPWF3/1DKkkUGu
kERMotPzvKY1OC/TYh22mZxwaIrVrpxs8UIxwWWyhSFVg7LSwbMdF2j1SAov7+OJHVZC+yVov/9/
8nStHb8yKoLZ4hXjJF6HsI3HX6/BUs0c8qx1xe9FDIvAgI2CYU3sAqhvXZh5ez8s8itJ3mCEMktW
lj+mEnn8E5s7wz++7h/2BAfUqnxhMIEpyG3j7czX054GudDPQqJ/XPpMYhicWwuN2reOTRJr/fOL
lfYfCh81iRcboKv9jpR1G1wGRAl+PJTRKsh6elh/fVygiDHwvMlSkL5/TtHyi8GWGFCF1fKjtYoH
lzV87k9IqdeYgoe6s61HJOjNuXTP3N1pxK5fleNkfcaRn3VsfGrHiruzXw3r4w0iTMT+2QHlH9AO
ITFWGSaIwij1dasfjFv1EsS2tdYCTwx+J9OMm+OoUZBs0op+DBq3G9xR2P0tqW5hpjPa7M7+SLRW
jMa8DMREGFmD3qlgYJjGGYlercW9dCz9jn48Fj49KKwDb3kJAqPExtm+VogjmXChph9T8U0EI1oR
/d8eDkiFVXtkedmQT2lp5j7Nqk5iWiifp6Xj9kYzjuiLGiKKbN8XWNdknw9JQNvtbO2Tj5oSyEYr
XFWjOKG9ijq+WlNVm7eW6fx5x9pOKp03SB8px1/wTizxmq+v3oUxmgeU66bzTNaC9psjkMHZ5omM
LaaFm+fsKzuad6ssMvqAjF+MiiGa2kR128g4cZtTIdmTwinFnpuFYBTaJJ5OVPQem6vwIf5xvFY+
nAEvguIkVx6F+oMbhQ+YfP2ww/cPdc9MQQxN/0PT+a7uOrf3vJWYqVYj2Ei41DSj9mOJqaqrlOfS
FKfkL0d0EABGKZdreYhvLrfCk6Gsl6TgU4rKDR2hGPTIkwPy5AfEcxj7KSnUw/hPAD0PFHvOntM4
ylCTF7vVqVDQTItvHaTddMQ6C70slxB79v8zZ4w5aukct7CqamuWV+DD3eSNK7aE2y+XoLVEuZ49
+fDt7+sFE4l3GJDoBUVl4qQW/fgnLTSPQ9gWRFBb6bobajH9YoHXMLOMT3iXYpsqcQCjZs/nJ0cP
PH+YGbfDcmXsmtQz/eRJ5Rgnuwl8BUP2jRtl2ENyci+s//o8wd3rIysO5puT4XBWlMTvVTrhd3uC
IZAZ98qTyMTfSCaR+LPj7n3rCct2/vOebWm88hYYFjCF1CBfts7N9mfFFVR8O5ju0AB5FsOgw28+
SM5K0G3Cev5gZPE7n91ycx1nSwfFB7HQGGB8oqvKPcGywjCRnCHxYw+DEw8OFY2IraQ0APHhJCUj
4kN6u+Crd3mVtfzMV1e98fdUUQNOzgGLcpO3ui9gpnA7CU/rBq0lps3inJGkpmOJWOk3oRYShy/E
f7qge7851f53qbuRHptzgGuqoU36x7kCQ96m1NRAwf1hxr5j4s/M0dRT2Ir6m/6h/PsaWx52za8k
yJCrACVmHM37UHCzC8SHv+IdTTJnDMWeSeJtRnak/N5LZ1E/Mn9aOA2T4XF0F7Lq5WGj+6NlnLAD
8+qCuDhySE51W3m1UObE8x5lVSNH0QDwvn1iWEHPAK0Yg6TwdZIDxjkNt9viWAiSS8LlVLxDCUsU
QUtuUt87tRGCD6bdREPGV7mhsY81HpU8RUnz0CWvzekf93HOjq3dCPsZGXz/t514gvcYuY8tsOwD
/LB7StGoEK8qd8QrkewD0PxtjjnCVV/TZe+Zps90gYYlMxrCJ2juk00atlmnjY4SxgEQ2qrysvYJ
OFRnDfFGU9PR7+Ih8vg5XtzwRL7Ezvia1gIWq46RfZSXuwQheR3MXwmnSMgfqaTld+f6B4JsqmT+
DNlaKZWZKAUnkjkEBCaNruDyYfhTOC35saqLge0OsFKfwP3ZdVkLexsw1BxCqCmQQ9929MlhrMK4
yDo5+/HYMYER8xE/7ZcS/QBQCUfc7deef4ioPqMjrj7y4H412Y6pb17zDA1KbwmN/g97/jyNTtzN
8S/vZ9ELba8XvuU4mCF53erIynYHYHLM0D3KHQq144pnSJbJ/TNwVcj4bus83GOPMVi2ku6b+Uhh
KS5jiBs30PMQh4ltyYQS6pbXrKpaVrOJr3AexmKc2RpMbsg1lXeBw1g05rMkfPs0PIgBfAZfK6uZ
gzZ3pX+2tFUSj5HC3Vu2BbTafMYdPsqKpuYvpP0zxPRvmOc20K/wfOwFQUXZBmQYahsa5HpEkHq6
HBGZDE6Q10V0oCXf5bg/j4LrMQ6E3TDHnNwpqGKpJz0Mu415lcDe58fFY2GeO1eOzREA4o9XYNrB
LP/2DdGdSfA4iJonNH31wuOccmPyEqMSlyw36G0ThSHQ0rNhmQ2J6OgIzTvP9QaGHqt3BEmv9ii1
iQ5NGb7ufUskjKF4HPrI8KqRn4Tr3GjJN76nnsNpvC0OG+pRwSKVLwcOpwu0IQe80VzirYx8c2qy
VBcYpPAH6rkta9GXU0dVHU/nM0iGQY1X9sohJe2/+tShvEd1GRnsNl8gRPlHM29YPvEfKGX00JHz
aXrOaSfB8eRgv8hJqGBV0KHifXhqZS9m3nm3/ohjB+taPHdqUxacgd/xNoaynrM4E5nb73AwMdIC
RgDru6X5RdflxZGVBOKx7JZz90BYHizn6MgNAtylsWG0eEPWesUvE8Bv6nDn0H3UXEZUNOUbCd84
egwbiuTUdTz5Q0yByvjRFq2Zs3hL7FYwPVnnUSf2eVRhiaa8Lvb7VKLJSXe4xHTk8o+RmYrZATJ0
fzAtJAbMZiAGl0fl4/bZuS0snSOo/7oU/fZHgDPMUYHNoJu7Wn15g+/joWl4WjelInjDritH0vME
6QhHVCMslsxDG3RMVeKlii/m7qljTIeNuEgFrxMYxaSZO3lky+guFhaXxTiacJif4xb2GEK06EFr
EpDJFmndB7BcAm3NqVrX+D3IEt/+YqeaU9mU343URP8PGZkp+2RNrcb4YFU5L5LTt0xOG4DH6GIU
b7l1cdZGZLtvNE8eEgxhm+goohIupNsyZMSpn48FScpU1g86pHlehPAo1Pm/RfRvMhXzB46d6vyj
dRiUunbNdTaPNIFaLaS48FPmOm3jDL/S9yL/9hVp1lXAJUz8JkyYDUxkzM08igCvwgXrX6aG1Tks
ZDiVfVFh98Vuy0ltSvF14cdJnL7mJfkAzkX575X5s+hQ2S0mRSrdpeU8xGyH1ZMvBu02Cc0ZdWi5
87nSmfJuvpAO1e+tBpOQ02XMWo9TALlfgWKFGghu6vwZNhXmW5WgJteuc/HTfWHOmzSmizH0ZJLB
mGjFAieNFBos14uKgcwrkST3hJCMxwogmNrVK6NPCcSozXOp8VfF3O1kt2CfF4K65XHuK3SwRJkp
Nz9W+Qu0C8/zRUwQiXDhDmEGPvSe2u7VKAguQdQQWs+SyubmytXl78/I0LehzZLxQsuF4dOEjLKJ
zuZol4Q3lke0/tnNzhuvaRdqBq5Yy+oKkeLo/DBfKquQUpR2lMFfnLS/53/d5OfvEEhKmJwIpxnV
Mp89ABG/vwMM25WsjrmAGIC2ILX+A+lTtXXHuNa2Y0Mei37W9c8kTz62OOGSF4STirseiVcSlGV5
1FlQeYj2GEtnAPLcPfVJlo52lYDlxBuEWfI2/KrxQZoLyu8NmaD8QAa3T6Sl/rVxfpwTjWghDLDF
gIyJ8vy/Qg4MoINoQkBGyt/VqCPSQHRxz3XQeCA5ZlQ5j7lJHgTZ9jEggUs1WIWTzILI2aZc0j8E
7s2YBEJUenXDk5cW9wTJ3uG0Rt8CpDIZmXJTFETXvQenSmcQccDDEtlmBuKEoaOWmhOidHjjzILX
h5C42ZlGKEwAeGHXK2qVtlRvwbW+dfqkEI4cPAaR6uBIhaGVRTJ2n2oXA/Ypq4DkqJHg+9iQ+Bvr
Ti9hyWmo3tiR2VvE1fJiPoluzn2XzCwJc2fF93alZvOkUGknCj9wogLBZptuXBUn5NZSqQtU+Pu7
OnOHo99s45qQ3d/GlN2LaY+IT3rWxoAL8g+kgzWpRjvSqexsnWsYQP95QombsdsJAHCus+uTaAX7
35ygcy0DACTo19BaOp55f9m87VMBk7yYzl78XbC2JS6yEIsN5rv7OdaZCTK0rHYq/dvazEsa59wq
W36Tkr7SHLAcIx1hssHI/lBsE1dRlsJroK5jkhzCH7NCiQYmif9WF4NcEWUn0JMuLFeO/qICDcHv
Vg60q3+dT1yx89fSFXrqYRhi6iawMF37jOd7vwdJvIItznZD8o4Cfzd0bGg6zBaglZevDegIHsso
exwYV7cctO7Psn6m252iuZ25WUgH6jWYg5ObnaB5XzjeI4nHEvVYgm/OG34Qr/1UoivbHWmRIjqe
17twgfct2lBtSznQr/TJfShrDMfM4M0RXvvYN7jEKbDckBbfRsHE2bc50IW+13xWZ9PERLw9mZ1F
BzivycLN6ofTE25YGlJd3mYg2P4Gg8UB6K4KG7F+bLqcRzblLejD3e3osH/1KLq+4Htxdodg3RPm
vz+FlRI/kfMnOCijoRyjUeOk6Pvusz0nYmYtYlA5I4R6K47+C5fa3yIHpzWsgq0Zva+0UzBAKZL6
MzPuA6nMfodaHs5HUhAhKmwBp5JBNbgeMbaG6LOPqCI1b+hsLk/0cyfmtXk3gkD02AYcKOOBpOtu
QZVfuyev5JNiYylzPHUmvpszP4jrkfeRlXlHyoa1qnYTPf/+8+UK9U/w2Rnod2WD1b23PJFqVuEW
0E6zudM0qW/Z4YluhWC/3lG3ewDlvWM7F/D8l3nqDgFoYyX2jwmzYrUwQmtbs9pvs2lY6Xa7SjDS
X7dmp8luDpG7N59XHWJk3IG9lDSEc6rEkn9Vw3a+9ydzaz2DhnUhn1F+Gn0AEx+CmhHGuNWKqpfZ
TNZRTqtP/lsxXIgseJlj19va7BkKtC/+omO6sqsenC7lO7Fwr+bKZ/QTiTfMDKn1GBL8PBNexZG5
9qrdjFj18O+E80AkKblFip5RgwVYtERlcsxUwv+8q+PGZ5ps9QvjwBnM0hLIlclQoSUUNMP9SSI8
HokVq0fjgc16tHm+pkJbTU1s1tDN6QwGRnzPGVF05B19znIf9FV4O1/Zvj9c6xh3R6TUQ0kI4Eh2
fSjOXP5dPRioeB8URXMxwva62k6vPinR7QGSSqoP9LxK2h9JGfrGoYcD5jBkGbgBBGLq0M2bFz8y
JVrmRcTlAQx08SP2DYcmtD29cTnSVFDlV/Us0dnNvH7t/SOUfSf7Lg5Cx5dZtVxLmH2EaIrWgDIR
261bcVAMdggemUfEKVj55VNZOWU/WzrTL8xF7aAzIL10xS3PmQaba7SlhhzgNlKcmnD3kwr/V75v
7FzP8vEXEiCIIIZqb/Cud4xfuQP1y7gPwgKEbnAISxJHJxUtOsXheLQXAPo+EdWpsoln3ri1YZHw
pbqvoczipVdPwr9vzQuPKDGUy684YMdXZDOwy/k6YtSoAKQwnKA1oyOyP8NE0ITAygfH4nUZaOIm
vrz6AggfJDZYU9ZYg0xER43cgrCe/KKAllPpcb0GdnDykNKs22Zp/9rHVAkl1yoLajIY70FNooSB
z0esZMteX8gaxve427I/w6U0LR86/SQYbNCD72Ysw2pazJw2mi4zEIrjOxhCuYtaS0a3yin9H/nf
mgnW9DyPPerkJc3J3nUIl6HLmWaxw26ZBdkOBz5pimg8MeF69kuDICyhRu2vRGeWLFtlbNigy44A
KoTkyYMwhRRXJB6m6uEktkiH4uC5RpERz9OUkySUlQRG1YtSgCI840bNY5Y8Lzoo6G2XJShjcQBa
vMQ4A9JGWTuSlXAFUTEjnCnbxw0meWiFA3CJBDkmuOOrgnDkEg+5Cg5gJmiFDdkci9/hG195GcJl
qkq2L59YukLAA9aUI01bODXB1unlgUsHB7wOJ3SVpzzKdpFgDiVVekyVhEXyLazQtqfn1UmVMou0
KjtITtIvLd2l95/V/fJoKNVKuI6pSwgPCt6zpAMTt/JAeH+dlvVXHtDIaxJaUycPx/QwKFtpUB9D
ur/agZCzZYsDkXYhA3tD9E0/3IozsGbTCZADd5Rpomt4CP/T3VOak8rJ2YzRQT7nFdtK/mky5BQt
YzJ/MIAc8L0vJa5tLMMRucomuH0NyXDCXbOFtrI52g8mpuMBRo8xqypt+LleXx6c70Hu3LG8N0xh
e0yqtfS1kZtItah4R0Ijqy5/ZMTme6GgkfZ1+lBFNvNCeczCQA4S4f9naEvJBRfRKHRkyayV6drx
K+2i67ZWfZXCXyfeVRZvBbqExLeX3k6CT0MUGpUCcMV7yBaURqdAvUVK0ly7OWEQiQ63ILoz2goV
dRRpqOSGjr5tp5zYY6AgXqUzqd0i6nf0LxdpZ34c/cEP7u2U6bFW+M1wu6283HJDEme5yGQfpxfT
SnYBNrSSJkfVKkJrcGpwC5kqaHgT/WN/rNMvJyUzeO+qPMWkDvYe3PN44sMwh+2gemG28WBlBUgQ
6RYh1NSKeruiPW2MRREJ7BN/50fjC/ofHqbXMEO9ItUxIYBCH3NLeVsAyYCsaZmnR29+BCXE69VQ
EUIw6qAbjxNhigiiOdFrQPDv2gySBj93skaZm599SWC7gBKHkSgBitlxxG3ts49/10zJtU3d3dQs
nS6nvFfiTMvZl1dUHgeX8sF2Gbomy8Il5A8as3psKnew8ga7akVKAXUaKDDJHoz6C6K++NRC5q5y
S5zTLT8J0WBMp9dhJvcosVmlmXN08OOEbbx5fAUJFTJplb0EYfgAKi+0nxX1zxpDpTC1VkFNR3l7
yI3+D7BOfMYTmKRhJH7jgmxab6Z2+l3pwBX2iBRAlPn95kZDT10kB1U+WijJc80BK+LbWqLXaO69
Zyqi1el7zd+fHYG2mRC+bRdK804NU8948oIoYcVVSmq1XvZo87TgwM+lIrMSCzZKxyrnxvfZSaPE
xEhAvSdpD149bPuwaJr1g98MXMMBjq9BDG1Ai0po4Beix8mXpY+yJbwzPYGZ+Dvgxzw9vz3cSqwS
HhkO7vSl2mTAbVZ3WIPS2N/QrC5bYIjaAFPgYdTPzNf+c4itfiHya64Vkq/sEMaBLQeWOyecGAFH
vGOFSxkvJpeb5ch1x+DPRqtkHqemOYwMSTUqicbJxDOV6k4UbtTu/9gQRvjoINaLv2YSyOnZNSl6
f41LEhFVZDL7u7i+UZ5UbfXG0VljHK4mAcmVv4QJfM4+MGVG+gDcZup3xluO1Yk3sV1hFK96VSGj
dQENnI7+LRLtyuQJxOyWPdXUw3V8sU2MKlja+2Djws1psucyewPrfLoOyZvAiRJflwaQFUnbyKBj
agPHsOeJHyfb70kP09VLo5F21SnY5uX7l/tEFEoE91q+lLZPAMNKKd51ZYtkXM4npxzSAh7cYCKP
N51BJq+owZx6jHRwFFRqsYJwZ+SfXVHh6V1a30+5ysWe7OIQc0mBPGk2JN4Xdj5vDu25wrgyqMLW
PCUje5kOd+F0/GcuhjGnkV/SooVffmRd9z7DSq+2NvQm5Eh0koZZFi5VgsOAOH5U7V5Avb17vmlx
PFGhxHjx4CWqC+EOZnUaLJ5jB3xmz8W/NMAEVjlGO2O/otxOxAkEB6Hcnp0Kcpvj2PHR95rhTZMp
mc0rd1j3xti6fGerzI7W3TW8etyU4+1E6gq6CFoBPcoU1D17a2x4QCVQeLX+1OSbeDtQHJToOf3z
NYO80/nQGMSAoMYewUvafzfoLHfWq0oExt2YbVhU6Gxxh4EHP0bzzxf2RNj+e/Om3/gGp9VrUrRc
45p7gmp++JX73cKnGbhbcJyJl9xlNP8k6ZVfMdSON6umHpLUsrA9nCc6RrwqMCIBrQGmOV0DEMJp
01GutfUQmXggU2DqPFeYujsmmuOvO8o2QK3QNEasTWB4kOI2oPzNZIVlIGI266tq3yUDasM2haKj
MPr2qeGLefSC6M2we1SbNk5QxHq+0ZoAa7tSElysN1cF/pIRjDCRscQTR8f4h2RbHNvKQcleUauo
RLOTD5viPhwGY0ZadzqZDPM4U6Z6zFQNphGbKOsM3xHcfj7REDBi4Uo299KCTvZBMKl+hfv1mOnY
Q1Pw6ByLw4N4iSS8aAbRD63o0h3tin1mzwG4GdeU7Znjn4w1JWrUv8r+ATzIcMFkbVWPF8NTJAwc
MqgpOhlqpdipnA7V6Us855Ar23kELCL4h57w4YgoVw/nr+u+bvwcWCMHARDG2MWnC1TRiC1yAt7f
pWnR2goCVminhOsehQNtlX3aAthtv3Sn2AfL1j08IgAKxDulgFtrS+O4GzmOJ6ss6PvNHQcO8UiT
rdoQ/LxSKML6GR4X79OGq3dvU6VpNjbXb/nsMgbWj/cDjZn5d0R9esphOddZmwFChIdRpkE07zuY
0fzw2asuudp16DXZefpR71zXLMybjQFd0O0/Yk/T7ncBDv9LjcUrSLiMrzowYdayP5vly9n5uqsX
JoeijG7GWkfFxGwUToGAek+ygKn+xsLYn+RHw8V4WICqGXiUONAZjhqpGXF+eHAgmDKStWZNGDnQ
s/JuOmm8EilHXV+tTakB0JZUjhzgzD/Xtg9XwbS+J/h5r6funo2gYO2uRO3R4hJZPr9Ae65Xq7LD
1CQMMFLHhoAur8PQQNCAEYhXyjRhaRsNUD0AJccpFyCnZZYOpzvLYuyepKaG9tbHqGD5XENy7r9b
HNlrnrtB1tJoXxSQucJqmOdP9gE9cMr0rUF8kwwrYT4156IXHumP0iugSGH7cW/cGZ7qgQejLw//
nJicdFvzEouykzLdjizolDkkNjChliuLV0gbQNMhCjXvKR2rBg0udK36kvECR36J/irzJ8SBKAwc
ORra+hPZ/lVMS60o7fWJCKYqBZqvLQTKdnXN6fuvCZZuH/lGNXcQ6CizmltcUSY1WNgK8OXUmsXO
NDdqqiUyMTcRzLKMKISm5mQMvPnBgyl7pSdskTcIzm1X6ZgQ4oo8fkv2aAZ4L7RhiUWQCmPjQGXq
MzKAyLrUXbvouSpbrQU/Yty2nQoCATEBDRymXL6b35FvPbsK8qdmtFwsi6iNeISmqD4roZ7+4OIp
HFtCC5VyUlDRj69joknIDWPaRtj3GervW0qiyaizvoUHOOyyB/zamavaiWc/L0Q1fE9iWhBVefKE
VTWxpALl52yKqS/cCntBMlrQ1KYLzG/AtQCHYt3Lb+3mOTvSjwsR4dZ460OLQ2HDRt3+n9k/dF3E
KV3HYRCRsb8W8j4tsgEMUCzIFt7M2yK+oLzi7sLKT7LFDlorBoGLyGE0SkKMunzhthSt4qtWW2SX
J+sbxIejCV1EPtfvrE/mcbW6+I10JisZ9B6fI/sNW2N/4/+DDvK4lHLNWFb6SAN7FLdl6JIhNx7X
5e+BxGy2m4nB3+/BX2zaUklnAg+jSLGTbLguaan1oZq8linpg/Xw16Nxvl5jenKpbvVsAYR8vvUF
NzizP5/S61p9a/ZtSwYONh4sHkUvNIElIyIQzqL3yU//o/SakzodWH58oDSnG/dyZ6PqPe5UrRx5
l4FaZtrTNy9CxNbx43pcMzHGx+qVgu67MeDNFZTvGE52DiFyxHWrrv5L7WLZ91mqsDvxnvnQXrrT
y3JeSn7uk25l6uYxnnAK0nC25tSnluFLi+ZaSKR45q63gFE/TqArqJCWWOnhE7jux26D/IQrznE7
7SLZkOnlGhj4IRnrVJi+Gdrj+XD7bm9wPtSzQ3Hb2L0uduTLCkidlOmuAfd8uF1e4xJfF3/Yts2/
a1U9OB96qnfCA9Xjl1SFjiAN8p9qNdJDguRSikZkFEVU8nxcYeRg1cMLFUhpPJQ9mOYZriPaiDkq
wLfejDCAItswS8pPGRD7Af5HiajL+tPYic+MwaNKgu68in61PSkDRS39B2LQa1ZoY0l+hS8z9vDx
HxalVPzPEOzoHhsix1LFXbzff0LMemzUTb1sabw9ZaAcP5sZGbCOBfLecjRn1TJIXihOvY7e/csK
IU/d781NSw2h9r4uRs4Kwgd11RpGecjhL0/kg0qQB5Cb6IEg3YLl9tLroxxI39JtfiHxT3k2UGku
YdLqw5ksIIEtX2H87+Qx5yzECwpqJ0R++8TcDLrUBx7ZGKMQt5WCs4oAxea9EaR2tMbgNj8IlslC
KnO52J5dAO/tkMrPriZTodjv60o97K+u5MbF1Nb4r8JRjgIUHCTpsuin0DqZLiahEe246YocWe3v
Vu3UFqVx8tXTKr11d45dy4jejIOWl9KutA3jU6tbg5vwbThUBeN2fBH8RBGR1Hf+IADtZpJOpxsa
F0K3dviJXQq0FeFD6MgP/kPBg3it41CkYILFflMqBsA7AVXNomwi8cxvT2JOGwSw6YWEr9U61L43
PMPZ8AazA8Tc5dPBLJFSD8AKCK3mF+jwUojwO/1QO18Xq9wHRVcFciHoraXHk+M6BaNIZjDDDvkk
E74tVcUjGzT33P97TupjZWOGdV/O5jfDB5Mrq97bE/MEA4G52zNchu0DvmrWTbsWm+KctpeQMh4O
QBUJimvklIbRzbm8U449TuwPyJSO8j5DNzKFq5ezdBhDPeXW52koiX0FzMY1cw90sNsn0Q5nlkrH
C+GCQO7N0iydNG8u769xsyB/aFeJzdw5L8Bg9qYwiaxlAnpdG3cece1zzvZgIQn7w/wojpTP3ls4
NPgZcI8mXb2QT8r1FACM+I47ij2g5B5vZ3fKfqipsDSrr1kaUD5BAJV3hMvdAWiTGfZ/08N7hBPq
PnUftfrs4SIXYfV3QMBu+bqx5OKozG/IIK81P+f5K46zed46ccUczlxRPyRDugrSivE1SewumHaL
WUyKFJQ+rNnxYX1LGSzO9+U6DzswQSeOxBB+IwviL0vrLFXk/CD5NQ4WNCcSSgjv4IYCDXJwF5ic
Vi0eP0Ko9pO/993RCZ0m26HK7R7Ge4PQAUlRoRluB3mhE0IV0xGOo89Uu2iolePBCkMOvQncAz5r
XdS4z8TaeQxOqB5KgYMsNbutzFknlWTZoFzsHE6FkQKKt62WfDty2ZCM/k+uVRpN5Zztdp76DtPC
Ih+UZZix/n6rfAn9ozwtajbLb2O+eUpv1FevZkFY7jt1mwa4PlYl5X003N7XNaEe1K3qotMFfZ3x
2nKgybPQux4XpZXlUnlOZpWxeLOhVARKtwWkDCXpkoE4un2D1gr6eKtwapvDhs2mIWMX22HJ/SkY
M8r5TtBw3RSIC7/3Y/j1p+bU7xb94XLCtRslvUfd4eiVd5dkDZoc+0IWOGHlpT8DCvfvwAg/Bm/B
/0fZxnPirdoooTKYXQooaQQEpp0m8kinBGp+SBBGcueTVstP56wbzbqKVnKZelYZXEwIydKDqd33
Rk6lBkYatpptl3i1hw5y5hQOESeKUXfO+6e+q2oibOsz9cGV8d5M3YTrkjbkLP9Xb30ZUtCjTPbe
C+s4jKmQprl6RYLm4jQXa2lLc1Q7PDtHrK79zcNj/mq5DuwnZ+fcfSGYSIrhgbdjPajVeXHXsVT+
4IE09N1ava0oFdkgOd05X1TE9QPeDqtfXC+S/kB7YRQzv+Ur+zAjxAD95RTp2dGOs1dDl+KTezPz
xtZI4kwgLU+vAOVCfSTDGoxy9RIAzq0cu0hRHOZzyOtM514Hz/AeacZ5p1d74mmL+HL41zfjs0Xj
IgnSkDb76bX2Do4/oeTLP3uqx/qEZzQipervQB4jwQ1NuudOpgXKj9afmRJFnOk+rFl1UPGZgrvv
86LobMb9g1tBdokYGS/8S9qP/HfGknWt3bNVxH1rjICz5TAHrKkrm452Iu1TdUM2NQB4SJ2bh5oN
MGKmkk1m/wtz3W5uy+E8nkAeUtqwd4gkkH7Q6zVHxmcLPXDagefbnoc3swe0drbLWTvu3dvl9R5p
Q81H/TpORV9PVZjO9xL2vaDM1RDCzGfpdMuq3im6AKp3eKNc8Enu85n4Ur4S24aMsUigBynA90EZ
d9k+uNZV1dSf9QUYt5s8JzHnvZ5ufiFNuSq4K/7l67qB7b8o1IOOBH88L5k/F+V5CEp2dY/9unK4
W6C5Dyz4f0Un2j1r3R+2BNf+hwgpuABkr+I0J9Zgfs2b2DDRdc9bWmEP5rw/OUIKWPJbBPYwoJh1
hr9K+oziIlPHcY6Feae5Cm8gC0de97PpvamabH5v7mj6IluLrfrjOZTBNHYG9sLE79x6fTl+DmsA
vBObAx0cbW+HJNuQWhRf5mbtAINHNmQPDIwkPo0V8fwPShiwNLs3KkwRu0fl0o0D7dc0EPY9m+VS
dYeTV/Oe+mTUHMc6TtbE4Y4rpLAUN7Q7mYVrkT14ATG/USXGxJ9UyyWLaudkm2hfsPLiT+OSQRUI
hd+ACpJYlrVL8QdFZCiZLXcixjc06nrLvpcK0Ka0+cJbOyeYsDvP0aOK25FD1KVdjUKbwU5wZk71
wsMHsIOKuFDzB8FDqEG6MMPN1QPR0WwY29fm9mI4B8YWBJ/q9v6u+CPNroSSa7rYjwlsWZdRXFsp
B5UhYHQ4J45RQtakp+X4axCt8l21Ygh0Jw+Da4BjIXSG2gya5CGxpxygmckYWA1qrL8uBVayRVs2
dNKC3g8UdsQSfUCdr1EoOawv9d/7oivot9RZ/V0X/dVFrN4mlJ2CsKKwV0Xjl6uxcFi+oZNFmUrb
IqEtpWapL+1QCqoHEcmlCYTyzt8X0tjIA7j9oe9YUwX/drFBPOLWqZ+MyOwmTg+FG9bVn1rBbC99
AYxC+1nFC95dvsQDlIOkhfSjTZU5Nd6YmkQGBYgCuTUVaxMmt/JXTCOTiNM7mWlT8IkoxHjEtVO2
YfCy/CpS2//H/taA+c9Qv4ykUB9spODLZiQQx+yy/TsKT/7lKJLKYhFwfWQAVKTg2acMjnlX1fJw
FWas+o5u3u0TgrWyDV9muoyPwUmCK7LxjWWVNyqQsjgE2zIWrJ3LHhs34o4Hwx2+OJEiUBwn5XLt
/RISwaeMJaq8LWhDnkD1cnpPzEBF88TXiwg2GXqhZYuUMothy7zC9Re6j1Z88z/w8homfFlTA1QB
57FbUlFGb9PkE8vBL/GBKSeKZGMVOsi02ZbHrml5sS7qQVBA100GWu8w4ujOFQE7d0f8OiINVhaZ
OlIvrATCMCh2Hu0k0W70HtHAtXtrLDrfbxMHYm7bL/9/a4W2X3Hv5V1K0DZx9+V9K5+wtD0Qm1gm
yLopvjUOvxbu581xibjPEsUK4XhoA+ukfYMJ7L7ENmx1wc0Ro/V1Z8Qqw80e1AoyTq1knJ9ZnAdx
Ml+ZnkGbP5TqBlfFjjT8/cVpUee1a/yIBZ7pViWCqwvtOKn8U8l2YY1rJvdbwJR2Iw/Wf6YVR3tI
9fIhEDUbOsBKBgEosw6aK6BCp+2mLH+YJCpLIN5y+zT1x3G1iOiADnySRkFDdIn/tw6Bf3lFEJ3a
gVPDin6WWyqAgpsFjc+fXDhxl/6KiDUhsp/+brDMAV+mhGIqQSQg4rtwj3MCJynbkIjArJ91kAF7
1fty9YyOOREI+YDt1Iz+sAn8TFjC03VTwubjMxoXqm8AouWqjBPkleGx6iCvHmBArEpNvr5NmIvW
yRUBl4HxY0yRtM6OGE0DP2eDnMPLXr71aUctSRFOp82Tjql2C8OWhUaDZcQxvjzghP0pXYdtXvel
i8UQQRblH4mRpZmoeed5h4PQCKz0cC2uMP3IOwwFL9Upydg2By6nAHJS67fCjg33qbwxcAZO5Tbe
8EIUw4defNzjsmLAwyCgmdHDFl3PuiBY6AoPhNhG8+T6aph5I3ag9TjShZgWVofQ9NyF8gz94ovq
dHV3VfSL+/ZKaXKJB6S6BufwPGM5X0J42xrlrtp+jfP+3DnSvuKequ8sdw6vp/PCqawTrSEcV2kY
oOBeN+nKVXBg7Xvzekt4AAmxablpFVYahrb7Ex2S805rBDESyzPbcVROjDvWw34PZR/W3pzAU0JD
P32FubZjppMSvfdOLeAp8m/M4VngTfNAl/w7w0xR6OXqJleszQmJGf6k3z0WNLO0Kodw/P7ldkRu
rK6aNGgwDfiID+l4d1mfec0XfttEbnTGwWtx7PfeRm6p+cLb6Vnmq+RvcwtYSi9jr3P3iWW8WpMu
QBBc3rGDeKAtXC+3BMCcMpvhNW3BURW8cx2m/SWfWqXgoVn4ImUwHe5UfK8Ix7YF6JXVZTMgQ6nT
t4bXk9+LcR49aEoc7fq/Upp/Kr0AzSEC0Ge/WUeDsHICnNZgYRWK5VDdHqK6eVFS+MYKiiS+/2Tg
hQv9ddVliU0yUAH5owJDEU5T8KOUOH/s2DOtefTBoAtRjfuk11lBKAALjsyuHMR8S5/L8fkv6VU1
wrDlaaprR3YkEXX8m8al49EqQHi9IMlCmyfR5c3iwZH5TTD6Y6xmw/Vz4BZ76XN1X2639j7jKYAc
FrCms2zbTt6RuTNkU/ovDf2vcw6sBfUFEFDsfJbozND1AVklbAsCGU8EDbC5P2BfWN5OEdZAvfRt
eBGJ0f2QgSIl6xFO+ckqh/fFnuI8m3rNaHNbKcQ8nZtwLj0dJSjxD3JiqPSVuplXFH3WarnxOppE
58s6mfV2Xae0WV6s/3CMK38qYMpWH+coOLH1SMRN686N0UDcYHId/Z66XBHbXYJLsl1/ADkG9xII
xdSQPWNY7ViSxka1dDzXEu8pBbupGo1UEs74TdH6D2o210F14o3h0wwGWLZjnX4MdsE+FMxjPbzq
f5UsMZ2yc6h9yznT8q0DsFuIwfl8+aXXK6woZxXr2RexQlalivGuEDUNtSOId4jrzxz2ZiIaU1P6
mbqot8ti+aAu15GqpjHpJbxt+YlKMU52v7MfKO2mohWq++Z4udQPlVFiYL7QK+00seWupSjppBYc
jP4pEjSut+8fh3NkPJ1DUDUk0va5JtjkFo3cW+zip52hNNPeSmbz31sTAxB/E4SrilQGb3sXzSAq
TIhzRyySKA+8t5pEX0oMWA7zwWLtHTkW8GSe5/lSWcNavf1mvOPLug9RoV9EFGLjg8KokVqkKgM3
O9zOiHhSmWSBrISTGf9ZHIoTCClOs0txDlDP4n5Y5FP0nUPoy0FcFKA4rpHVghZdNFxydy93TH+v
HAQUPj8tbjY3WoGSvC/ul9iHeDYSOQSjHSK7zdeWHUNpMjmuILhx83Hf7hEHHgeyYxpKxFyKWwuX
WqOV35lP1EVJMwHSaP6b1U/rMMWzdly54N7zU9NpgIUcBnYEiIQRJ0CqndQ1nJoo8PIpW4804J77
WxgqrBAXB03i8UnFvgsN2uFleggjXdJ6fto6VLIBJrRBZYu80uo/EQ7Ft1dpugQy8RgeWFkxN0Ay
8/JASszEkgWI0K6SEcEEdCDNf7uCse4Syw2XO5pbd5Ca0RL1mcMoWDf/1kgEAcDruOrUBOtU0sAQ
JZueVvk2HcrocdGnhAGKNJ1+saPr9BtFUQF1xgkK2oRJsm4VzWc59Xs8+2jz8k+NCJsFUTkWL4MG
jwqGuJOq5GRXGkShV3Dw4f7G3GXbVcVZCO352xIq2ArUHy8fRQr8w39OUsDJgX4Vx3b9C4lx8UkK
eBdsM/8gyAQ2wrOJb9UIZGoR/jiu51PKx0w7E0ptnGYBfx7cG+t/yPHUdhECvOGApNsksz+qI4Us
lPUzr1RD4tfbwMt13VJ6H6qkoj9+sPfsDJ81BeteX5K3SrmXPc6g6ZSEK0yizsIV9i5kEOyMIfmE
5hW42lzV3rQL3Rx5jrkWA+Y9t/1UrKB6V9aR2i8bTBQJPD4ndxfjHVbUcRiaQZW2smF0T/T/23uk
NllL0WVlnO7Gq4pqIZCMk5T/PbQkcsW7uLLQafZPGhSFIKKwcfispkBKUdRz+M/h2VylXTonF2RI
64S616WgHZZhQga3TCURhXZL0eUGJasrDMc7pC114IS77EyYNxsHqzkl5BtxkYy1NKBHKiseDC/a
6yC0H3oD8teoJn1SLBvKYts0ltbTffl/e44P6xlAh8c9Lghp6uhxx8bHlG6+kWSQoP0evjW/oWPQ
mSWlo2NWfPq3fpUsOTwo12JfS9QWkM1KN2AIth7V+7sBnNjqsnxtyx/TInOloM01wKcSzh+DKKbp
aukLiUUloDZ4j8qDFrPC0zduxOwH0c7OteCJPJHeoziIeEn+4NBmmURGMorJ8bHCfptPi2SpKT0U
2DKIi8nA9dLsJvxFiHMSFqRGjSwrMpMFgxJXM+tqS1qm/jnQlg1FCVa7f4+YkSVDsACrEowIspJb
6Xhc3nOay+5pmm3J/BWcFjpMAi5EFnQh1m+aQvvKaYIzNuPhlviFSjn/lpjDLhuRpu5EJfc/Dwac
wsAS422HKmZwR6cIIXwGEqQhNa4OD15HrFRWIoi3tW6a3C2nX4AjgpCAZeOTwymBMOoU1PfHyrPh
nSRFo0sxv4QU+VOndi0PKUXuG/JLa1s5rA0JZWCHF3G/6e6dFO6eeWvVfl176y0t9xu942Uj/iIX
DuyZi3/r/kshZ0tq/S+gCFYX3+lFsG8AAEChX2RmTYSXO1wSIqNdXPCFbZ09YFkVs1jdTy5wV7Ih
PlE6AD5xktAeH9pOQHW83aoBIOw/LsiaJ38wu5paLmj4uACShzV1l1AXWa0LJbmIkwdubPnnAszR
NVD3aABKVwWA0/wcI9ZbjV04FNFAcQ6WvImcmUMz1ItbKyoMgSz8EVo88yVJ647wO/usnpon4TwG
Mw9yjbZ8+BLRnVhRF23GN4uhcybEQs21geMAdxUtho98dlBpS8Y7x2iF8yA8+UHK5v0025Nj40tr
Pkr+OK9zyqHS5GUDG98uryK6Z0y+NkmX6B/AWDlu9DWvSUe7WJOJQhBsvsa1HR+dXXvRvYkrkzOK
YUC+Xg7uwwK/4fDgQM3lHbqTiIFKRrMB0OD1XXe64iv6XP9ECz6GtPrrnNDROmKVxRNd265+Fr1q
CkcYxnGG/Ovkivls7eoqAik5a7XhvD3efUoQRd6fHS5Ipxh6En7pZ/PNn+1p3pEu89v/VSXRJjnB
bY/q9xDjvb77t3aNeW49vOu18aiVTQNVFPh5kKMdy1ei/s0JyIEmueoi7bpJLztK+VxN5QxpqUCO
0XVfS3POiP3atsJ2oCJ5LV6B/lRtV4bRQRbBKm2HwmDy6x/pNKAJVWo7OFoYfs5EPNg89W+gPjwE
SBcCuyOxXZuLvPnQWutsdrjl+ekBhsQwsN1ufkExSqfCAlnEldyaoGeHldP3eMpb8s9K+98UgsXS
gamyRFWG5YZBn6OmoAIHJlLcfbX4DRoRsKHcfahjoqfDxP1Dc7Z7cHDGzeURV/1RUA5AggWVBpPr
4xUP88D3ObUb4sJeE1kd4Hxw0AmMHxYUxU2FyvowJB9EtCbaLcgu4YvihVh2VGsHW2TW6sbt3RRk
EitC2+NctYBX3O3i3Qb60jLu0340i0Vv1ZL70uLYZQer2fx0CkDSnjkdWqIg+2RxRL63niEaTy1U
hZKU1OxBlKiw7WOggGNRL/sHyc3ps/lhhQPxPbIaej/afqgz84xmd1+xxoJLj7S+cwN1bCXJg4Yw
mQk5lF1UwVWcdoe4i8Pp5/xe/k5VcwVI13Ds+EXZXbMy2vttIc5jBgke3S+A/m2mh++pfZCS3q0g
pQZUbuh0RmKVtMkCqeAHNNgKVljbS5T1E0bVQPefm0enztC5yWMr5XDXf6yDY2zZppEJPokiJJ0/
S+zfokNB8OiLD1Oq1fLpEmY8ctyZKcWBzgJb2/q3Jy9V0HZUCP+F8Yys9cfsaaKNTToqTZ0KqhcH
NQLBRsg5xst91N6FIRCu4WMDqKQc573Ri+rfCdU+PmQ774Mf0aM9kH0Dogp1CijSERqKBZmaCXai
dKE7T3MwsrObeAO3Hcf4lesD4rcjq9ruBvCgRHNR01RMX9P/naKbx6FnD7/NvnkxY7gFq1URKiGs
8OPDHqrLHDw7vt3L4ZiSzI0BCYtHbGFq8zp7ekjyPoBZvpKwdo+5s4DjR+ai7lNrEfmPVDGkCMc/
17t7RiwxwKMf3QRTFAyNCc64gtmnoTHKa++yefxYGLsilCVt1q0V6Y0N/WHT2SBXW99S7j7f6Fjt
5N3ttop64w6NJvqh95RPck9H2V3XW4OlTImEnkpydmXzCkVGwxshi1sZkCoCAjlPrIYXbHuOFMA3
9kuupqmz5DYiASevFty5kTaMKLgOwuUyrxY1CPdsGhauLpX4dlmlnc3dKheoqnhSnX1/QUmpUC6V
l1uBnSgzo5EYa7IYFTPPugAIqrIizipGojaZGgIaIDObKBWKiTMbpDT2xtsVh1qwVlSy1m6X1yIF
akZAoN7CnWDXDuh3Og1kThewsB6j2Uq/HAewFVrGhabuFoYBviBk93r53Q9fwwQV7jyL5ZP+NeP2
7rpHcL0mAFDw//uulUi5CE9vaVwjbjn5bcKUpIhtWvgFyvBPwacdKzF195degz2QoXQCZxQTqSCb
3+BohO+++axmFqHe/sVd6UxRM2wOwnxR0hgkvN+XrQPFx1MwlUUyS/jBmgkheLt4zAbBRsKlLp3t
cg/UVJf+bO9QzFKEpehPVJYAlJxhVmMPX3XFd+tKkZI/1Ajqy9CH1JMwnxlrurZYpd1nXZ9aL6/L
moEysqEHNYWOCadBYqiYQskHCrZsPZQzm8rurwm5WZWNDdHCrcA+PcPVzdBmOLP6hTSb+XB4CWpU
vPeM0fm7VMjSmhAV9rSXw0oDwZBB5CeUNt2uMK5SncWJg8soQqniBiNOxP6RFpFNQM9LupXYCgio
SxXQ9yiDwoQqj8UVwI+g+csimInzFWReQYowv5VrOtHbPAWI9KJLFHzw3ffFjzZJ0BJ7ErtqSuL3
yFqoPImOhz73pMYJSSkJ0l5dR8K6Y1Hy24vquKKmwJAcggjR9XniZx3mJXe12GgiAZ+dQSWdBdxE
9n5UhctzXP0QGjImlYQYuTCUy7R/WBB+zkLRrkj4XmxdSoqYKx0zD6hDb/jQ/VmbebZIt45aktMn
jJBRmpc1arz7JRCW2YckyE0CjgTE+OJHaqUYDK5QF2nBa0fHnjnwHRet0qFMXjtnzvZUeZhNhgcV
JWesOcOW9zzBMBtO5xLW0hVipeXRJZEq/45BbyKsI3TtvXoC0ZKs0JiNRI5LERdJ7Cm7Swv5D5k+
MokZ1M0+I0zbBptjwLJyGzEm0wo79SWVG/OvmQjJa+mtRT1V7pSK6k25Mdu2fMwqJaKhViRMhZgw
KRLhJwPM/8Trf1tj8jyRH7sdeVlHomcmsXswnVbEkTodmZ2aZqRXBoyFhlKjRf6M5+vTFmBu/2kQ
ygmQ1ZzSRDm7ArHPRMV9PT2DjbJOzk2GH6MNLl6YvyhZkZp3dwmxj5Qxl0FPjUCrK9RXeWJmmVh/
8wNw2WfI2XKLF/R83/T1GfqNxmS/pCMmuAEMPXlqMhRfqdsmk48fefucqlEzihSobgR6G1K6fnGu
2OsKAGkj5hTVahlb2THxY2wjn4bp4RLWUaFKrVV/OQcePph3wba48agnH+Onj239/n9fSl9kY7f1
qgzUyUrXFSvi4XXeJhtlA4zBhPxIwlNlZoQYwjPlzNsDD03LRcnbK7y62AyoPsWXwzKT4ynvzu9L
/hvSxhnGGxTnR1g0XTLYULxIbRvWYuxCibQlzErQ3fbF2vPjKsdro9gB18hkMPpC6HdNA1R2Qa8L
OkQ1xlC1VICmfSsoi9/TiDUZrWbuCnQXwYv+ao5tPoTCP15A/xXdPkT2Yl/v6YrGa1Z5ZXW6l7Xv
/xQCAgCSWv4gyiEQXIFbZLzItbsWIdBKnmW2TKMiMM0W9Qc9mWFVu5nqNc6CMOHcOe0P92j6Rjxa
BNiqdzHucUrP6/kt1033DFd27ISvhLQqNb+LfIC7UGnJP8oWbIKw9biX5ppnzLEFVshnSNTk4fKi
viIB3UCWCWe61M3iN4YmPOWoA6ZMbaTYCtRFRHcVAF7R9PzJuDtu2mf2Kk/jB3wCrcNmrYsTbvAX
QDL9zvR30JpcHXFfHRjHcGRW3qXkieYkNCXY2vow31fNtPKHlZ95UeH89TrGU5ptka0l/aAL1sw3
3I95d0BUYzCusORxjro5qc0W45sXhrfBJT8NVLdD/axEf5XkGHcpNrB7Et6CAbu7xB/4X28Oc4DI
XmWv4Q6qOLj6yr4gwJzbHwRBWjUrsVK33b4eGNGhZyNwmFQUjxAQVTFA5/hv1E4urZPPTV8XeSVi
MJz3g7uz6k1yMs2ceurW4nmzyd164Syxz/7SJTJCoVyYnUL2MxUPmfD3MY4y/2vd0BRv5xRB359q
SpQkZpXtfn0+RszIMa+GsMu89WLZFHDyqXPf+OuRFZzcVU3I8l5v49vhY9OLx54uDfskvYKNMwxv
LJUlK6lJXJq0OmMSDb48ak0bVy2nGKb8H2Qqmt1QytGAUhOtbbl+tdy4QvfWFvQ+6CJG7WnQ0yA2
2BOsCsmGQfsJW8aZiQpY/b2CO2Ih+mv5HessRPhZNx0RRYhDEGL7B0YGkUwALSYy2P+q5LK6Q4tQ
NHvNeXklv7o7Z9+9HvrZZU48h5LX3AI2RnDn67yozhLCYUeV94ZosfliUFONXroT+L6OJ79ic6+G
axhY3dCEhlQElsVyKgJL2aeF2gsWtkGC8bHqsHsykMjBJMC/f6wCUjYIY1ABvctB3BidpevRcaym
2bqp+Q5eQGRTzV0Q8S8SlrjjMdYvEFvD/mzAnaMDBA3uauqeJ1AmjFiEAT8bR4UeuqYgGltnsDxL
3uawNiR3Kq9QAtDZfCJvvg5nqPRJfpNfE4BFdB5vLdsAfrxsD9lLtDOjmZ2E6Mtb/JGD2d5dR9KU
KxsC+9ftd32C9KE4xh/qYAAH34dh/RBX2fwZ0bU2Gdn5I9Oh0naXR6wh6z7KsVijmjWkThnmNY3t
EGJyFxA1A3qH3Fe1103phusMNnBBuSgSPpMUSmGmPzyCb7Ww3XZisEO/ouRvIFHQHwPO8j79B0p6
lPSI2AIBADsm9Nn0gtFZoco2Ud8Mj1j1TWpKDV8mT/ww9D9kHHeTcjixAmLVoxbJGwVGt3/UhEFs
F/1nivCXSDkDbtd6XqX5vivGdSOMQaKA8L9ySa67rQ+afc1OWbreVnccY5/n4yAcaIsDAb7HgigT
R3XF/6TgQ2zLx7xMJ4tvJDgiz0mE2XK+BT/WK++OblIaiDH16kSprg2vbmbexFHIpQ6YI3C/QGoI
n8eexXvzpbmFO3qBQJdn5myHRJl5JUyBnnCdJluouULEIcIBBBQMGFs9w/fuFNGzD5okCHS2NZqj
flbubCCOJirZKDG539stJPszxu5yNqZd9EmN4ImBIxv+hjjLizEj/6wdMlOx6J2CqeWaY1DKjPTb
m+M+k3ZMQMoEJvTQ9zS5BUWcmEw1R6gsN+g77O6dGueo9qhumBLXodvb5p3Fy4nbvyEujpisamfm
ff0uIcV7N4PQKXtSkhgNwUsDPFVJcmInXC/T3uVrFs+b28Wsm1/iRWpf2ci5Q6PufaRyR96pQ3jM
K0N2Eiv1u+nyXDl91tG04JdDQN4GvRMdwFMBmKop1x4Z05NZvqkXjXo9RczkCr84Vz7X3ngur5Jz
HrCAtRNuqdd/ow/vCpaRs3djzJQhBhVZEw6eadMB7DbE0KE91B/lh7AsT/R8DiDtx4SebKo5oYir
nFYrGRvD+Lc5dcE0T2j3R3pVdN7o7noVK28vaHaus/7NWfX5sJ78HVon46BKORgxncLpi7rBo4gj
ehiVKWwAeBGbFrFBpXKq8jtrUBQxOuZr1n1o9pzY1unQ8CUuJp+QsXebkMeBE0b8ZfUgBebgYPdQ
9MfQgPTNQv/8mNBI63M9C2UihqJUwWyylljE/VMAxXAXcnW4TLFvDfmtIxsX1f7vtDmGjo0wNk0n
Bh/efbkBSDRZBs+F2px3rlHzCATBMTGZ+WlSBLFkGXSLkv9lsfqQ8k2dHDWDUpj+u9LHoz12fwqC
SamhqNG/VJTwwO+H82n41GMoZD8xEtoqjA7SilwkobjDJCi2DFGX2WfuIE7v3BtlEPY/FczhwRmc
ewQn7OwJoKS4gFI+hV/N5Gobvd99rmUn6mR+1JXYxzyxGKsZopd8TbDi0y+VjCdrG8KxXytB9Tee
8hyBSAH0nyvYwX7BRWpHh/JFCbiraN4KwEJlm6+JtzVBWHkY8H5CxioSstkpboV5Qe3ov17VYWe9
twmNn3BcdYJ7v/QN0yZuj+E/JGoQoB30o0hBaC/ZqSoML5WtppbxYlMrsQIBlAnFeCEY36PDbA37
pop7pS7pewvk9d7Lqm0A0ZXFEz3ZDQn6K8HQeL5DRhO8BizUVG1GkgzTvS2nduYIUXQA88D3jMEV
o3QaVnmiwtvur7ajMYK0xnNI44eiWhdJvoCX2xF4H/T2P7+k7DvrEZ+Axrd66V915xhBh+WieQwo
8VAHKvM+B2+AyFbaJv6IYJtCqWN0lJ8Qg+EUezTSgdyhhvh0ePZOWubHcmz6i0BkOy5nilGjktWf
97wDx3xLIntd9XYmD0aUdNJt0xnK/wCUdcVaxVIBixtJc3bQyKcBEYGZ7yM6hjBKiEizsupYX79Q
JsYPvXDUEH90eYbmWaymBE9KzPCcqh+SpdbLGWSZq3dx9kFStux7VS64UoKTMxydWhfwYmR76KYT
5S2YAcRO42NgrIdpfPesvcVTE86+5+2TJPVmhAAE+1FFXWzHMLJxL2MN8FLLN0ZcHLv2oef0fqam
ccLgXhXOSwHTWWLBKVGR6XXNfl4sbh845jxA8jpwLcY1JY9ABRq5+mUfqVo/hJUBAFP5PuDWsCDT
TF3rKgU08Se7D9L1+vnLOuZRVVjF1Sizxux8Kqtl1CHVPMILzBzW935FSrJYCWqudoQWBr0bf7ia
TcMURDjg2CKYE6i1Az45WhKTqG8fkwTzp1pt54fBV8lqrU9npBmfdjFfmt5wsZ0t1Rl3QxG9D3iW
9Ji6CklBfJinnDs3F/o/XxZwDdnkjhq/OjQrhIXeMaCm6B4mF6Okixm+V9wE03sbXcqSrYABdoLy
yNexFXGHCi43cG1x7Lr1eRpx97/+v7lyHyzX9n0m80Y6HQeTfqmFiTwuBIGzfLqR9PSKuCiabu+L
kYAg09QFAKOJzFGmbPM/fdt3XqiltgmZt3kC1Y6+ENNSBEoxDp8vQ1OSRXxpzOcfAA4bEsd3FDAO
jlwz4/jtFIrYohyveaEGx+IbskadMtSRXRQOsFfPce9SNOXMLHJRyE4vQXTpYcvMIybDwrrAjNgM
Xv2E5t+LqRKsTwwpFIWs2u9S2MqNn23AFyZmGyvzx18KgE5HvWamwnVcYIdH9z7ofbakHebuAZkk
onE7Y7RxFLp3guA6Ykxj3Y9PL/AjLj59lMC8TeGQOR/vrgcFcsCPFBFI3P3BCJoZ+UXj+VBrvtGL
9mmxVRDjQ1syP51n2hUAlCOZnuf+VmF6AtqIQPD85jrGl2i7UWYlxX/m4q02xov1QMwit+AFArCe
0ogGXHgIyNysHeFxtuyv5LMvoIKIdHR1qKQn1AdYHj8WVNZnUYYBRRO8CZL6onwM3lxvO1UlIOI7
IURs7+iKl6iZtvz2IvA7edFCKsBBdwZbVFe5XNdDoxHh8vaY5eMf+mPaJfoxZXAirSEwb461djLL
oBxiM8JnwAYo7wvKE07tT6jPMbDW2akiB6XL9CzP7xBVepDJPxS3n3dP7eWkQ59I2nWJ8bSj2yWf
Tdf1WzXUhHzz4U7DEi5dLPAxfu/yCKUGuWUFAAYBYydL9ExLXA+PEP8J4N+o99xmCrTYb1HOlGdy
Nli2w0efGhgUdAop2WW9lP5UwIHVH//misKRzAgRuoT3OT22QTd2C0rKClykQ5VHzLO6jiYF2XCq
Nf6mwhgz/mZoZgXf4J4R90erEvWrqtclYyfPY4PavVfaqGLoykNjbyEoEhJmBwkB+2dZzCBlRyvM
mdhJ1edcenPOSL0l1z7DM75c5GdGouvO6YV1LQLDu88XngYHtE5btLtPhYnLEWuNN6coB+vb8PvQ
vQHKoD5+6ymiw8X/yuLXjejRldBbPLfFvi2gwC0Fq1g3Fs8zohedYxMjTqQs17aQl4isQZldZ4q/
MY884I+5GyYDMMGok1nC7PHma4TNCiDSwx4sjkR32UPC22IdepH/BvL2fNIbMidHcGSySHIb+XBH
5C6l/LyHWlFlzZKwSBDQEmvoSsc1HH0Qb90N0D5rerwesT0+RSIuTqE76XnvY0lqVAZqYH0UDPqo
MeSInDtv2/yMMQl1hv+6AOc7BIF/0ARUlc7gZrBFqZMUQzb+/gXukRqmZdC2NoB2mNmX57UDZnHP
xUH5uJU7+AhQgxO1imwRlpzRdM2vT5gqyncmg6iZTZyxdOMkVKWlGKmOzfF+AzBmd/Rbzgw0nxuA
TelpYaery8+nGtayOTs7t6ngo+ndMJkG7nZHK1h296MxjXQegwlXDubxQgx2LLGopiBw4s8Gf52+
MuBnJLq91/YwsPd8k78xVCLT+tyKn4Sg3egwXequc4Hj4d/iSCawZ5SL+eMNO/Z2v9QepjqUgDfo
sx0pf0MbDZ9dKosr0ihTl32Zayxjfkd9b9luHUcShhM55k40E7/fV8lc/+TVYpJ2xfX9/O7cTyX9
H8S5Hno8fHV4qAAKvkEt33PF/jlxjbcxvi0T7IuVgKVBPQkS3fAIJ9w1q/jJfu8nNWUUZ8ce/SxE
xO4NTVmiqWV8VAx8twooBcae8dJikRNQ/CmDO2mZiWyZprUWRWJjs8FSWeZcZVToQJPLx8+IkYGd
p6ZgJG1T909sTfqIPznBptSvPACY8Q6DbFnui/sbUmQVcOkLnvHNS+YQF/jn5BYSkD8Z9RpjzP4q
WOhCwVgKyqCp9/YwdMKesSmUS6H9RkHXX6c6RUka4GGynjj2mQtEAHNmZYRYq+23ktrjdLeWVHvq
vqbwrFCCMZbKNeMcAzQ0UgKLYNRsVa6KiBQzOlEtmd5aUzRZCvmfAH5OvHAr+XXXYwfjnW6z9Qtl
rvIMnBCiFOZnu8rgTH29gm6nQdf0Ug9cz/WAGmNS+iOhWW6xVD21NG6PtbLtTG7kiamNtaq+ubdB
zySEE5nr86W+2O/4zX4FimWR5Dent+on5UOzrfVmPdl0MXpYUavGF1WKDPrZ+jAu4ab9ZZ9hmejJ
wsPMreq/X8ejyIADS/83e70F7swYpghTLrwGZcNNF5TU3YylHe8WdavExk+UWQpP95fl4Vejl6bJ
rOuNEv5iVFT9c2FyWfZ6i0/+UQXabjNsZV8xdti0YWbWkqw41Gfr4FppPteERHHVHQgllpdQRsbU
1qJxB5TTQxjjIrR0k8DRMOctFxAwaaXN+3w2Z0ipO5i+xDvvx1WXxRvoCBtwvivl50yMcE+wvA7z
mpdyZxDompEYu0OSjIZpT+yQEydIdKxxcccLM42cmybkigrT9YsVriKkUuCCjv8zHa7+iDPb1f9D
yvlmzYLErHqA8CPVcoHsWo4rCqQZhig11ejqO3sFnAqrZfDUHexqcaOi3OJFsn7yk84ruLcDNXuJ
EjMms4yFgmEyrZSuWHXU6UmnZ8G8P68mOHJ6tvKVMy1JPzv9EkzRQNNkxnPY02oIFz+bGsl3lvnT
Exz/KHmK6W3EDoCT9sYKg5WJwdOZ/aDSkxfDKBB3KhcWw+16tPLI5IM6SsYOqObYiLjtL8/DhCvL
eqDwICRxjacHfrVknVGerWkrY7V1KHsC57I39A9KWJKOX4pY/JbZ+4BOF/JA9rBZBNPfFNQwflWo
gOdpu4JQgaY39xQFs+fRZmLMu9hT6EUmjGcfws6cS0pSb2SnCdu7Z+hYfyWKt1aTiNQ47MalIYmK
H3It0wR1UgomZYlAALK2lesVgHHXb9ldUomP/hkiyhMRqCIZ3pdSPK9BbZa1WscuIgv+bXb7jZU0
14JFfeWtKpPgLb1BcZ95lzswdwestds/mv5Iaizw5Hg4g1gzVXfL/EjvTUD+hdyoHQ98uFhMMU50
CVGcd0RuvNYR2KOg+YVNbPhlJz2UIuKZ118BzPF4dfNWAMBbsCBok30SR7uoXOOvloU0VftqyKQU
6yEgZpnu1/XddEwdj2gXzNiS+y8VkqTfYCe0xsiVkhs5SKEzhUgFxmYNOeaDF04swt2w778+kFA5
/iKNNEmutSOp/Ust9G40oU8xCrMG3JjCkZB12zJoE4fYCw0R9ce+O8DZLWz3OFmuK/zGfYtRoCi+
cJeCPhLof81e9V7+Veq2wFwBOTvSXG3wMw3lmWTlERSkKjptANRFxBoThsTVvOkp/4izjBP/1O0r
dIvQ6Gtk7g7XepFJoj12NdWbskA6XdJVsdD6p4JC3v3iwrUlZy4AjV/HYba/ypH6BMGppqKD8WuU
PuoeJCQ4aezqAlS3dsK128SNaL+ns+isyNyC0iB6Urq90+xA0mZdapzBkCxobwzY4+ylcOtm7QDJ
lXeja2kvW5LOYeFRfeks2dxqcupI+cj/aOGyEMYB6WB08AvCBKX7wjLIObXfkTboKM1N2H92YMXM
AZ3fbe49ZsaIZ1p5N106/QbY4R3iNaNpl0Een8JFIjGks3njz2Hk3ntoxcOtO+vNxAt/udj8tm8q
gTgnMscn8tOU57LtJXaK+i50qjP55Px1TzclDHYT2LrnLqgBE6BpxdIWlONRZnwY5Ns4LOk8Ixza
aVFth8rXOCH34iS0noa3Yur0UGijzOZtuOGliVbgsHZUfEvrsTK9QDnQtob+ViFwjPWYk6pcRfhZ
KyxDWli0CZ+JlWafFHi0AVmyDCC/MrHpOve8wDh2bx1SZob6IAghBE+7RlXff3P/36Hnpgh/ehjV
01oOGOUtgBCiQKem1TY0deR61g5t9IBUCQ7kVxbUK4AHUl6GrbhK3E9XZTFLOlSmlgxmhBUDT8S/
fWWmxglwy7DTOa1m7zEpPu5rj9FWlYrngPLJCMM32ZI9BTwV+JS7Asv3W3EjyToLvcVU7KfRKc1t
Q8C9EcPA9XqvbHZcBAGhIpy+FyKjWO8c2U2XrQOqF2UuglV1LJM2++mDobCmOie9jy+WGtLj+Js9
PSdUsSS1sBLGBO64AuhEE9dMR/NorHKmUg+ntjqC3zBrnWM7NgyOrjV9glqSadn7Vcq3pV8Mxrxe
dT4YO+1eTsbTnrJfVIjulzL4UFQPn7KlRsJP9WhsvnNWx/2OABaSVaNRucvwobUNEJ50BxKVF6OL
JA/Z7PaEwUUvALep04IgldzEzef7n0gT8pBfDRFn/fSyS+DwtEcateqU17JlsjYly8KZaBYaB6RT
yPvdpkhuagQ16YGWHAPhAx4O4gliiZAKcLyhWEWm0Bo+u0xuw0iqgabg9yUXqGeBvQJ+ddVtsmTw
3pn/qJ0INpcwQSs4wNFCHh0llXdCCULC/0RuGJI7jr+6XBP4kuCAhlzTgGVBbqpwUJfcpVd+o0mV
tl8E/jroAHSfJofT4hF+sUdHA9YXFd1nJSS8F/+Lr0zW5K2jz1nuDD7Ts8WiOXyaELOni9M2g+BJ
5NSQ54gxAnLujqix4nanhmSZAQMJ1cDk8vHkc806aCv3tK/YQWh1MytPOElyLHNsLOlUMBmoRtOk
T5kCihsR/cm5awAdG06pIzSfaNodhwCUsfs1TohT/6lknMFdfYiyeJwg1h1DIYvQEmVBYr5rh1UY
2LFgBNs2YWJr/j1JdQ1i8XBLRsaQFXg2EkxFxMiUi537xcSYtTN3pJi9++Th6Vq9LMDX/R0lmD3C
8UHVfs3HmlyzYlfwfRcB2U3cy5ur1ty55Krsejo/X8BKbIrEDGEo+StsGvHyOyY6+onxUVvX1Ov/
Zh1D7hOB6UwuWoUM1ex/MEgtbjIvvFuQA0AhOxHEQSMvDTu3/DxydHyjV+kca4OrWIpCNQ0O4i0a
jN25V5gRW7BBd3cPop3ws5t3dz/AT6UiwHHHt4CAyzL1sCXjoUMI9FLtjak2j/jsH+4wamaZJ9MF
JnBhyTrNMFLyjMzvUqiWybkcn5iRZH9dmznAJETpIpUrohrSxn1g+dV/IQwsRV8aY7z7dYhomwLC
0OJlVemLj5kgtUSWC9a/3mtt9RCWk5hZpTFgV3Ufpz25aeh5drkCdgCoLo1GZ7lJDGvCVRueSMHY
NgBDAWBGeyJsYGpFGlcIwD/LBbWC5NIgLZJa8gbU6SAUqg0bfwL4EFjM3ldZJRLhhphu9QGgaSH7
wpLHeqOVvgzhfkn8efEV4lPYp5WyxLcy+WQND9QL11/ejeI6SFbNHcGJvTXAtbY2eVKJA00s8R4Q
4+vSQCb1Px1thTE9UxCerLia1hNQZeuxd7EGza9ekNFrJ7BgtWO5myWzz9aCk+bqvhSNGcuGnyGu
SuXAchoy1rEq7RrJ+yVHxWOaKp/ezBZEoSi9Y5+xEZ48NUKlrtGENxVsBK66K3ULRcs4eQLvLXzU
TN2T0BaqLT1uALpPLPEUWEHnrMJdKdMalQH+3CVwf2XaJrNs05Xd5D6zsMuOGjcN120pqwW3KCMO
eL/yOe/BOEp9cenqM1TmVnmdTsk1Qte2uhB+Py+4i9VUNAQVXM8wvRAnTPPcUVa8aGlNMk/BPFjs
IKsCKPYh6SRgdV0afPAYQBQOeWu8272FqZXieJj1F3RJf7hT3Mn19DP9Xm09KXnh3xGa9VFQHgHH
4aGptagZ9Gmsq6LWIJ3698omPBRCIyUnfRsGE5o+Zdn1Xka2aBUOaIiauHAFAUDYDR8bgoFYYJy0
PW+uM/9UXD0tQBE8Lrd2/KNnpib78A/HgWg7/duGu0ixvr1xvaCYEzy+SAvOWc2py/h2oe/ux56/
gG2UkKxTivhYSTVv2GI3OdorydOTjYo8YC8zJHQcYmG/nsW+tvrnMoSlELD9ndP4gOVqUHpEkdy6
j1kyUnlee7QXOvohzydwNVrsXZrfKcDrtYkgCyY3rXyxB6upw7impmmSg9QcjT/pqky/5NG4dXyl
DDwROzgl4csy0wsREU0LZw5F+ajn3JPwQIuc3oaU9ajJGg8uxo15+Gvkwn0iT9zrQ4j7fwZutjYB
HFWDjguw8zVN1NUqFd1TZMCVK4T6NvwJArGEtS7gAs8Z3Nuid1tL+aXAS88OA04qq+IetHMzKIjO
U/f60v14fidTCKUX2C1ygPOxKV62vUK1x2gVQTTLcIK/N9JEHpfN6j1wltx44bHFLr/301bzbUTZ
Tc4lj9QvaGL8A+v0YBeZCtPsN450IVfVRVa/NIs/YwR/q+JF8Vz77P/XtfElKnLHR/ESvclnGwm5
ohu1hc/UQ4J1r8oXFHDLvFVvtzyrIa5SRjMd1OMZSSZobXPjgs0cgaJoMzikhMxz/Bvb68upevga
uvGOdlZFuhLDqaUl6jMgVsUjTRPo7chIXCHzLFRk2P+Fq09rPejkXLRea0Awh1ajjWCDCpWyazbx
zxL8iSPIBTw5+mZ6DFddrzHhhAPkVSQQAo6ICT9UiWFtWS010hoAFfXEGEuB7RTmTcEQ3dIpjFyB
FxmP5drmoKfBZwb8qLKG53oegd6LrXDzysfZ0HrFQc6d1rNYOoUSRVSJpld9k51sSkqyBS1of9S9
or5KXLokJq1OpWWdYvfSkV9Ef+YJSI1E81K0KZ34the0Z5LrBZOqOoiyn2vXFSiOB4h9aVcSALfY
2JFmKsHUY/D5QENDkQbSP1X/4ECxAkkn8QszyaIBlFt6fx0+BJk1zIDOiiQIm3favgUUaU7EWnFk
0GkkP1mTLRo5l4yBbLrYQInS1DRbIFrc/Q8ipW1RnOf7zvzwBwBNktH4xPW5dnYyR4qIFa9lj9RA
5PGbtI+bR+sMYSQr7nQivkFwKBw5VXhcpwu0//htdFp/FpbcvYkNTEUT0dgCItyP9S1rhD5UBmhP
2Nu46iAgEKLO5UmS3fs+YM4+X7aGK1dZQHFQF43OQF/VIg32gReg2SdEw7Td2w/W4MgQg/Bq37c/
NUPxwbyeWvtGyEObDckGHgYs8LlqJg1qZOlJbCMfBDQra6qE7ixy/pel1LNkdCrnhuuDV4g1JxS8
pZVO1rrOnEPf5ZqyQu3iRYVmdM9COoszuhub8B2tt7Mu3zKOLxzk2wLOlauWL+a7kruk09+CIt8P
LjTUwCjz/Oz9gxmVTYmGPTEw1OYzKGM44vZ3aAv8a34Q8UXCwUp0mex9I/wbJkTV0rEbbJ055qlx
RR/pz96q3Dfo9O1ylnobY3CW6u7GAiibdJ7lAJwEMkxiYzkAuaTszWp3J1jcIppf9yjYYQ7/pOKf
Yr3uttOg1b/ju7NanNe2DAM2KDdC6O+LMUmElFZ7eK88pBifI7ydT4a6VssmzYtOkkTKj7RlH4Fo
8RDwtMZAuo4W3QOUkA0B3s4IuUdMWny+anJa92Np+8pQAFC/sxPQGFqfPkEBEw+yatIV2pe5KRIG
RQK6jRDWuaIZJt1vnUHuA0wghrKqpME8ZHpsFhkmND5cTTokWm1eFzTR0jrxpnbZ0nQQNrtMWfKr
6mmdKaQkAnhbqhqvQa7JwzOvo0OmlRbrpjvLcXPRsP/vsV7C4yxXHXY4mATwT8X4cNMX4QjGzzvv
q513TBoKZ79ZE+/CMahmKAtPYNj8PYVPO9Jq0NuvtHMzzXyK34qjNVsHTzv3hdLVeo2PZIT1oyxI
FHzFTNw4nahKzcdYdG1me44usUfYyRgZ8qmc+QZlsqZnhsS6LxFFdsOX8jUxYo6ct6VVREjZ5qqj
OArScZadLpIHcXbl/KIXbGKtah09kwvA5fsOO2Uu6UYHkJWRcgXZpIP0O7Ub5kQ+0thU5L5UBcUu
FCSycqy/A1hg+umGZbityw9EkcIgaYtfHb2YU1w6hGawiHoL203Sd+T/yHnNAXvRDV+OvyEHE2Gw
dFZKvItf3CFIiN8mDhR4NmBVlVhzDtcLssNkFgesC5Gu1jcRoQb7mHvhnOQ/SMvHAR/jXgSiBiq8
Kd4SA7C8pvPaJFJVwr0t5gKJ5BNM89EUuJwAEHffyQUKCsSPvuKfWmQCZ8yZJeiMU9r7EOfMSJ/y
V0md/7AbgubS+gaFzofTxBRxlxF0wQzAnIUIfGI65gktSv1upXMgK2tKCZFJhZyc1xRzFSoECelK
fZK8lNS5m9xdzmiTGqhUt7xhaljC5T82/tx6nrXffdn9iWcamjslalPg7thcoeA+Bi1+EdO+5biV
NYVx9zc89ZmrLeqPZdGUUhZ2hPRURWfgb8AQ4t4DwOkNgRx/bPNSWPNJZ768kW+IiSsq4UXeItOR
o+SA7kgGD6PGEeijIQnF43+KgHxz4t9QIBgSntiBsPafsrd0D0it5IauYQecqL5ca9AqKO3/m5BY
9fi+9DFkR+VzX/i+lj3+80VlL47TL69wR7/IepwzEH0V7Se4gcYCWX0PPwOlhefbkIhKkbc3B2S5
hq5TFZA6EL/QGC4R2+IZr98jUNFIm6hG+14944K8/WNJepCT81ROVrhWQuo3Jp6SNlPRwHKz2DsD
3rc1CEu9asZLo/kudH6/8I7PmOBza41/PKQUtrIMVyPNwNdtNH7RAT0kzt2eI6zxYGqJ8rhKeCuU
gysZKnwKGcuvaEZdICcQqId6vkGIGSBw4YwHS7nXr+hh2c7VzV9+5kLmhjkeIZqSLfqxaNJEC10X
IlRpiJx+lzeRbBNejXMRlMjvw3Zs+VRxCtd9SoZM+z+hZx8gZKdJPFDszefLBx8w3JvaLobIwZuv
AkRkhA1h/Bd5sLdzJNi11PBCzzaQXwdPA2p0yTPCAx0tIW3Brl4asxnGbFBO61DCroWAR8pPzv1h
mjvnt6hrVlksO4X7lKBKRCsEwWcleAONnFkQ9/+NeNkdzGIHtBSZntJ5yLasdFWgVGXSx+cwpiAx
7I5BcnqFQJ+Mfe8GtBKCVHIm3LzdjRHop3xh1nrDbqRRGt1wT7ur5zaQolGFYR45UHir0bn1ehCe
LDCAUI2799slY+zzYa/bpubdoAuuSkNhbRpXbnZX6JVUiGc0Lr0WlAFhE1UXgF6+Gmc5Zyx3Emn6
O//0FZ4egxn1jKuOgF4fJ2ce5LZKth24Q55yD1oIk1dCsDicr7et/zLtuAM86AhgoV7PW6XXqIiE
H7k65whrQxNIDkOgwr46OxxuuRoe/x4vncz9XO9zihwrK0tzkxBHvtwiDCIbG9BUbtoeT2viRG++
VjjE4fbZ5wEAdhgH4aGsGzaTK+CZlgUXGy4YwhCh3ybWBeM+JwxLdY+QPLRvpJ9tCGYW70gvs32p
trBNYD3ZjFjk2Po9pik+ZvApyaW9KJEUlkb/nHYiJS04ASpMuLhlHLqI5xGBsq+iW+i6qaNBvXWR
3w4L5u35qkIocRRWKaGslDqxuACebd1Hn2k3rtncXK7xki+2Pk63Mr6kR69q6rMhkOpGlPA9+fhx
IniHtOeMDw7gNi33bnSo48fziF8vxEYfMK6Zy8G2C1rpRedFRj8UmGl7V0t87a8yLxIgaG+HHP5J
LR8EYKhuB71DHLvBlj0/hk8ciiPFhfqJoUfArNdYnKgpbTVCeP1uHkVvqwG9EUXPabkqTDyARTT5
4jp+k3H+PHEnXZzJhnthzs+W4YnM1HzgLrlz+8gKQCfT+oq0DHvUxPY3TbyPmltNIRRJKo/NYpS8
I7XVvyUyJpIzMVReVAHHFuBZ+h8nzCvl6JV4+076F3R2OLpnLO4TAmf8EnGx1GDbJyigmdEz8Lq5
uS0mwC+AWe8OFpUMHm9wMxI3JLEQHo8J3oxlkLVlafSP2rO/E9ZMEozQu5MROBv4gLprvlrOxJO+
a3hmcZK9Mg9l9yveUMJYvP6QS3K3Z1bJF++lwfOcTL3alUorih9Qn8xhYQ3rRPg1w53L74U68704
xhsxgbi9LHDoI5ebi9bEyrji6H+mXSNhGn18d2HBpUZjQeTfd5Jml39+RRjzJ7hBPhACvppqwaEy
L/c7NMCCfIXj3aTuvYZjkRJF7ebex6J0iZchbVxSQSWWEOVD4Z3bIVbLoqiUn35hO0QJJpuSOdp2
J+J4wwZL4oZ8nPG2pl8L1M6pAMTFb2O0tTPUWFEdBz4tWL2iCsFoEy5hTkxha14Tv1SKZbEvs+V+
1oljss8nWX13q/6mobFyheN+CdxbrPnR5Pa5ek+ihgmdmeDnC/Fnxk+p45LdLt6PfCAEqLmrQpPq
PUYM3lVWugjuQ9zOlBh55+NniX+o7g1rTKvsG0uSQQK2g2dkCFBDCwFTEbGKh7nd44R8PlRL22Qo
/YKi+kSzc85lzdu/82tBXgy9UsHWJhxfiNolMBqBY4wpwrxFRnxP5sGbX2uIlkZp1ADiF4IxFFXE
cqy5xyYzhJfI2yxUhvUAuXJoAB6UNltTikv6BmiOb3Dqm0qsD63NqxlwxzNTuf00pLvgIJoRWcUH
Ob5iMVaW+8Ky8iAm7R73rVOyU3DziotT2Ofy30cAPU65gYgmYAUacCV/ftSbQRaE9GE+PSHqeLuE
9mxgKj125NJjIk9ru79wSeJTH1kxMGy7w99cZHJoFnLw6c6jgJbZU2DT3mTr9wGvMZFvjAlZl7To
6aHxtpOrjFoA0NXpQNglZ0R2/qYqVSH5xoHx6hBzipr1ub5o1tlfyQTg8H0xLxCztP4XmfXxlg0H
QkPzqh+JSD/mC8gQak9mSNLjReF1/61E3EB36mu1At0XrAWJjmZy3OSpIO//UPXgtAZ/IejxjwaT
1CZuqwb3A43BYN3yy42YwjaEn+Kz5mVXjhsPa+Gl1zvxnlF4OZ3K8ha8aBwAt+NYLCK6/RrK6F7m
uhMUO6HXVSwp15RVu72NvQhdWK2gjX9VchDKM0ywcX7vLl8HGuXLQm4B3SBWGbrNBE9gf+XKV/i1
U1/Nle9GygCHFfbRQ9V4Mt8q3M92ZwFfOC50d3Y6FTf5tys/gxcXifN5I2dyfXoDhBUu6AknAmYp
9fY8e1DaSyAeDtHmWfuxxy9gD0W0GmZr4z92NgOqMN5MtaDLblZUHYuSc8Bs0YEZi8jPDkDW5NgT
kWRJ2p+H/TcumunKSsH4D9OXmQR1VmZ8KaPp83ntmdR2l3adtwDds87FptBj6jnXnYAMPbrp7q+W
6k2uhhWq9GsqL08P/f/7mP/nvE3Bo05QDrrf8kJjtHe3/iQksglAv2rWNOS67KpRNYCiLTxlGPZS
2da/2ou8ckYVJzn1/PeRX44zaQpZAda0osypBXo5ovKnw9YqCYB1AB765tgNef/+vEnRpu7VVuul
UL/AIl7zZ9PW0myHN+LwI7a196DIJ7z6lwbdptyrltSX6OoucjGsL8OchLiGV8hNplvMjtT0Ya7B
hj0LwZ24tUSQSbSAjWK+u6I12uIBpd2pSpJOtXUlr1gd/9YxwcUHJOyKmMPsd9M/J+BDX/22YFOH
joRRxeltbAawRKUuV1aV2ur6FL6StLKKaku3PcVMoMph7h5OywSCp2dSjH+Jpz/pw5O3vXZIE0bf
LgJnDbErMXobb7NZ42uiXXiGxx/GKfa5rpjAc/G+oapu2tfTAZYqXgaSL23atI7ylr/bAKTT0Urc
HKMra31tfJqoc1dSls5LsXh/G/ST1QHWC9uy0550W1sIg8TRIsw2IJOotaJPsG6RNf53OVK1y3oP
88Kg0gDIwaRy8PhPEGA0vXaJhaLLn1IPiqnYJXPMvypwE1rBmygzknhJmA/KqYNcHIlPWXlCzjQO
SBsP75NPliLUwQdcCgHOLDX6+qwTHkCi9A/ijQuRqnGPlSBiU+6HqyDUSB/1dEIBBytq3GccI678
Cr4jWB2eDqwBscsm6v+VuzqFE4117VgQz3udOAa71Ql7t7OoLc+4IBm55OSfONfRT8HmC0GYNcDT
Qqo0uFfKZ3qzfpjh+BqBpT4xeGego9VA4GN/MVcVbV3EswWvHDQBW86f6cJARvY0+h63sywAI2er
58qDpZ46LkJS93qejh088APaM9nkYe5OhOOcORG8KnTSajjuSAbq1z+49nnXl4W7YQAEps8+l5pj
fdKMsz3h1AIv09P04EVkTSOoyK3x7hVnEew1/NEBHVogu4bwgXYYKaGuCgfEAnKJVfHz3WwlPoIc
9BEfpJ4CouIl6hsAp4nRH+KlvFo3pYzCDKzewz2jvKEbaMybpuTYSYVkRkTw0nByUPNb3reSNDfL
xc0fP8rp4RMnP66yZHjF6tjZ98WKEJUaxK8M3LUO+4Cir6roENidxiivlgtRWdOU2x/wv4ypdL5i
EmV/FWYf8W85Ar4E41a7tYq4wuCdKspUw3pH5Aiyqx1qDy8/XS6TgUG0U+UWgmJhJk3irxve6cL5
38k6MUXkri1aCPQ/3H8zXMONXRUt2zHv0I0fRkWkIXkp0cbCScVFNMJIgNeFe3jhNTr9ASChhmh0
UYXvJwIWjYXUAAFS6IMIfRFqzyJi62HNy2YuH5IiFpAaAB8rUW2aF496C3UiePYDBeftG/bhLs7T
ZUoDNTQUo9GlQQr8NM6F55y53hsP9RAX4hIzOnTFmpRjC+0efQTpCh+g20DHcMcy6mYa+J0jJx/V
FTwbd3D1cGz5m+Tg47LVewYUaonODar4U9f6DYM71DbUgCKgoyEShmcPdAUycVmdxBTxQAMtcVZ0
ptyEp9Mw2JjI+fYcnkXo3z7n0JjfH875+CgLzyBagUk4fnFDxQjMkwH/LoPfgGSyPs0B+o7Ar5mA
cNsWeMU48JbDaO1idrDNoEPlmxK383hr4iPVfm7FKnfxVEqs608Nmm/IXDNLFEuFPpAAsViUN0rw
ITGqml6+JLo0y8xP3HlSDvRzwTZ9NkWhoGAlh6L61WZaaPnwKEBLBgVNB9EygLQ2GxVtVEtmugxK
d5pp6QDTsHvHEUPimu7roSvsUkLHIj0YHfY+7nWTDA59hNEFw+1Uz+YSt+hClqF8bn+ktFdWzfyh
hkFeCtN68AER+/BF4Gk0CPL2muQLun8xyAXJM2hWYt2bMNe616cibLaZPN2Z3q9SRgZaIfwTsG6X
d/lcYCnT31L48mvH+y6UyzUbPGAbbTEEJrBBL8rHx7Qtwdkwvazg29o56H6C91jZ7h3US7qushq/
MuILx77zaMxxrrq9nGiZHh459idH8DSJN+hcAR5t5Hucu8GsTVKXkJYtN3SM10SFAlySCgXoIJVD
vOoPmVTAs/1nkOjwljgomvIfsnqh7L7fj1J6GLFYTgX0vXgqUdBXprkmN8ETG88FEceuDwPy85eI
ADLQi9dM/+E+eRkj+PbmWEpDBtI2z1+pqGU+qQbqd100u0aLNjh9TaQGgU4Aev/T1K84z6bcwbKC
/xrX0TiuXk+L/cmCn7L0AW/pYjJdCUrDzqakQZxkufXM9pLedFqiqO39fNlbaaUKqbfPCrQ1h0CP
WwKZF/VXCCLzJiClKmir4PxCkuJzq809vNiQNPupFzwJcifBhIYsBx59G4p/ZQPWeUww0c/r95d7
z3USCOijxRqYuLpW2iFoG5ODZgfzkKq8KZLKQip/1ybxCKvcMVMueK2l4uwRmywAUvhvv2R9Yuq5
SQpl92HOSiw+dJoOuxhXr/PMGYg3Js7S5tq/Se6/V+aGBRNCMkersCNJrp2DK9zqhbjH0gWyrvWO
/dduQ6TL87CD9+kTD1gaEPTFjtvW0cFHuAMyUufRz2UD9Ns840NFKlDzyzX6r9642kR8FQ4qwRWu
/90CL535JCaW3Q6q66LFgPzZ8ieQMpCbHP8RmqT1viz8m4D9aDKGP1Qxoz3wl/275z56KGrtNRTj
ROHJvjLWaaubjhwFCs/eHTYdJiJDnhCv5X1eONkytKfVQrPEbDsDlvG3+n39SIIxq/kZEZdTY0Dk
RTJd9X5pKY31X4aOzsYC3NzJbaU9hkM/9OT646qU7r1DfoVpp/BZAJOzwD3YvF49ovm0MtnOH21I
Gc0GG9Al76GIJjunLYrJMTVVfDDpURBiqOePaZk7g1HXrp/bHs5oNgze2Cm8ySFAtpCxLqJz183y
JICOZzZafI7iIbPUaOqBYTbR2tbnhimlmboNVf6pt2/1beyAzhRT9N9uXEXqxTz4HTGHsaGGcyAV
XVS6ZMlAWZ/Pt717m8tYqAWW2Roiv1KNQhXii7WqHiDqjgPylTHtqrnzpw/HtRAR+voJ/TlnRC+R
xe4BNx8YluSqk2Txk1Jrs0qO74TtWJaL4XlQJ5lKnsikcUZm5dA4uJtNJ7mR/2wvRvPIeX+3u3e8
dM3K4BDz11doAmAiwwTCzXHSLQjRXCw8+Y5m//xgNivpnliBy4QMLba+hY11qaXzWyHKKRbRHmWf
T6HO4Mi5wsAfOJkMIGI0inoeTbU+H7yaAeKi4GyzlIUNQnI5FI4c4iDEohTKZ9YCFaeEGAs7BHdn
eGSF1rYlxIMntUJ22sr7l16dsylcXAwCMUrnyS6eRPaWfks+4KtZ00G15IVNahTupypcrwdUPfdI
8rqKCdmiKVESfqEbswFIjQ7CcgKWFA3FEq3rsqzv2DgTvoV0YV9j8Bqq0OdhzoZw6xvNt7crBjL3
f5UHdHFYlN7OJMw8c9hgkFgRJVCUiCZG1BfVutNTIaYUTjgLkkaXtmlBmScB05dKuc2r6m4vF4MR
pllki9T7gnI8awoSxSE7HP0CWmvPzivUB+mmLD0fLpj1D2U0KlX1f2jblexJjBFiTkE6dXPeEhKn
xdg3MiNYyD4AynYh65SUoi0yOqjpmvyYSXe6u6vg38PHqaeeUFgvmj6AZMkWrMD5KiZZZwerXmPr
RnehoyrBo1xoUD4UcnUsH0fsaBTRBqLOpFKPdOx83shLfRIFhxOcoEt66DPpKnJavyvY5PEpi4fO
aIQhqjemcaRlp/77ee/9nPb/a5SvDy+/vdJde2Z1MqHtSTCfCICc0R6ZUPUfcC6By602LhnO0Wd7
NHX2K+cVm3AU2x2h2WHNLH4KyOjxf5zmVep8CYgsGeOVbikicGcC0InbM6xEcYvrGO8yPDY0ClH4
RV4S4pj3zZkUX/A7JJOCMjqZrKhSHwmJ2XeFZFPp6YxIDdSmRQIIdbssEzmBZlezJ7jig2Taf00j
6o+8AfkUUEYGON6cHmq0VRX1as549DBDErlNcSNI0+siX2a7U4EQQzfcpKrgf8xgT+K+R4R3Ia6j
m+N/tQrwwQ16Gp+B3XV/dUIOVNKrzG3Mao4Jl+YUpp99oDj2DE5XUmwoCsxkX1C1hWNtaUufHnpm
xPtqbhKGE+4dB6TWeIfjo88traViosK8PB/qUo9l8aHIfirt/5p84vIEQXwbWldZQKCp4hL9RRER
juyxbhUaShG/iPy4onXXGDdL+O08cX+PzmVLM+1B38bOP+nWO4KclOnfHhKWi3g+frAreC8HKjk4
2W33Xn+xqcoBltJE/EMcMsLgjkNj/YB37AojDWsCP3CoG+YcIUCcuivrfSDMqSrU8vFsdYp7QkZd
RvkHN17BP+OhInAzniw8GqBR6s4wc+tjCwQBr2OVq+4gjifpR43fpfpStheSgs53vbFVaMSvzIz2
HEDJMOhADWTHCga7q/THDbYHQIL/bmQlfP13Wka55EkYJXiR2GBtX7qxHYCmVfvyKcqzdcejJnZk
3vRrixzewtHSp2fEn00uIAX6KPlDF6igtmq1wug0AaF9OQSEM/RLAPnrdn1aUr8HWhwsJIOS2k07
sMZlQZhHKpHM0yogRB37JNVQmd7UE6GgqHcQCuHMjJH0KCzdTe8c4ObqsNkaTrQy4NWN6NXucLWG
BYQcGpyL8QSvI2U2qwqcSW6E6PlyafUoZLQoLg43Y6rjSv9WmJJy1M4WyKZMWcdcQZ6G4P6/D7z7
7+Cyqf8IUCjNMgak/8Es3SHMNn/RLz9aaWFInyobdejqr4VDRXDiaSAUdXwz3WofLkwGlOYVrEIV
CMsauE74t4UBVm/rUY46mouDGEW+Wrvi1CpqxufoOGae/0HDfNQPtXBuwrfy30iIt1Xxew5CsF/K
34i700prbl6L3RSpR7H2zYaMzFwQYKizoqQlABrglrIRPTJK8pLcAw9P2h4cFL55J7YQXO6n1qUb
m+sjJYOUVQ+n2hm2/rAtIs8tddtmnrc/IzvQKk84zOrj0GzwIuMvgSciAICAvPuXpBW9WVumQRrJ
8krcZBfYAVlfWRVoJnjBT7QZiHgQ7Scggp5TFLDmarXjLLxkh4m4URkjkj1Va3INk42C+VMMweA/
P13p6Lbad5lj1GuOMAvsGkFzBtsZq19LiQPDZKqxsbFwDKHlU7e6j7C0bGFF76wSffcH5glY2WgK
9Y/bZ1GNEKWFyjFZC54GWiiCYpaLuhXmIqyLd5chKB3Hqf9Ss36dSlfPCBl8hbS1lRIQVS602xpn
W70bOwLf8hGmJKIvCPov1ImhB0rcMeThFGsQgneoG+9ilANgjHR3pQl0B/3sURwM6FSER7e2YluU
I+3XZ0ov8/LSQTJFv7iNdXqWVB6sqod7M5syLvbyiD3y9kxkDc8Ym9oBsbxrRYye6E5M8kftnzp8
FRBtESGydUhhS7g7P/cHML18Uyo5rc5UWo/mpScGrSQ0UQ18v2yv4EJumtkeguzYNiXq+C7kVBpO
qkdkYeDVICmwxhg4zhN+/f07a9ATMaueWXDzA+wII7EJ1DqaV7Iw2RaNnpH3x1sLq8yKEFm5QKab
Ad9Am7iD2uvBIHDntcpIv2VO3m+gZD/qiEFr2KVDG3qX2T1hZH+QWdeGLHBGYSjqAkXZxnZl8IbD
X488qQJTnKwmVXgRORgP7i0tw44kqHI1TSSTyaNbujGR8ZWtf9MbedwVK9JTdHu2A7Zef4pQwhym
wdBezfHTRvPQwvW5ZyafeY146vSDJyEFNm2uWh8XNOn7CoFvV9n9rG88N7yn8F8UQaIqgV2UnBdX
+wtzdzDCynFckjkqRS8aEXiSN3Sjb8+L/UzQIrjyoovnVGt7NuoYKFgFyEPcSku725bJEsCWxWuA
ODtyE3EhSseQ2DBlu2h5s1QKRQXhKx1QMNtUEq1l6yc17HfHZL/ba76hclzyqdb4m7OscULjPMe6
tQ1Q7OXGx83TxvOluVMI3QF6MRGAXTt6uxV6w5dhZ2aE7v5UXYTfWxQ2wNl+KxiOPCqvJu0sQ+L9
k3dfC9xV568JSclpGA72CEgQ5AWRODPwMoAvAL9C4+nTrO+H6Tz4aZAoLDqs8maTtDuqeCpyv/dj
DLOD/IP8ua1XmdJxFlAOpLkhuZ5IUjoM0EYAqB5Xj5K88VJG7nlYfqK/iP7xqhFk+p2/Wfuks28A
1at+Z560BAhUI3ggm+ENXomwK6gGGzuRB4ucH4GkPaNWsZfM6t+7UjvN6O6A2q339HgSkOVNA/JT
dHLVza3NjLymFi1v5OcQHpa/6qPlgfpC1WjbEjjfXDDTPlwg26ZQoOp2mRQ1ic/Q2f/3NUhLyWnA
iZCUxWZK+ryrNTKT6tsEjfzTQmY3GvJdk1fX+r9+sKUxQccLIBh/8qssSN0w5WLzkAZgsFJ38UAF
hDgD+MAQqOfLvweSr3Kmps63YOP0CMNWuuDfExtzF8e2v6jioVAD3QMiGHL3re3vzttQHUf5Re43
idDDwqPYVReK8ij44H0uthLabGFgywH/vd5Ajvm/fObmjBPCMWtQy+ejBaUcacTWrC+ZERIOoGbt
9KeftrkTPNy8NwxTv5qsuMErgFO3k05dpgbPYgn9WlDTT6Tt2GvwvwEctknUucmLAIzlIgz8Lxo5
i56TUwfsucFcIEbZc9BmMGLexWGBsaTTEtgPrh4oFB+swXM6OZC+KVujay1wRL28UBvAs+wztcF5
6ZbTQd9r/L2H4CFT9A2b0Mc0zz3R1l1SKfdWJVUteC7pelI1jAzQH5OxGJ/k6dQeoi3ZiMv2jKE6
x5/S4XfWn0R9bydLKMHt+nGLvv6Hz3YuP+eRDbPTiIdmHEnA5ZcwKn6aLpcrQf+XBnnSd8dlB9VU
StM9IhziuN0Cxpe1JeaCRFV0qhES4W5odhOCFYoi94BSoQSF8Yoqi9hwZUyfEkSCLMKwQcuJWWlW
gM9YNA7Q4OBJOFiHMBxAAtNwQtd5GpI+JhtfTQL4zmZnfc3FuVJuMsvWimAgRPN9M+p9NavMB7Cf
8OHco6w0NvPcd6mWh+2HKlkjVJkwv6bTTJHePuAAZHJLykE+PwQ9hWzaNxGFcPesSas56NbLxSQY
QPVx1aic3dRED2TuSDt9JneSeduaWGd2n08pVnuLg/GFPSJz9wg/A9QSasIgITghZFrYYFWx1KSj
MDrTJ4DrQpAjK1B7FYBJkg2OCqClshdk2R51Uofb0nUcouFA74nw82JZv3k2SDd1xCpByTUcqDSd
e4KI7iQ+gyn1JGaX/3t56HbQMETLiMP5/+WqxbyBrF/B6eOsWttAmN08LK6pufqUjjcOryHNdocU
hMQrvCAOhwnACtlAlQNYjJip+7gaZILyup6vlQiRymTw8FFuj9gFVl+V3AFQ/rLTgmVhMboTk4aE
qG73xX8ycFpBBJn8gdT0e9P7FockUMrkTCe11kvX/9o5EWP2Kt5Orq22afFIub9bDAUw3tEhV1fH
xY0+KpwUitfjjHUhubD52EDyz6F8IG2BPRbFqnL/9jru8NIiyUMxQOhJrhEwgFbQogm88cGCTd91
H00stuMeLJ1UjeSq3yrN68HaEyZqErBxJ+EW0CjmlDrZ1GqBg0IrADz95eLJ0z+meacwebm/T3cg
5Ikui2J+eovcrXPRYRu/tCKMQosAkM3Rz2mVVtvhVRyrG7OZbZSTQBRR4KeJq6kEFCLbUnlsdCvo
qzBCmAaAs2pVVCDDpiNfpO0D9SQPDzbDRDzU2GRSfy+7TiQ/tsUVkWCiBnzb+XnABVB0JZD7hmid
yVgCwi1kwnzxpKKuggcqN6UR+DaF87MEn+KXwYr8OOvEejGfx7HsyNwYLqnAVnt4AZRNAiSNqyd2
F5wHc+qGlw0nPP3Ju2oNVENXZj8PCd+X791vAcL6l/jVPcTBi3esMTRNvDxq/9qOR56WSWM3KUYu
Mrq5tybrf9nUu+/FiDc4WjYxg81085nf4OmbqqPB9CW61A3IlH0C2gfv/tGvt5uD2wX1PyaNsMU+
QDolKyLwC5G05PzsycB8xOBXyJthYkLUNV8uyuBKl3q/CfsBJ7Nt7iKUlLFQDbeXokLb29Bg53Od
HO6dqYh8eqfkScXOAp0wVGuQX734hO08BVy7uDjeeljGZIfULZdu2yMRD8Ii1WZUdU9bZS4MaTUD
F4tmBaIwahPyIt98zOXEnCMkhyltZ9uipQEiSUIPfebWFd6MmbhInyUScx96ZBCVke4Sbf9TlfoT
gG+f1gqlBnSj8D7c2WapEyvE5kuv8mMBWxZ0RZ+LcK2LEX0meKPFx1DVVys6BW6CqCKJJ80BmoMJ
tQllxtvv2avsV2X17xWckNeUFMZ9CdpOqD1J4d6Frh+l9nUpoKq20Wn0NfL7LumAUf0X+eD69WNV
htymSXPGoQnikf/c3VhsYpZ1j5ruRWKy4uT5hnE5uMJ0VeuL3TxMyJ8WH4elay/9+IHnKupCbcB4
+StxKBV5VaMOCur8Bsy3YKHOAKlkaGjc5Jwh0AU9xkiqW3F4T124yLDDF3vGEr7HS/UZcbYiEJ/M
/131rpWq/5Phv8k04/ntGiNKK/hgypalFPe2FD3lT+OelJfcOh/GM2AnoYyl98zgYhleYslGdBPU
pJ9KsZXDx/bGyyNVqowoBYdSl7A1rSnkJ4ea85Tw2PvPsbzqyGnAVclES6Tvtrh1fc9CArsvHIRb
nwr8akt9vXrXpUWpYMJohBwU82kxLNZz4yssE5BriqD4E2jHUY6kzG0HwWryzWmAOH4MMNrBdJtj
rCsQFgdy3VgUCah1FRRpC7m4RIyfq+4LnOERK+1fbcEyVpU+mYb6BvMh9saJPiqyoVhqxnfo/Lt0
ZGxntCD1GmeZkgbI/u3UBUCQB6DYZ3KX7YbaeDHZc1Svkl9lDnMhnSN7UkNNmIifQSumNjG8FcCA
PJC0PddeOI5marEYG3MM8NBEVeXfJPnUCJlaXFCFg5IVdnXPVRlxzuu53UdpwAvRgD6UbWIwxA7k
D6uWQPVSVsWvCNFR9tz9N0wULxMjQpU9so+RrGtB70P78wDNkIU6+yJk8sd5r+ADKzbD+6IFsDyj
duXNsSj379wIPrMoEQun5o+NMePHt9vCriID0r3772jGVLr8HW+hkkiWwQ52TQk0lsknZtByEi5q
hl8Zp8KUY9zvXQl0Doj+9h0BuagQ2cF1JZxLSs0MUg8ov07LS2d8Ot4HB0mn7wAkiaJUfbDrdTuL
T9AG4j5h7MeNH3ZcuLtvahZSfuzc4d0HR1+y1ZxnXOjDYXbRGQTh7j2GyP3DV7WTRCRWFIPTAgXm
fLXL3Iysr17bMbGpIQm2DjYNfiIs48O+o1D+qMIWgmYnxqBipEihU/jwQK+pqO6cJDYq9RcxVS3s
4tJl7jmUdeXykH5ylCaA+xnMeb8T+dqL9lZEikF2AIApnV7i72bTHKL4PrmS8PFR0ROCjLeGx5d1
/CEcgJD2PEgOdYLj1mSSOosQ+oCje2Vc8rY1oE0sVOPYGgCw8Lo+BVj+A6EbRtRz66XAx0aOV5Ob
GU7gV001lyveO7dwTA9pH6f6ZszyXngqHk6jsNFmReZkLqCNAXX8zLjD6szhKcCy9L7k9X3qEcTX
SXfktC7nXtpkXQhCDKdsLKTkHT6mvzzWFZMdlxLjvMzmAL/GlFYU69qQAGVWaO7qHN4iRzIiH+GB
Gwd1wOc3RFkT/v5kCBsck175EXRrdRFhO9SClG8dW1YL6b/Isywdsl8FGM/3VA9ZheEKNUa12EYT
xnvns+XiU+lOTm+lHJHgv6RmV7AhNGfY6cN6+1PfBWmL0C8Zv2H9/nxOLMGS9oi9ki5wjljq0OBc
MVk5mpT6AdPztDDkCt+PUleS+15nz9shNR8TRaZ2Kba0pYsm0ZfaAr8WsgCsVnIamdV7fT64ogiZ
/iDKkJloPD94dABcfi/1hXScNLe7+0Lz/vXjEpJXb+rHCNEC26ZtQ6X/cZlrP7T2fzOBqk3R5w01
GAeo7Eh1bhzcCXItkeZYTiagir7UJj6t9CiRdYSMBq30cJpQF3k6ms2TEDazOnjObSw8A0yAp9e6
zxsaGnXPbWWEbpMkdem/SCPIlFQPW/2lFn/p3rruZI05egToRhmvL25zNwfWodZY1sZlyLKlzo0a
eXCpzm9A1xVTGd2ORVJXbRrTcApoXQQqq9Wvh/9u8ehtZ9XXUW7rPGaCoAy9HJQ6cWKQ9LEVNdrr
qTPIHLVCK5TbT5X1rh0XUQO6D5n1rwEa7Ci1W6osaDTGVAL5bttbcigjyTA1yCXEieNW4kLdylgg
wPnqSFAWPTwtDAH/J8Z4QdPwP2LWvmtYtrqxFpOIYmCXOQ5I2a9sJnKiGMzMEexBNm9M8O38GZXz
VJhpXAtIKzH0gYlyiRKzMMaINdeSHEFigAkIRmXBMUPVhq+YgnU99ObNW/OmgOGggf62BzsWabMw
QTY7Wse6AtqNN8hYtfYzjXpmzXvFKH2Y8E7UzPCob/SNaaHFhcaiqQR2mGTIBw2I086y1x7DI7wp
8RT/Eh8DMlj4RbNYj5wUV/gbKaglrFZyOUcauXV0n7wouKS72mH111u2L1yHQkrZDtqI2TEHC/mu
KgvsA1LrZ0osUgOvTSxGfTXnQMR8vfv8OEacgvDT1s8iS4xxj0JtKDtkEk7uL8T3d74gNRkT5D2H
7GxSe3kfBKpIdTXsX1ktGM+qZ7iIAPhv/ugtmkHctKydqWy2NJfux5vuJMQzDLqmPIeWWg1rpzMO
wQZm1FnQXv74x93hHvBAtCS1bO3FpP93j1SXT+1ABo6rFiZKfKxsXhnrv0yfrcx4b/RhmOHfyPqk
5usRkTcmFY7HzmR5gNL5Vh0vIn9HWPd8kizlN9XH+HEkmf6RNqJk1/j+YFbu3ms2ppUpArUZc27j
2407dN484ZWuQVE9AXTbot1pG+8ONClrFU1fWo53FQadl7prxLyISEg2GClGVpGI2WbabNPBUIeK
Eq4GDACgHTz2Ey42BJVdH2sLdpuzxYx9EYStOY44XU5Yiqm181vlDTHEpItKBZdCULfLn7QdxiwP
01xK12MpcPvuaEgs/iXDnS01ybxx9zAXEKJoCXn5V+gyE7rfwZubUI/fVdft686n/e4ePhCptyQC
6IyK9e9zxLF4xpuS5aHT8z4Vg2POno3KYMwACOPsxNnVbN69zx6+npl356FK639e6/BMT52EJSgF
lNXiCvZ6Eqc+i6h8HLZjr98T2IDoXh8VNnlafXA0VQvWGDiwnJt4etbamQQoqOPckz5BG3lcpjP3
D8WbZSC+A12nkEj7gX5yQImfWkBM7NoO/1N0iNN/VrHUz+VV7X0RSurM9mWzPOBsGixA822ODL44
mpK03PkUWrAHdd7OUxU0ji4rPgQsiFav4h7Dn55qBdF6T67w2AML7pa8V4uRGS4uvD7NhA+kfI/y
r8/FR6NlRGcLQvM5iFLDGCrVkcS4Bt550kNJUzh1ZNG4RpnE4u3uQTUXkOyCcgMPMkYJvEs5YNqe
TI7DE/7M5AKNV6ynverHwpc384n1QlNTSPGrQJzE4aPEXSgfSlfS+Y2HJw3RAQNvvcSFja5vXlqx
4D/DogEXMKEhlkfMiybt3e8p2E7JrzEnpefWtDOyDG76S8MPrYsuG54jz7eaiIx42cVhf38E6X3w
sQkICadqGCPNAiaCmViMC9S0tP+bSQKqS1+blRKWr2G6lfNItsde4zIkx8eOUryIJyOR7pFJIEgl
h5QyChYOV32tawL8ooOJTrKAOtY0VoYDUKu1MGGr5p6WTMJwwoRbjWIHKFovx8GSfwKeCnsu5ZRG
S1y1GZUOtSpPaWt3XknnodwJ1N2NsQt5dMPvoJ3n64gdTrMjQS8vQ0vlYG/t11YAra6milWiRolh
FCbom5wTRQzzWqPJ2qtzzkekSthEVtEYmOn9E7gaqAM5hH3MchS847d18q8LSX8waIaSBp6rBcSa
3Q1Q+jWtGKi80Lza7qzWMyw+uuB7YQFzffqt7Lpo6OlWSovjDyMU8XZrSh23Y0QuAUZpolER7ClC
/l3IUUpyqdJQmGrlAhW7UEdWSQBms5nYUC/JtZ1eqJOV+ziCNEgSlTOeM1MwaYq4TbmKGRPYWe5e
4BGCF04gdjT0D40Z8Vf+yjMIheFE7QCZY3N5z4LWstzZuNNCfjAKszgiAwWcKBuWMXKQAGcl7HUR
QqpRxT3XTpz/wkGoRqRZRxG+S4gCixJSC8g6fBofQ7BAtOjZ0hkSXBHoRFHiyrcc/huqnzkMGuEw
xWd4VWlT8vEUuM37R9+ZsIh5NT3UiTzLoBbgAKvJXDLxbbi4Ungpl4zPU5PjLJ5sHOodIYo9s60d
FEXKkAwnkKCexPn1yI8KhzJw3f/Tf86Y78HBaxRII/Z9whp/Xtgda85YHPNHY0rAVlWkmr6R0ywb
iXiMVwfuRCUdhVCZcarP3b0WKVJJSu7DWvuSi1nTrwZxp8vqAeczrsh9m5IsVWBbKmG9+mKQGJyx
F/7zh63EdSEzuQUi9rFVn6JaSE1tjdUtY3UMI0EI2gF9iYGEXJoLLsiLgTVJk6GPJMFas8y9ijMr
B7VreuvZ/mST5C73ssHLohiE13yc/nrMC+/vPc2ooMcR0nQ9dvta6kofyqHWg7S1SazywZkLFJQK
ClRyVI7YQ12eikneySbPSdQ/PvbD9qONyqviOIobruFMJD0aoUTDADTu37ZbsNRqtZ3hLx8AWO3B
euThLx19FVg0If21efrTOpOnThpqRKFqUC6rMOI+1wI1Cd+nS0qkYuBeE/QidC1ShRrxLQhqFUkv
1MU28UFnA4JnG7ZsXPZssluMPZHfhEHMmhR7sqGkrDn+ADsiuNTWYwxqdWZ5ucD4CeFFU0UeIvCn
/vVDswjDh4d6l5taxm3mSTfU98VHwkgsOQC8d3+YZ4KabHHNiQijbolodMyTT1vzshjCXZgeIxJA
cc4zvPdWOPQGmnO0Oyz9+CQWnRVeGrp2npipoqEsKVBkyIH8fCAn05wQxhWAGzfAOusXHsawQXSN
qtkROJSVECoT8QNblroaIkgGOi/DXo0eVe33PUJk4bRsNV8FyqkJfVWflUCRegMKOZf4RG+0x+aq
ZvJzD0Lx44PhoMX1VLZC6pCCk88MhQpnmkzGvRQeuBjbbVuBT/r2YMFB1BeW8wIi7tmpL43TtyG3
gvAr2V+skvWoZl7iZTCKl1pbeBr+Y5aVDapx6SMFxP3znUnGZcuKV3Wr4Mymhxz1RwfycDZA9pMN
m1xSRqznlAq+g3GDJx0hrdkta/7rJGN64Vh88aDA3ehgnrdcPvye/X2S8OwGxWX5TYVZIycMvzMK
AhXyfRl2YKK8czM34U5fK0jbYYkR8IDlwQ3JMA0NItuZVBtQeuiBK9RLn6JM7wXgJRMFrU7iQMYi
6rSNvrrD92uV6fMfilHB82AhaPK0OH111xb7zK9MQgHV9c7U/5V3KPZIPP06c2ivOAwdesQvlzE+
kad18e+9lIzSkZvkAQXTG6DFBbTSRoR1+2IWfYZF+nqLykkJMf6EFcj/zlGBe+4uIY5DCe+76tcH
GQ3J4bKvvxA2Q7WqKs3NV8IcdO+EGmB5gsvk/ShSERs4qjJVdLLGE2IAAHaHaY2EmgtBTogCwz1N
WoV1vk6RnF0qaZG30pZO+geJTuk4MWmicFsw78KzTptg7rzlX6eQJV1zMHfzaX1tbzT0yEHPshe9
VZEw8tkaVJXTHL5UeHOwistfCxkWJpFYX/fOEQ2jx4WR4cwz7bnQ0lEsK1gbnBPP3JBEbpoRPl40
woFiLSfXsN0IFxLT+Q+fQXH4N01mlfnEm4ZB3twDuHvM117Cz2k0irZN67OU6rUN4MjnJ0qMLqav
s6HTrGXUqyFWc5WYkJVM0qsUjR9IdjoFqJyOLSRPagPjvKxVjlunkyootHHmlWYKSQNx+q1VIXkw
c7y3z0pu0JoBIg5PvPxb7fOLyE6PoE6sKqGe/2AQXw2mlcAE146O2BRqLXBOUJE8O2nRSuOBt7CP
UrMNFkpt8UL4gwBvdBg3XPBvL3hvmV1hsrN73H6lq2yeF4GXbkrDhG3nL6xJq6dEj8dDG7LpujP2
r5k/02LyJbApalgtgv4V5HvTWkOu0cH8egsEvM+912peK3V8VPQpoGuyEkdmJ43mclZ//7AekgML
3xhLiGfnecenqXyfHRwYUyAh/ilNOdPYRBheoQC4aVjm9oHqvOOgvvKbTA7f9vnOY/VhedbMm0Ba
y+7N9UJv3LqmNOck26B1AW3TplEhxSiRQpZ2ZR0x8W+siJWwU65GZHgb0yA0bfT8bQGpHv5skqQV
re01R8KyF29B8CFYdDSbskDO398q4sJAVjqI4MyhfhvIqDJhqHUBW/cFZQY/y1tIXaA0DFRpBweu
2K2xfYD4RMrvFXEQhzU4w7jX9cKfdGvVGizklAPazodZuI0QjtSJct0VS7O5ZD4b351ZkJMZIeGF
1WkuZYwSMCfKqtdv/tCeUrHGrGZORgQeKCEFYrjR3YSYRV4iaYrG+PUxUZfv4MZnWQBs7OfyBQYA
DuAZ/dw4zHZKUq3kkJEQRtHuItpugn9xfM4MyGYYfQUVJakcIYn2s5PlTUaKiqvc6gO7nBajur1S
iUBneF+E5Kh/ni7rHCyd496kZdbNFlISAcCQXtGusJE3u5L8WzbslcLtDe/gcG9/Slns8Zdw9m2R
AqOlfFj1e+Xl/I1i1Yk+jHPdpvr7eXvV2SuL3gCcqULDtUAUAZk1g+1Y0q+IfnMcttba+Uc+gDGN
Vt7XAW1ZRobF1AT5zSxO+j62h4T+flzz5qRQviKIzDpBCQi2dnpEVIGFLqGhwQc9sf1/H1cPNXBB
88esE8sjnQERDcRJFk01B44C6AIDiUn6JfhcprWyxmDTPjbEavMX8vivq2DVU+tWIwBgo/GdOX7s
VcdvDu/isjzoU65z5Eq45/AJZf+vLOdaBeQYZE5RHdaTih6FiSUzNnmlwvr7Plc6WFzEU3JpqViA
sKgL5OrYkSZPCzZv8OwmGV2NvhB5+MgbXFRm5BCiTfTrNPkpQiDYhFDBv0jGtQKzUygAxn16w5VX
3Fxhs0tD9RQTOBg/ICHbPrGmsAmIx9CVWq1pfAHp4gQp1+oMUc0gknRTY1KYeNgY5cSx1OtmFxP2
O2sYyo+/eGXhj2sAhcueBy7r/J8PFIIZTNev1mxpsIjA8+uBVmEklxixUOlu121t77nIUEydMynj
Xz6PlHHuZ4eQOV+emTpQ+vetGSmyYprZNwaOyq/TMaRPYlMsSDqS7C8QYYP3OygCDc8Jr6qvBrYJ
oI3n0OJMlgBjwDMSK7raUqFI1pjkF2UlQw7YasSI+Aq/510oZg0C/7xNyBOyIo4rLVYMt3GFJCXn
Eq46OQrxAOdiabbvLbivPnnSx7wwrfDq7CPG8PHEJado9ti6z0WT4vuJkoSPCPoCaIfGhqGZEnAP
moaG2oqHV16qpsUiB7zYUBFV0+9kQGPtZ7D8rmA5EKwpiNe5ZmOmGZqFbO5nQL/KwURDV4duXxRa
GpgcBGGXski/FAp7WRBBxn8YvNEGpqwlDwSK5/ekKaMl+Nq4d0vFHRxPMc2iRs8nT9gntviuxAN1
fmvscxQ6RzwX55xLFTt++N5/h5sNnbizum95SQ5E8Ir+XKEWJCixG4HB0rfdNnLE2Q/1KNLcmtSf
o1lWQ4gqm4L5tDwwdwCvudt9HcKrY2/C7XBsSQ4TbYFD8FNcZ99tRtuM4uvztSQLNQ3iRtChcgIN
4u075vBzS43XkNsh7DgYxV0HKHbrBmjzz7nIg+7dNRlUYwh81a7UmB9tNFYGdcml2mTTg56UCbH6
XWmGkX/upzAwVaZFMTcA72E09F9ToEAhS9hEU3NA2S0pevgLcm0CQ5succSCST1huWsSyQutHHnz
yWH1C+IUvhVAfqI5CSNjTaNTLeCc38Whxk7VTTVWDmLIERtKCnZ4VT83Cdh1Zr1RTG/g0P6P4qSV
lo5NRziZ7mqpiYF9ETCP32WSpBzNmPhOIUXS0M6TeEckzn79DbX/2CRcnCAIoYJQw6Zpw1IukT2F
CbQ52T+hus+NAvWscD3cKwk3skYhL62Tbse13/l8BUc6ZTnT26BdtWDiQs5aKjrxSI+j3cLwwx7q
gGCRMq3cAYxe6TiOw66Ti/F3FGpQqaqc5GV2Z3+kHAaQ6gNYaKqoA7apCSRCopM/+hTb+wZNRQPK
lfiLnQ8B6FkgBmXjn2t3uFIrUqc8fgG/OoFjE2phAXxFz+DURWF6UpLCXcqiJnbspX+m6NtM+5Pc
wM8CCYCJjkSSqInrGI+WS9F3VP3VMUpcRLp3SZNtxvMTxVnTVoEjjPQ1oTLUG8CEf9ELcFrbG1X4
m/+njIzmQAFlGxhWwsOHHHRfP06m2f904bBuW4/Q/4WPWdfHlvRxwtY+Wkh8vDeX1jw/pz7H/IVJ
qDdHeNvJvP6xyyXG0WToSUHMX1IluX/uN5zjOfqZzm4z8lsHXx9K2x65Ujw/W8hPNwXXcEpUZgBz
GgWSjku19C+4+5aLZ8dDYidYzgAbKIIs6F7GjHNbSk4R5xGCjEadVU+7tMSA7Q2VlgejZwUegXzV
eAthEWPixUJr6ECYlUEfkjTI0bdlpwxg2EuI9LyHHgMHPT7C6X0QbZt7JHXcZ/Yi08tnGTxMKe5b
BDRsP0SnVTkwu46ylc+l3hHgeYwnFRUL0pWy1L9gH4fUx3MIQzE5DlPBDGwZ/oHe7yYh7vLtJP+H
bo/2FL3iEXfPXRvqLJCEZbC9mAKcKCazmi7nnAi9AJysUhzxDF2qanlAKJm3lXbJy6wAxSZSl2n1
GRkNRdGOL24xTVSZWvA/rFlDm8ZmfTq34SNXiUKbv5iBjmI987O8qY/9Jpl1PYvHFdlpCALqE6DA
vuMkp+zNuzOk3OZJLQ/8KKwV5f9/CY4fjUP+7mg1V3rujdqOBvL5sQRfuXutMGIN9rYK7rgkZ869
j/g+wWV1t4/rSGIiywgFJL5kZOBOofNiudD2OdXf0zdj183SshVBB8/LZszGVqo2ioswYII6Mc/q
vJMgdmWjCuWCDKMIvAaj1xI/qKWVbVFgGUqXbRCgWfIQM3efnPsfGmelS4St9qCy7PY8Lo82M4m9
BL2SKxsETHYpRSqdgpPCf2G+WtG+jUrSaaex9TNByN36RafeHDxad7cgJdBodCP+kPNTDj8DJwyy
K5IVo4bOTff8cU/b7yC7hdrwXsZChVjJ6TXbt63rCyYf0khGJl81lbUNkGiruCsPBeCoZlbqhm85
ZMxVg2XLmH/9IKve51pleYwZsigqUVPASe0UvplkYPCfCmy/ExDmmWCuqxAiwtXZL+5N5J/tuWlq
IFgZ31DV7YYf8+C3XGNL5JPWZdcmtbBx9Q4vXLZA2n+a6NiFoRW5LerlqrD75qMHRzJxoemZjy5S
AROVuVXsqA+qnCFR53hcucGScZihX9jc8Hh/wuxdtLOs393Z/IPKD+2CYCiA8WJz6oAjUHSwJ9od
YEF67x198lYZeoZIcRBoP6p/OCqLRicKcwSUPGUtd//YHVMCXNhnNu58tCKl3T2jiF4eZh/p9EeS
FkD/Np4OcQB+5AjcqpQoNogRhJtXja32p1RGJWKjqL6g8vSC0nF8sftbOZJdXzBJzen5n0wfyrPw
+5BEmh+5ZkzPlL8d2ksLBXlO7km3EV3YaoN3B1bE6WpKopLX74oVpAWJknT5RaNh4+zbh7UxDdzs
VMnrY6Pu0fnFTOflNLZw6nF+c28RgrtvGFABW58dCsOAievDkDGyY8W5V2Ko2GMflVzPff0V0CIs
YJy96KGMpRJCzF4PXMuOp0zvha4Fbb5/GigaEAKcwpmhkRwnuz4DjydTTcJzds0gPD8J6BMXADPw
d+U1+Nd0tEgIu7+v6FdpFwQPsNESj8HqghCN/i98arVJzelNYFjtQx9MHzAr7JJ669wGzj95tIs7
npZWVTY0BVvHXoK9h1OWqOjZmWZ6gDkNWawk9rJjdTwYAhypBUcf+HSWDegJkQbeMQQ+KqqDxtX+
8T7m/JOOWSfs94VOGLe1SGymTqgBI1LmV2DVQomLglgGI44CqDlb1wxAlzSfGiFY1kUwF4epEJLD
2wfuFvYct7QqXtangg+IpLRLsvfUjln4roPmxRZX7oRgojYwry9vOlKIE2xzQJWZjUEZMBvyiIv7
Qiqg+NCMZL2dvWm6xzJ8xKfFPJTTtjXL7t0t44casbC3/VayZ/jhXz4uJCJLShbsvl6GyWyPBMAT
Qu6v3cSLwgPaXLITcDiOwrggT90xh8FjOEk8AOscHmU/kYXPpQ1Z8qbU4YRkS61Afx+B7do35G4M
jARe3AlyIlBg6S4xbJa6XFFoDMGk0xDTPQ0ug6+zKFRPUMwzA3f2TNqVVdlmAbSZ4bPQpYeKWz2K
L6x1sL5XYkx2DaxuQJ5gjDwo4fNym/UdlPT5x2SFCZibZ7Ob2Ca4bPJMADpS8yBVQkin+lzqGydl
Q1GVkLYR6pRtj0UoGm/x/zrE6SwvS6BZbJmks8vEYT36dzwXL7ply+tDftzf9SSFkVn5RAzUonqf
XASFrwDIgzvSmzQ07H5mjlDt1RjkTnWaXhcxHF/GOzhvK36XLbE2n9FreXsqtgM26NFEiIz/qzy9
EFEkKd1/YhGBgl5HFPdvlVqni3JKTqdzaRNOSZ1HDT4VESJ3JkGni+FKefLll2/LFnh1fEdHlhyk
oSbpuh8btHLFRUIW3lfTtGr2VMqiG+J1WFaJziZ62S178Wmgndz/ZUXAgg3VKhuxedbfhNEBx+MF
bekqSE+oLcGJmQVApKLhT+Fau44Vaw2Q5Lebr7j3Kwtp5mElGTw4kLlWO6tx7KlY4a3y9ZNGHRxL
i2MXre2vlojWNPSvfDgWtnW41hzxWAl3LUH+XBOTmNGOj5yixmIieHSZ5YGhLRerKVAyMLsHiP2f
VGeK4fV2jfY/OTes5z46Z87VrebDoIamkZfL68oRHBTb6fImjh9JXDwnYxloc2dZE5R3boWNsno1
s10rQ4HASgOLadcmbSgi0+flGt9cMPDIJ3B9lcSgwJ955K3MfK0OuMCM1GAkhJnH632rqWkkWovF
9qRqn3JFKQ6dXGU/lY6Qv2DJhvhSdxB3kTEy/gh0Pg9N2uqMQSvcLM5xlBoAu111ikPcctUBwWx8
2JZD5S7PgCPYZs2uUHus9wMwPCR7pvJz5651irQriJl32uH84gAnhph3s3gsd9GGxQYzcQhnaWuL
k8Z178yJ9aHnLXjwJn0ioS2JC0yIbAuu+ZewfZoBLFumnWA5fYVRBdpAnM9dYzhVa0xUg9Uv3MUd
7XdN3NKrgBS/3rytOr5/3E4eq3KD6ZX29oubfVGj3ZDKXyW9Y11neztY7NH+i6cnQyZ7votM8nwq
520zsjj8Fm7wRKFg7/YlzhSHQcDyLDAfS4vVOYOIKza6ljPFp9ys3TwvkFEf4xZSJh/jn5y7GIan
LiJPq5HhwQTDQJ5SeYzJUJI3fyLqKvvveCx+X5toXrWA7rR15vye7mn9un3F06RiOuJ/Tn6Y4GqF
O/HTIz63ys3hvlGj+hDU6Qd5N9qLRNn/jd9Lks9IwQkVGTI1uT+NQAkjlUyjCKLL010Srvo1RlZw
/yJ0jxC8eCLM+I3bJk3jMtqxFmDZOGG2AwjR4pOe82ZZLeofs3eJclYyB3o26mylPqoA1MRkOTAM
w1l1fQ5y4HS2UmVrEUdS/VWnvIG5xHwR/J5alKFojCdd6kCfdCboCa3bxFU/89aYiT3cG9Q+pkCc
V43HMTitVx9crKzw7Oz0+x1n1TxY+O8ai/lBRxszVI1/OlBBo8yIRQgfdNilvMGRL5Fufm089c7P
LlkUOVKN89oSNzKF0+1QJAQGsfg1b3Kdfyt5snBHgic3c7sJSNOkoKOgxQkTQwS26GoOiH07+jlM
LYRLGlOzfIHwpXtgHXHU5yx/O+I2FHdAd4LRKe4Pb2K6LBreefWk58NCV11Cig7X2M+1H3Bfxcf+
CBhjo27ZyUKGYjJlwyKfqsfIgmmvpsNpR38oO2Tn+ocLVQpoPCIJFC6yUAJyfeneh4WrXO/6lC3u
I9GHX0I/af/fr1vq7Eepawz5b+WOaXqIZT85yV9I23akh5vv/Y/gMNuizMX6lf/UuMH0sAqurqna
GL6nOQIZajmklIowSagzW2s/xcFet8gDrKVVxM6w5tj4WP92e2uIfo0Jydwk3TGJc7P9/YUc2V0R
1lFoawiWF3Sktmy8Rfi7ITOb9dcZyZnqe0S3UvV79nyCoD7JvueLBqpF+HI/d5mcOstxTVRzwgWb
g+GVmav9Q1HdBc+cXh3EMe3lIxMqrXWuywZ/aIH7oDJiRWHer3C20WIxDjFmLa6VMDHsodvQO1SV
VjuAgezRCs5X2A8IUGwgDAp+3sfxukc0TnXc6BfYuStWlbFBzeYCiuENFATgSPy0T5gn95YFoPvj
7Hi4P+mUatpDPNTHpfZQ23IcIAA2YkiWLIkRAQ+ahYTI8OS5JHFT/Agn4/XfltyJAkGnEaC4HaIY
vX7RbAErYA1MmrOo4yO/Dr824T4ye4l08apVdgp0Enc2E4QM9+KnnxT8yyvBYSQzzv42NLKbN6Qv
CshE2IJsQ9zLbdZn7cSf5H/o4l4BC0vhE89sJulmsEE8MSCqQldDJMrcUFUiG5vtHJDKO6Xm/Ehx
QOk91nm99pNQ1gyonfgm+7IujPCsMpdhAmUqq3QqwNTzxeJ5q0zne97jSMvzkOmwkr9XnOnmujkk
shuQ2xtk1/DX8bxnT9E31VUiSAsurVRuhhfYEfBpvXPxxG8GtnZ+5GVCH59xUw9qNr235GTULMoq
jzjeHvfUsKTRbOH0f7jv6V8Pt4Ss2Xpvhn2nkN4xw9i4hm/oX2u1gd/pmEX/VoWF7vS7tCSnb9fu
M0GmqeigxBTDzoTGJGNybnufABpAaOizIfLST+ogpYSTsJDeUiZEpU5CmjyGLA2PivKDJKRwDVe8
fb9VksZDUTg/rc9pc8qYwouDGvz5J6br6YAC4/P5/3reyniIw7qSW3n4fBaCU5poQeBRRg1PACom
FKe652TN8maJ2G2HhJbSCyT41DmS8rW8V+El8rcsUDkkdwyaqvS6x7WcbObZtTHbpa9f1UjO6S4U
r0PsChk2v2KEW+pcJrJum16SCZgB3hw1jh3EuIsyXbWMSVQa5BJjzz0ncSYII10R7zWzOZwzMIO2
EH+eojq1z7B9Q8taM6582ipoyZf8iBM7vqu4nbLELh2sDMKoAikRwY3VlQMkMf54Gmog0/KdSxgj
eNryK13HXlCzjQU8vCjhdEzL9fioHxeppWtAH/sIZtqXJ4S4Da+4dczmx5Emj4cmn3wwuPL1M9gv
3KkW4FNPa5Dilcl5YvNelOzqsSe+ydbIAbnVvrq10yII2gUK/r5aMaWYzAp9tiHx8FQkTHyvlCc+
x4p4iyb+YGU93mfeqCAPZjn4JPS5Ds+7rxGCZsBPUSumteeNAtWC2Zor0GXrkOmdyA2mdEWTWlpn
8to4B+G8jM3vynJGNm8aQ1VAg6vOpvjQsXGfMuX2QVJ2/h22JWgnasAuUtlpYfDbo0yDX/s9pNOC
hm14UC9KhKjah9MJhDd5nFPCfwRFgrnrayYaTL/q0/s+kDlY81r+nZB0058YRfn85YftxYxkGoA/
7rNIEF6W60sfS6UgbopYpr+ycObU2BSFXp5es/fmUxPvgtpuAQM4B9ydB+uJqEE/0if2fbqps5kQ
GexmWTm0e1mgOph2R5TXXjPMkgylMoWwaxD6EBwx4P2lw804JrdeGTJ4P+mZB3yT8AtIiB4VdMMP
esc5OLNr51JRu2tCt/R0vEv25i0sQ74VyJJlHPGs0S9PDzaRKGLzwp1DE2dckrT9CbCc3mWXsfP8
Cd+GbaPQ/8pjPrkH/LIy0+Y7hBnjzDXwGQ79QmbANhOPq9xA6KAPb4TqFMpr4UiSJY18gUbWI9j8
eeOmdx4Dwb7iaX08PvocrDClL6pVYSrtIUMwCoTbTi0XUUR2CiBps08aOCydLqhPTjzvWRZCrXGh
DHN+gl2Y8CLIJCh3AnwdzyZDVtg5d7aDi/gbsD8OzqoP/5zFeQYuAhbEJ1k4pdR01fXBhboOsHEr
oPpxLxqFnU1AM6lbGFftO88xQqF7yAMqz2/YlIYMiWIFUBn45XTSyvjttJHnM3p+GWo90O6U1PU3
ME08MfpeGkBEAHKBanhvXPW8T179nch3ZzUcewcV05jrqOFeGcge/XJq5lhOjQuAPup5SLJCnR35
xN6R/5+J5QxcbegE//LGDvwV1oPrHqh3InCTbdTtZnLsi4BvrmEoxJ924+yQbBABjMB9PHNn698w
ofmrggmVcqZ+bnwHHvp1ph3fS+xYhtsmN4MgoBR/fSAgc8f/C5qLvTZA0i5rAIcW5usXZPsYandG
Ar8W6IMJgd/0upsnknjuYHDeW14gms/h3qRsjQ7JoF8JoFF/UFrUKbA+JaBx3ZZgw8VAk2PrNZEE
Rhe/bvjkWbMakBUpb5v+RtiaNRjvk7WhyL/ovMMzOv+1S+NLOdFKJR2I4LjUYZHX6XX1NcIUxNqp
fHAaZb3IiwNAdpugQajDNLvC7PtJp2fPlrr4NvY6IHDlxY4UoNX1bEIJvFjrtGeCFZAMydJM1BQc
QYnqbCmXWXSIT9QQvWNqXMepz5yY7ve/EcRsXG5kehQgcS3Kwmm64wcIHsmmnu2b+T6p01Oon94J
lF+jROS3dtSRTcytIcvPebdMo9QckIl2XBWIIxQDP4FcszHGBkgNBXl4/wcaR/eglETVb5ALF2qi
ukluF2mzPhmNU9Z0yQ+UzGsScnTxslgnQiHe/ktQ6HnIaZwzZkWhMqNnxpRsbfikPQRbfRxBrd9h
6NJqYmCUxdYALoPXhkcTFIEa5KNJI3VmxABNu/DfEUvzh8AggtOBzbsY+7UKnD6HGhVpgDJ1ehiv
OxePVQYxslFIEAsOUOCEj7xMOztkR8aOcUnvsU8wBB+TcJSeHMRAK8oAOyuqY9T64jfCqCNkMtnP
AQqcJl+NcJjLmdbtBJtF53TieyBhvwLUZ2Kru/OCazaOKMkOITnWhMqXSBBOt0UkbGvzK+1FEG4b
RTfdjZy6FYgb3xnEf1TX8tIlE2AjV3jNfwlAOAscXrDc7qhCIhII6/BJo7OPXSce52s7TBJcjkhA
7TL4Sjtw8QkbrfN01iN/WuQZiROqDxGS5Qwth8B0nU9WaalYRG7zhxwtyxg350bt52UiGUSLsp6J
V9roluhovffhMeV49ccGSLkoc5m1TQwmCbMRuUVTN43//pW+rrXmqHc8bi97EOlA4hjr/dLph04W
NrFvdDu6lCoZrHix+thA5eu2vu2hcrs8Y+XT6sV8CHJfkH/V5GqnSzciGXBYoIi6OlY4QW9mHEIY
6lgFXDhTcBD/RyJvtgqEptirQ+GbgSqUb6EDoECXjIEI/qNG7aonM4kiMt5gamHK3qPgVt6cdtD6
iF2NIRGf2Zoscru7QfTYTAFMgT05n59jpAaVlX8wONTf8C0FkqwA803K5VAfloCZHsGd6j8tNYr4
zl7/mvbILolZkQPUpFELVg8cswUKAdvBAdSId+dD/ac8q+ws4wIlS0JsT7mh9AXJGhpHUkArFrrO
OOMCgzQFJOM7X/EKqmhqcXk3+Qda1uzCG9jd6aNXqP3h/E5OHp/LzzzdmlUI00AtUy9UkQlT0G11
Rqt/6Z3IFURlAy7TOBNvPqyVlWxMul6EdNHeNqJ2YScXHsAKti9s//BGCAXv7+y9l3M1uGSqceni
COE1U5fZWwc13yKVeDW/egiTSecuKi+rPZKERFaFBOq3IEQ5spmQJ2K+q6kxjyYNJp/hIgQ+P/hu
vuP6Z5NJJfGR2o4KFnXJg3y55ZjbKkr3ZbZ332dH2clahgZM8AXW7HnUZyDp3dcm1uZx7EfiOugp
9iWRXVKz3a3KK9Wrq6YqeOMdepaiY4zW3cjHPxfXOVhbIPFI1/RmlT2geZEec4hQrQj7t32ifO0U
oYddg/gpxSBUDRnhLySB0vn3UZCPV7MM+qTHsQ75jjmW3VEN42F2oukZsOb0cVPomIzcpFdvETHH
9d+3JOY9ZvIiOgj8NtDpWL5asxz/K2GW70MPhM09WIegBxeIhiY3D+q9xGPJf/LIQ8wPrhjQVoA2
9xIMuXwe426i8NoItVjf932rWgOJZLbnGWqDMJsZCCUjKpmba/vFacb51YnZQTnfiYNte2Dw66dA
Z8V1+Xx+/i7ycPpZr87fw1oZ1R+SoWBP0BoPhUa87bJYdQqfC/ifajJ3/J1qaFJtdrcJD7xgo9ce
51UvGFFQerCYz4mIbcB74V76LeEa1BFu2VRLteSj8JAJmE/mFnLOR0r8R3kscdjCTjeopNArILFp
ZPftkn/uiHg+9QNV0qpESx/NBeHO60XkEJBBNYEk+7uj6S1xFmvYjEluuXBgxsisfzNgvvRyytDX
EDpQaMrJMCUuIJrs6h/lJ5GsMkNPY5YtmBzaEJjSVmApkdONezFU4gn7Z1mvGcqhfHFSIJ90Lb6p
KO+oeKZRT2xI3LWuACYm1ESmeBfpLCcVAXtn+aLklCOHd9V54dm4OZigZhxT0J36HHLV2CHIWFfC
EguWpDYb4U7/ald1Zh96+vwUuqZz0cRh7w+5PqN/lLiAZIhge9uUvIKRCtga3F5dptPgi6F+BzKL
WZVO6OstyvRMUdYpi1mHo1Rnz3ntQoxot8pvBLRVm9l6V53shz6pBr0fOec3KijCQo5LOXNENvce
ksTYdvBiAIN68b2qRmYS40UNA+/pL00ajaPz8LTpI7CPByWgCYoopwWnxcWYkxNwDKmjBgZTKtL4
KN5iXATRk2ji8p1gPjzajIkkv0YuSSToS49npbhMdeKmJNiAT2YvIV/EQCmB/ikZ4OczXl+7S2Ag
kPZRcN9zvcCCFOCSPfpNIbC7lVc7B5PCysBEQYIsDptApmxa808JJrQvN9RX6C28ml4pSi/TqzP0
mw4twTP+ERLff8yD9zz0sfYPXHjp88OxZZeJPsCXewuMHGZ4ikfFEyp7HfQVM4qqCZPGgrCgfBfJ
m6YXPeniidZRxIrZIELf+Typo6nUKzwgtQpQc6OxxGSlHEhI2jzoJNHHeDpIFIgNnSucnOW+Q+4j
KA3GKd6pkWyIOIxNqQbWto/kJ7sgCqCC3BERR+WgR37J6apK7xL1Wv42lf2v8huN7aavkeLfd6I+
rAlmtzWyJTjSisT046qPdNqmeDvT8lGtyJDlmSWgKRjd2y+oP5qa8Qr9GZi6s6K3ePHQhxWkvU+j
1b6DYBgPdh4+Z2JUApSxeEGUFrNwNMY6ndl0dJsWlH1aAM6fWD+mR4K00eZPEO9QoroAY/LjUicl
jVNyP0tdSIyXJGr5+KdDbCLJ0VWg0Mk9H2eBEyvJ4rYBnXs8ajLc7HgTvFEOlBzirqBWQKqmADaz
pGZdBKJdBZnPfji/gnlDh+vSS2DKR5Sjh4am2yIQg1WoVTL0yPq3GQ2vdrWNQi3vshTm5W1R56Ts
3vo+QTQbT4yiaj86nQwphYVeIQGglAQ/IWu/eS/tgAF76Z9q+nwoqlDSwgffm/+TGzJQiYYg2TwW
dOx3M5qd1J4BJoO/jNH8WULWK12snTjRYFE+RkdGZR3+7pcD4C3cO5IJ+DOQp2pJ/bA6vJWAZ4yf
TiT5KygZ5qT83IBQ5BX6a+P5Tj+KHQIglycKeedL2VvRsi1mF9FADaLb2aeJFoAxP+b9KV19OKij
Hol2dt/Nk4CvQ5vSgIWjRz31G8hhzkyuH2dRKI2VjrJkB7qmZX+Bwatk8C1pR4N13OEiVWJa5UZk
AFZyo07O2MceUdZdE9LQxrpB+F4+62OONZbrl3wvTGGeR1zUrjFJJNvG4pnl5+RhTAsFrqsJFbIO
Q5Sp3qe4+hItdUSD9nojjOzIozspwkZhR/KaASfw82nkhryNgMl3Hn/UwIaaXK/+nlDobMY2g4S8
MJ6LEewR5JxksvbfkMJbopaqQgKGMyOTmDQHg3o8UiDvtULqqJpczXH5ez2OR6zWexkSTknFBeZL
7Q/nMOcLtoIhBGjuRh/QLBzRkXRIwudFLZP3GZVrbf6AwEPmUk7bnRPMV7q8u+eDZgSwMniXPXFW
gNI8jO2Lg3aCIgiIPq5n85MecVLrdUXPdoANPET9c60l822y5Bmka9GNByhiIdlP40HIES2+5QF7
Oj9tGp0PMYPKYIsE5gqHxzLmy5EIdcmt0+JpEi4MJkRH26E+OkBfwVmiKDH0doVlqielb1VOaG3S
LcedScP/QlSmqafToh8JnHsF/CzVs3hIFvwWbcDprk8Z4Pqw6qY8gKeTUm8FY0QnpLqy0qfopZae
JGs8y94wKHAwsVvlcqk3k0cSrIke0qClRHj4uxxa27k1JApRTysTUjTB174mODO2Qt9ZL8pSDe0J
YTWjMwcAP3jYOW8ijEo6zkDhPnzXC5/YhHFdejXza3n6KCiiFwwjBFoo2fyH2bxn0WToipJAKdNJ
gO27uPAnK0o9+L61QnA9AQ7/lxmitHoCAGEUmaeLaLVVMGLRL/x6dIv34c7LKG329eQv5puC4Km6
WxQ1S3rxl3q/EkXdQEf3mXNfcrILXqiaTilCpKkITCrCsE/cG7OHh3qhk9x00tdjQWjPa73S0kTY
RH/RaDwg6VN+TSZBEhCkkgZq41EsmaVv8sMlYQDdjrJU5TZh3vuJAV2uhh6oTZhvEeVXqF2Du2QE
PB8uupYsg+g60fVz3JW6rRYE3FAmjI/OUpWfoB+AkilfZp/zy/Pi47ChKSqEvBVI3i06hbsRc68k
JAjiMO2bTcvjqHXoytsL0twpiHxJqXL4m2Civba8ZDhlAkl7LhTRkzHgxuWG9Zdmyv9kc72IZOKz
f1YcCzPcG/AbQn5whbTsEwdUjnBUfM+0BdUjEZuDbMDpZ8Jy8hembC6V6LpW/Euwx2tI21NkFyqI
7VnibpXUkLShmzxb00AB+rwcDw3+56noj4hC03So3eFefGxhF4MYppATCjONNEFwa26xtHk2CIj5
OQVTZ/BnGE0qaJh5MILEn/MviyqrDvAYivb6i4TDecvLaGPixhvNoV32LmylY4YGpmJL0VJEeuG1
qDFpSLCcRfWLKROIzTEoGUwCw5YaYTTcmCl5nwcqsbYJqL2xURfaabSVdq9YmzfDHAxkG8bQUMbZ
oivGdcKykhfsv4d8SvBrRQnRo3AS7dNsEpfW23mcjkqh1UF/PmHioexqiHVsBjKuzBjjDWrg8bda
fPF2SSPPvBmA19a4pEfzTyuRzRgBkxvI4bwZIKLWYqzQ4ip3dxJlZvTGagqamtckGTgX2CjYvfRm
XYEfN+5kAVYK3Qp3LYzJJrYF8n0mP5WkHhrti6ABWnFePE7W7qAYBFs7At7qsOGLOIgyMHCujPb5
sGNqVDs36XmBMwkxr05HeB+oT7nQRLzwxz5kyEJ7xbqr5/JPFfMW+EevxOGH35CCIOWHmexTAk/5
OlY6buxiIJ7VrdfwhJr+HhUoPnTS+6BcTu1SQAErm2DD5LLVveRnoVzgn3Px/CcdRzmWtumLY5HZ
pI1pgIIqpfG0vaUSCSGr1RKA7vh56x/k04FuTIC870zKd0AbN2X0FZUpgtqbX9HqykZKfvgTO8NV
O7VJ4tjlFTK44WowRtQ+H7ZP9brcrvOcqLGbsvdGHTKMzfXaDQIJtvY+sNahIoVkm/rYLX1p2IxI
VQf18CUzgaitzXCuAVG6EbfqHbFvd5Iao+QgY7f6mpfH5sUlZ+hjklL1LdxmiCdRC5maAizsLaae
Zj9eRm0xEnsrH/N3PVuacWHQUawTBn22AN9O4uD1ljfsuZUXML3RE9XQIJskS/ZO8LbLGH5CbqY4
ANAMVaeegd8to84trH+zyUoCYxEQczr/rhq+0fuXa0e82/2948tdfAN2JEcytoPUrwmK8rGUaCwA
SmI++y49nMX5bETLOHniAnxXAMR39dAOWFJNhm6YnWjaDz5Q2kPsVoi/dIvZUacX2THCxFqMqpGn
U5wc2mxG5ZVCzwpMLQzYuOjnZsXC6GPl9nurCxQZWhI6Zc+90mcbeKPu9sCWXFepiUmdXmApqP4O
tqRi/YTCFaXlIR8dfrxDqIHEVf5b6LCgrkxATruzALTC2EW0BQq+DJlzPuc6z/70Pd0yXkusPTJX
FIIAGur8atijW8U5PnOrzeZh062MGgnIPye3ekmL/LO0URaaKTkO8BY47zGak6VwUGwmMJiXvep5
ryXaHrPkLOQqFQllTco8P5nbWd8/IrVEl+tekjjsNJyoNX6O53z+UsWnAhIc5frO4ruWjR/hZF++
D7BRgWpzqQys1rvT5Y3vn2HmpGZ0eO9Wehx3irVzjTdUzqDNeM8FTqqyKbU+/CP0V6+8+LMgbilT
Ypy8TWEur3+mr1IxLFAbv6aGkkJt2+YB+UvCu6ndQg42+LpkWSa3JqNvBkkMRlq/GU8wH4EpBVnu
A2d1K3Rl5aBy3Vxmxy7B7YiSECmAYHi0bkWRms8lawMLBu4l6ePHq+veitviZarJHF2ViIH0s4/Q
G95JNdKi+9cciRW9C2D7c56hNb/f7/NWu7wz8eSPL2WLmKAa3edfVOxg0rlhCHy2Qn1jzCpCXedd
DhQ2jG52FgO7wYcD5UtVWlLYR0RB/b+Y64z7Mqlu6wl7T+I8cwvNUzeBf86ERHyCkOg+AILFEImj
8GHwE2CF6LAhBQyQ+djH/dqvAldStze7XuUhRLA9dltCgvkWo2OL7qzJzzxFD/wfJHLA1JNgK9DR
3ldc2UJ01q2hSXNyS35WUH7Axanr3rNTWR0sKNeQQ3Q5LcuoH4/RLO5r4EXRPmMX6gOSphJIhMC3
kbw+qQhnk2jEi7q4CwD9ZLKfHKzCr4raexaFocbEnZZoF7fdkYsF5wHD0uWX50Zk1lAf3F3pXCi0
Ol6eJRGiMKcUCzy5qLBrf1ugqDbk0bsUK/F+Yirlyb5vT6rTTQRQWL1HjebbyPGJrX57xDIo2c3G
bncwGTzBE0GAVtJG+rXRk76g7epr+lJgtvGuIp35rdm1FlbGnf1XON3YvcLT3fLxYvvJ9/8BtT1D
8qw5uyqqiqBdVd2Sk5BJeQM8aSmUNLcMbD5MOBr/MlA2S9iUs8DR2T+iLChbq50aAqOtj3RJ1U9S
eRwbSdVAsFZaFGt1xFv+dSOXgv9GEoeax4g07yLz62Uep5r8+nQIX1B0TJYXRbUiEt+sIP3iTs0h
AkxrLCeXLomZjCD96ooN8lLs4BU7zw5XM/CZB1xdwMxsSp/X3fAVCteSiI5LDguLnbQysLVE+naJ
e3vronskLAoLZgpdChz36Y5ZQj0rqxtAFo+sHDh5okiNWIJXoskaSOpzaoZOTbPadgiStPh2DT1R
w11M+c46yCEbmKtTGlx7ha6YSyawsG9E0LOAjLf2mgxmisI49afYqQmlb9pUkvRfaRdN/Y8dhpZm
7nUkwmlrORuMGYjEcxU/GY+M5Bs9bUb2PNa0W16B088/7mwav6GumJ1Jz3lQQlx8hfeIfRQKsmmF
m5dREp6PZwqA1GZBAtazvS3pH4OBgJrhq4X09lRCt4//yzkAcRDyu+IV7bUQkoCB2PyfFIMZWVFR
K2Saske/ysqL/C7bA173+RjVHnqa9tRJU1ahR2KAhCcXCNxaJy5InRyg4rX8EBoamJcvEqNavY44
sioEpI0/H8rcmTUAB7FyLtSZx/2+c7b9JgvRaNtKAHKfBVVRyTcMAwO0UuRdvAVZ46HPZMb0j5LJ
7ur4539Ga3W2kZMuthQ1DkqKP7BRnrLnnfegAGJ6pS2zygSyRza+bNeA5cVf3PsSo91ymJ/kJDX9
6yvP/Pvw7mU+LaODKADX8/uZqo7l7D99vyJorKOqD2bJs6U1VsKw7/UjX7mrE+f7DDGmtYu8R+SR
GAPCA62gkpVnj58v7abkqRVNsaQLfMfWcRyPB12EmKfkm3ZFkU2/vPjoxLolOrG36iN3ZLH/77Oe
Yb8pV4le1aVz52yPSCh9Un6LI46QEwqCUJeNSySAFv0CCBl/LJepNDPc3IP/ZzS9v0k4qTpkvpUw
YPzXGRP6eHxzZo2nOYHvCVqH/DmfrZAt9npsx5Cle4h9Yc5sSaMXO7UGR6vA6Ti1UrJzAhyfc3HF
GMd1IyO+49681yT7vK4yhRUNhbn6LArw5unMz5y0uA/4C0ZigUHBDL91xqBOVT8ocXZ8o0ZyfSQN
JU35/hXrnDMT0KyDfL6psFmaLWrTaiCYlzM2Lr9ro9NaViZBOpdMu34G1xopMqWm0BrwD1mehJqd
d6LNX1wfiBDQAEux0EEKIb6PGHMuyE/mJvyO5VLfQly6oaRzuoX6hrKflV4ZwFjAStK9Sh1riWcr
X7KArUZOtIIlTiUftcbjiJ/IpcFeQpX4C7JYhwG3rJk1ly34L50JZwacb7Iwb1LN1ueNyEzPwDwq
SGu8oZ3i1rFBUG7xWa0rzNE8FkogGU+54oZ1v8JSmidyHBAVtO1RxY35pU99/Ecgj5qKZpBnFqjL
vZlfc3dtD+gZSmbCGZd+pMGnu/yDtwqNwP6a+0AttlfSHmea24kcp7nk4OjzNI9MoZrUCvyiQuFx
lM5995ZHCpOlEVJfg83Mzk+MtxY/zy3M4n9ZUy1NV3wtC4f1Au3iwX1Rst6bEF+lprgz+YUSM2Hj
RzOEOUU6jwywVnhWJndmyHb/W2d7nAekto7fTjUBlKYk/7FVClMCMfM6Z/di/uzG4Zor8xMhlif3
pz8CzKcnqN9RbMJAHeaN+a2iGYNzx1SLqG3wjZBoiICRXdjjInZnksZ9qptI/ByFHCKVEy9QfUnr
GQirjjsIiTLhJdI5QzfKXCUWqfj4DcczDQ9OZl2u6KVE8Xh5ZuQzQH4Ecsmo4/xU3gB32QYGAob9
mrWSmrXS0rv3I+MUkX4/LXkXCfIoAOvIOYBDhvSAEIJA9DEtoxfIWC9nKmTlMFBMJdDcx22w1pO1
LD6+hg/0hT5HWlnfdPhcQFvNpjemG/U8WaPOAeQ4cVgQFWY6ujgMgX4VedUMD7ENfQ5Bdewnl90c
LK8S6He79nebpZYUmkNZwf8MadiJ800NqET7tZy0njjFuRB+vpY98vD37bY9W0TkWqXRrIzNjIr8
cm7IogyVz58jW8XLzhGgFbkAqRGmzjcfBE4LzkrHx0q3EJbaFm4yBAIpTZWT2vI5kxDxe2uv1GGB
8U9g6fT3x4hnkp2LqfAlyFpnOuLQdPnDEqUyALvfL6DWKg0UGnsZLZX9fBqrmFxS6PDhU/FjKGmc
vFGAtp/N0nCbVIU4jlHWdillfzt0hB3iy6bi86n4U4fYH5qd3iTuRlKceJyCDXJgDVouMRM5bkS6
K/A3TZHEqImb8Mnivf4lsAlKzT+0v6lLyCaiu1LkItMmNaUx94bIzAB1Q7rRrdIUPeu5cSX/mt5m
gV3H3VKRQFKex+X8em2+OJTCef45I1dWy/yK286H69zghvLyk1d0sMuHys5C46FL1sYNKdhHhgcm
WtqBmWLgfQjdpFkAPTAXjeE63tFH2x9oknvmkVi8HWxqw8cW1RFFIb80o64WMRmVoFXNTCYMS9j3
gYZDa+9UWCHtcTfm9rvDbtte/3JuK0KDOtP3hIRy8IzMi0+oTiviGcmw8SS64HDw98vIG+ORodu8
xTQOYh+Zp9lH5Dc2qMOd/QlyydR0+Z+PGWfLy1VoKEdoIoj8PT/y1NHO1a5SiHhIyMZp3noaL8aN
ug5H/JO/kuh+8MuiZQHd+lYzXs/EoJnzUwW/bHaVfnI3lLlgN+iZeBQVl1pQ5AVc43LR6+7cFgJb
N4jtx3tRow4r8m7a/gtkJJ8ereyllrJ89vd28qbldQSpvLLMzARFhQDX2xUy/oeoHTcMhiL3VxCh
+BamO0WCgnFx5a1PwVwqt0R5j5BRzf8TMJIPfIBwO0EFrY58eHLzswD6prm7aXiOgReYd/sSNyQV
MkjNIrxgCJYk1D1EU+5jNMZRnGbO5By/Pn3PyrNn2mabUNPknedF9ze/2HLk0BbE0tJiFvII/ijT
1R8yzH7fNQBUeNmkKt5G4XLWU+SdBWYu7f9znHokI3aAmtEFNWo3dVrrbtZcc5l/UtGLiT1EA4l2
9+4bwwTHcGGnk5YHQx9ZFmPFmYRD5aWUk9/I5tOUz+KbFl6pW1bAaPMJxJDxaqhfY0f/R27WOWat
ukvitT6huR9g3Vwn5sQDohraImOF/ArVJ05kbd7g9QfAnVzlHHvGi26yJChpou3UQul8JD/RR7BD
SILDNQZx9PwHLmKIf0s1NpjQcsocCLLiW7b6bGPmDrULU0WtOCDdbr40jIgGFRFDiCJZe/AGPS6K
FGYTEgSD/hr6Tw4IFJngrcc86g6zImL+mmXaUWSG5WdHi8hOeIoqXMEsPWxmghaC/CwN7pJN2j7E
gt5g+ECGusCu8Cug9cI811Hf3dgjjVoBrh7Jsj7N+x9iIuFV4Wveu5xX7O4ycqyLC+QQ9R8iwhB0
KScE/Kq/deosejF1/3GOJ9YY34A3btKTM+sz/+QitVO1FrLEZN1vUZIdi0rO5PSKUJN5s0wvgEAV
HTJ5SsUmMyORT368bj3ouLzP7w6Xa6Ju/97IqSlnfuxoEcS6sXn40RNGQfMnoI/+MdWXgJPfQd+H
rG5r0prUu/I7joI0Did8PVvEercq+YX/HQlGuotkC7+TvJwgQtz7vexU7IHoUT3AGK5R3Xd+wrUl
5Ox0O3fPV8tSL4Xvp0YkOetGbPsTLIvJ2vHFMaiA1SukIydU0XYi2CZ8lpEFENLSO7iTL61Gg0SZ
d1aZdfoLy2Kdw8njmJe7H3eiKAL1WRHSwQxI5os2yntqXkb+q4VTnoL73LOh+FRiC+bPpzo7j2oY
RcI5wrDzxf0+n65I1xvDCk/QMuxL3rBRD0jsdHVQKibjC/3tx5q+mMEkqWG7P3xa2U9VhAWIZrsS
2S+KR1r4PGLyDLmfkydkZ5okQHS1ooMiPyddZlTF32QBJACn4xBxl9E80PDDxLdk5i2HwPXgpG9R
8GyQxlSFBKiLV3YQ4TWzCHcbUffxKtmN8x1uN+ygXjScYSi3iZdYaOg5ePl2hUwDvb0fSPjrAFqO
UDuGvRmEZHe4fEDC6p1bUS9inn13KJXtz4HohzqpWDW1IcK0ofiBaKOzv8LWl9TcABES7iGF3mrC
kxzfz5oAPKm8wRKf/HYJWehkt0BWNb2epMGR4gNfDF01Uwpj0zyh2XtqE4FoKpXKP2WtkTyWhNoj
x6X0Im/EZzRReIVdnhuiq3ZMmJ3KWuNAguRwCmxY9+0yUnBgNBNBIUyofzE3dFDyfVYnwHrRS8MM
b7BMsIlHCYxFU/wUi7DpB7x4SkwV6towFzcJjX83DpXpgUIvi6rNoUn6KkylIR72zBaJGkYBkJ4I
FWug0Sn1eTvQkA1+duwHL6EWAJw4mAVYoIOUuUmX4viWt2lFv5XY9lKiL/BB8Ht6kcEo3Rd2LFq8
T1H07ok0xBnaN3oOg/enc/gM+1XhkupvSO4wzSaNRYxm3vm9IJDIjESa3aDdpsNXfdbBtfp9RK84
kVWsMKJfZDcyhaIehz3vaYpBzj+2yVWSgaRV9bcB5r10TC02zn7o/LjqrMIKGUdKbz+6G5SXhXdx
m89cT1euH7K2BAguPI8vF8+NE3vZVwADTVNyOoIEcwgD7tl1KqqFJ58hVOud4D7R3GggQmoQlllK
QGG5TY7+g4JTzcoDEXaswv7FHvAQjBuL5uR3HqX/li/cr3qG67jPqVKgud4yHk5Z+TfWBFjpuaj4
RgC0eqgdUlD4Ah5czfEQYMbWtzFYMotXwtQk60+0hvre2AVBX6oS2kcUKevZNQCkj352TcnesGWP
oQLPSGhKVbKGhIGWiyCXi2mfjfjn45hQHfShHrn/lQIRHvRvm3n4geXJyoK1YfTC8AUvKzTflVeV
oos5uU5fLlKBD/GUCTHmTcY++8ldvCv42Kcme8XUdfmoLn4n2U+DcsJL/XXwNpUjlmAjNlLP8JYQ
ErLvbZa0wui5pMMO9b9p7D+wx7V5WAMB/gvJPkeWs34KuWfoIMzqYgHAMH0ygJEzzm4Our5lkIXr
PB223yWtItLGgYlanSYEDp3zGltN+OBKwDgwiNbYFyWb898MBcBPqK/WtxvYUBOsXUgfMfvzz0zR
m1eizvXHPYvFkpPgVSYS0TyeGZxvWFicI0skiPMlo8jrV2t+Bk47eOMKh4asWIvWG4WCiIuTBGxm
KKcKI2D2wf5bq8Hwm3RUpOKJdNoy3fU+lyjOvkHVlh+NxNA/Xa4GjEdSea3px+vkmNZ2KNU/ugtb
+y47zMlTFs6Z1h3Ei2VTOENKeFS9Jctacw72EYtH4TpF05wkyX5aj59HA4zjA5kS8Rugeb9V56KH
Ox86/avrGPExVbPwIM98ArpBlhzVDeYtIRbemGlQI656IRfovfBxnaKZKpt8uf8sb2rM2vzCc4wI
H30PqBVn7yFn2Cl620bv6Wiw8NF+y4s97PEQ9KZnwoLLvnpIHLafJRB4yst8vuGfHRIOeFhsLjDc
6CvWGqLBIXLj0lE6Og24h+NswzH0x3s1yD4qrHfzMsYH4c7iflIms+qTRKGJ005uqFNzf0hIzBka
KNkDa/eQvmXgdogXAtQDpStb3zBTCRcNCGZwJhFXtUgw+6u5uc7ESMHOfBsNe5wn417qSWIa8cU3
1EHsGgpjPPnveuSfgnzQHP9sLEmFR5QlrAogQsdNVVx5V9Sp8Kp63k4OHZ8cJiJW7b9sL+q83hCb
PQFg9jWT+G9Di2WtxsbT1R8rMffD8jZc2/3dAOsuSPtMVKgnErBE3uDMLOKBDODO0cFjNNN+Aj01
HnxWM0XKhaBidnEhSZu77VtU+8iz1kBViFGdBhRBufg7Dmr3epDBIZoT0jc8IE9DEDnxEcwL1756
ae533RFt/DAxcooRfjV9USIdyZLUtYpDsj3rXLIUBeq5OG5N1wSUn1D8Z8XWBuorB8KGvtHNN1lG
SKM16KipELTyPiakZzzLLWzLO5n8ZNqcVR45kwrc2pwLmO0m7eknhtxFi3EXFaftx5mK56pKv+e1
n0MF5o6NPUtEhagG26C98Y0/ruMlzzm3t+sfM3EOVhjI2wZWZwzznyyvA8YDR8x03IEPCz1xtyFE
Jctyc5h8wGN7iWYKd8/vy7KIqh3I9Qu5jxal2sfWruauQ2M/hZLjSkm03LLL9Lw8Z2PHrZm+GVEX
0PRvkGdRvWXM5qLtIRxM5jpqcmHQ9kFBY1pgqffIqYll7/IfZStBfWLoYMxnlGZDqmD2IDt6i0gs
21VBwtgT6I1OsrgBx/+DyWUfStPugokRJsJxeAS2tFhgqC1DNcNya0VxPhwoFpgAPhSt2YqE/qkn
nc+PU6S3i+VMtzXh1KJRWSDEX7XfrYmvqSwNUQQudJaSkM14gF433lEsZon/YwUXZLjxvGqBym82
zRjTnii3KWJwebVAKF/iqsnfjeJHb63FXjEBVsNbNR1VCCQP5XjWJ7pDN0zIfmsy1Ol8QrxlZGo/
XhsRPapruURoZQDth4hptlbVO2Ol5LdUGVG+7jUeu/BthOt/L/iawnS6IxbR1SvYH5whvYY4WGyH
wogE3B6/+7Vt0ZFkSzXjku13Qe//gn+zgk1cHeGY0wWiFD2veRR/DiVOAWM6KGA9WYxG/MjvHoTM
FXWXLiZJLAFXlWvEgNdIgW7B6C1ZBAA8QObovXyEVJJXVL0wcGpkrzeUXE+Kol9ftQKoumXHnW2I
xk3RIguDHACyARGi0H8fRAH84CKrPnr6IgneWbXk2y3oThL4g0lriY4+9iGSBSrnqwzPnSRWtTNg
cxDkw7KmAh4sWRqvvSEu/1W9cBUMLyDUApa1nOixy48zN693yaGzozBOSVbQnmWjjn2yucqvD2xj
VRpO8VpkoL0F8vVGFl3nBhjK/PK+BcaZ/AWUbLdAeo5fFkuQpQJuGHfZw3HMAhUtTsoaGx6iF6cD
nZMpzLy681o+u5Lw+ldgny2HMnLHBG/SSeABDMdfdi8iqxEEhpx0g61iJJPlc9BwztYldFa6XhK7
4upYdt79Nq+cdJEdQB+mhRUMEHG/LNPu0gbNbRGM9vPQFBSe44nGA8QR8LpDmM6cSRq2LTv1P+nE
RVBB+2tiELPYzKgc7N+G4qZKT2uHxN5QCJ9f75Q/NDT1xeCl8mIsnKbpEB8mVKCVb2jWKOsFh1fK
daQViauXsE/67vU8M2m4LT2fRAIXnj8hH0oLSNFw0C2EDxj+VUvRqIcYba0YRNmF5OMc6fEiVF2J
7SAaj7LHwTwvdLIwdfBDQI3zqkJJ6ty/as9XYP/WX2L+Ij8BqxeKGhFOoE4NF6qmK2GwBkO1nMLo
4+NyYYqtrZI+VKl1xhWlJyaBPelyTHkP3ssyQN1RtGbbzNia53xEyMK7VQR0p02LDfw+wWUT+96i
BQnoB0AjesEYpf4zSGFzYfTszE+f/rEyjrF7lNo8e409CENct3kb9QIGvqoyVzBDtiWcmBgv+nT5
iuMs0KctwBNoNt1nnjIbepGtBvlucrR2rTHTNy3pOY4uHq3De4eztC52g+u3r/j7AyPvsate+uJq
qoP+k8J82Fs84ZuvQb0uSOlgqS3RMf25GdcEkjKhZPJdIdFC5mrKon161hhkVyHzoK6xkwgRgtmi
zv8Z0NfQDr9OHEOL9jlnPU4FAhL+KFaqMt30IUtOWtWiJOO7U3nwrYbfshrtn7/OwsExIBBXK9WW
qlfsUrIj8bGq7Xz3TcgoYciqh3DPvZpB4pv+rIrbQGPOHQxXiliyuALaY6LO3INeKQfWGGLj1VWI
8YkwZm9OqkjMDsrK7jnEoPOWGNmieltNHp+6HcJQdYkh7xhZ/eirYXV4WkY9UGlJfbbRwxD9d4We
OwDHVdPus4K49fxtgXuEMzKJX30Xnc1dYceo3ZOqbbUd3TYEi4Eabtku6p4ggRMraqLQz+InS9XK
qPEedPlrk5qPaof4s5VkXuKlZIqSbNMYsVSaGk1o2+icV52bvLEhcmoXu8745WBY9z6q08hkXFS1
Z9yBPxAFSWQitCkhMQVXHtlkH7wZQ+JHSCxhH/u5eu9GUKJJJOBsu1O+o24RKlNvSWvuD7ySYH39
jRg2btvARRlyzOqc878KA7IyR38kyidy7c+iZKsLUaLNQf6JqDKKsTs9wCsV4p5ET8oIS1o8NnTj
xRaaI+w05Acgy6O3rmaxF+xHHaHyPQx95l/kHLX8gUxTwLDIjzqt/Xtqu21GrHFH8VwhLPncoFT9
eXaDYfPnhjIyTfUIyUYREprrT7WiiIAyJEC9H+ae76ccjuavJffDRcuIjb8jjZF0kf3X7dgzYY/3
by7m9PTeysKkTsyi3uAUVmoNXbOf/Tc07eqSGgnSfErUKXkWZR6h2B7YiiYysrhtgd05Sr4qro/f
tPp3r2/e2UDGP1oy1O4ml2Ufqbpq36UJVrF7jaaTX1+i3J74Z1l8RNWDT8KxAiZm9aKBJQ9wgvX5
i/4kThzt9btbovnB9ahfhb0+bOESWqIZbBUSuLyhXx8g8+US/bV4BmRICdDSU/B0im2yiV+rNE2P
LzRqyZBeuoSXZXST58du9dP5/6mwoqSkX+UfOnhYUQ1ryW7COt7JMHuTeUfZOxtSz/fVQbF/jg/f
k2QwkJRK7f6+FnQ66YQhTfNEvicQhvbahDdwDai5FJ6v0Nq+ocN7f/QkB+sy5SJM3sDliFx1peAh
aKNPDdDlUJ+zgi2DGc+q/FcQG9H7kQcFsDTHj+dY0GRfl0jtjgDqnsUq55HlcFw1zlFLnwnC/sHr
gPuhfYWz7AwBGiyk9Rt3zP+lqm6Cmb0iUhIWFDlu5z+FeCj4rg98YRDU9i8BLE0//OWneJI2PCWa
j33QKEfdlTYdbqRH3CPHixVffyH0ltYGcwpBZSVKUBKkQ0knrLFQOaExJ3cIugVmyeCKJUh9sCvu
poxRIOBriB/ThGIu3wRaVFoNjAIpDwE4mTTdPLBoJR2etwc2UOrB5SWpgy3SpZMeae3HqCx7FO2p
iZnVzuDHKdBnRRBxcBLKzolXM3pQxyaDkw9pfVoid/8lbQdoxcDS7iak8xhiFFwjlxxPo9u1j6/u
rh0F3Cb9ieyk+Jbk0+1Hm9Ykgn52WMUbXxzqZbNTtvcD5EwEo4Gw7RvLlUrbm5OXHuRX4L8mpvLS
9MCgJBT1qLQuF8si3kicU76jy+0sEyylJ57O3FRtM+QNrKR2ttuSopUWQo/0vYrnNdcDEn39BwdK
Q0Zmg+j42Ksx2ROPqmTh8T6toZrBBqETfhBp4BiTBJ5z+VTjTZE6T07dTz16uB31jRluvrpPCLCt
R1wztAtgsRvuzgiRyMeRQezZtDv19wdOfh908tFkKud8ddWzWzBiPLcvTvySaUP/KllOU0CNdDcM
pZ0Vaps+oGRVoaqftsSM5RXJniGp4jFKBNr3oozZjnZW25BEhlpQt8+BTe8lBlaXvGYug2FnixK/
TfkvHmPfe86ay+s7n+dW/KQIhkNVc9Q4u84ZjmMDs5dk0Ry3Z4oWqqfLwTDkrGiignCK3fRjjDh4
jaiGe2exxOIu/G6J9DBjKDvh86HEhyXuqOdI5MI2vwfr7It2rzoWYBeW7Jw705++5qVcMMPdsunc
5gbVANcRrjh5K4HiV3QVy3t2Yoa7r8I6LF6ycqwUXF2RQPhyQiVS4CFcmoiqvU79aw22f29ExYaL
h8PIwZxU68r4QwiEZM5oDZ9XhXUwkgXdzZmvKN/+vSFp8o9svPkLlL1Gtd3rH08YTxghPwxKo7zi
oL/kF+Ywaw4piCBJtLnUlnT2wCuxjxq7O5Zpz1ctrwjSi0mj2PTlyxDh4TaJlEpTBnXjkhlZQpEd
zMu0yAC66PHOmKMcLjTv0UxmeaKNjCygwgUCJ/K/FWp1Ruc7cq3OC8a4Ip9ROi63Siq9EhG14XUc
seAMbLzQB8KufU88AUed1MnV7UAoz/tgq8fsD3iihYKSK0wcXKxihVznyI+UJK78S0fx5aW+Qxac
M5nSMOQK7dXiVOKrlqz5p8UzN6NIlTZV3LlyAEk0oTtwKf4YUUOl/pSQ4vmtKIM5DPheodxtl+L3
yVz7vuQf6368e2IS8CvbwTxzxb0LquxWD8C5NrYCA4tspp9IW9nDU4sGUet8r38NTToHvK7nobVF
HQU+8pB7aPomXrxWTmBChgzSnm4pQLy9K0QYXKl2cSyz2yAzzFYLHM0f6z/C/rbB68FE5ASoxECo
eNOnX5ysMtKUu3ko+2ozOl2DtH4soeihBcmXowjn0tUszWMy/47n0NI+KKFcURKZBtetUqeM/HTz
Hx+Robr7GRGgnXnlDb/5QwImg9uTAiP86Z6a4EjwEaoxxT6t2yJ8KY4EwkMYSjhyjdd0laVI28jy
JtDvjuWiiUzjHs+oir4Rjr7k+yIjLsN7JEMBdcEjwwzNAIWqHdnLyj951eRCEZIeUaUv+etfvTEZ
HLOeIyTTg+6T6+1CqSzdf0CvHf0xMi0tiM5uMnTh6iBS+LAbicTRxDRViGOd6hLwAB2tgpHqtptv
cZ/ntgf02zXV6FS+gNfippDO16aQtkN67nh6E2C3w8qdOXae6JIDsLqjuoOSoTTY5WsWE0C6D7Xd
OmW6+OK5Lj5zaVpJrw9aicccjYDv7LjH+5StxqimkobfhcGjKP5QGnWg6xZ0OakSHVAivy0DYhX2
dhdGA6GaxBlAcflaqgjr42PDiOvUN0Og1MXmOppIyMRS8S+DUxS09Uxtl+5oQ9Uxnj6OU/v0o9u6
3A/jj6NxwEv/LgbbRZHkKdEe05/Du0k+jZjXD8qw8DpnY2Iex/GiPr0drNNoItRda1RRcDL9BcTz
PUqVIvmX4z4NOHbnNjoNqhhcYgJ7knxGfuO4YXcuLlvZ0kEgbY9ZjG/vIvJXBaxjx6Cq54TrSTs9
csDO46R281Xe5jbnlmcSjrVMT7ITM2L1WJxKSY7emJs+VEa5ypD7L5T2jxw7mTJHc9dG6O2jw3XL
o6cGKo8ZS8j1YueQCLObAydgu9MVH+292f4G/X1keDnX/SBVv6PORrSdkI3qbwTGDXPkuO3bix1s
rxeovsdwr2a9p/yU+Y6vzXtDReIuLh6smj492VVkeEEx0XZDezrqXDkKWX3lkKvb5NUeL0WJ67rv
wRwpZkDBd6dXh6fHN9X4xSOa50Zkh92jGfSxEFgGFqgRHKf7Uhz5VNyoCBZy6+WZUxxXSOLOeRm8
CkQbsxE8gskmuq4+PXc8I9290CFt/CXDiMQtFq2VO1Oy1P8dUtjkYF7E8kBE+i2KjfQwcDfnJ8NQ
aF7ypmq94iO/oHoosbic4CW0vrj+sErp3Qx8ve4eklh2gJFYSg0a67K58I5oroOIHsOFO2Sq4Yio
b+BDSP/O7twC88GDQSk6iUgltrat1ctbwprfPsBgiGzxu5i1r3Dmu4z5URndM3h+HpxyMx7f+G+u
YhURNQfMGD0Fq2uxbm9xify06gw37Gz4aT31sX3erjkvWcjNYCNnfOR5tMR9Vg9yVKhbqWwbhj7g
exLfPwxXEz7FtaRvKCBhBwmE+iFrESb0wRGIH5rmrJiYs9sHh5YGjMHfB+gyT9zxcG/zhL7mKPym
jS4uwlXEtm6R8QbzEqAZ0QFf1J45pdbO9mBYUu0DmlTxmGxtYwtmZRGrq9COH9KTcrZNgjNR3uBw
QfaZJA4W+PJfPf15nmb9O+Km3FE128DT47dWnJU/27Fw1HZrMyEd7t4pnq455KNCSBrKqXdIiyQK
uHGWhMW8Swfy9CUJtiCrgHIBOidMgtS/Y5Bgojqw6NNBfnJHgQpcv/HdyVi123B5t9rbMlNBsx0r
DFGYhBuco4RhyaWujRwo9z1Da8aWPsarvJVQDdH4ze6+wHmnEQG/apgD3D0gF75TTYi06ruS+oZK
GxnUxXLygbTaGTaViLJa4odTALsFF+RaQ/z+y1L8Ndk9H5tEzASEAFvnv5UYwvGEIOU60ECdlAKO
rpIEoEGJASWyTlIN3uzOLD02bsCAJZsbTIkcnpGqRE6OvFY9EmwFbOPLG3iZgVs2TWAgHIPzBBZA
B8mX8WznoO1eRmMYu04j2VEd/4nMEN3SKK0D/13lkyJi/RZkUeJlbsDtjpYRyvDKYl6FF8DiqVfR
gA449T3QIfB99KOiMkQ7R1OXSjL4EZEI8niWvMDYyPvI7ZUvupk4d5vJYYFJy/bFXddbAux2X096
NIrhzK6RJuBgS07EjBlbaDSz3Lx1wv+yU1QBazyoyqpDSRszyjJnA7aY/wGXloljq2qoaZduYgGi
Pu6M7EI42aAI3014vG9uijviJMdf8T1gl/8Y5pgk2bJb8rqB2DzHq5Z2S/emdY9nSAJEs0YexitE
WcSRbuPi8au4UaWJr4NbCsqp+eQm66BbvoVGnPTO0KYplD6FG2Zpb1MPx+E9UNQx4lP00phuI66e
ySfCtJj1l2HYQ94RIEw06gB5CcjVdAnfh4qWgQB59r7ncBuchyoPQhMWfoXiMDdmuqFaQfqASSHC
M/zW4sdtZN4t9qzATdm2F9MFu8D5yZ1iBzaOjwtyBVKJJ8vwRunhWRYD3TBFuiO91pNZBVHBxMaV
hXnqmoG/YqdUDj9qzKiXqC4MbwXJG8uf4t3HlJZWzIB0+NbwLTpU9jg0Gm1ZF1cq+90PWy0VgYox
8fSqelqCt7We+Ny8+XssaqlUdvweZJSni9trmttJkfHW7VFjKHdbOVajAoKcq60Lars3TKNzxK5n
vb2qaQIyrzNpqlTfewhAeCrJtZLA17SjwTgQX40BwWmVLla/FclLS35osXfq8xPlaD4XAodKny9e
k7Ufmk66uaWkjVWQr0nzpHA2lriPVcPqf5REn2IiFPrKS53+Q3KwZwOWfQmkzj7M/ow6BbyRRFGs
QacdFVqik9+Pv3kE0v54ueY9uXR9YmWoQ3EjqJ3fCNloTxcMJxo9YkDBPAlTUG/j1nRdRlEVmJJv
9OeiWbFKMwOdD9QGdPoX7uuhV4b5dzF2gnsJIYOHLDYFo14MK7/RjCUdh+sWaC/VOAiikOY6ZtGT
Fypgy4ryqCLqsfXVcRh1kkpVyDQjJAIjDF4oYpBzkzysgwzI7rm/v0lo4Z/chcFh4YHhUj3/iXkQ
AOExGUlZGt3ACOszo+o4D3AFHM04lLdPBr0Gqv5KSiAqj5I+Qhu6ngUccBOpgApS+tu4GUusyb9O
/tGCYuvMPzpG4tNdt9iZoyY/o2IMFCOfCtDudTYSr1gEHm6/90KAIFytM7pnxvw2SpiQo7ziO9Uf
snvV+OYgFhhHaAe1yNT1mHMvAbI/GMcvsZAXjq8iawkHvdK9C+J9sKWNgvXr4N5Q6LBhLSrcYsu8
vyy0lLLmDWgUkmkNf+i1S2L9VQ/hCvoTSFKAb706BQSUlCVSVUrI8RgHygg0qAh8jHvFTe1p9U3y
5y4Qad/aOdKab2GvNXrGdvydqe/2TrLpb9x09aAMnyau9W4twOVJmWGPnH3jDm3DoschQZskN0yG
zGmAdZ2BIE8Uk81D+ziWUJzwPOCcSVLflr6UdcHlVJs9tc1C74CwIatX0pxYmJ4kak84dbS729xd
e0ABVF6MK9UyuStMSorLgY9zb0sC+W6qu2BnOsw+rPK2H90EWDqP+m9Dz57s3K5/iBM6KqwNkOGE
ifDpTOzfivBUnxBeG4R1Pfw4OfEIUwAATi1qm1axVj9L8KxHsvd+2TT6BZ/MDs6cEOXywk7OkYX7
rR8jgYjCCaXs3AAHe77TT5CbBDvsN3L1obRNKuV02fnWcVP5HrgTKV2kFWn1dYuo7oNkBDcA47bH
SDaNbLTzDRBQ0bP0ZiwLQPvOaYRA5PO+KfsUK4m6didouTo57eCYahmKgHhtHdEMUrtJJE696+ub
MLarC6R/w7663pVaxq2/873lD3Tr+8l124fweX7hvJ7fkjsrLHmmPckhBolN/U6yRGyOWL0v90ry
3UiFQD/3pefVyFpPoLf5NvEDXJhAaM1Gs/V/6GrNUa455ZGO8TAPKZUGnrA+qiGYFisB0GqJI+T2
w4Zr1nKsSckqfi0KOX+qP1LkFTsbTwsGTuqCYfbY+JNE646beQAaG//eDJoV46GCgNg8FxiXiKkp
xkO9rnZTfeOI5r/Cu2IVMaYZ+t0gFDDoG2wwA6I3aDddBHm18kgoX0c2JX1Fq8MRSFNJ5+w9NR/E
tMj9Jbfoqv3SwWiYdBIqr/bOsXdJxYpfeA/lKZX6hoGvjBp0e54HaUKqtruisYvhjwjAdLRHinDj
2J0JDwu4y05kdMY4g6hlLcR8P47m/D+KePqP7AlLGlNa1BzHUC8PhaG9Pr1/KYMHy7RgonlG6IIs
vPDt7+CdlJUdscThPaaazGwsOkBBykXoQ3C9sbb8cekZr/CovQChJSctrbWp4CWzxgmUMyxLiBBh
bJeT7AJDD30Hh5vF1bQh3YptyfJSY3kzTbAYsukv+Oi+C/1Q3YBapJKZXSgxEYNg17Nvp3j20Sli
erzdRC2bySqP7GQbjnKzKkmqvMuXfedk2bLtwV4wbec7irtCZEK2rceAVbeh9HW2EH+nO9wl5AEE
ugC3YDB0BJp4h3wkpVPSdMg53NKxhQ7iUBXHJtZ4eAuT5iN2Rf9VUh8smelZbWp9aswcT8k9uya4
camONuHgr2sJf4EWuFsnCKvcq4uyixw04DrN4Px8BSZqgR1VSfEs7o1bsy5K5mI2R3fnz9UURRTw
JNMN8Zt0UTDaOEQSWCzFl3Y0kL+viBaBsmADMhD+voWdP2aeUaWpxLM2dN34HZk+PRSHTlo3I3CQ
m4cDklW+g8W509J5f8CpCamQbM4ZdYwR692o7tNXpG9dA0mdTKdArNdtZpCvvAYX0v+r5L2YAL/i
wJD8gOMo6KAPAxdyn5wt5qM6fqC/xTJKAaaoJL78KDLJh67OLjBNlam2BifxDYPs7MRxXBE/ssFK
NSae7oIoiS2X2ZBQKM5SxO1Iz0tY3TkhISA3/ZZlODVqB8SkMD/usko8GFci+63BSbREdeVcu1Nm
wFONLF404tNxciwdgxn/Ty4ZAOTkPim0SYDpqqDf8WzyL5baWflSRr9JbCTcR4Qm2ipqUPzj4UWS
rNAo2fZuDjrrUy+AXlMSESle+nR3VFQZYUAUujvvXsNdAjjPT+zx5Td4RaUEDifhAtTzHeI55swa
qsacUbZclQn10QmDWdgBp/xIzAltHNpBhv0D81KVpPiHTAQ4h58jAKZKvmA+D3WOGDfwCGpURCXW
RiZJsOzrOOAjfxGAqHDrFi+tNTy3ZXrKjKj1HFMwX3jMud77ssiuLDXOKk4TK09SkxSw74wVlEfL
mh5/QbNwiFiuc6XegARjVz7XImUOvWNHEoM77OlbOpLGfRazGkhP7atEI1ea6ne1x55fkeuYO9od
4yGRBI6m2kmkVL/mkyKjhTSLYxOCHJcYLKyBmXXK7bkRyachtKFjPiHOyy2YXWRnBo8McrUmvGVm
9wGE6lfgTpoYM9PWYS2RXFrYZkthb0wam3s3OLtndatUu13bukHhzetJ0UBICUL8UHpVScggQ5vG
ZH8isxjDgHI1XgBU/GM6WPrBF04JHG5pKhe/mbzdM3pTUBGOEaxqt74KYqOv0GI0Hfd9CSO+u5UR
Zr2bdPabBpQZj8QE8F0t68AW/d6WEgrLJEt0VszFjl/UQKdMYJMMEXFCA1PeY3L3Ga1t9nKmTzu7
opwMJln9h4eUaSLz412kW3P4kpR3EkBgmOyMKFAdpfnotwz0LslwkLCJxjtItLJstbLRvWt3elOH
zDFhFxCqgaJSrr3gNnZc4HiRM/rms7ERiGF5WKuzkvXZAoXlHKaSAZ8ywmK2LC3cqenZTARXbvfw
+GDvfJHNP9xQcP3aQVB8Dnr3U+u7JrJ8Hi+pshWNhBt+p+DM17xdQ3DsqbNSlT8ufZ9xaKXr/4kg
Avm8Bx8XESeauqg2lc5A108ELmEF/g2lvRkNjtHJYR2VwV17m+01RgoqF2TO0//ea0R1gjeA99px
5BEhbAXxorfmdB2AIXHt4sSOBfoNP6LGo4C5RfwrIlrkjY90nHe3V/a6/yhVfAWjG0DaqQ8DXVGl
Mpo4A9u85Wo1avLxo1cRhaMNsHHFvxzEn5RksFO2WvYGcf/IvDAKjKEEngqkFiDUlHN+aCBE5760
Vak3rYhgiPCA+IGds8UKe7t244BO/fFEwLBZDOv7hCjozjAmwqKxkzrJq0Xtb+AlnoearAhn7w==
`protect end_protected
