`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gFPxhRrTYv6VaHVPGAiPVy2YZ6S6v5BzuhWPBzwrubAT6kReucnryQjohV6YcQAEW8yJvtBp1Ysr
C+Bb5OtwkQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZrUOXlzrvv6qQpYJjywdImSGK6eXCI+MVQlcEaIaqP1/0j88qHcz2caBn7ko88g8r0vYZDYOxV5n
bwj9ewbJDQQ9ap8inJ+mdTFTKMPo94XSVrTA1cg28DUpjvYCwKrTbA1ADYh7RUYFbkkhMydUo7LD
lH1Uea4TZeH7p9fvCAc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KbcSBrdjT+GWw7UD28rW1gOX3CWu2vBfC5H9w+FelX3uG1bnT8AS52Y+stg85peQ62PdcFUi3fwK
NXs462r/hLo1nXD5F7+p11ru4OTbASkxrndcH0xh437UXtMIGNy4kESqx3cwYEQPIPbRIRHzo9lQ
H9EeuRfgapMIwrwKfCXh5gP57kN6zZB6sonyIx1xDfWBlHzocSUfgxGgT8hjIANluSQYpSfuUlo+
dEI3dEYoep/bAM20bt7RM5pEkOJajAoAtlMCTYREM5sI9ThqVmwHm0PxWocsdrpPEQovhMXL8bOt
27757RGtc969a11Cl9CQkDFdiqII0115hijMGw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PdZa1nRU9Vl9CFvj4B3l+BUQbX3f5MtNMaAyCvHevFovH8IDhuKgsO//TZN/V6VMR5YKx88nRmJO
9ayU3n6NN6JGyQ3D58SFXa1a3OL55wVnztwe1sdhcybNUAinICFBWGz/HG3ewmeUDTJCH6F9JROD
zSKXdw3fVdzQHjJ8CBI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFmPg+ESJU/XzKxI7CxC31/2b9ui3jWsU5VwZ0xzon7uYu+V6+oXRkduShPEbf95d7/36KCCl42c
DIZ4bKmOA7sL2G1GDfX2uAXELrSU6RP0dLua5f4h4uJ51pxMoZ71Og0jK8qBTgKG5/XNcTiuzcSx
J7dExt5Zvipm6MezAEpMNhoncMZMfeEsTHfNvBWH6oe73a+ylanQijwvhLoY7BQzeOBhwqx8DnjM
9rOxboLIf08CAVrJMdT5yb+t4+XQyBrBTrAmlnTZ5Wd7nODE0b5llIj/BG+v00hD030OPT1HhKY8
8XcBy0JYRhwIxcQi6EWvXDTos47nlnr5S4eXhw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25312)
`protect data_block
WsmniEhGXJ3yqCpRdXxXvQXVHBCVfysWyVF3k8QSuZ6YigsK4kMR4qE5nf/mJeNtRJY2aLF2OBGd
0fMDjYvvmnhYSIUaXTPyRvdL5pNXUwg6NGqPeYORyTrr3FhUZFU2rJMC8x8+VNBXfryKjgSsYRo+
XprjSdC+U37oB5nie0tg1lL39ddWX86+q40fB/w7i+x+WeY5Vd0wNCNbfuQ1OgH+91jml+M/aTDI
b2JBVhMp46Sszd/3B4EMqjVPPBd2hpLzVOZ08ZJ6eqwGq1Tow7xRA7LbkkXoW0hCHX+/RDw5z8dl
Szo1kMNkEt9sxJ966h9AjCRgoLhU9qVGkznnDkFjegzXuEiPgdZ8d/uewNDvqEzg/232xukRxItI
n65fgbUUtksx79GpgyESxHnd8WCixLeemS6iwD7TP6Yg0Z/W6nM2TOtyoZYH7FUMOr5AATS3dOQS
t0zDGfhQNQ0b/VDvjushi69x4AqR5IOovXaCnlZT4P6SEGWwbLrJfib78o2kR0O0d1Ir288GdO6I
WHT2AQ/upAGsKqPrmwHFgo0d1gpL+rl7qKP9WmJnbnJS5H/CLHWvU23NWq7KXeMKAglP6lrYYa0S
3jfd6U5gVP0RAh47bnR5EbD12i1Zl09Psf8niFTs+s6w9fnmSY1pyd4QnEJEvSrv5ToC7e/2vIfz
XGgver81zQaIkh4Oq9g/rSsgPVG8ZoILBycqktG7k5uelbdLF/QXJJCXtV7WzIWH06DmpTYsqgk+
TqydCwFit3yHs/sKIcBTERNCljmPY5Pj78MlDfDT+G2gHtY4gHjdNDsU56C8ybaUsVW4d52xQvlb
ga/PBINepdk/FqxfQKehUJiqSJrVLgQAcNCWyImMZtmsgvBxW9EYthtNLYirz5N1zHczzYms2F05
2ll+vYkQz/zc7CqRh5bWnNZNfpfe8djAWNWwPUMYe23SBsm83eHZ9xtP48kB0yluo1ooXe3+teBF
ITaIgQ7qEk4XCpiV1vMM7Oy/MQdLSn6cZlOK2xkUCNSLgZ02ZM5BLwGNUZLZ3kyRlmo8mvSAu7Kx
8BjQZ98G7DfdXQXmkEI/U1t9Vx6pPRHUUrkEaqdaXt7scDc8BjwtK1jzcq/QRLycX7zy0OFZgqwV
jGjHUTNivoQEW9/aTkeQTWJeQtc01Lf8zg1FEdFcMU5E7NfKQfi+ntQ3QJI3OAtbSvZd+KUjxwhb
60Ax0EfSpdnyi+Nq10GL+463+Pn0TK2AqeACXZjCVAin+5h7ztt9cnlWciMwddbn1ofKCQ4+D/m1
CrsaOWN231gmbMeCMEZ1u0WqGKmsN8dlLh+PbO8xkr/W5kzP7nJqnTpiIW7cPEQCu+YMIyS1bi90
hGk0qLuBpQS/AcRgMAhCPAl1e8Q81U/R6VjnyyCkizoe+t0Vhgl/WphwjEvgIYrMgzj2MkNvtw+9
jImfttRrdEDOtPUpXfiOwg5oGMGFVP4mejgmCNVMe+LERtiOwSxx/DlDl+e70xrmVdowfKP96xGX
mIXshS8xm79r/QTtvy9Iv5j0+ZNKBnmauqt776iapWbJgYTvjOwlDky0gBrujvIb9WB9hIYC8Ttv
mNnFGZ6osA8F61S4Hjd6GFgQpMTmWPk+olH8zPAet9nKTW+IvZ3xu8EDivYifEco19Xpq78ZndxK
2OgxDhTA+feKCM7fCS8Lrb1dAhhiL98CllJIiwOplrmowvdwU+FWIMd/O39vvYaFMhbm2lo+wRqY
IjKFvehWImIjIbc4QU8nvytW4UTUnsYgtiSk5AnGS08RwIMO486qBAF3qcTBH68QFnZYjfhKOKOi
4irERycfARU8D0Tyl9cHm/TdUMXVGuN0gUEVfSQYPp4e41Y4t2mR3MOawyJkSoGmCMaCwSZqs+Oh
p+SS47uy00aRgr4tk86HJME9SZKHKwZCvkTZWYFXwCsbofMUd/zTLf1++2u3ffbkGTlQ06TbUVhc
kxpMJVvSb5OIOqg+bD/zMBJpmur8rF+ZkdNlxyUjdRG/Hlt+YhCQiyPXErVgtJyDNkYd2iZY5HAZ
w0zRRPUt0QwFvR1UfYwpujNwCWXi6rYLBpNE8sU+HmXZNuXD+2suDPTx60aiCVj3xzrx72wxS1RY
zzWfsWotWcGgoey8ta+DA7fJm8GKsYeAUtZsoWnzidDW0nU62vJCZyLNMB9v4kBRwce8Tyr4/KeC
abEhe+E1+k0jMZg0Y7NHXXRtQC0LRL3a+OFy4GhyYhk5Gp3GnDAlgJK3/GO50uhd9rnRIrx2SnSe
M9GFXieoo8anJJ/4+mvYFDqIHl2g0nNxGTHp6HchRd0cOuwoqyHko7Yx6OIt5zDz01Aq7QP/HWfF
xXtj0h2K7CDpnDQJlsqgf4fJCvETryAyvczhfulff1RuqwQkPDEvvxbDvowIG9nfRLcENw4a1/cg
Ho2iSwAWWEDuPsPcCxOwTqyED7igMNUisLl5zG8DCxcKcX5H4EpAuqgrl83KeZtumPn0ULZSYlxP
xsrNiQkl84LF+QSn7WOIEgkMDdz6cTksYwbhOJdnkSJaxbgoYLdpad+6VB2iAGHUcrTWH1/R4tIk
bIXJjxyUFjGXxlSWW7KCNRirWpimrxQvD/2nEB9s92mku/Pf60jfWrAex5tHBeFpjnvDGEnimedC
sNp6mbBn/zXjUuDOL6Srm2GCn92ffojj74jqTbYDX36n1lrdxUimFXWMdE5653qlMQkZUfbKyEyt
A2g9twAKyRNdSO9A7L6qnzPUMCTGRuaah5KOBkK5snoxd8E7wlLtdi5KubRTKIX2mt1cjFzbCWLK
0Q+QalLqZSOe2AaH1Y5V1drTbSFFdK9oxBoS/asXC9JE2h1bJ7RhvJY1lJxjLpgubPUhaAdxR2l/
V5kM8Rf1akBlM4drKfWdiwIkR73OOfUL/6atdvpbV6wtydRzOiX8MUOhnEyNMCFdoeB2k4WFan3i
O9jZ8US9u5mcNr/ZAGl+NL0WHjrvRWtnQHkSEOm3zvXDlvMzcJ9SUBtG1SmT2mHzz6PINjWlqix1
yoJVcbVRSs91jeAz7JJo3LMZpa3zzvCB/kvuFk74Aqoce3P8MbIyXaefmrXwm3XPaOCSE6xMxIkb
8bKXiWCkAqHVil4F2wF22qUR/yCwCQKaPQFUS4LsuTggcmczGlKN3x4YpYgDkLjDtTRS/D0AOWa2
KAn+NRzi0SyLXSkBRZogn0bHluTp/rDPsLxg/gjrFrY112AXtydv863yhoEVR2G0c7aH9FWVuMWn
vvLSQSWTMLMuiNRx824OVu02B+QrZndy/9ol9zlL+DXJLm2Zb14b6GaS6Zkgniu1znsLaX2rnfF0
Wug0/GxpT3YAyBJvr2jlPQPIRItJgdhgUPfArKHT9+0+Fo3/1qruE+m0QZ98hybsN5lXfOoCOEQO
fY5a0g+Nws8mAT2giJ+gwwdiFXyPqrNUw3hevbd+dXss3mIl965bpILKHDISl/4XCmM8cCJoymgf
U10A+xTkJhAX5KVbNp41Ur0LVWarE3RqX12zRc9yHZus6hjvzmZTpgXerQe1SboHjkZhpszu87qz
mr65GKNS4UJUxNZYdSEH+jhTGByASgd7jTUpEPXyYbqi0dvP6iCkUtL3PBrHF/z+MEG/YfM/yqe3
cFwDpy/ZgLEKPi3DvmNSThLWuZJ3iYc3bbzqR4pohVoA5z/1+/+AuxQfQzoK00p2RhgZosgdN2GS
hvh9yZIYk6ETEUXxILCqOn2iintLuNpGrbVIx2gTVq6xxPicZND0pSV4lnYv1zEPSZIhWDsCV8DJ
f5TdHfez0UPAme73DmNsV+dglM5vrClLXl78K/dzcAsK4o8wkeyNqXPbdBIOTNupr99T2ml+NRt+
4aHc3+WgpTeVfTA99gI+r7/dj5RoVHqDq7/zqfyUWdg2fPKkpjfMyXj+S7Qd2h119gOwwBHnxMR/
vPouSWHM+WQygi1ldHGRh19dZdGB3fKGyGBOgYMVJa3/Amc6FjclaBgfgQSe1u2EJTpz/KJKFUCo
91SQbo/EW5k6PZxwe4qe6YLweFZaIUNRj86B7rvc0oXXYJv+tHJrqNnHwA3f0toAHPHvZAEIzp9x
2sfhqa7Npz22nQvFZTvKodgCvUemlLq31lao87BfpVHxojkfx3UFWDeG2Sq/31DihE+PTfZAzTbZ
RZFMOI7P9xoEAiW9KfDspx4eh06W8gy1/S+oElBncQjB2cpj4gjFiX/63RdmxT919z5V+2AKvqTH
q+YgvduijqRngSDx+wXxCXl4U248RRFZy6Q+o9zbr7yfLI/Mr8b0nMpRuRovdvfwsANcrTpH024P
lZ6Fib3d87U3YitGVT/cZNHeEq47pa8CcxClScuoYDrpEf4+Hhz7/yPT+8sITTZBu//OKDZ21wVi
jQy8Mjqmo73Oh8QKOdJyzDhCKBg9igxSPOz1ccrKsS43VQNonxxOpwAhTlTx57M/SyepmrEIQ0X1
edsox2aRW8hZOIyqHLCxVuz10hjTPrihNSS+i7KwQc9VIa0Q7wLOo80maM34oqa9ZW0x2BZXO5sX
uNgfU3N+46Tq40nuieaHExN9OwsqDL2pwAWYM91J7R6BLdD8mtuw8pH3C0mnhl1+X4Q+U+skK7G+
4ecErcIf/+BmSieepRwQQzjYaZIvy02gyctzhM7M8j4J+I3XJbcPorXwyfIjKD81sknETVH9Tpby
ADe0tXAzBmKICzwuJXIylVrH16Rmv3YWaix6Ple45l9m/xOjhvPK9nElR5B66LoIP7hbAC0Ghinn
KqAjMjh3WZdPnDaHhzm42wYBecWWRrARTmEhNcXtH0HWsL7gkeHWfxGhA4Ty4DUJk4Hz7nX9+14V
dGyrlw05mITynLKNgby47eylEjyiYnux9Y1vktSwFDpii9xNCMsw8RDK2YoNI+zbZlTzmzgESv7U
T2tfWanoQm5ehNSq7JkOOm9n163Ti3KgTkXYkJBXGdbH+6nu5T2NYcasEeRdNpOTthlBKo5uWTSy
+1X1sK5g9BVMl9mu4kiZS4UlhJzWk2oFL50oYstVWKWKBZ1wkeXP6ErgqLjFW6hyJIcGDrSqV/0w
klF22YgeiwaAcOIDV/yePObu8U2wAN25NbNKlOYBvlF6YbK8dz4KZpFgLs77bNm4eRktWp2GP3KH
XoH3TpxFl/5eeJ+fsuB/TThb1Kv83I2Pql/xpUrX+oUa+GFeU3i2HFpMBu7RbsKNiVmsyzxGgGMa
cpD3zQL0Jm7Sers26h/gp+JocJz6sI7lQxQkiLUUjz3m22jkFjF8pKswDrNNMrjepSmDv6Dl+kaP
H4bKpILkHL6gFoD1u21bmIHPSbdC7LcMoUQzqc+vODBqyYlHkWf0fdLLi78TN1WIWSk/4EnEzBkb
4FLnaFBsUjw7NwB40JQnQ2v0IidHG8dpdizgtuAlfdjzDTNmUF2/NqhKy4yFFPhAVJ7MOJxHZiyG
a+NaqXuelN/Vc25TFQMeweR9YyZU/ZZcG0NtWfd2MntCFvPPqZGya/GuoJKdNVDPqvxpscbTZGGz
y4OLJ5DcTAg/TFj3N0+/sJpmJ9B7zLcltxmUM+NFdPgxapPf9MdFKAh4a2VS6sYxUK8KIHsLTxZq
Xc2ZUBsI+dmds86OuScoSpDUc4QRQiwv0KLKn7BHmIcXo8ixtgIO8da37daFJM4Q+egbKUfJLiYw
KaUWKifWqxOUkIQCOrUK2yr8SaFk+N4WT4MCDN9ay0AtzAQw4NQ7cdUxHTB3u2EgcEPGCeZqe93H
wZrjkdGHMUymDk2jvMJPiC8DvP3Tm0i7oWBv8H/eJe1pxxke13MgtZA2AJWdJ1sqBvZrglBITjzm
VP9FRW24cHDFCzCVRG8wWkIVTfvNO8peJTxl2L1IgpwTbzxtKdQnAd33p2U6yMQV+DJyclkL34zK
TntzgzZkg9xqTne13W5uYwuYwXNxzKMwu6MhsFZRN3zl/whXPVe850aRuVfqe1nidDYr8hShRz8w
ao4I/Kx4au49IY7UbQPnIpMv1tVpO4mAGC6uSE1p+/sQWZgKFjW59jR0GFiRAqdy9uVDCvQ2UDxK
HYLsYjqaTZ6dbIt8W5jcIhKf0HkI7VyQsy4AuxvjYJILli2uc5QfpnirJSASybH0pAQqWBfBAnBn
k8KmtYM5kRI7mvHwe7yAXJw/Yy1cpZxXU7T0pHY3VkzZZUcqCe8AlAEw6/6PO7a86KNxH+eh86Ro
37WF8nauffHltlTOZh3PG1Ls8tqAlUgCrbb3ruzRxiVeppyoUwuDNhNleFUpSi4SagdzzgiDDCIy
kMDrOLbHk6jkXZz6tNHlHDyt4bup3Z5LiUSdDYXdDDxZ0b3ZXI4jHdH3lVWj+eEyKNHGI/S68xdB
UEFUuiMdfdvSBVE+lgvi/88fp3N1okU9M1z/0ruuQFYJXfhMHHYwuphrhflgaCuDKDh44ICX6/Ay
ISvkgm9tZ+/TfQD9qmIJhBfeoBTST3UNPDvkhP0zT6PdYJ86zVeYCln6qlKKSdJ1lC2oarqCEIa/
Ow1F0hwJ60iwntkwlx+q0fzbQyXvEBj/FclRJNowB0LE0rnLFAxkbPBwh6RXgMkqAY5drBU+8o2s
FDkkcwclOLRVCzo4kBXWZa1+4nmLiKCuGCl2rrEqnmph/MZLpuvcyax/KwaO4Gvytt/v5oxAy0XD
Y2KIirgAItFEZzuMJguPEb/+Ln6TbnPgvdK+ZEANwwNWwX6vPyNi7dnRPSTmpn3qEpOV7a3hh8vD
0DugwIaV0IXg3lUijc2xyvdTNoPv5Few/R/7uVCgA2Et8Icy4g0MyESnhwHPfMtyVai3UpI2ANNv
CZt1rQtowzaF1tOPbg8BHedllF66MaDY08Wax69IAL9TGXSoPOJ+bO6+1M6m1SolV0OXf/PNAigy
Tj7ENXKnc1aOJ5hQyPibn0+AwoeRyVRExdhfnp1dZBI2kUkIRMXt9wU0BprVlkAJLyjmtFv3z10R
k87zU/G4B7en2qyw47j9SMt0OFT/hV+yvIH94o5+ljHv8gNSA5lQTSszaCGFDqL80qoTdUWDlQ+k
7yNX9xla461k0XXRSNNpO8xYDOhOh3wHY/jochoHkWzMzTWDI2UQQSSzbSPXwRhdX+uoWdB6VPLf
d27bBMdFumMm51ftKz9XZ472gYsjnBGgDFwsIX7odEWmft1uBEIx2pKl6dcfhY825CYTRo0uKkVs
DiawfF8tmUzw/hAFbvXNEJj/lYn4XiVKLe7KE1dVXqs98xunFnzXZ8I9FyGzeTZMcDDqgElP9DPp
lrr0PxDWg/LqVaavYVecA0WmGHyjDUSY7bVsuAw8F1y1ueBI53+Atr48Nb1Ehv8VHKjVaSwRrCtJ
xkdOO6MlqyhWzNBKKV46LzMq3upIV2Av8r9g+BqGapvLl0F043LG7FPW3mWMjGXq57nOFH7A5SRL
Wa5F4eVVqQu42f3AXmfZgCw8tTiLrBOFY/OjwkIOX3+UVDjx8dZgu0C/pOx4cpbzeWXavjJpSVNL
ZtXrTzkvhqlE43nyCgIW9QhS5DFYtUyDfijJdREN3/WFc8POZkxOIZmApmdQBs39rXx2wqTaeOKk
a9AECNfTU9dObLWdcLclq0VE/nSNK9/jO6AsUgN5e/bAualV5V8wfgCRssYahDXATatRGqLsud18
RPmxIMREpnPdqClJlmw+pk6S+vDLb+2U7L1FxxVOvonp0QspcO4Il9SSJqWOkwYvk1e8Dp3bfNcC
0xeKdj/H1twoeHWdIcDFM9uE/iIDWHQ9kdHunx3P1UD85bIsVaAE+mbBe18t7n8ztSSUKdPnLPtG
OBho1F7hCby9fw/RkgObAce2DGUspuDy+JTFh8AzKwnYDurMqA74quSTRh3M12rlSbK1ZkGfp9cH
o43xO/8XbhDHo6hEB2hctkB1SoBMHMt5XrzdKgx6t2gVgqrx03UL2BO5oPMLkbBYEOuXm8snFJ9i
I/Nlz9Ceelan8cEIsoRJV0ppKI2G5pwBlwKoRdzpW5k5yBJ7gEhpwkRqqwfZMcFtV9rHfq8v87b5
vBMXeZHdArvCWldE31ZRFvlHLvsATJ8QSUn4BjoMP+KpYh5JmlgiTW+PXrol0z/7UqshVNDaHcw1
z1R5MkCLL1gpgtOSoyDd2yFjT4DLVS2/SeZVDoL/4p8ZUZI8JpzJG6M57B9hsVymEmobT50yDmVY
yszFrY8EyDlIHB15SDWhDnLfw9AtWVY89p9P8X8SkJmmyeDybSWUx5t1A557HtzqUUlqtgo2q24h
kZSCOyNnb0dFVn49eHEwhdeVb9MM+hsVFbVUg9p/otr72xJ1Ewtbm+ubKL0bJch+zK0VAHdatZTB
F6SXuRtcgswf0IVsgB8pSgbb0Jn2qGdRYyb8GUa28bEriE7Q6gndOo8PcSQ+4IT3EMx54xhWhTfV
ebHKpuCgxxeRggLVijnuoSlR50sJ0G9pPYPohtF+148ZiyUOwhdeksc5evatIvfdIyntp29K3Q/g
HiHKwEFo3KKvFXAJkWsVFcaN7FWvDp53xInK28Ng4bMKyCodbt2mmbywQTspvR+N11mZrOmGpA3d
N6lFiNzVed6CuLONd2rrQH/+1D/r53gewJ+tqUHB2PGWebtEZZ5Z5rlRIqjOPQ1VaknT6nqEYAyz
JmI/+bud025e1s4yto9XLa/fYYfWJO91kQinFRlOKzgmXz+JDcmT0Uic3n1LXEWfQeBee+qisN08
eJAyWw3Y7B9NJC7pdyKorcdsuGrAdNRGnzIgJ1g2UtdmaiQXT5gPakUnzTEMCKWYA4HbKMvDWGK2
o9DawqP0kA0eBGSkeHguAvp6G1HITcFNau0SctCQSAH8Y9o8ufFlzxc/WreQvHprUziCrmp+E45n
WLhx8Nmj6pevBrYRll1IlJouuxZYLu36VauS7HybiUckWTj8NDS7pOGaeT9k8tMsF3UGUxENls6a
L8cSPXJFmxZRHrr+zAtD/U9Bi6t47hN94ycerguxrBRJNRCicAZ5++MUdo3SyyUYndiEBlCWtGuD
7B9LujMXsPwhAVLf5jgxRMGLv9SCXVJgRyGSPp2xqk5WsxRXS45KbMmxmcopHbSw90kV1XcSeQDq
MCeiWLkviAgElxRKS8ZNTeHODjWp2hnyfTsgSs4p5jH36kO4gbcFAa2vSh6yGQTexUnkpQbPG0JR
lApjNjuIMgico59A9A4nIsx0NFK29loWSHyD7UTa7FrCyuyGhmIXxrgNFQSbq3cN9l4ycWhc1loA
W5HY4B58tKpDCpbiK262dyOdVXb2D79MpiSAiSXaVKk6fm5mOdZ/SJlAKI3erLuG6IQv8hehOGtm
Ad+59zYrlUZzqs7CPld67exJPoUSO2W0PwM1RcZ2SGGjbBtr6KdDiIOIfmKvLAmer6JuG1lYTUpw
IOKDWKpvpm+JwkBT7mQE+Kew36n/MTamxy3fWP6D1/w11HtQys2kRWVpNeYhz+JlCsWbRVxvYIFn
xC4l49i/I1HwDYHkF5lU8LHX9LrComDajJwWpq1O0hqUHJc7BV5MKUwZpfmr4VWz+ZgROuhWbqQE
UyW6I7PNIFS5r8NDihBa0Uv3d//nwp8Pul53LUtGYGhJn6LZjRy4N5jsDatumoA3iuIuC/3fzK8j
TeMfbFgFEFymTXyearmM6zhZBFEGXm8dmotPtqI+O6GLfY7opE0tjUGDyMlfc7LX7suDTZbHwQDl
Y8I7gxaqjeFjTR63NVMWIroGFSDeTT1vherLXwUqUBTPvFiMdNPVWee12XWPYOSZ33G8aIy3jpd1
XJVZH/mGOSs1b4pgNntb6DSp0HSYgwdNlmUrGYyo844Qmhv9cfN3GLlobyE58ucnJXomhHHDsLkK
tnU3cTouqkeoCozJ3Xa29M6OT68e1PzuOvu6VdaLyVRcCs5u/ZfvXWt5QZ+ThY/B4CNMVWuX2yH5
TV2n2x8sMmSiR+lo8SSQS8VblyPl8zRGRNfa7AdicrdIPed2CN7+04yjmRSs3OOMii07fRkDLYrZ
N7XUpwvvrUYTeG2vUw4y/U1qEjFjTv4CZwGMd7OtgNfrgOQTSrbD0zBBVFfBLnH4AvnROBfYayeA
+bsn6wi+ppj5vFPmw3wzq2HEXHRCI0S1ihZREyp/68W7yAQj1XkYgQF2ka/5VS9feSC9VyFGMUXA
0AZ+lfgZ6H7OXpwxwMb7ecTiYfaOYWfLbq2oKWhq/Z/zzV93tkaxkDslfDEJjBZD/Qvr1Gud5riD
XxYYlj1bSOJ71F2G98CziHoqkSYqW6p/G1VNNjttdKRzkt68Hmap7SlTuRxScIcmBMV6lEovV3UD
WxoVD+pCs8nOOim7ADoP7CUSGmkfZwbUuUuZmhXNszW6THFmkyGqScw/F/Gu8q+Ji30vw1nVNhQR
lY9lb4RWAiy0rC+DXLqJjSVxRqqFIiV/Z4sd2WWmq71Ygs3lcH2pBGw8QNTAJoPIlJKs0vvks5xO
cO3Q91WPYCmbrafipNWwXi2frMrROO2tqJO64yyf+DK4bJdNzVjnHz3qXMaQ2r9eUaZfgbr1bqLv
4iCUxzXA7DBjEz9FbokSlHXhfIYdPAG9x19twXy1UpVBLiW0LH/i9WgoCmbf7udqTzfmjjMPxKsH
RyloFa5qDBq676RtttDJxYP2jWdmylBsl62aaf/R18yfsUzlan4nZo+cQUyksNgAlAwsWxHAbcj7
wJlELr9mvXpNvBucCjRiAPVRjFPIiReztuTRD7wB4aa9TbWDnZ4nF/00OYWP78lgY1Zz+0gXYRyF
Lm+LQ0MPxkb04ZsyJnY4d+j8Z7hpQFdwxQnCptYbB/7MmBvRt/Fe2GGGZCLPbTAqK4ROjQiVhm9m
OSBEdgRL4vqDmPx5/T14w6BwCbSkUNu1vJCoUK/6d2MdXDU6I7IjZgy9s17b91i3XLL047qUArVX
lqrIw4BlvDLfjdQK7aXcHkMSj2iUiNO6g5vROWy+jmjMlFA0aL+Y/Hqgo8+nLbyPQKd7NmvQsv+u
xxriBF1uW00IcUGh4ESTlH5v5aahOsC7DO5odmeiZ2KXjg2ml+8owbo36FGCS+nF7wek8/f+Z8MZ
XkB77GpMTB1irRQcFVJ7Kbw25k11WiOS/MX2U5km+VHxCqu4FNsX4Vm1ABcu795WwWHFtGFvWYE5
WF4CA3E5aiwfHbPkX3fPix/tvGGJp/pJl+UCev66akqDyAm/+6vKm/owUCmB8nipTcjOd8m3135/
jLEIDSf3hLe5Wn0PUMI1jfSG6KwuDszbjq6ZkdoFuHlfywzuLP6T8WG9DmKsKUkox+0tO32ujCps
rR7V7g1m1exi5yGSf2pP7aVm2plCtf+i3lFpWzNsyJR295wvCgp3fjumTprgXfX+ybSTmCe2JB4L
wRggydVeuIW04FLdSv9GtaVJPAeF17do/cgEPfvWKeV5YUvfoYrX5KNBn8PkFBvCQkoVxsGyp+jI
ygg3gn0zUbRMbfkPDBDkur7prMV31G/+ijMrcIgwf0R7c3diOEzdXZWhtuHcnBQWxRgscGjc9PG8
ICmuIBpoJs+SB0t1+4qS+6rHcOSLisSujir7aLihJxXcnUA3FFp+uh7tdiXNJT/MTX1XSA+hC3EZ
yq1+5/sJxT3YikgvUahE03zMsDWp0atI6DWJKEDaIs/kKoP77mf0g+s0gh1XmMxDHtmBohgbbfWm
j6j/An7tSutTr0AT7bUBXVr20Nmqr/40TK1AZZ2h584wMYMCGU4F7YCdmv22liivv9EQ/tqYQ5P1
vFwWykV19cTVdIsTlyAN30kYTyT/f1xbbKcnuWDI6AIWafJUuECWbOf+C0dG0HRmC2zopqjBb8eu
Y7adYmQjnBevDOkfR92A4QGLSQg7/fYAhUIwu+/Fat38tk3uqnuLWndC6keTRv/vzxTLIBWc6yco
hW4lFqCsoLC5IGdXwlI3qTnjDAZtWzeV28zT95twJavJs3adtnGI145VfSr3k5IATO47E/Ce/HqH
FxEuZDGmU9WHOHCGHI6fiC6sy/ys2Zyfvb5dK6qEPIsU8cbWSU+37zGCwqFDG/82krx6toApiKgi
oKZ1L+ixCOQaxgebjjzhVkNTkbauksKSx67U0TP35cQFMEJ8B8nCjnpFjIgjPTmj9KD0NzjriqVU
2CLHjxUyAUz4objBeFROZZa/1I+CtkAGM/r3aYkb0tsAFBh6ELZslF5O+0YVC+R1/Wgk5M+ZJh+R
V1DzjO1m+WDz9Uqb3nZPNFXxx9Q57tbdwj34L1RHNrU6jgLYMGggvKArsaNfrFXnICXM6K+Fe1y+
6fjZKOVtLz0oui9+ZK+g5pyN8McGLy3MLN58c7zLUlwKvg3h047MR6FDd9b8rAaAVQNLNSCPaRHy
LgwbvHoBd3H5lWBcImSbyPrBoF9s8Q1V7jd+MiJgb/t7K8+uTXlBNdwPBz3zLRDdjxC0yEzZ8DVO
Xp3R6hG/TAIJOtlOHyKKiFBtcYiVIbYg6OF9tCUqF3LJDCAqzuasUCpKQIKt01rBm7uz2U9Pfe/T
5q/ftY/GhG0zccfk0nOphtD6s3x5TkhK/MEpGkEONWBWM88lveV7VJAKtiNrR5J47hk86ZSPZIx8
ZCczDXEpaI2gHuI+54j99tsRU4Mp51LT8q0+NLAgJP/0LB7dsJSEfoXVIRGg3UXxs8RocHQHtEsa
evzrT9lgjTsPJzghBYl2qBMwt7w8Xs4LTE2xxAP16x+L07bdVxLKqUeOKNYeyAA03ghqZ5yct396
6ghSX+W5mKA9B9PiU/3VNNxECB04WJUW3vv4KAXAaOEJ/GU+PFIs7GKzzFoqcosdqpxcY8phGB35
SzOCTpcdNKqdhWCrxTm0y5hd5Kffe6Jw6N8tkhBWUTv4renW+BQui9OYkeaS/AI021XlyOjnFmAs
eszlpo9MIdvPXYnI9yFUmb6h8WI+MuRrqgldMAssc8ypjjyI1ZsoP3ozs/aGpSO3mWPph08KmL+7
SRonCvQZ6yeJdprHZEZX0lGV8a+zsY/65BFBEJHY6PHLSTw4yQzDE7JJ9W1E4icLkdFtU1ua5lxp
Pif9CpYTAURwG57XqgjTiTlFr4T9DRBIR7MyFo7oF+fqJSInPve2QbDHA7pCutHJ5BmWSj4AklVV
AZ7kphSzdH0YlZOygKWbjvduagwlv6vrAdrzvmUjxEfQ7UqPxZJ9QkV54yjznQYxgmrqmi789G3i
jdpU+JwKdt4deE3yuBfTUXE4sOyQs6f57Ux88amYncIhGMSz/jkOtV8nv7my109RyQ8z6C6oKufl
afDYqwOJMrVNGen+snSpieKzXgIEjFf6Ezc5XduyXOBOSaLqpgAgVUjNQ3DXYJuRvwmdSfboyfWO
NA4Nhu4jMc9eX+XU1r7JhBqFG2PtgYYq8Re7gSzsFpk3HkbonRUbuqsenn3PLirgRLuGGWD0vPf1
IlXY/QTvC6krcSvcRypw9qtv4+bHjyPGJx6tUZOuFs7yiW0MgMKDUWSpZfyu3Zy62CafG7abSl6y
+PTla+eGuHXfbmrez5QT1t+rgikqUFVLcXp9VdI3/FXp/kIqFP+RaLy6OCmUuo7ErtN5wJQ7jDpn
tYB6m9LGuA4bbfXabXtiKsCYzrKGwu2eyd7wRkF0QcMP7qTqHv/kUaRw/ToNBzUm/sqb2lUpwS5F
k3T021KCgCH2N+KmjktTR5M+FKHYlePoF8a3kzgDo1IX3zr9SwmEllSBvinoDG1LsGd25yXanG+E
vCeHUf+GTerebIRjzdjMyRyke+JknOJ2HAVmLPJmJsZaT7+ApfyDgM2ovdbtpiHv5rndCCg+DnDm
1+HUFMrt/Nq/QNeJjerp1bUL+Wn2lvIZyyM6ovZpWchWFpZ5tnjQosWYp7cIz7HuWwOQP5RNhGni
3cc9BxolSa2HVjHCCOBS8g50jdOpSpscZXg1/IpcJDZi7QUvTUY9R9rXxrHHDYBzxzGOzD4dHLT9
Fc6jxUTl30W+erlD7CG3CswwRlNw0vU2G2VX0AYZWDOo7W+vt/mUbXcMSPDkC3ZwiV0xBFIP8U3l
3xlVh7yM0R6ba+7w+lxPSKpMcR7yixyBVxYg68ckDbGn4naNjAnCEEnm4bZHf3+/5EbPFNYUv8C1
78Bx8ru8SVdPiCoOzp7lZjHhzRz9t3c8g34qKk7qnj20Hkufgwdsl6uFgm6UTq6Ee0eUBOZIJlrM
l2YlzKVBcO/l4LW7oA759Uex63Dpbt6caPMGKKoi6rLa73HBH7ctR50135Oh14XB0WVuBJcU2/Xs
vOxsdHI+AbrsnqC/aaiQjsC5Qp3nBdF8skOtKI1RCQzSgDb+8Y7F5LUesFkbxhKh+cTNnkz0eIHq
2wkZC/GZIHbtseUP5sirzCHJ5a86ng5hnGGpV//vSz7+4NLz03QD8gDbTwoM6Gy6DVh5xyio02QD
ZXmbW11RGgepZbJZYGqB2ywsHKw2tQVRag7ZXO9Za2NyLdcMGnOCE5uIKppJErFj80hnu/uzMhKe
PC7dZ2I/8AswafdEMNsuPM+4R9n3FVkrW2MW2ky+PR3s0KBwiqYRq+gLCDZTwicRiM3cPGY1nedw
qDIqyXRDMfaDqQkFXc7wPOg7j2MMR7bsiT+mgutvam4Gd7KfggJNUTWlaVgjw3dkmEyEjlsAnrOa
wHr2ZgStWUYciKWQc5IhxJpU9SFDOYA36WyBjV1qOPhzmBZ8N6lH01BAUnsXHFGLo1RdW/cP+2xU
w0GeihIlZlSxS2LW2AsZPrTaslMSZ21324pbaaybqJqiV8ddP66hT0Hb/vjz/hHhfaIiRz1s8tvo
2Nqb0aL0wENCjcoGC9RRGj17To+NPvVWcHlTvhQLHhpmE/3sbqNQRAHqS1tQ4lDtVqhTbRb31pLd
gxU8s9A/qBVP5t2vqnGpwysRhmJ5LA8kOdywPIBGKrhC/UBEWE/eiEPXZEzdRsxrWccrxOVHid3c
IImQ+9gskK00B3Y/7U2gPAE0KQototD6IlBRAmuwjGvjoKwxv9pZkhysWn8RE8CB/jcu2fxsPBfD
0UueXpbRP6kxlfVwZ1Z0HHIaWZpPbTI+vKOF0os8F6dW2/tWs7paNtt1A7c4V8w/Wi6GimsAKxXR
kJG6CMESRZfAlnrhfiOGohJjIfuO7s0XBjMI4CHJZkoz2C7Z4drwy+6YSzC9z3++DZq9fIOervXs
5UJD/cTmdAi2QWAF3zu4m2hR1OO/H88An4+whQrK/v+01NSoszhcI8MLcwczMUlFXmhtPNlBgi72
3YI2fjP0sy/OpLd5vj8FDQmeM+11FtzaexeGQW2oG8UyHLa+PvlbCtvFdC9VIoJ5yNbprc8BWhLa
/y96/b9Qy8Uzv3fK594hcaH8zM/I2+p3JVQIq0t3aBeXk3IS/czxTcZQ/FwI5IbkE7RYHfwyBqbR
pAuKhfakq7XU3g4TFFuAqRquUEnQy4qbjIakP1AGWKqCSi6lFFHn/UF6sUPmyRNUGTbTelWu/8g0
US9L/auJ7PPqEATbrVOSf/ZHrzYndl8YulfyTQ7cLSakVxoFz4AkBuI9o/RukVKwqovNaJQMWd8c
fVHlSxp+CGmMbE6tD1SnYS3DSFo/OqX9Nnv3Nh7mINeAk2effMXcLb5Uq3+xE7sHzFrpwgYRHPwn
FT/s132Wdw2soSHl/k+fOtEPCnBCCribg481B0KNgOha7WsdGASkTSG1KQqGRoOvCcHLZn0XHMK8
X6YlDjhgcMSaETuqURK3E5EhSW2vlgDL/xhxfzvYRjjBKrJKVwGgxF3vgyaX/Bs7mE+GYA+dVBgn
SUIJ7/zgrkbm/wuHuUwA/MbtvpyJWpav2brnQw2DOPdjVjgnwdJZfhX2tY+YxQdB0A2TNyp8Kpuz
fE9jXSKyQsZ+tl8Qf5FVTiaPfTErfS5sthlhAHbpO+4soHnqiXcGUTzD9HkQ+vR9kDrEc5hoj/tZ
J4VZtCNv7/2yhpkYrBRsgDxJgM4LGzPGXj8k5WruTLCvheZkuYj76UGnf9gZartS3dY4gbox/uR/
XKwrxfBiNgKOrzdwAQsSatcKtQNESfg+tHEXHk9UAi0t+NFVDssRVWbLq5WoOmp2WfwO6mOK52d8
l1FZoAUNaGQX92JZETEqu6Zde8Lo1Xsy9i8+X6BsMEx3NVO5N7jsKDR3uTpDr/NJw+8Wdenupgfm
uHm2y9rzDca3CkxOPlU//lqtdjU5xTKqN6E2rKd48px4wmv2JJKPg5K4+rgm/hyYRtq9RBQGb8Sz
0pk8zjTc1bEOKdZ0s6+SdQ2JRmLs5AsIsf/oYz7FD/7fIxfNlPS4wRJj40EzywDOz8YKG058BJ7a
fY4rBCutayY2oN7wRqhTxw+mm9SBCFI0UErt3w8gpIiaSTHSvcjFFp/Zh44U+wuZrp0QX57MXxyn
SnRcqTq31kQHRx7ZHC/GwMJGy1fcj/sfnZp9Gm0I+aAdCvtaBUIZgJ61Tp/i6r3LO4c5+aVOiUx9
UlaYHYukpkZQZjA+Wlv6MPYIxpYV7/17qCNXxCMc93kCdJzSq2oOGH6iADDu3Rz+JaRAiKiP5aEY
XpZ1tUbM/yfuYqPffcXRS0dK2sMOl8tRtoqaJgUjnzVHnq2o6eL9ig5Ssb5IoSgACoEW9T0Bo1n2
sfKhnaGwWHM3QiUsOPgAYOkIv8KBwnum8ijJGGf3ky78PPVoBBlS6C6HijRRLcnd9AA6gton3tXB
7vaNR6dy6aPi68+mA38aAaVGooqppNp66Fi+DLScDsq69iIeZPCMnCsd14HrJcUsn8apiQlYfH4k
ZQepckCbmvi4OJjtyvLX+E3MWpldj3wj/JstynI/0fliHXh+jB8WoSQO6+Knuecmy7pi+IDwZrQZ
vSUTNOmLjfstoc0jSpi3oOTUYlcY+8KGwoR17ivcWaFtYhhCuzRYFCQlcPeYBX8NX5NJcHz9Phvd
UlAL88qitYJ2ZCakuZEapJmMuz0mwc31KJD1Bqlkb8JyxUL3fqvrFhQi25Yn+ax6fzXkmgCA4lm5
H2aGVuKsipIX2tTaQotY5JVj04Njhucwc2gtecr+gy79+j/PKOOmTh7PgOrmWmnCain+TYOUipDE
7eeOBtn0PZsKLCClxv5prkTFYC93AoUOK2pqx9CUbSsXIQ19P0cKLZztsBEtCaX2GkwjshgfOX4A
WpRus6CgqViLTgXl8juxsH2c6hdnDz8tr7oAo3vvOvbqBG/g+h2rQCOaPMLPpXSlexIj6eQVOtGK
mW3+wHCwu9XrVhLUgD+rHYLqz6vjDtfpLniIWw0cOTEEjdEAQRJa56jCI01NxnZtZztnKaUYZK1Y
5mVELXG7bXfN4BWBEB+chu7u+QagpXuy1Ke5epYEXVhjW0QrH8oQ87le10XTKSWt19V+vRfc7Vw3
gKU0/5TyUSWGw1rVZBOcxxSyP5Bk1QTaqP287l5xNyc6i5NcGV3txTLcoicG4Wr826L3xmS6zpr3
bpQv+1WY2pnfLRW5jZbTdgPFQb9uAemwJlOm1GT2I0HS6ggYAGthIYxd8lH0DR4NVL0yS2dkbS8U
gsi4TNqkX/aPjsw6WrvEbpAVKgE6nKKQ6tjrEMT/gN/Gq2DhWe0WqqiMGppz5BBTBoFF9AKeSgCL
aKKG90fpSwPPlnSl/anx733UyBI0G6i04LVW+7+oC0MaPI2VIwajmf3dq2UkHl0E6trFLzvIwBwb
VuzgAgQ5ZI7WUcvBz7OZhxwMM4oPEjzv2WpBZ3/5/4z8ihuJUdD4Vy/IchsY8VPwz+zIjkX570Ac
vS+R9cwrdQzyZOFr2aJMWh/3gJzAbiQosPqten4v3hlSP81a1FVKRfhCcbnyly/cqLbVAoFn6+ac
I0L5teJp0JO7v+ifmV+yyiUgS/YUotk3Eo+CPS7Ap/2M5xqZBrUWIvugjApSa3GnmfEUiRWLwdVo
bA3E3Ik0+nCGKDmP1L7ApH6p5Kxe1qv2EaLd4PhsEQZMX00fE7h8QaSDnzffuzt59m3Bax/E6BqU
P+ClXMl9gwQaMwcEResZeKwwLE0u6F6gkdCNsO5hRCw+eeJZhxN9zf4HDInHQsrM/6m8K+3oyjn0
jDkVQqnJPDII+Ibb9Fu6Gw6yR2Edb8rAiiJamGnQYKW2IadITG1IRi8FgaUjK00fuR9Uk/fWNqb2
CIC72Ig1scJEjpzZOuPlSKJjQvkZC//asobAjTyBBLbAcqkuRsYGv5X8GOZa1rY+NWrqjGlBTA9E
5qPbVs//LtwTCD+vpmqhEqJSr8lZSxl1GJyPtiAPJozDgiZGvTLBQHJBlnJJEjKSJvfVMK4EkTO2
6f2NWkEMULO/boDrhv5wRr0jAaK+W76fURbLp4alZwYW2MKSmbynSH1YWyTiBpqrRWSMAYwIDC1N
DSC94eR2ao31TwptWkG7bbg1GHuh2Ju2LToU7HDe2azSKj/tjZC6NNQMpnnO8EJTM0K/6jSLIZLg
8/VXqov73AnBmvc6cldYvttc2Buy2e9klgrUBhNv18ubFZmukPBI7D/2HDpgliG2C8ikUlNdgEVR
UyOMNW6us7vlTngqdI2gkmz2p19jHRfVlY/PKKRZgNjwj0pUvTVRfRX2cG/gUhKO0wsedB8A33fZ
uwfY0mYKCQ6azPcIgdLxTR+FBRMqU4HmUW1wZi7iXSCUxxwTdmSSyL5MnIO4m3jkWhWT16ydNfVJ
V/HqvIvPO7Zbh2ZRV1VlSlAh2aKfISolGRa+xpvTS/l2gWIys3nycIVXn7g/665+vlbhaemiOUZK
HVPPDJEzE55N2RQkR/0Wl6R/3Ql3V2lOCk+H61Ya6Uqp49JLld9QCp2z90wnusaaALOvhONSJTxO
jtDlDDu3LFZVSHEiTrhSvv4pAFZ+3ZDPFlU/UviSFYWof3qBLyeWxTaycqT535sy/pgOHtEAdvDx
wq2QoTfwdSVLiaxOL5adO664v3glWDXgS8F0snl7mgCSUPnj6c1nXf2J8zhcDKlbGfonGkQIRCQQ
oYPQ3lznEjn7OFYtjNk895qHhaObWqCPce+kp6DwFLXyrbURJ3/9AFgXn2+YdUIB45FrEl5YztM1
zLL/XnRRQolJwVCoUPxKVq0mBnsPd0Uu29Or28SWWvFvPiuHjxLU679zjFZjUT8kl0jwWGIfnO1y
vkqM3OQXY+hmo29OtvOlOrWdnF6csuzc+/hd3e8xuX8PZlLVgTnjAv9BpG7IvFZAfNTyHwPJmtvD
73kHNBsqhZ0SvNOjDQMq5Y3NJ4VoVOcdsqMisxpzXjDupNj3G3xEJZ5506s6RxP/OFbinE2nkXVk
Uley57WIRz6COXYd6T6Bu8bQiER6WU1xF/Qu7WV5QydphK4SazojXfm3ywGengP5a3YMZmtz7ylu
b2aemYzTCM/hzNMVRbpVjed0hN4uVeekrYdt+VqAgm0GVXLd3sA0o6LUy1m4mw8LN1vBgsEvsYmH
f9A1W+IdIPxeH8K6ZfXzfTnp+xqluOARW+bsAcAPuYRKzaWGRl3VGlAc1KTXSaKpYycpvL8biGdi
LUt/GE7J0Qjs4lAcFBd9eDfbi4OyGMKG66D+1HniKA3I3qBBGkhra3EQdStiTJFvNb6ZbJ4WMzg4
s+S5IEZrZtjBwwLiwEUGsETPm7MAdt0t3GXwGG6vM/NnyuMrAHqevFt6kMSsAuH8XVm6vOgTN7RE
ww16BWyHfCdU94BwSU2KsT/gbIyfJvue2daHXreAjpvzvkbqgNkH/TVfz0vY0tk/+eLhM/KMC8uC
wxbXcOE3LUhHAXgmTbQr1JTFgwAwFZRydi/oyLm0ibmQ0VXr1OO+ygZNpWoEK31YtmXo8KJZPftR
3jcfGJ+rwVpHfjdyGCZI0C5ELkJ/VS3rOvPWx9BR4gRp3UxD1+jP7O26SeqCrRSlrlnCjt6RnDvi
5BrozCvtc0VBFSz/7rBagKqXL0MpaQLnZAWzahFvOH+/jQRFs/cwEpCU4nU2Fi+LOXWWlsyjZ6mt
cJvTUhZmnVcc33HnwapkfCcIlgSsjlY9Fas03hnfB6EEXFbHCUL0CASILDLZ5XXtbD6y0JbsPRdY
vzQ9nJOo2F0FaxxvK9LuHLgNW1c+y1HQnTuNzkhtqHCKaRKaIaXJOJmDhrwQgu+TRY+Pfa6Pmc9O
DeW0ayj6VKV6BD7HLUkTTew//bze0Ez+PtIYMj6XyUSBDswSL9DWp+jfSiDKJ619I4WXU390c4I0
CTz6pEF60x+hzeBr2JU9CbutDAcfnD84zEd+AztOwFd96hYe/48iM5WHsbItmYk8jIrw+bZFGR5m
xzq8wvYFG3GDsXKgX1gfRuB4hNnsa9mNUVWVWcE49M5xBwnMGkkytvVdOeewM7jzcY/xfZ80lei0
t70qc1rIkAEu//jL2E9TNs0R9swSibaKzn7TxexErfdDnnzlBQWeYAVlLKYaqYsWwRNv3PhtHLLK
V1LEB8BzIAAUWApXyWAeAyhK1QwTprlduNW58GmPyZsrYQUqiqx7jWUa9jRx2Yjpla83H31r4sO4
GDmRhcHkAGWCn859/4zScHQ1R+oomk2r9OepbJBKNORX0IZ+qGSzJwYc9xE7Fbg9X6GBd9otV2eS
ExXDjFW+2fJRHecMPggsPeNAB2q2SWAgH2pi4/ZU8ooAGIx9Hfh7AIP6nlsNvWIGx0pSk1ia5BQW
XZmEEk2aRmQn3QkuYxJuZUC7wlPYtYa0JsXBBUFHQdtu6S862MtrhYFK7+BrK19FnOkFco8XFu5g
3XoUVa5OU6Y29sSQfL5+oQDqCtYPVw1FDRSesJzCBsb46zKgLiXf9vQIDfR8WbbW7zsHmXQrNtLO
gWozfOIp6clksmO4EjCfLUhgH3yGQDpmzCDYiSvyaLWYeWwbSsAsGmrAFwUV19/k6vn8kBVgkMNl
h4G97RZ7B/w575BcdF+mqvwHULesgZ+1WaVStxcx/OHOLBPLSaDcBKbe4/iEt56vgGlKuE1lKAyV
zIue7Eqgjwwf/FA/yPonScYtvervUugwnJTFGIGxZ2AuPqN+mepnnedxdh7GTEvbxDjsGuhtc3oT
DwHShoz2DiX2G1g1Iown0vvLuF1R97hovumqjVyhcpv6wavPOAN3lF1dbbYFye4QXsARKnNZ+PXE
XJtjSu8JskDTLYUYeyjVS4vAJGEFPh1o7nP448O0pyk8vD70KeiqI7hAhQfAqR8KiWW1DlVGgjZy
BTMh3mC+TxjFWvJGJOFcfi0v0uClYljpuF8wnLMu90alqHeH9Ya7mi4m3QjDqdAhGMhULv1QDUG0
gUFfktuC01rJ5OyQVQ3JXnISw0/ismyq7hNY/eux8/LniFFkbUOLhCUFWyzH91thednSNxnNbb/d
MQIznAsFqIc9UvITZkFiw8Vh+KTVxSq6dqDKbMtw0SJnYxkoFF3B/BVS6NS5SBElAQIWA9Jjf/0q
1CSGAcHkEwGkqhssY9vrhh2xriAWHodwc8BJaiBVV2zU5kHRBYqxKO9h39CdRUxCuks3lEqudELS
/nOlIX2CIpQuM9QVnL5ogkTIiDfR846HztUAS9Vlzlqstmge5AGnlg8mwydy8SdLntLKeyzRpLF5
2IB+SupwH5iuiBsfnz6jT8SZwzt7dVeH0p7OyOmOno3/ALQ8bCmEjJAGjHnc3peVx3uP6V8qme5P
mRixbS8gBH3hv1SEiKA336WGNtfLIMcvthgGucYkTkB2PKYTB4u9n1WgZPx2dMqHNfvLxRVzCrn7
EKJdTip84WkIVDpGLTrV150z/pSL3gN7XqZwHP6gnqoPlDiUWpkJuD/Q5RG8noC1EUHzPctzsl4s
IOkYyk7cIFCtOHNyTWOlkVN9CFTixD3JNLuxDIPKKFSeKfwIzCVLpUyP3spI1ThYJlv672Lu7jS2
F/HHOfV5jmSxRIZ9qdDR2MzNSyQ7CNQMADvyrLWf6U/nGp9YvF9oXiTFSLHqvMjAz5TQku+RPQIu
Us3LqDno9Imfghw1vLeKjRGuD/v1AC8UX93w8ZBa1fqKWtRO2lrQ/4z68fqRt1gsW4lBUkZs6Rif
TPFXvhxEXQXCGxF/hdkWaWgDpfhiAHa1A11FD1o4L1yQzY+Tfx8l1O5OYOmpiKHxuwSnOgVJyTfL
8zJCg1Sb/6Gtqt203aM1ezYVJCE+H1ppHbwlAQLNqsXpAi+KXm6mnF+AD+NZI/2eOJwieYqMAzth
pamlSxpzwJdh0xwkXk0YCY8hFOm5kgs9WCVD1C3g/4a86f6pqeRzCVVpsqALkwJeJ8HwXLvN19ED
b3jQhT9i/bTnMB1Dpoh38FpJ49iwLOq1fu6jf6b473Nqz0xYf0kInk4gvZpWM9P3RUUo7B+xQpPR
8uAuDUqH3Ya2QFTR6ZERjYUcfVuOGiGsPxeqxrR4AijrxtpTCNse/H4eCWkBtENy/PBcICAfrBld
6m5yWOlCU7YoGC6Cttr8uvUpmRMSHDEN1BMoSbPB3VuFVp1qt2I3rIroBh2lQkEkg/LuBWWbW7Q0
BMlCw8eekcnMP8C8KjIi/SwTNmsmzXLylS4MhX/w8+ThS9YLT9zv/P9tAnPVe2Ybr9qWO/zkU18a
fUhZZI1Z/Ok5HSyPvge26WTPMWqe11vueBaY6P3d35HRNaJMlonNWWsPoFDGYsGgXwyd+/Jay9Qy
zsSgWttHxnv+ap3RUsxa8u9gCl9zckIk3AUBJBktgjt3XrsS1MbhP/fPEWoods3I+pdWosSr0vVo
4h5dQrMKw22Ie0zU1yGunu2BylK9EDzCLKnu9p2qNZsL6HsNb9ItH2/BozbydKHdk1OKRQPq2WAQ
K3l1dD3eh0gP+ndSX9LW3rhSqMSd6qjLp2WrzjReipW+kGSsdEmQntuHKSt0BGOknLiVCz72vz34
2AM9JVB5if8jXP0nV050Z+snNKy8jPvwrPwj378mqJdHKys4AVU4E9m+0Lh4spM0g6I+ohFfrsya
/9jk3T0/JL8oR6CjBata8/0xahZY2S27c9kf2COVGnxYwAcHbeGNSyFxU23329cXiv6wro4Lzi5w
G7R9h377nASxnJnilqKOwT/xPYGuw2yrjheplY1zZ4yEwKEiOxrSmdsLQyRuXNMvxvGimjV4RWiG
HdwixIM6bbxYcv4rqQDCBdy9obsOlwTvI8I7hwcJLMA8JMTmnJqDL7Hk44TvFm9xvG/pewg5OgUl
Whh1+o6MDfc4nDMDlrmPMOdZKPgWOU0Xqr0s05u3y8Z3DfqIW0h+es/nJOUTcuksbiwMrgi/hmiF
jJCx1I1PDF6psW2vd4+CI6cZJaxXCeaZpH6ss51nDDsZwdzZEYQOQ+iD3tLnhb/b+4VeKGbjcsxA
5DTCSJVn1L6HZXlCUc8D28mVu7EtbDY86++H1brQ/lvwAcY1vC1i5LwsyzE8IpmMocdzCw+zmUnb
RmuUqMSnIiPVrp6lovol3bx8Qj/LfhL/MXFjFJDLQJx/dDd8GKcX4Di2JECkD9adRXFZ+Vo8Kv9D
AnlelUcM0IC46KJHRgpCsNRdHQyQYACFONa1b0S3f8ZxjLKqu1JS0rkDPjVI22iejUaHVMC1DLxh
tZD8tIxHxqJVhonGtRs5XSLh4HA6ePEyu5smApuwPO9Wtzoe7RyuFUNq9Wr5dt6TY0IFCqilvt3P
ibX95RYV3PunAG92Hro3YbR2d/eaj+rfTCJp74iaSHlPLzaEWR1GrmXAmitjyhVBUggeesnzMe8v
mUr0GDS8NksKF3AlMK/lcbuOv2F1Nn3ObZcACUvYMGsGD6UZT+U+Q7ct5iWokFNwQOhcYrQ6BAuq
Bm+m5FkSnI+nB1wu0BoFdq5XY9gAEUttXFyDXYEbtOwcIBoI1HIEIFEa3o+UgWPAHDfMlpMfcpUr
dmCD0fDN23nUv7g/jjPRv1bBKgBzBIteHgdMWxow7WzVSIw1ZqwsTB78ImneXD5s2sMMd0mqHUbU
fmU/mPA7IMp18fT8+tNDtU08uozfB5Ua2VepoG7XGBK1OIlJTWDW1EFtsN9w6SwSF5U1V0FWivUc
uDvMQxaWZjfUCE72/qF4zUTGtLeRFF3rM5MAHZi4/mCXeVzi2+ead8UHZAVkkynUqhfW9cAje1AZ
GJqBRJ+RN+oPRHgW7/YlneRWHgKDt6EbLLVpSx3IJEq4EtxAUth7XRPdDBUx3ooGylmTfY7Cc7qp
/Z2c2rg6S+xFRgUhCaxssOVkAvo/L8oTeQNzLahu+cZkqyIKoE35Ad4WtB1iR1dVkxPzMyIKgRQB
BSMv3Ysh0hMqJmyqwAVUkCHC2Qx9QIo0/XdQQfz3d5K3etQN15B3RxKO0Mlksnub4StCxoReH0j9
7ErAP6e3/FcJ1JSb8E7LVzRjkveYscIWvu3lIf5U2UbskaI96V6H4UXETDWp4pL+gdfnr9Y4iHeY
cufy9myAFJhcVmeg7T8fABHkB2G/s4TJd1X5PmFdEtHKDQeGyIQmzTs9TQWeYrYeG1gQr1S12ZOr
BfpvjGq/MXhepoTm6kGhRfHxq8+BLGZ9jHafDXigqMvwP0YB71P25utQM6h11mo8FTmXTH8D6T9Q
jdAhoqQugk2BVwpl8NKrsVkNALoOCiE3/BuE0UnIBJw7NE7QSzGyCl2Qq9zK6jstc5FFKIPztrfz
vk+A0l+wKmrJBNXm4rHqkg/E1NdQSRt9Uuci3xEbwbGa+ZXUtxWqNccCzlG1EQ6vUigP68PgR30B
eJRquzmjfb/4IfRp8KOxl9Os/1/f7X8sNWarCOYbNEJc2PJs/OWK1f0qmunqL4NdnesRJEyjttG3
FjYTs6n9SiJC53F58JhfMpvItE2JXwl2G0sv5sWk3rhsEr6uPFuXZv6sgqrUUiBjoppDQS9Y7ixO
wdNY2wDw5N260jyKtVZxHz7ngPfptMcO978KXVuBk2cQokZ4Nyb+HIDdNfUIXAs6dUdRPTm1fcOi
2/cE55Y6tHZKHw+wbkliwXlIk5U5Zx+G1qjHIt3CLIO1m4I3pfuQaE6qOrqh1ZPHvJEhCyHOW1RB
FmQonz0Hvdg2LxcZa0tPcqPCMkuOF36QPDN1gAunUDc40JsWYlu/+wbwI9ozxf8J66ykBxNFL7+4
urd4OyTWFP+atT/nGKHSHp6ul29Dl2fWJtVdIzv0n8VqedEhmkm6IjTO/w0OR9NuJosSB2q6PmcQ
UqITa3CvoKeIptZu6K2p2pEYRUmxXtVfjZ0hHN6NfXf0SLh5X5OREpK4MAElfJ1VXY0gCCe3ckT5
ysc8sf9jGcu5hMeipJJgBLOuQOZfSwq3uvk796I16oO6VQiW4JT1d1360xy4MMGdWFoBxPOAGcZB
xaOsuf/Pb5KVYZXp6SmmY8R+aGd4pSMPnD65DZr/Xi+y/1kQd41XkolokkJwSJ7l61QPo2x6rDPO
iHukUMQmuFV/rDnYhBOygOVeiMkHrekJbaEE8EFPQb1SILbKYjzc7Dzhg7RwOc/JOlVhhpAQ+S8c
JisvS9tqiLWEF+7tr/XWSj0CGxnXUvqvMPPYEPsHK2A2i+PFSZqXFO9OZj3jiU5pHvVTfnt3kbQC
s2fudN0iUz5NgOOqsofnnGViNA8s4jEUjQB0h0MwjBDmA7eCutRxmXSzRfjbb3oCnUW3bs8Mtzxm
6IA7HpOkJzOssMAo4ateRa+76p0uEHOb3PJYtAhpblKIWa8UA37a4qTwv04DPtdN/EmwMb1FZaJU
skNMaYgS2phr4Pm1cClvLw04lLiOd/I0cInQJtV7PDfipY+ITiBlNaaaykqg6c2BSKh2BxGLj2ow
t1EdusCtToSxzQ4NpC364dTg7lKj2wAjmG8HyopkkDwA0sUxa1MTyY0U49tJqmN/Pib5pGsh4yU1
ao6qS44Ykof8waknmpfJiHmNFVoIzVmDdgnmUr++p7HK5qsCMPRFMx/v1QVb4bM/M3j+5zmpfrYl
1WB1fWQNcKCanZsidepMsXmlB18VwD+u3F9ENg68Z2UMP3ldNKE1aBB60XEsOHpTL+Y7wDlG+mjA
DIa83EdRbmcF9zF+hPCsE3e+7dQ1EWJ1yCsZjSz0YaKSuPrBfdFnAnZguAF4gI2BTK/9TS9lXlQj
LSeBd6vAJKMNT5wtG0L0/NnsvcguGzXEpPm8UZlornGk2pIDZ8HKQTFETIRr7uky0nomHFPUabG3
KtwmARhr4oblgeBE2TYOiRl2ZpmSB9o/s0wNWA1UCvyurh3ZgRxLqS2NUo9dFP51mOTtXYHZWmoH
eomn31+jXQuQ6esz1qUqK5PLrmr8613/NY4Cvbv1QLfUcP+0ETmgr50NyeSDuf+dOnnwNc2KmJ5p
gO97L0XlBIk4gfM/4gP4LFCHXYXOVNTZxL+8epB/EY/S3j05H8/6E+C4BPyp5hZDRwi16TtehRba
G+9xVw7mPCFnhl645ALh+sj92KAmrh8TMz5rCRyH95on9cdi59W358Wq4z6KMUR9HTQVDRbhczCs
efZ+hsZmBHGZSfZo2sSWlJDqZ5BPQphN7pSRJd0CCkqTTzGYkowW9jPKRQ8478xyUcNZo5EMGG9i
j9pgbAnEAm+QzpqN1EwEKuavsfZjFm65vG0OLkyRCNhSXUgr0v24XEy74znp26nHoKR2fAiUMOrQ
8hIRF0MWf2ddI+iWdDu+dTnXhqWCrdzctIIbQKIF5oqcHi1TUjMhAjEynxIixzuWW2txxqba8iCJ
THySIaIbCocCiURUYT2HJG6iR6OlL9JHocbMhuhbKsMFCQAc815JnXfHBq/WnHkHdEzyvThyxA+n
Y0OCCHdrpNnGcBT0l24vTD0+hpzDHkHpSj9mRaNTOcly+LwGp28q4c1NYCG78gzAIvPWSGEi1Dsi
+/T52PQ2CkMQdpMTXbZ5RLUUoe3MUXCLD0RPtQoUc8DZ1ArtVAzvotxJNuvMA10ZPKI9iAforx+T
lgmbbs8/Olp4FWdKCuVczh959OSYXJf+l6PbsYtn5Z5KFpNsVmutiSy2mvngBteXMK0Cl6EdZ+ni
GOSNuGM3GpjTY0TQYmpgzg7MxTwEgH1hVDXJq72ovBseIW5J1mCmbUwTVm+Vm35ZTAlcbyHKGgHL
5OJbZ4LyJ2+9Q78CvSsZpySbPXQOJ3vwhJ8bfxTmtMjhOBX7mlDOm2VcgAgj3Q/VWy9OjgOFZjRa
UsppSz8jkWRSsfkPSL0d2KFsYuCLWpNE3p/FKYhGGCBUaFehTcaZkeeQJ77ZfxXjgineBhYJOKDt
uzkpKzdX9AVZNpGmQfTrPsrtQeYV8zhtnMW8c+uV70pXcm2kiD3rROiABWzYOUtdkkwQbwyGYLuj
xSKZ93gg0Q/xZ/uI9AM+lA7pXkc0V6tx3FEmWv/dsO8tH+2LU3FAQQC5zOLQmKo8WlR9sMAJeosB
W1PzvBv037DFLAIBVjd16iZFdc0ky3rRiwG2Cb4Z9ISpGQVmKK3oYoOyLgfkS3xIjaYkLy6u+b27
RT5nR8Op3ywg4wgypFmhq4FQ7yO3hTa/h5DwNb5ek85OWFhktkyKCNh0r3d7UOZQDzA9eErJ0/G3
z83r0w7wUJLrF/x000cNwsdz6a1aQqyzZ3lkMJsLEnbUHaE7LuTlljPFtL6SBKRWpS4m6cxeAN2p
PA1EJ1RlKidZi98ZNlhRjH0uGPxmMCdSpQoHoXc41PJYKDsKhpMKlDSdeugxiF3QdiTll1t19BF+
EY16mESMtcJgaL9pljsKswVnsF30KclIja5ZlbmlITsd0JApA+zASOZnEnWJ7NZWXv9viI2L05aF
XYsG3V1jieFZBB6vUxwrKcgLx+SmeBiXKQEiU4s8zI2tzh+NBf/yQARbEOwW8d0t1PYsguEa4nJL
WPfiNYIiibN+II8m72XiFJQID7gS8BNNaCD/etpXy9oXFLUevis6BrUenOfJB8zj2egZ+OTNjabK
5THafD8/QDhfbhv3H0QEMH+5q2pXUvTGhfDZDeCKEaoNiB1fUB7EHS3voaFPz774VJVoPNyzVJQg
VczmpTi/5ggm25MrxuZAYGhFuV58Zjf60vYP1hS6f6DbTsl0FY23PAgsc8Svc4OKUfvBiM146RH3
uMATDeP4rOh3kjsZ2vLgo51kfpTLhPP24jo/15UAS/h2QX9tj8D0MjCPEPejrUcKpOYuhZh7FE09
v3wv8FSSX0nyNjXVqL9ACr4xE8djGAdO58NOKGBQm7PJs9lSNLkuwXlSDGcNlrPmW1CajCBskTSw
E2AkMhWqgfPeb7KUQbR0T+drgiyg97s11uRo8o+E4h3OBpZKdpyNkUPfTf2uTBStaC+bKmDEM5qI
ecqtgJ2Fq+5wsJ+pXu8i3olIsiNwdyijeXKB/GfQkVCbIrc9jZmmSM16rFDEHTmgqY8IElJ0h5FH
bJ5vX96ex0mCjJr4J0s2ebm3I3QtYVvWDcR92r7YbunpTbza09sBz0tMBnfttSXX+98Z+E1y1ZOp
/KMCT0/bR/f9PrMThz9831AQhOkqugVLL3fkFR/s/ezBSVE3/K4TRqWfojwBKxlPl02Hb2NDI5co
qnO3HUvfg/L2UaOpVeCmsFegmIWnxsGNcKDF6MKEsfY9mEZWdUGUZxVbohygItwCgNVI2Bjm1CkW
byCe+1U2vhloNvgvioUrMQZwWtCwA+7a9NzXdYxJt9Q2ETFpnis/xgc5CMNCj+/u5f5DP/5FzxkR
WMUilpofiyUhoTcQ01BgTGTtCT98kSJ2v2VAb+JLmuoe+Lk9E8dmf+qUGAOwx3jp8HrMwjRADS36
B6FXv2LS+AubQOVhDdLbQQrthNqhcL069dyiO8prOUs1+zZaDTHjBdsavHrUIr6x48RzB4SIwxtg
/I/psna6kiQbYEBSXnVRaTkCVdg38kmDo7T4ahap0MDtWkAhxisO3Yy0s3tgAVH51sZlN+y+C9Ec
qp7FzKVOKtU7sKgIvZiw1quZVT3ZmH0Xc/BBwGsKpmktkblko1jEA5uKQix/cq1yhBS/LbquBmZs
jv0yt46qTv3tdTH4uzYBjk9+3O/2rJsPzq4MNRTSFR6GBeFqk0ZlkqYrF0PCYApTO6zgfU8tDY24
PVBjdO/uAMRrG5IHNp8gr4MwXnGBgl8dp9Se0wU8wQdgbMTftWkCjpyMTUx0ZJtOHJVCp/ISoofi
nfVDtC3lMlWeAFJrXPYO7AE6wiSb7/o7TvXP343sL6siKo20lCy7j9flSUFQv6dnJU/OObBYQHik
qptJHpsFNVn9FE5V5jMrue9pZxHUtXsDUe0UIL/zzAie7ghAZrAsmGosLSldOk5we6LgCGw47Zr8
7arrNBAGrkeMBOjhf8oiJpCxyuUpNV4FHD52d/Lj45eSogF8mgILzA46ELwuxCYQW9MOxWwecgcW
7gg/VVBgfbMYEGAl1zQtDy9QrSpFVj7M5rPrP7hFlfyLjWkKxJki31HyeYHbYMza8fSLUfQOcNGo
OR+pp9h4fqxyHutwc1MCmflpjxbYoiAIeteC6aO94DygAIMb+G1Nj5YDf0iCV1UdJB4BTjPCjflq
YdowIbn3hYwpNul2wpWJvxaoJmNc/rRFNRuv6r86eGDOghHJn70sxU3S1NdFxkgrSsFqVC4d/THJ
mlUujpLrSTJSGjTmaUIY4VvAgSqaEx0/hUJ1kPtNj8EgTRDyrblCD1cOY/3B+W5vrwhivk8o8P0o
lxzahTz7gvwhmlkNCU2Rwi8BJog9aU/L0MUrDRb0YLD2ZzZKgftrGJRoODOLyTLNtoD9lZAooSzA
R07PJpdu9jIOVxcotFam9moaKuBqgVupaKB65tdzUvriF50D1Fd1p36wEYHruuFT3GLGo+GxghH5
dnA//pDlQ0fMu7FAwhClI1MjRmrtrYRp+7L/wzQf/hEmWfB+YasAs9OrgdbaKHRvyl2w/H6u8uuK
weftNUmZwE4CnUG43LVnmn9ToMt8nh7PgdaBXdqhbchGmsAun/BDsUxBMiKDeK6RYR/4HagFo+ps
AmsNWS5ZrPAM2SIMbzLlr5v3pfTFOJAU7TZh0HUna3WCmfXZHEmhkrAZEju9G9a7VXoDqQKdAFlE
laxbXidL+o41WJG8bR6ZYHdX4VqyUKlWQUDnZ0pay9rOUmLn7Sr/Ef8HwJXQN8etl/0UrHHcXpJ3
7f6sYptI/GgfD/UVSi9Y5b/BgfM4waAvGpLTnvjc9DiNx+iKdD4VXDSWqW1GoQ0qAnkMQvgCXpYf
g8kbwPSQJYq7UxcHHGCjxkS+I4iIDWXNRu98z0YImhEWTDyW2AI/WVZymosHsaq7QCBgKPAA/jA1
3HxAzkgswqUz116tIsk8d8NwZbykY3pgAJDzGvpbbZs4YXLd/hTuSx23aGcC7BV7EN2RrD69g4Ss
l7FcoMOWDKH/5VXfImMPk1G4CSj5y94wjgJehloMLNZsg4COjtomlJqw+9sbdTbYgf1e1tpULSSq
Xh9ZpmSGJF2PZpSDHve4LmtkVbq4Z1raqCnrCMvp7kO2JnISdNdrWTC046uKzyE2M3V9NhjP1Axc
QS5q1duE7iljDhZ2gWYaGugMh9EoCvIZsCyz+rf5qWeCQhWpzE1/0cMNgDBpJXNiXNV/9FndYHKb
m6sNJN7BiARVebyzieIGdbYVipLrJKVhzcyNCjnJicgv6y8QuPxZ+mlFpyUJrEtQfYZGnkNitFQk
Voou1M2GZC+gm7XdoNfMk8ZOsnSXMvbbWebuCn21fE8d0Y00FzNModd3Ocim7VJZi2lWNorgHQMS
KkPNeHHZKRJ+CN2a0a2c38SHdEiZpalnbumFzSRDRrylYfURFiRgvhhXlWDUV6wSOq/jt3pIgQfV
DlvKvQwg0y6+FzFH7jltmbBAuuzYrOUismvFRcIvBept+nc/SLufZfCN4HL1ARX9s+xX2EVe9dRc
/MKMH4R3lS1mXZYMlZPw4Fl3A40HYBAR7dMeud+LdsyWfESBf8SpwObt4q5oJBOIi/Lp7+5wPm/Z
zjvzoHp/ijN7QL8XwiC38ZmW/x5Zv5T3ZoNTC4dPh4nwFrF2jx9fV3IK2Vk9mgKplWKw7I5DJ1zD
sK8Fqac9lUiZIVeHY/JdYcY+pUVQQYlOkg9M0NUxAqkWjwPoWGhTpdjlQGScUgB52E5YqQCrjSZ+
X2YvLvP95wPbvB8ikX6dKZ7u6NysilsV06mYQD5qkwhjqAAaybKT//CFifRq1twsWOd59PkbLR7Q
DJNQKwKIuZZ6Lug258W8JA+4WWEVlbVLqmaBoLgtFHygBfn2LZ1E3bZOOwy4lyCfpOv8w8y+6sgF
pfXGhZVtPD6C/K3ZZedtIdewAQAC0GOxMCEQaBcYiZGmK3L/BqzWQv8cpEKrmST+cs9uhv/uDWHo
gdG8DlIeJQFYRpgj/ciJsw4fZoruq8b+l4VvTZz62ITw5Dh8Vhd/sVBBjKGxaISOi+GGcqa5IWqy
7HYkZXRAl7YwDBP9BGe2jgcpgvwtsWyBUzktQSWhy5m07ZGAiIgi8v275RS1755Pgip1G69csMai
kCartcXxZuEoK57qPXjDIN1hc800TOIC97b2WFNRtxV3sgibv0w1Yo7qkUsM3cpf5hWwIJW2DIB/
SS2D8WcA7aV//JmFDC5FJRaExXYZ333+ufly6PDPvnXngcOJDroeuPhKW3ohLJ9gV7+4fNREhjyk
mYer7hq/HhnkD7YAOATAs1cyYCHEoPlf7Eal/XSU1KwJY8a76yAStOpIOGykeOuhwV/DxzkzXXBe
G74zVL8lL20NS0nIosmJ3CxzBgA2BmxskFSqm3WJYmNwdMOz8PGgv3Ne+csXV/CTyZYSbJG2v9SO
UA2sIYW9Ar09UsL6Le4TqP4XxSVySZt8MXuRBGY0AKzRkwnEHdDiHQsaaez//UlO9eEGa69cP2Tt
3CqOEWG56GaooaNFKpy5javkDWrrm8XNdrPP6QQxWdZf8/PZFAMxcQOeWwwV0k14ZpTjOwoReQx2
s7LHBpG9/ZQLO9WFOoE0Usxe+4pt3T1o9Md/xYdhDOt4RH8sUwznKifXEOej5VViU9BQotBiTSR8
QdAaSXNAdk8HcH9xmgi03ZpOQBT0QmFovncOgA5XkJEf7M+hYBU/zjP8wA8nH4K/EHJKe623cJV8
96xVkQfhRyKc4Q0uYO6IEwvAlSFs9Eou8X1n1DyIFfmxdZlyMKvTEuwfxs5q3c87INTQWXn4Q+nI
B0DYDx44mKE8MlzVX83nzcHv+elgEiyEHSuR41CHKD15dI7aue35gmC5vwc2qzMXhkpvNO/A1tsu
Dahoe0RAxdZhY+9gHJWtwP4V/9i0HvW0RJSgmSbj/5GriBG6/lEJvP/YjjlNmD3U5+8l3Ldq3tF8
22k0qPjdh9pA/Lk7rdev+wdxaftjQOugqosppEE6LlWIuHBbpYHxw3cilga+19pJTijZxbSxlZ4J
Ld26jg9DvOU30CUjXn+qq9i7XbkOQJicBXRR++dMe1tEmQg44kGdOnnpWhxRZeX3fCrd//4EwccW
+Yc04pI8UNRMRuEQv8AmcQOlmurPQpzMeBjZqCo9Qvy+90lZlVWJ221p720gjkT1+jEFVCOiqJ/I
aEGMsI6KE7MwgxaYD1vdo7czTH+/Xf3xSiTjIlXEkdAw2VFHPjRNjzlSxxIH5NqXfoXjXrhYphuQ
QQz2bmrh6QbQp0ClEpabTaGWoTTy9T1nE3JuUuE9O2MGY+dM+w2pJfexyBxCgdtsldZxfVGz5jzI
C4DJLuqzoqocBej7fYoKiihxA3gpLQWXP22dRTDFXL+e6ionH08oNJ+K4i0B6Hkfe7ICQOMSIjNS
UBcd6WtF1ewDwApTOv47p+OPnFLZjeBrPdybLmRzC8yv04iN7wejSqKXNOfA2Tr597Z7H9YDKBXn
u6yXZSuuF+hdIS6xqJZOuiaWiz3sHy71z/HR/XpQbNrEdzWt3nkX2sCd/FWWf4Pn8Hdkncg5Qv+Y
szo3XKikZSihzSIY+D4TWFNKcyqPxjYhB6IuV6lPPcE+IjIQBWW2BkYVMH/CQMtlJh9kw6/Fdmxt
Hc6lpsQxfVJtkhHmJzXUVLBkkfePH+RlUDgJfPtGpqMvjYIQGrjEfV0ZdK4OOueS++glycjGk+RQ
+ZViiic9E017ah0S7pfvo2jHZzAus9oGANKMJ2FFeSaqTE82cBBbMh9arVdzDdFhuDLV8QQ/r5+j
LWZeWgduWjqV40XEaUG4PPM+DiQSI00//uTPxO86chqRXri0ZmLXK82mTOfe4TmKQimvHjA7NiZ1
Rdf89QerYuAcFXXCgPXKDtABPrSatDy8Oj9hY9o+e2cgfzittXgGg8oecF9US3RMF93KT/ob51ZX
nuqE6JaAihQR1JeGrcgsMsoRpb6K2vZrUQnwB3TGr3FXJHPGImjWAdta83wv3n2AYd4d2JlpKGvx
fjtyug+/wdz29oTqm9AWJcFWMh6IzxRRDkrzk6PAJUv5Q/JNMkc7hyDXnWYPQe2lL55yGVwYyNz0
XpuksmrwTv8yHgMEfZK5W8fCnkJaMRYJ3Qxdh+BLWNBexs+CDEj7H3tpCJq7dbhpfJGzO1Z1F9Uv
IjbpvD6oDiWp7s5gWv6f8mb0SpYoWFbiVGpf3bsV/HjZ+Nc3s/Wqjg+5MR/yizQJbPLTxVg8ifPR
j4L0WoiPqhlNjuCpRJxqK0rYPXour2K4MuLC9vUJpV9difZlqD0Pq+xbW4AJzEL0asJeWQmBhMCf
B7Aks740E0fDOLA3HWut+eqX4Zo/VoQ4vdw/zsBwwCVtBt3EVjYMi5y0N3E66SaTkuZOwCyQdK4M
uHsDlg==
`protect end_protected
