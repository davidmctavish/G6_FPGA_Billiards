`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MVrW3iH1zuJGrb0LaxOZfWREd6ahohJrHPBC6cTQIbnlTuiKWK2HW0ixBATydpMminmUZ9o8c+hL
+ULE6mqtbA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Su+fdr7iLmwio+vYILVk6UZsrLxKMznntzIMqRTPloyj/ktq2DNEtMc8inYpZ3+1DsJGMqZH8Nv9
BXtRouEXu+ut8d/KMKq2ZJeLfYegP6vkuSn6VjLDTTw+a23UOy0KLDVDzVYWNwlK+lL7cNABRzRO
0EahhBqHzAhZDH5KAHI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WwPlYBbDXDzenyPcViY0CZW0dq0KNuAJu5ErSb3mBnA31Uo2qvHMTmC0G3+N46Xq4PAQW0a6l0ud
PnISnEa6RXxphsziPFqlRUBpVq+OfS0gfWagub+83hZdpnZXV8txo9E0Go6LeP2ocguMYy41URR/
/szX/Q4SInrUFRes51lfDKVZ4JkuuBDBDdTyd7kxHXO2S4TFTFCanM1b3USubtDwbqQlFmKkJ/ig
0lLLFdMWm9hSX9YUqVg21rOrrNaKaVH/zXCA4218MwImJ1nYkc0b5qsJ/Ve3dAaXC/uyybt0RdvI
T0m1xAAPkaZ87ZHh1Rj+KJE/ynrneGYe0Tye/w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mm34ytP15m8qswuPYaEJSWzGavW4BWN24CbEdOE/hvrU3jNidCHc7b6fSurzksKvieXv/sLpT2hd
gu2Ack21ma/huh9SRIVydqiyf67llpTVTZv1rckmTcNd5C1mDHhX0IJN+nnLtvoVGzsTvrv9u+pY
zOx5Fez6UuPqDQWrvuc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Mf+ouAEOoQ8uMP084TLgBHEnQ6wgksNLBmRPsdAzZqKs/imLoMjJ9o27nleGH42qT0oTlwUJ1VNu
t5EiNghAs2wLRz7xPAcXS8WgAQM0rg6WTqFPUt5uU3GZwCyf5DzlmO1FI2V+/25fYLrsYf7lIIoY
xcOSTeqXUMjuP5/3F+mS5+3fVxcQnfwTHi+7TauFX9+TCuj0Cv/GRB58OG7jxxlQxy9AgzDC43KV
XXlL+wS4c1W9svCkd4LPS4uH4lExwK28fcoVvUE03T5+k9bVo6KeNhcgTId8w09ITLMphV3GTs3+
mNlKgeerTpNzkpZq3VI3LAjIHwqzzcgvR+5prQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`protect data_block
yr4vO0PzksD2AvHywoFSp7onzuwObCWm48pkrXcb3xGgis8E6HvE9tg2q9+AlRsYn2856UQygCIC
SAvPlpINqPkOlw2uBbGxqloFrc1ZlmpepzHLMHS7mNaRxdmwjKYMSG5JKPgq314/X9+90lPUL7Bb
jKrrK0AkIDRscsAXIjglQyizwYxEwig0sx7sxtmZhBVM8n6Z9QhHvZoh3/DwfDYsOm8g0Tbbnmxu
YUV4Ti+9IhrLqEyqG40FwCSZWYELY0x7C8mFohuOAqsou1oTVx2P5KTK29yTdPlZTaZpWPipnD0n
u9/wX1T9aTOpNeI6YFgI/EwGbztxrs6TB1eF9ILXIE9bEf1pOT8zHplukNOW5mtAx/BvI5pT/nc9
ODJKGkAuSRuVw30o3wC3UIEWnGcx6iIYbLXG/4g5aY4mrdP+MJgXzKu6j9tQwXAmjCnBroebAV0H
wu9mslgtDiIUQAGS/BNJlGIm/7rU7HvXdgNWYyZ/EZ132C2sRk7FZdcEkLAdNXIKleOdESM+YV+v
1tX795yeTDwvSFlY+6emSQhx9MI1+c3JkfJJvoKZE01/WR+l/q1pLH9n4tnA5r8XHuB7qIX2s7S9
VMTAGpEyUz9OV9gF98ORfMZQ8b4dpHxIDSY5CPJlfE4rq4KrgifKdEDpvEIAt4uYaaswVzEhlf0i
PTKpLPMbgZ75smiEQExoBtgJP9vaxNKVvR2UHrUFz08VwY/ovILQ/iHf939ZMZSF5YVbYcGpeO85
VI8rT8jlP3C4QqhGw6dSAXahPH3VyFUSbfPx9efzbWhBE3RdTQKmcOerMMs3c4R0ja4POp+xKLJ6
LTTm3aWJT7N4igQEgd4sA3ubCBkWTu4eGPAHtlsOtb+8aKg9EZwZt0dtuQdai6GRV006EgMlU/4K
u07BrZiUpxtDdMj4NfXrB+JC2OUbsvjQgHJDzNdhYU4abI8weZG4dnpC/wx+7vuLg/9QQBwP0auU
FQ1cF5NVYBLQGxUurr9iuBgqpQMPU8ueimfItLr0qm7qNIz7juPXU+UG0JAVwY7aXNnzfJWCDaqU
GKn6dYBxRBo/Dkoa3tElZWLJ2Azm2tbaTSMdk9NWosRleKcJQUKF83QhFkjc3a+FeJITaw6KxOvE
YTD311xHGN3yOKsXvb/v6owI0J7EmbGgSobPmpNhRnpuY8nJC+jAz8diT59MOnbm4IGBM7n29xOI
VKgMdRtr5QKkleagp4eEBz4RpPXTKuWL3pHAjiPDZMZWgSiPd6pYoQriI69IUV4xAGUuqU7TG/nc
B6BZAm/UsYxw7F7PO0ZieQPDklWtRq8KQ24+65mD0xuoKbae+iqtQYVojPFY1lEozznyw83UbiJf
gH/CpWo6iByHGcp0knKPHIkrFyFYJsF5gg23Gr5jgbSuhzWSynEqANgiTQ+n65PLOE/91AmO4ayX
2FQXaGazpfmkE639R4OKv3Sn2b2N02VPrImC4vIZlXrCzCjgtnlx5kwHt+qVg+g7fGRqEQno2BIU
FAXUSHDTtu0v+uR0E8uJvfInyazLwovz9KZa5H8hgoei/NLjIJ1oqC2CcPZMvgu0sAsCVH9cY5jI
72PIxQTLDBi4XzqI+OHj+13dbmaKi/6ufY+X8Wm4uwE4qZQLFKVYtl8G2lLy3/eUqRzU84ii3+T9
0+9kEpImxYPOIvm8BV6mJqH83usAOC4lJAJxBmXdzxiSCENa+3PLVYUpevnB26HcTxIk0er9gtxg
vAWtTDodcAVjQrgzVXmTzEI8DSA2vZbfWSbvtP/D02H3s8D8i+DOWS6lvhaDt9sTkzJV2DPs63im
zyO2+HzhTqqpcDM1hufmIkGBV76CJKW/MfB3m69anlWSV++ETGMBGIX26x8Lpn61D1qjdjpDsgFG
wfxZ8qtqZdKbYMgt0+pLxXVOoi4P+yZt26NxDNaCWaIP2cT0r6D7oYUIi8hZm3gWYUc7pEEnc0Af
y6Mh7KIjB7/+deGoyvRtsAc0XGfMOeA8wWumbF0lWORvM6HlrGn4a6ddKzbzhx7rpI9Lb/cII/Wo
IgyHkWgNh/aXEpieP1a8o7TauIiMsBKbs6u04bdL3x+y8O8HC6I002ZQvAxKnLe4vbRWNWlVE56g
qanEj1+OCyNiPsTuk6eQJTHs542Qje9DmHNXb5/xfQkw6KtFcdLGGqwEFfHtVT0gyujmCR63+ajF
BDBSOeTH/uAWUgNOPgnQ7A4cGN4jmNZMH/G2OZ9r2wzu4dJKMOPOLYetUiyjELEvc01Oxf8IbkRC
kjOMSTBWZhJb4U9/8yRwqPRe1T8zyA2DNEDHItoOy/pyLDnuV/pCbImZp8QRHwoGF6Iqf/0kWotc
qiTuMTlan41HXhSXXJ6zpW+eg16pSyiNFZi3kNdykmMMpaQO1WTTVaY9l5mZgoGbPLdVaB/8gKgb
92Tv9yz/1qdJIgmBEXxh2g5Aax6N2EZhArk9ndUU3FdtPY258YL0kQHf+HO/7F/eVXWVivB4JYEd
OB/BgbBG6v+jwRpFnPhHBXkx45JVDg4RPbNZbGLDd2Yez5VlZ9dWDpYyyLj/lwW5bIF2HRfvQWAr
IdUokjYhD2F54Nlnh3jTkIYfLiIlvlpxz25bIx7iwMMdRxRPHXGrPSl6G8+CcqeMSaq6KEnlwlh8
XfOQMvfIZq3leJnAR+53zxdb1ilUo2DkFuxHsnydBOydf9OtPIUqXhtaLismSsRPXt+p6e6akyqz
vBKlaPgDJXaFs0UQGnkqIGtce8gO4ZN2MUsjqOJWMYBk8kiY11MA0ibumXOhum9z+3CmVcadMo0r
CqtNq9Y8O9YEpwoC9RhI0tP+DSZQnCwFYrPW4tBN2p4aXw5w9E9onC30sPrSABOlc6EePyOZBNIE
beohi/H6JQOli0aX7AzezINyNL52hJlMOoLyCpg5NLvE1XhfEkaXpmhvZdrLko2q38BUPRorSz3n
bO2d1eSRYK9eyHUPE4ptPTqQNeo9bzkrH32cMCkyYFEKo08jYlgouV3figgUYTCrpEhirGz/kXed
UY4+VD/lYaYLltLeDBU9MgGlCb/rJ0XnMN1EVcaRc3Ma+0g9bxCbGSfSV64AsFhCgCmIGk4aMqGx
XJNvSOgrQgUiuaj9J1mzqcthz2tGcVCxBXpVgWT7W2zgkn7dv6lZYvZQ9q6KTW4RyGQ1pAG35oAU
i2/YfuxXwabYBSGD0e58Ww1Wlj4yvjlIBVZ8Fucex9yLVC2M/I1UnCtHYXmfU7HRLlhB4LLqiq2m
ZoHdQxu2AmbprkkRLa8lqZr9eZin1wdIM+E5BXZVitamiYxPaPWNz3w4s7M2O+oFsQIJcyRZv7+4
WBU6G2YEFFMZ6hkVuAEEhjh2XFt02pKsn1lEkNT4uFcmikiIDGvclUaDWUk/+8Yp0WEY/Cd3VqYk
JNi1+sbln/amhPBFZKp/4ny+ekaaqMYO4bJO78tbNi9CySDcCNBq9uYDfvtBavmX+J2TM3+t9+pg
1VDSBK8LNVW+6RLA/KWu18Ct2svQQ8pOFGuuYNlZQgC43zAqwFe3QnpVdK7Vh/fKouTicw/zV8HG
tzqCvlPUX1vGwPZqFi5WcfAFGeRA1Dg/65v3ZQJpNsq5WgQKeuprfshls883NMFUcjP8kC7+w55A
+9rCzJCIPW1uPXP8fOiQveW/xSKyfQO67xN93qq3F8y4oeTJ2pGk3jJREJtlP/OZqEve0Ecnn6lq
M4KQCZXO0BoZwOfQZqPeIk73Im3YMpBoOVE+t5HDFeH7MGfTjrP/towXN+mOFZCUwHqZCHU8sjPj
zKV5xq9Td4+qkZRh9Gq7lD0xBNbtcPFs7Ty8UXdDWla+7z55hJlZspxc2cMeqz1exFgk0/3bRJ51
Qlue/RLl2cp+s6q14Xw3axPX/gCNJyfG96V1RoleZIihVXfxRo+MA2+Okw4T39i/VUEmqpuLcs2q
mKhozlhBlw9jzAuQ5ZCFQOmKwaQ9aTh3/exkY6jLqMss5EzrTJl8sIfWr9ESaZZGtIkP2aqiyio1
X9S7HWqgl4XOjAFPxrcorhP8fG+gLdOatE2+njkRnHMQNAyAPdaCx1OQGvSSQxXMilVTrUJBIaIp
fo8he8TLGhxM/ulP8apIky1Su4juMSvepAXIt45K014alaf5XYEmB/SUwH7QnVPKfiZYb1JSo4UR
fUi6EsyQZgqBYEbe5S2aJ7CYYRtHtY47US7QmwH1oN4bHzXAuDAJhP2NmhXUrl+zUH+HGDs2dkwW
bjxKwBnN344+WznEZBz5k1D+LbAg1qxZg02xTTvNTuhjMb3HpxJp/v5Atv13Gpoumoq8U9nECZSa
/u6WjbCMUXtK6GsJE6th7gJmH95/bz03IwDj4g2HfR7i82omQSWoMgvHTXszT/y3qlsDc2PL3xaF
CX2af7tN3vZe2roDoa+ITqvO4T9XMdDtuA8FagijY6erFATW9D5yfqAma354Px3csPIN9gSuf7x8
VwqjODBHreCu/wgUnDsCLIYZNwJIwkRPm56pgOUMnz37yZGljZYrCCa6VWlLSWlRgRI73R9i1Wzh
axUSv5mSLA66wylyJJtG5qOmRtam2UV2uywkqKUIaMjhfalJ69pASXIObY6yRKGV3a14PjSaa0aZ
vDz3vALISaLSRZ7M8BuUWu4I2Jbdx2E6kNGOsJ2mbnZItrd1gRgbCvzLvQYbM/qVSlwci78NnHr9
BCeBRR/+fHmQhGlQkas9VV8EvksF+7XX3AtVxF0IwCSSAz6/Ffjjn60OTcyfNJ4uV9T5YOQe0x0R
NW1SWKWDOcfgkMnktfMSY9fOpLeV6VUAZXrwnpf39FS0UTjmiQl+g6C+kRrMFQIM5nZy6nClNZyW
/L2AzkUv7wxSpB3is/6TKFo3YtJSx6gXPk5MIDKKj/Ukheb3Rfy++9kctgCpsW/ShK11Je+nJ/8i
MQceWTD3jY0SikfYkqHjqKO1TEAWL0yevcopX2nt1HT4gJ+ylgx0cM4WZ/o5mlr7UkXlmiBc8Zf+
TJI9Z+KjG1LPmdcQUeaQNPly14cNzc16v4ixHgXobHPyKVwRoNt8DI0lhFuLzx67c1Oy6INsYFv9
UM5/kEaZMyl3H3VFAr8IssomcpaJ2wU9a1io4Lq5mReyDXhvnbdPRAXyDS3meaSD54kxSgWMaFBt
SeglSv56xUf2r6gdzCDiuj7XoRVk1JoPlFAozblVosCBZ4ha4BTKH80/fzT3vlf6xM43HsBO/pi1
WBjj8LUE++UpObJ43B9EHpSY+XwAL1mPbj1oOKkOsOcF8iv2fWYXMjN0h44UIj1xkmqi0x3B0wnT
iqIfD1pOoEKMhcyRpm0AhqB8L2L29rgb9fBd34JddZPZnJes2E/Poxi1w57x5U5x9d9cQt5QKv3c
KLVESWT86p40dj9y+JQBeTipdFjH7Maara3i40a+mClMargCGbtrktPeANRS6ywx79FSvK9Qr3Vf
59T2KikEWiWLoQsP6KRuEVfPVdm6PEHhRqMo5ULT9s6UvfBMSEvy3DVrsGW6cX0iyivrIRApoWds
OcML+wH0vckhY0GAOx/C3Mx6qbVdbvdUPSBR1dYeBqzOsdKIebmIC9pVtwSHb4nWzdt/124QfMKz
2ULDYGH6N9E2i8mOuF6dA9VCm0zzymWhiN9FI5muhp/o7zJvWtG+O1CKAlVN7CT9UGBkzgXNh5QU
6X6XSDsTueAKtLNQRIXwJFp17eM1BFrzs3i2O3d+4p6spO/1sX9tyGzyjkH7dHB1lwvw95jLE//T
1N4Xva3NOO/qG0wwnLa5h6IlrZWmU925nUGJs5FtMTP8FZd3HE3IfOVlDPYEoFY+AEIEO6xP3TNa
GzNfgZ0LANbKXn6c7G/eoi1vfZb4ZUoCF6y0D/rqKq0dQDa7Dij9NET3nkxSgmR8acyjt4Bkun4L
edK5/+DRYtEivmJODJ6klU3xoUcl58lKhd08OrVQt+oeHhqa1gnmfniwTMdmQc5Fe7mlrGnTrdv9
Qg/rHbkcMI0JQ82Tn+rMnCk8DndjhWbHag9qQCc0/j3y9IBmXOzU+88B53hLBKodT296BlX1r7Uc
wCuf5OOVaGZOreH5ohR+32EtBNU6yS95d/nER8hB6yH5raovHFslk/pWAaYc9+ZcghFtxXoH4VAE
NCidCmJju1MG1GheUopdavc9qwTfo/wKEPqRy4Zq7I4jlqMecx+FK2G6HRIaKonlAPwnkiaPqikQ
CXM1b7LsgUpRqRcaT3H7TGPFv6Jk17Ua9Sie9Ceomg/2GT1V8Gk8cfUKyq4wINOkfsa+8V9xD0Di
63s068sl05EBLPQjqe548VipEnhRiVtbo5LGxiBWuguiqhA6DyAySRNAs/eQSQhKKe5KmL+/SJmv
jFCLJhmi88iyzgNuNyAl8GclfKZ6muoufjvx+4sIpn7AJcJfSysuZ73XMg9Ys4k7fBUAvB1CKeqN
N4dkTnhnukISOs7H+sV5T4bHNq1XiMu6sKb4IglCEle8lPFCsSzkDDEVD4XHcUj9PCrXmZdhlv1B
7a88091NwSohXkVTL70bUcWOdzwlRdKHFI/wq7qh/xNiCDujNNwf7OH4lobZIfKXq4XqxWK1ZKAO
VspofgF4nH0KdqzZnXQHFgVw5qSqjBIC+2f5EiDMRVR5VJl47lG9QhQ3PYcv2OPtqvr1hb/p4RSH
zTcISxSQu/C8GdQGiti6SpxDh9xYm4cStJaqXSPh4dUTEui1awj5uUV8EP+PpXh0/VqkfhSrqwfX
B8SxjjNcq2BeQfYE0jC/u1JbojodI0MHMDhXsNatU3qMmWMbz6+Y6E3GgbnVH4yj/8y/rEMW/c+g
IN+n4qXX74dKVaQt9azUbkd/hXl2Z1j9whJrquAF3Z6IkJdxDxj9z87RJsyCa84aSvEDFj4sZdKz
6GYjA1ZOa6i5bkkTgY/75/E/oI+zOCwu4yFw08VMIcu+fMU+SpQUgnzP5AelEHMii0GQdHJwUg44
64OKUFxCv7ylGuQyd63v7JhetfOYsw8bz3yhlBhmfitoTZN4/8Hk4sqD6mEFzrZtZwMGz/lrChbf
cWa/ZxzgIpuA4c7MTe/AzfcTjYnQ3EQmKiq6blmq7og/IK9rOaNnx9LAIR46vXE+RDQUk9ogt3+q
psQEMy4HorxEjC49J4PW3Mt6cllhKhVbFlt9Co2NiKcCUAwSHi48WANULKn1i5OEeUl7jzTMfovB
Wn4dB2kjyRzcG6Q9DFH9j8wwDmwz6SuK7VNQjUCd1OPln3YzeVQAFiUZ5HUKi06coVAHkRAcgOPN
dUw9KdwF60/LCsO0TL3ZdxwAKP8lUfaX/UnQjDSlcslPl10r1v1OibkH7LvScsYpg/y0TBiaGdcN
UT9iqvfyJJQFHz19xjE504STtrwOnM5V4w8RbX78D+7I71nI3tC2XWUgXcOVHRjMhldet41s8Cvj
UFyBm7MklJlXdrHAtKA3LxB0F9rVO5CBvNlUXNA+yuQIs7/8au8OhRerPysiHW1Qs17yo5dvM5id
8Gfk9I0=
`protect end_protected
