`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RsG60PnPR+fjG2NYmg7fxbmx3mPAjfuPq1NAQ654sl+5ZVpiFNqi5J8vVDUTh7SxulmJtapLbrXq
C9Y+RPyCrw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LlI6RcMouDios2m0ErNT2qZHZwbOjC4bxD2nva7mz0uhu1nLiHVCoFKwBIxaZDKWf7Y1pvbbmE5n
0Z65NVdj7IW+noR7UPlt5MWHsNqjq0VssLCcn/xNCYuXCfL5D1V7Xg+da6sMcMhHUFEaXaSAcboi
mlxo316c7KaQQlNMxW8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qvz5RqoJgjVXCx+EkjSYsR5IxJHJl79pj6PhAklqakqXQggZYJSNa2PQXH8d5d701AGCxI5gPR5O
Y+JoUEE8V4EiMgzO5nE0h7qKAMPVygl+ETVJnTtxENFYKyaVLdoUR106WPjCoYOUlh1hbOXV3CB7
C677hWF0bSmj6bxmctVNfH67PaY/aJ1EFKuEctz8hK3pOi6/qkBKRrJaR3BGDfgnbK+2oRDcLCFt
DDkWMqJj0te16zahUZ4zf6Vz5z4C26AvywIkGWtg3ZkyCqRXhDuQ2zwVxAcc4xHyOR8GMU6vL0yl
c5hfIXiIxHF+omQXoBBNVNwqnkDqCZiE8T9ZiQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0TdqttMiFGueyqz5adRq45agZAFQaqOSDqnrYesrgoyjsEbUQ0Kfbe00ye6ex6TDDeSkX4x6jz+s
0A9i5hcHmTl20nK6IIZ4v7G+FT7RgFl1QwWt08xGI2FX28p7x1YFX+LOdIqh6jcT/0Us2f7frBtY
uDw2lCS57SkpqgK2QOE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oCiutPVE/9DQhtu//ymudMkJggwZWFU1GThtJymmbdDEkRUvGctKw6YjdHNCn7iceKrDt/G2vlSJ
lShxdKHPZ0m8AtcWhOpw1j1e4qZ7MfSfhRRuIInjdLRHDCe9VpKWsnDDTnP0HuOw7xX4PXhb8o3Z
uJWz8ff4ABpiIyRB0L7o9v778NjjzfyEpOylXq3kKvy3wZlS7R2x4lKIufrQoDnMSomubnHU8iVT
xyVzvXEYC/v+GXwkWEmDIArIG9uOkrlKD7963MH7GxKiRl2nCKVxhTw6N127QXfJ9G3DKGSjWbFh
T1xP5OPoTLJpWhtt8AVC1K4ZAL44uFacmmwGpQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6640)
`protect data_block
NTb1fMByUWAoKNbYXO3kMd+Ba/Lmfvcu3bonU/PzI7apxf+zr+1C1oKqc7J7S0ZhVNUiT3K1nGMv
w1NhPyXa1wJrPBJcMm8606w7YMhB4UndJpeYmH3tD6IrxihyiKbKtZ+h7eFRbpAvtQcRffBme2Py
XIhbCiJLlfijsnMwKlcOZBZfriiKj5uvo/bFzL1AKcOFJkeAgIvLbFgPvkh0N/pL8hE2GKRgLRHj
eB/++WAqFR8G8bR8F0LPdceeZ05a0aOTrwqUrEUvstalJVH+/4UPNpHZ1cbpoibbKnw60PZPkhh+
kqqeu5WOi4rbHTnYSuR0evt7nXXFw/mO3jCdylQPDcxn5w5JKIixIhahQ5MBScXns7JLl1bd6MnC
vAHVTiTERTJNdmn0sHqRD4PgwnVnBqfHIDYH0XVZzq9DdCya6SMG6OQolaVwp0fRWx3Ukq8+VTj/
JGNGJlZSZRM6lY1a7Ho117G1b5y/0CI9gc8Y+wUHJknTg0cPa+iipDb133gjxx/2TYlSPojXsfO0
kedW4FR/FJbEnLM/e1Ipdf/GeivtpiGMirY8+IsKFiaRMAx4sa70Cub62FuKe6Syrp/MeROnoENl
klsFffp551vsyg4oMqdIJzx3Wb/77yGuSITbDYMA1gyw4OyIi9ygg20r7O4PAaLWL8KTRxbXCm2Q
kXv1B99zoP5TV5M5YWm+ByziNQ7KOTIwHSEsvlv8OiBR4LM6IqWMwWpZdkk3En8G47b/5FLVj1yY
/IdDqYVDZOesX6Z5bC3L7p7p86oq+kWa2DNEY6NLqHCrqj1PhWI2hJDW+/SoIM+lJJJx2tkbPPx6
m1Jz3bcXPPJuAhytp7gzV04pacIYNiFlnQ5a7BebgUQN850kDK2OegaseIgzf36Xn4EkDIrD4QJp
gpdcYQxAyLP61lcew/JxqPyq1ntD93OuFpYW39wqgoITGDnhnEy6dSGCKkr1RY6huS01upsOdK0P
8gKxa8kHyRH83EPQa6vMXzSZtjgoSrxBGTTKkCvJNfsM7JyEu5sf0wxHs/D+uTH9zo+xujfxyZoK
qxJcboPmP6QWpsJZZB1MimJxk39psM7CbaS8WRGZP4YcGfR4pGVwv77/lGSD+EZ79WssaCqYrNpS
3LNHZyH0fA5828oJm5NClIhzsDm9wV1U28lMUs06LA0Sw5UVr3In5hGvN9zmG0bDGK4/Apu8bKfb
ozjv+k43BU4UK/mTiuGGyTGGYZ6qe42CsnNkDgTzLaClxzbpfVxZ4AJLHHcA9k4hGyOxQL3kt4IP
V5W+jmm8jA6mToTyycA9ZMjjOADSf9F1rm2Qn9AZX1tgFTkX/Nas2Xt0dWRIDmjpXwdHdy/U2n8v
MVlHUIBC4f1TLAs3Z5AHax58BaXREN1HN4nzPSb/N2TK2SJpBl5q0zKddjSoK9QzXQaydtG1mv4A
vk39kSox7AGo/sBUCB8TVauSapun8i4qS9h3ahG3ztt/NOoogC5jAlveu7URiqnJP24axPCcP4Lz
1bEBLnJu+xKqlAx7ENEQ42TVA3P6QIx1SATnKfTqHX1SET6HDSR6gOf3zs3U4GXb8YmF+HI6jRMc
HoMN/X/Y5hWxc++kt8e4+LcScFoExfZ+xfFIRCPEHTVq3Qkn1OW87AvWIiCqgs+0BjphuZrigE4A
JObjT1lFpgsCMIJHhiq0MfpXJ970vhfvzO9xCfuK22LJ/bjlxS8Bw4ttVFPTi/BWPsoLoh981KeH
+DQbFoeStQYQo30xa+c1YAL847UPnmKsSOt09mTYOZG9EywGmhv2HaZTbXR1ZpECRbnyAA5PwYhx
WTJ5ONmor1HTU5st5FwDDQp/VunDOM6LBg/gjsgOjGobozj0MUcoIAZDrGdsB4aGkLGiXSACERve
oMV2wPJFgoGwrzAQyQBhB5867OJmwGFz+EzdCzqCd6HovlJpgG8yZQr/wD6XSwPNpv76vL1vJeax
1X+a3wMJ+mh/gfW8s3VEjWmBIWygI/VOv1E5cXo+OySB+BpzF0VwnjX9AXOCUdSaTtuwraq36cm3
ShdlUZEl0AuY96RrhdllTGDnjB05ku4yNnemkeL6VgvB5xEhpi2B+ncLbngK5LVu61Je8O8/3H2k
Eh+Q3MN0wSWoie8nkECSSTWfK00qb6uZfI2zZvxssZN7rU+2hXmd/a3vXZqFxZK9Fv4UIDxUq2P1
NHk2Y/vs6DlyQ1hpmDPhTNTxWZSGklPkQwkrvNY546o99EFkNxIYGtxCYbvYQ8EvXJpdwjS5p1TC
VV0IIUJCtLT/oQarFD7E+VmCcieCR7zbJKf/3DhHp8cIphiyuzrq11qlISM4GNRhX89bam3S65S3
2iTN2VpJexqtvGZIFRmaL0DiuTm+BJsjT2PGfjaPcEl4YFTXy3CDVQT+zvoZp2Nkm8A9tKUZrUKC
6Zka4GvJgxMcAj9uoLhCkre0De4bn0u5ITdgojMKfADzLEQ4BRBjYD8slp8/wbPFJCpU/m9hPCLw
oiNY5ObUdP+ri3vg9k/223NNpfzOstHtUeJUyhUQc00h9sflq8ooMP35yWWiEnTZRr49p5INj551
4QZo9GQK4AD0eg2MFbLPN63jV8uOmdC1bd1hwC8R0mzW8Opc3QF5lJgR/UAhU7l3A043MFFCr/e+
OVK/2vgyUkK0sJ0ecjwTw6F+hXbwEgj54XT5CozLziGugf4+n1cQlDDnRpZCIIRRUz2i+w5CWuKm
M6Mq/TkKR3x72lj8AFZQZ2c2gPwL3dRQsH+O0lCxLCAO4PwksVpfXtO5Ack+HgzYddPuyDKsdN4l
P11kqqqdTO+InmdkQ8K+YnL19sKDlZMhBzFdJ1vvq1sgCroFQTxKAcaP+yRpxtedmVTQABADc1EV
SJ/VXj3bhMNi1dM3/xT4G+NXLZPQXalXnGgZxJ7b/8rEA3ytufK0iccWjLDXVccKdLo+eKja1JVG
SWFuRgk1eddpoUX+LNbXgE1Q38vlN4cZ9fjDYaxVdGudui1Rtz93xKmTUyTIKpKgur+9B9qDkdvh
OCSNPc6XIC0uYwYhJ2hztTr7rw9XrebGhEM1I00O1xfchB8nbwnwZA0uSBT7b05Zg4mribH211PZ
+jlJnY5oZfkXkhSSV7BYl3uCqwdCfL20dN6OY/wzXlujgnEKh0b/E2cETRDT4/Xy7y8vYbN2mP3n
KEl8HhNBzHrc6DcCHqG6uAWA1oPIkWiTISW0+fDdHsBOnA3vrIcM4yTpp80Iuty3WxnGfPfjYf6h
X0bpBBSIc/RKt/iVnqaWAPYZ38cXQKotizUMSzneE7OVNOm/HSI31zCGvCXrPh/aiYex6NZmQmtT
Qn23tQx47h1wfs40haEULTnq03EnSrDOmZS2HLOWBWBbhQkYxei1GK3hX4+xEJNemzPGPpeHBf4Z
13FLwqzE+EJIkmEp6wYVxkfDl67quhakM1z/qxv5nm5otQLySEIrW3ISfRaOO4oj67/qL42IqBRb
jPTWpk5A4Z5SQqJLC48lvJpxqV5rLf3crOQmgMy+QkWaMntnZLYwbvOKFJt2ltMYqAx4OR4O17a1
mHUT13aRopiKYIRxKpSCdXEtfSFo59ricqmIi6Y5mFYVpz75jpOM8d3GJIsnHMxyPPsK7aI3Ini8
Ee8reVgD/illg8xYQ3yDfabQhT0l6B+XPPK4uViNDEP2wrouEfK4qqR9KfmugtfF4zZp0bYqyLiI
QtSAeKWzbKbOJ1meVYAn//lJvI5rUetdynWrgWH6TeM+hwdC2oFYBiJVE4i69VFtk57miEbafIQh
/C9FiZ/cUDVwCWvihJikbkFqUL8MGPR23MuDgtyLK9SEqs5d5yN9h+o/UVARa4nGXeLU6zAXbqqY
RLd9ojPgteXYBV7m4R7oB9216uxBpdacU0lSIBfeG8YmiIWw8Tv+ZfZld1gel1hibGGu22X3zJSi
R2sISFAgkI57R3t0DvLXaZIkm0XA3UHftgIxof664Obtq9tK8CpOhM1vYU+hyroVVxPQHgfA0275
xrOytkiuASwGtsJGHmrelMkjYqsfoLqRNievjdKzMfjfG51G1JmGugi/+RiQXCfpGBCTTGPBTMkv
SX8giTOvrePbsgBwDII3t2Ypu6HNgWzrR+bweAfzfjx6Rf/lk9WD0Z38lpFVvsRd6r/P2kYJifOj
2aE89U17S64Trxo69JWJJd0SDJdY8D/ETu0zbisa9pngOnGn/kREhpdjWBdt5mAzsKZh+Z72mMVy
dva714hCjOTSoQtmIDIPC7wFdD0tkxOSLTOTTvDoUUPoHtZadctZvOoX2KfbfpCdfkmlQEsxWKT7
C8K3865S28uUWXcDMzIS5s3NSoCm6dAuaymQcNoFH0AjsP4x5nmkMopd53GbsbLLl7aAxfjUjuWn
xOcno+fCQhdb/oqqqAHQHppzsskSIh43TsJnqIGM6LmeqhkpNild98GpamP7MQLOueEfGH2NjT1e
okdMzrjhjE4na7714tH4cFcVj8RlC+/9uTZ5DNzrMAwNLZEjhdA6aqOCV8gOigaIrN/fS25EuP4y
2v1RCa/27L8+0J5DrdeRkHQKr2JkBIEvaQ4xWF8AfBR/IjubU6SPuvg/a8eqheJsaUCaFLZqJ/fu
SCzYNm7AXrFGT0kalBqxdxh5C/knqF88M9Bhb0bc8o/GQtgkjjNIAFsYLlrWobMJzmeSjauBquy5
gjkLDIT+Auu6jy0iIosdxTwt6e3/FTwpWSzjQ1mMQkTj3fwYjHPct9uMFbC8LrVSAUndPvvUZ+ve
NdnnKN8JFXNtgypFSIt7l0as+ObR3sVH65RTQiV/fSxy37aRvqLGxEhU+SXfS49h14pKQd2Kjbcx
k19pQP6UppD4kifCfrmhqa6k/IL8XU7J56t8hVGXwIXC9eYgTkOcQDsIZXB0ezDPF2LIMkDU34H7
kBayhHsZ/s5KWu+lkkzpZwVnyPzHGzeOcEOuRg+MBtpixU9M5/4HkrkR4liFrJ5UsoIOGMRv3262
fleJ2XIwkbfy/A9D6qS/kcnwCXt7ppFPIflmtdPbBQQEEmyv8m9dyOKXzZSOKtWkzv+rfmALFkCO
i2HpwQ945ieOSrMWgSLkWhZe5QZT8B/qnqnxjp11ZDZrUW9kpnEq9Mz/FNOgXERK32OdljTTAweP
47jOAMjqBJ0/R12e857TXG+VoqNSVBdkh4XJyfAwVn4djJyojljCpEdXRIwQSdIQSHDOQDgt/MHN
wZFkBj7EUCV5VVoq7M98BxRYoDCgqP1l9VYZsVQe/cjBLfrOqnG0GetAIQpRza3LbBE5FAK+VoIT
7OqDpUKorLjcfrqXyx9TOwyumnTDxNygKBBtKsORYu//n3hCLAHoeo2RMx1KwlRO/1ojrpUxh0IM
FDXwSE6BhRRLAaJ7ZGkQcfZYY+AaXKOT8/y/rsXKlpSuM7CwUqWpq1C7KYkzV4kzeDzlLeN3oPGj
DcIjIiT2OPKr+s9qOPUDlx8etP5MFc5BXXYDl60DibJ2Q7Rd6F4h9a1h2VRnWZuUQD/Iuv19iGya
tLlLMJw8WQMYukPbyn5ahl6DhMykwx2nK8dZE6WOYdRj+OuPynUd6Q7DyTgZkIa7nf1xqnUfNy6W
AekmBu+Gj4mOJPZkRtth/vddpQHMwkPT0tkIvwDsj5bX05oNqOEwTi+yfgBRv18dFxXHM3/IAEG7
MXP7V+KhjEFk8WTkpzzUlEGSLUCwKMpflyRxpkM0oYUOBRmYgCR+SgCPChtM2JAx+LvZi/3qZdV3
hsWJsKPchvOnpRFMQtjnZ80E/uSejCqwQ3fhhtanPGSSxp9QQdrHsw3FO/zsBEuPnD5P1rFDrAKt
R8x6KUETcx022ZIVGBV3qncgaj0gLFGYZwDshb+pYoLexccPLfu7PMlxwECNs/BlgN2Gm8HhDaEk
WxaJFeS/QL2/t+dpLLhENV5F8yJzLWT5eMsRhK9WOPQHdnWLRifQZ0Kkc2PmF45YjqdG7xyf7Kcu
DvTtKorEETGqsJEJAH+TW9N7HRVWou6uKyt6w4LDpAK7U+MKSfqqWZY16/y5CCr2u6c6OWfFNz51
o4UGQZ+CpsVJQUCbASfbThM5lqgVSwBhHQefTBmo5yIthGWn+pg+GOYp7xkWuMPHL5Ly72I2NXhA
Szyg2byiUd0K6TYFYI+FOxr5gw3zEt3G/5KV3W45E4XZaxH+0i4dnMUmUbGm43q51/l0GgVioYIi
wBz3ZH4GYpN/+Yo1DY1BBG84EmJqD2s4pKuJG3Otq+URg7ZCuWOGzmBcViwBzARhnF9d3s+opzqQ
jdynnGi7f1bIqipEBJYiRQNHzlDTiu6D8Z29B4iHqWkFiSwi7aABMhXwR0cKhm/EEthX/ZjngQ5q
Sod7bVieuPpHhfP3Yjg3tP+BZ4vA3cfhFamIoBKR2Mumq/qtr69MyEo79cRF1nI4t0EYb8d+veTn
zPCIGvxNTGG6wTBMrMa3FqByaMRBV8Y1UKtpZYuiRu8RJyEjV4KSX2rRwF10LRQAMGhiHQm9IvdH
VfYpuAtVEeZs+cfeYp76OuIM+QTZpX9i3WmJsZ36x9827rQyy/26Js0DMmElbu0N18JZVyZmi4v/
Q8kToAhSY8D7biR5sUod0wqBe5V4khX5aQwoJED56q4h5IHgp8Z3IdzkPsY/aCbW3u61Gaf4rQVT
n6IdY6EcbKrdRd9ftCXewc59foy/8tIX9y8VeHVleirlGWC/4628LtlAJuGCHuGq8Pv48PzgV0Dc
JkE2/OL2oScEqmxl67q6eieZA4gZ+Z5oaTySpXFNM/D06t+BEz1BpLiQi1J0wk19NmtILZ4LAzyw
2eAPNBdnt0TlMo2xok+lxmUN+grXqhYQCJP2vVOdYe2UlBHzjLK5/NtE6y+/ODtJJX3MyG4WL8G1
mZ9X+htrhVFXVTafTAy/kQ9a36dK12QtXA4Edry84R2IbDPkwOQvsJ2eU6laQ2w6fMbR49o8tw/t
AyUN7JBYQmA8HAC+DgW1355Fg/7DMHAz1OqVgyXENLgPP4KMRaxNAzbvgUlkV62LKy1QfZtINOWu
OGuA2dZ366jITMwYkMVDtuVTbrxVAJEy38vQbkEm1PNKc+sN8SuuTOo/zQfLjKAxW8tGK/C2t1W/
hxEEBEW6fCaxV0iDbvanUH4tgqm3wRGvHfzOOk6anJDpjkGGYRrEetyiajiI7CaNODWLvaRZmYBA
on6vlynwwyRhJSFwHf0jch7GBC1s7mPfb5rbLzLwyPYqapDDXuwjsR3mjbwelAVxKUDz+z5nmVDL
mnBz1c7APPQPSkCutR9lgQpSZmhNRUK2ds9ibpqz1EPUlw/O7LPknSWFTyuZQitJg1uieBHNfD4Q
0Sz8myfLErCunORUdKLyPYW7qQQ3C8ZxDz2KhEz2HA2aA4uctVuUDQYN6yUCkPNt96PVkYgYpTU9
OlCFCNsSUD/Xka2We6BzQCzakFYv1yL2y6oDIKRwn26kpZ3rU5W2vqnDuTDVcZWEND4x3dqY7Ska
0B6PMHm/cO8DeaD3BYFfa/4dpyEcShRkIEXWe4PyymBGoBsMke3V0xDpO5swz4YEamBKhE6jJLz1
vxKftJJ5o6qhYCPQT1irnJKJkNAM3v0+WRjg8GLmKKS9jZvw0EOzj2hcv3WgZ6awWHQh3k7A4x47
GTghfnTdRd+N0C7UnmTtxRYpz4F/pLJvfYZb6PWJM1PP/jQWw4HnzlTqB/BAa7GMjJJ1L/m0s33s
2qvJ/SoS5kqN5CvSXEvW2QYBu5M8b8XISw/8a4VNugAxjSR3JrLL8KQAH47B2qhyst2Q8ZB/i11k
5/KAhSlx+lzJwvEXM4Y4w5j8Z/sYMfL8OEDzkKXFmgjww0zZZRvqey1T5A2y2XweBhfmHlDr9H/z
gmVCRxlS66JVZN13pVxayP6SRf5z7idU1Flip4WDWqradVik4mv9j3mBjzUvbm/FMlomu0+Fpn8+
tHo6RSgZjI7KytYXRPl45ktofi+h0EFBGime6Qooou05OLcHdL1dNBOe963B6aP+eozFT7PPmRgX
5f5Vk0UNXTQVJWB1pv7BdlqCTTCp4/B2yldj7ZuuD54/M6vFQ3sStxdzCP1u6R4I0e/ZBXU3gvFC
erPrMPyiotBG0I4jXbSfKSdEhGLWnB2Af/ezs7IOsg1t+s1IhpT3P561+tYS+/S7SRuhNTPLxqx0
Z8GApTvdI4SZ01Lhse74ABnE+dTL/ajpBbV0ghgE62Db2ySx0Y31Sr6QQKSjNnjbrJjhaujgyk7w
8Qn1btaOdAOSao61uXEXCWQt8M+4m6elg3WMk4tPAJ2xCxnO/FJ6e2rGuPAPf1uWJXE4NjzaBiyo
8Po/FlH836E7qO7G86Pt5hWN9oVo7JVNf2WOJsAoe1/MGf5q3OJ0IJcuevtcHFk/0v28CaO8S15l
+WaiJ06yFEOiBgf+alFXlruyxeIhWIGuuOFolRaU+I2buxAlodibvq7V3xVlBRKQWfpbFjIAcJ8j
FF4rzUbXbbUbXzUcUE6RN4pGD/oMc27pNYVKo/lGemUNKSAjq/t3zBHQca+xHByT2XL0pnMPyRyd
iqFT1mhXb8HINc48yrKHlshRsnheSOyLmvkmKzgXdTITNlHwmHkJd0vehVj05BXvbCXCqUy2tqDF
MpkAwswzulU674CXh26dXctReqqc7vUXZfaSFQI0LYqklT++5QfdaQm0+bopFJfSG10g7ylTemeU
YjUFxiKc/4O7wf4fEz3qjReZcEWXF4Pu4lNDL0Y3UBx7/Y/vRybWTpBhliVFjM7cjp315+pgWCLm
aigrqYO0zj7pi8HArKdvD7iCZM64TzmZFlZnBw==
`protect end_protected
