`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GGEdS9Pi7MLJxBTcDN9C5AjQJ5qNPq/VYl1vIRZAuTRezix3jresRizOOYoZtQoddkrIyj1KLx6j
1H8H5lIa3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J53wVJ0BT4U8EW5aw8aDy403OSY/NdYKHsXgTxyKZExrCRuxGQUG3REJlJ0OZe9hk9Z4cHosBwcf
T6lWWe7gGg8pNY83bGPBmajQS2N1/uQmv5lyfeIo2Bptq6ezqgqYW7Qud1kLENiNWol214kCTk6n
CVb6lnm8bCi38IAmc34=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rS7fIuclhHntjWuxfdNwERfMdRaspcCGH+NGRJJJlZcFbsy6DlE8p+3T3q5ivtdeFuxYgHjI8Vqn
ZMkz6zNKaciGEy8UBsps9L4h7c/unSqUwWaCiwmgrmNn0oDwqMlaz4HEUF04B0+3DYCuEhKBORXR
C+pAMsBbFrINzDJ5rBO8mFTTsIlj3/qRK1bud331FEhPvgV0hraXUIVCuO2MPw3VDGaTwDC9aIag
/njvvDMUjY1e6YFPc3PKjTwBBzG08lQvPYAGbrDDFW+sdGHxPXCVbns7oweH81baT369yBxguezC
bRpqn/Omz2a9N/2SCxgeAQecFob/uGGijii7WQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4EQoHLxFvhKGMZBY1DwaQ+mYJ2osIRk1rq7R6pp0JQ8G6Tw1Chwov3oCKZEm995TWi4AyD6vNOjL
XccAUz+hHpRvE60DLF61TdneDOsjZbd3L2NYwPwg5S5AJ7ZrnTJwAVYwvFlzhW131tm/lurPq0Sz
8df0btXRylGQdpptJbo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AxERoGEMba482M0C8sy3EKLcFl069KmT5qDaJvThv4E3gFb0sCRDhBzQjiHiO9CRsB6zBsdyeU3w
Y6fgDE9YYC0V0pTV9ZsG7c7zJ2PLwK16NhLbcG676xDjQndf9jPtlo2Pw5rqpo/oGRJTSGLVs32R
11Q6RlxpXviJ5RhtaKGyKHQB8u1MBEnTEXMJrP5yJOlRTtAEDCicg71rAIgHTsep3LjmeIbmoXGB
sfB25uvZjfeV8jFOx942z68+0Bggulirrc0nl3ermhlaR1Xgbj5lFqbZssYgngGjd2tfdI4/WR/P
aOwZkVJkuayTsVEBE2Unb+GH+XD51oao/zeNCA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35776)
`protect data_block
Kjw17PAtobpF5df+12GWE8KhTyUys2i2wi0lvOfOy/iXYBvWHPJWXUuChtZYDnDSRRfjLD/meUWq
o0kKqvCrGdG59fqbB3+8ZH1QDSphqj++Bqk5aMyjWF078UFY9StI7YSToDI9B12Nh6ImE0e8qtgZ
7JfJBB+QleAZjKisXHxYUK67J/820L3PeREF0Tdg8Af8GxFBDvL/BNDaVm0yN8EBJgahnuagJp7j
eSR89deiZtNryIfYi5/7v4RQn/L94Jc+ilhJ/2qPqmvXbdI/C/sioKhYeK1fWHuPiPKNKxLbaFK2
wZ+a7PjsyTBKseLv3ONaaHfzNE4GZ0gZG3wZHbpqovwuLgRoHcRK9e0asbPoqL45MKZiBmCut5j2
TXLSTscxt5ytKOB8pQPrBxuA+CYwuffvA/NKsPs5Wy6G4Fs2q+hHxfxAiZuASidsPshZ4M0fES5s
VyNHdfwzDSIXpdAEppgsG4qMvT/ZZKrn0ph0KHET51DcERT5AhcmDPxCSHWUEjiVdle4lViH0/x+
yTRD1xnOV95bVdnyBtTfNjSOc9bOa/RfPy9QNXAckGNVJX0+UX7iQgbh9OzmGeFBdyPuDY4ZSTcY
VaeCnz2sy3uXgXKxN6BlFHpVZUWn299zEJk9B7taCHKmq3MrI72DOPf9USv2+jW1BdOmbetVFtUR
6VqHmHJD2r2WJT8wmnbpd90co0x000S+f9kw0ezgEhkOyyma/EEo3/UkCofLU13D2Wv829Org79D
46FrFV5NkBckj0MrPvbQfzrJtfeFSGOP0729gny/2MzDUptrEkXL5TLdNR+UkVz5U5RRKfPJBIMj
GOU7H/udL2bmlDqmExRj0lx8TSXUvGn5epP3tqJYlk+qjCIkTMreg4RDfpP3+UZmhOcTTc2odvIP
4OlIFcMo9fJYmNaQoxT2fY8Xsn+JwB7K9KPpmveOmG05DCeazMFoFf8GWcT+ZATKPJ2i4TR57iCT
Wo20bAOA/AA+8Ml1tE0qR4n8P3fWa4Jakgffh1XMwBmgLtB/wQmMp3GOdGA5AEzSj0Qzc1jvjVEz
syJbOMoiEidAmQHYl058WYhjyS73L2REFiTNpIFAyLPhXijWFXAO0ZkOJ9IFPIqRHLr17omkVSey
dZrAMIAXnRAI9kyd2h5KMQ1ue0jakoh46OMrwq7XJfwD42mifDInFdmqTPs51T/xeYMEHMnE1yPK
zvRf9d2A5++e0Chl663o2Mqs1RaEjx6nMRC5Nb/KlDlAi+P9dU9Le9qU/AWhkq5oCQ9YHYeTqIU5
CoDBPPkcNncAKHjJUoIsfVkU2f625iX6/D12decsPZ/1hPOVNFpqd3grX1/K/EZqzq9vQ3Mtwbtw
5G148uwAsW6ENWRHu5E5tJj1g47BYFbBpEAPvugJw9kBfkymhhUr9z17xKlguvo+lKSS6hBipXnT
FCRh8kes9CI25OUNBiAn2l4G2qfyKqLNYFQMgyZCj4x9np/SP6fZBIGfmxkNgxtSi2VzYR/Tfkd1
iZO4VPkEDGoqG2ivFMFLFJgH4t4kHzoEME0Wfl38PAKAWHVYtLi1Q7C3XcH3r8c4VPuym1F6Ew7c
l7N9UXYPvXCFsyLjQ2PtPow4xvwmPtzJP+PWvUoNGD5b0Im0CQsnuQO5LoSNb+cjwI6xFvDfs8De
1dyAB8DQow4ODQDqEZKKw3zlzjn6xbPhDSBYhTgTqjPF2f6Qxu4r/B96uq5M/75U7FGlPgbjwDuI
0MKtTyGVY4kES1kAeoI3DdEuyUaLELDp5qgZUkdFU9MO8QEQXL+EpNfBs+tlbNHiUfrza06Ou0TG
YmNoaOpajgPVxVHfWAkIpizc/BZ5wpfdz8PJCfvx8nN8tM5mYotZwquv/V6lMpPbLCnTSsrb9UlE
RMHRQZslrCP3bRfcyOzbkxYz+U9az66T3MtPo3hCE2/0vqkZIWa1uiiSWBHLoW0SEkNqo5jX+M6H
Tfby2YdNtApwCVEFJOHwDeQylkOsLRTVISr3nUs0svGPer29bU5dVyBiQWoCIdVwGcolFiOzEeTH
Uh8L+WqBkTxrMvVzaekjGhw7g82gjsioQ4hNnGQl8+EukNLu/64EaBrcprrPgnm03Xza1qN8Xy94
bQqTXDxCM9rWoCZHrTB52RfiQYeZFT0bK8uJEwJfD7TPccB76g5EN2cw2mKVLEWFv4PJWwKBktS2
dmAfQsF8gC+7LDfQT6Z20URsvIMOfHFvF83zg7ea9iKxbfP4EFXWk8bPmoV9CDU3z5gZaAasYxAv
TKDwh3yohiXpDu8ZRdTuF44B2amPeVf5LINdLObJt7c1+FbE6mxeb+aMzMAsk8ppdoRKDAx56vH8
SzyYwxw8Wro1pOCofC/8OrKL7yfbIr1B2ogxjKFoJE5kzlsdwaPVGS9GctaWS5RvI3FStzpizH9t
Ok2CCUr3SEV1DiwY5+P1VtAz1quuiSENDdJcOJjtrGjrM78CM0sR+rexyr1NpPJI8YrNQ1itSR45
bYulbyMNCiErKLwFMF3oeOzRbmyWDGtYTNPcUTFFqaqQO+35heSj6z8mUc/Lc6/wJDBTl7Kh6wPm
wFX5EVRnlQSXwvWw0zR/ypIhdPq5yeYVtvqt5mlOyijj/PJtc6IHGfsxWbCDQ9QuYrGvdYprtOp6
VzOc281W0j8XS6sJHP1bYu6LUB776s0mh886+qXNWrJXJlHlCvI0le5roU7JPSTSID01pvMLZ+wX
OFEi+Ebn/eiu5ihudeVfCFmtRVv4sPLv5S12WMHdbMgHdQRkcBLggRszFSU1Q1SCcTchxzUSGMkH
/ado+DKDt7DWVFACQHLGWEVr7vF/w1h6uNZSuu8pOFDJgrPbvS+FzZG3HJbO4fHzbMNgXnbEUZG6
NGCsxK9F9hhdcE7a8mY+HkmMpI06J9SQm+dVltrvpWuNKwVRQZyOdq3cWE+V/xf/MUTknIK/0v7f
5nWGB6NjFwiRclJgAf4Hl97O4ySFAUcIsALj4EX6f/x2rC5H5MHtHBuQaBvQflnfNDonyN7VPx9v
+ScXNexCo2jWk6mmygGH+OIU9ape33WJ35knneHAkCL0QZfD1P6pV8odHBA1+N1FRwQEJWKyKdZA
IfOdf60GwPrRay2xkRTs92V1z+2urk72KotQGZtiE2r2YLRSWMQdP80hH6LzRHdNxixJCI6jOM2/
vzaiFKlQjRjgEPnwdY/jHAh+O9636EMET4I2u0dxEvbw4ZVGSY0hB4lLmdPo6yKa/W3e2IKIfzqj
EeMje7OCWD5hrFfCeVeXf/lYqUrwC8PzNat2Nc0uGahCFClRZE5Sb9tT6zfBEcbYznlLFTMGn985
pt44EclzQbTzd5G+dpk1q40QF9qDP1A2H8w8tiFdX0nJM1h0HSuqNVtZjHHnD/abeJiuhxSvMNx4
g1gGznIYLu2k2kDS3TvTvhlrDsDBySxEizRMeb5X4lOY/VQdMf7BnNjyrwgzpwUU8FKo3n71/V6/
L/fuxDHzERBYoGryUonl1IVvSJQjsG7ltr8WqOCSUP2yGJsLJKk+w4XmnPjyE1tryJGDjIoQxaZI
PzXz4q+mZjONMhE1ff4xL7Hz6iOablmXpE+nWJC0CBNedURoDPLjjomuOeIEDU3pBhf++SFKx2xG
8BQNXDiYDGzqZVaeIVMVgkO6rk/FPyUlVk34vCP+I69lKAVBWSlWFzgmsrYj69182b6/GEqtFVxk
Jcg68CSAKFFcQtrIDfdGeogub3Od9lQxCFtX9rh5Mtej0zjTPzSgiq3uTdpPitR1APiAN9GgaZVT
aGOWySUstfj5FhrYGMj95ChcajBvk/FBqz4rAVg64+jcnE3zJRm0xGEf+dL16R1AWVIPc4lMIYlI
7gXOQae6KqO4W/B148JIH+3YxVKlDCX3vyQkmG3qdm0LjTkDL9xdQEstM7SNAeOgY+oiNUqVDq8x
NMu+rVKZEoTJLcPf4QwqF2H19WF/cZsIOqsTWBqt0DbaCfv/bWJ6jttTp6ayFO8byJqNooZ8bAP7
HfXSLvy14UsThe3kJk+1Si5AN4s5SVo1/811dqRfs1gg8EcKY5reERetmdb2v4j+jqQWbl3v8C94
LKDaQS81uXkTPH4mDMCTe6ID9/yfXaEgydaKNpn8qR1lg08swkDODe4kuwn9230zL6W8t0XJsOPy
KtFsKzGW0f4Ey9opa37XzlHXL097PjUcuDs5zPlBmjeoFJrYNfXVojW0ZFX6F9OesacKia8dDnnQ
kFKY8yjam3c87z31OnfWVkTOgz23i+d8Jqp3FRxOrTPeSw1LDUzvxx2/iDued/86GPV7QowQuMX4
fe8pUxTBMoB1XMbtAzghU/kI56aTsy1iTPurhGsYZA0CT/elpBC4DwG+myj6eAV3iPJ2l9WrkD+T
cLKqPr3XNsOLWSBUeoRLVPLO+wiUVMzGM7VbifrU72gtiCsjpDTbtIamMVds8LNnqxL3ahJeQfn8
LxnQYWiTZKiF+6nHiiCHb/f2ifJamb3aSizMMa9CW7ovf96jSHNoF4URLe35s/mN0DYkth+CFSyN
GPEgC395UhRbtM70tFuyRA9A2et4EAtQvC5/iaq20YMQsVS3lYQAvLc/7/apCZoKSnRJuM2QT69M
gBfXrwRb69GCX9QNghP0UHGSeTAhCAErBZBxpnn6TKMm6sKc9Jp6uOQ5g4VW4HtcJh1w8Ehpz5VB
hxsKmweih98QBsJbg0z06ECv1hLNs/39ffpVhJaXACDHi3OM4bhDJAEar5M2YAlKjglz0zvtTihb
9O1k2XvUiUMzocmqksLqsugoL9w3TD1AhYZoBsnIc489SdiEjZSO4BGV9W6Q/oytjGG53jw1bJjt
lafUaFWRbn8R5lqNeKwdz8Kdz1MAwoiOFYrdCRi1GSdHKHIojqDCE2z/MVVUCaYmTXX/xJeQ2Fys
DUTN+mqv/ACmNwrSPw61UNwIxQ7EGEwCejhZK+q007zv33wX3wvj+BebFq/QmGxvjY2r/r55vxmc
43aSB6qwtTu0s5/Y1uTbBqSZHtcSwpjx1ABsXGSi7/jn5cY2bctyMb2qLHP1+gtNcSnB4Fl8HvCQ
eyxuwFUlktsQq524vNuayZyxa0q6kxcTsPJTMWgZZAHNw0kaFS+JOEiDRxm1SxMkQ2AHEW6KSim8
AQ+hQRUJC3YaPGQNDLbAAATdrDiAp/HOM6bdtDZmUUMc0WvMnF0nmCp09dm7f5qOagxwazmMyElI
c/88p+dAhRmd83uzBhMqy5kWDP9v0h4hr9AyQqUWNnFwsZCXPm5dQ+uu3zq2kaDRlhxN9SlxNyCM
ZlvpHFJnH5S04/KSyXLLgm3zH5QKV00S3aJNyMKOicwFfNzWxm82JJ1UcJzpw3dqGcHd9Czhzivz
vG7V7yVWLxsA9pwno1qqP3J2fldTWaNayplaf2VVizgBbIo8n26EXRB3kGIZaTa/f7hiIW3dNYS8
jKm0I8ej3bBwLuFAwBdDV5beAu+SEiuNlXxDdo6fvEFoIfU2zIisBxwWd/rzmwhA/C2D9DW0Q09R
0PD9Q90YhfIQYEGqsOlvwJVQqKt0WjiUBcVz7PBU10WNOHb/+5SDjcOk7Tx+2otceI1XwoahieJt
G0dfyqqJjt/OG5w2apjWhVesJCJGgYdV/cjbjASQfvY/ACaQutvkEMca0RevnU+hA6NGaH6BHbOR
fsalxaYWPyHU3UKr+LNwqCUplpDTH8NAAv4/uT+/Gv+bC3oJY+vSqJxPNbLepOnOTypOMJiXKho5
ET1CMrqEezbPnQiKiXxIr/0PLjNfGt8j3zTUo4A9RcWH0qez/41t8clB4Slkk4P4YS2btnJrZo9R
VpxYT3nDP6zekI8Q1c6aGaTbD5V3WQrUkmnMODFfc1tXbTd+5jkaLxSqXH6ykdP/LOhFKey/Bpym
lJU9PuFNAAAuo7ht6onKEyMV1SmvRjp5JqunNjDYhSmnACrBe53byQqPssmfMYuTqjm/gzLvPfuv
JshjbyhCGBFtRtnspG7BZwgeA1bVHrgz0lPcSmQYBrf4DZdXHIfFXOksM3wPe5/YftvO/dM7XQDV
6WIV5c2SmPqK+OqKf+1EXcXoxwnm/vg6qdGeaBjkkqRlJ0hlY5W6F8uTrzjohI8i/Zfo1PQZNEdt
p+rkWc9YJJXBpdYnbct+9zRge306FkM2Ls3drDz7VQezGAddNMnZHk4AuvwXenh69ZLm0EMaHgnk
oxeXsi8g4SCugMs70oJbPMsSNcbT8mgYAmUDTHUP3U+YlgSFKInpy3/B06mLIcN7RvC57qFO1CPm
oQ8+XqfciCVWxBOatAqiZeT28KIqqkctDQT3jMGro0hfHvrum/9/lHn5kVLxFrQzUVDwltr/kxev
rDI6o7nJXeIhq+P+2IWMXBfpaS3Ll4YeRQIBlEChP/e7X/q6x4diwvDE7++R4vClgvKsW5jcBhIk
3M56Rah8IuYHlVtA90CZ8aPwY/gA4FBy/6EVEl3RjMYhuSAixIb5PcmtU5yZ8y5GbcF1RIFBgCex
vP7M3b92poLuYzgKUpV8tRkkpmZ2P7H/sOSvyk+WWOoleblc7h3/HXjQFiJHzMOwHUAMuSr2UZgU
y6NrsL9U7ACRaWUMaNR2kKB/LF9Uve1K3rNVxsBmRoWyaKMFz1eSrEnddxPAMRU3o9WPXRTX/WDQ
7sETIgY425Qn1hmclRRmUpoeh8eQMGAacy5mKWIKOhDlYc51tnozIJtKMwQlzcf4Iq47o8XBjr99
Nu4ZXw9X+mN6qQcnxyC2Ote78UgPyrpEvDmCKJtVXb49TqUMwB+0nwrMBB/xlJGJnJ4YSiEVgZLt
7KQF+MIYfJLVF8uzLk9Md9t6nAFBnjXnzqgiVa7B49g602cEwGcItIMIxiRBCYaJ+l7fei9s/ao/
S818qkT7sj2jlCnCOHvRNBdI9n+y4kiGaUDkUsHi9OSjFnOCJWYaqz57EfKU2bxGZ8xgpaHgMYPr
uCi2/za4yIPXbw0fTLuI31RoSODSuxVE6GTTy7Z72wbdbPJXC5rv7Qr6HHy0TJdynFS9LMuf1hPW
HKpBG4nzA6m9miDnZv6Er/AE9XH3gX1F1dRjhwJmo4GaYXXAWVyHKI0mNL+vcMVg86EtVjSELb22
T8+AqhVZWlhB2SUDD0KcqVFGoUBAPoLDm5eiOFFmJd1mDr4IYqkf8R/qT/jUfN0TXv6WgF9ImDWY
7OqTZ/HPdeMJyxC+0iccxGxBeN1TpilVBlza3+/dAsmaljJn1izmPS/qG4xiFbc+eoeJswBMe6e1
5l7IGOpRZnqdxOgvhMYpQrPTzzdcbcnLBf8sD8MJo/2cwBWB1DjpICXLQqy4hyjcWqgNPhFZw5Lh
BBa2KyU+pEsKZKS8gAhc5WwhoFemNNVrn9CrL6vP1iClCVjcOeOgYhEW3TzFrRICwDhkqx8pQqjq
Z8v3zWc1qQlCdgC7h+ZiQrUljXToMzTpIm7Wset+Te1C7nPcLGz9mZ1rW9HbmNY/QTsK5rxzRpq4
wG0cK9/K+HYyQpb3Q33To5/gIpm4fX39ikgFy6Cpl+ro+PrFOdEt7GWeTweCyYHUEZXD1kAhIvDU
2l2iidY20imEdR/BfkFJwZ3Sd0u/oWILa+xSm3VG/8WhsFFaMwUlwsrbiZewjF+5U1cFcq2U3wvp
3U9cb4yo9zBDyp6UZZ50hidErVwmx8MIYqyyX7Yh2dyMHRvDzbaUicBjVHZTmO2kP6rShSytAaSE
cdg3jHsVwN8Wqk9AyisVia5C4iuNAavatJsnCzHa/EHbXLLi8IL5HT04OJ76UG5/zW83rMKYrNM+
uPQ0oHR1K3vYn/nW8o/0iVU35yiB2DYUhAWKi3T43dn3RpDTtAEFGXDR3w6z7x7iL3SMRqJwLqSF
fpUn2O1BQuW4NimptHqWPHYEaODYh90qJJyZujOFpUx/2kGqywJC19VPtML8CUyjjJGVf6Jst0A6
/sqkKzGrLCLRJs2qHvEfIUou8+u+vzWjJyHVZT8EVLP1J73HcTFuxM7nXD7tsYiE9yA+vQIxrIMS
2ZP5HocV6o19CmDhhs6C0noW5/JKL0RERsTZ1Zox5ZrOdLaT7zzB+yPjiiPzPz9yLR7Lrz+AHwQd
BdU2kUlpNIDUPuItQP/RbJwY1T/9r+6hV5C+vVPgHMQxZeHZ87WgHMEC3MlSnNnUqvchSOL8OPLm
ouEc8KEP4KZ8LWcGn0pGSn7WZtIAnX+o7FBn26GxRpAZPlSTmuCPPYIW5ObEszRqbnM0S8s9ziJ6
v8KO0fJHtf4/8BwcYUn/ltn1PiMIZafK5G4kiGY7n/+eGY9os5jpCZTaf3s4Z28KnRJ42ZcF0S/C
bd55fB5bN+pRcS1Eq/uLnVsUXR9WgNtU5u+GeX0N+jyt7VaRxcLCMZBG92IY67LG3l7ShO3MizWG
usHbIUtrlTyoVOD2NZOeeTZYjlU4ziHjwpt8IVkOJqXi8IzvZeMLn5IZxFSc40FDDFt7WqhGsq1g
7aQ5cO4w9k7/32yHT0bIUHgZVcoij6IWMHlTwXqKJFPNPOuHPrMbFojKEZpNh/mK8kHY/Z+COFGE
VrFGaQ+bX3epH9LLWgpS2bOh4CmbmyLo98m95jkxb6uJk6KQGEVH9XEjdFya9AkN7/nKw7eFPG8P
RfJljwrKXHY2G3O0ic/e5sWW2ceP9wgQIiS8WuNZdDU4kSGCL1w8DEOde6dCEZIBVe8TeJ46KZL/
1GJXQi7wXYwr3dqBnFWA4847YMnEve5ZwJS4NjMCCp/cjVhF2dwTRNUPTIjFEdfUaPt6xEZjsGmH
NSUy7PK631C9BpITe5b0OenU6tdAC7tMKymHCskqRUYQBA8/Z2k2cgh6wZgmw1r3uaHbifOP7puO
6JgsUA36WJlX2/ThgmiLgcRSKZ5V3ctqeNaw+7F3MbsIkPhr9Z6ITlWA4HxIFwAxZCIQSlElAdFF
geHRwzCbGN94+qHrmm97v2WENjsNTctKvyBkSwSqSC6Cfjes01gaDJfZH2OmRV3M7DjnkakhlUGN
pTyLKoEa+eVTk+KUMkgDOvefWuvukBtWNCj2+CrPq+bmBkXRaA79ZKgDVx0tyiEPpz7Iqx1+subE
c94fI9yTVzE5k5e0d8KtGP3Rnr1gfsnXNms5SQXusTXU4Bn29eUtrKiewia8hDq9IPiDcP21OqKH
EuTKlUysQSxpsAY6ZjEtD2STJwStcGw3A1eXzxGXj2iGTy6l/GfTjkU+owHT3jfr3T8Ww9lMmhpp
V9Zu/KAN/nXx2qDLuEgcpWJnFxOcY+okv5/HWli9P19NLxdfFLSnAlWDS0K7lyTWVkFFg8V1iLTv
6q1IopkDCeoiLmHAI5YvZQBp/skHHLhKB2laJB3ICjGatIqMho5fl8piLXo1eWo6hi2A3A3c3u6s
abMSBg4vcalkcIAD1mA1EgmOX9SuiWDO0XaXasDwdSqYyap3uTpyxDVfquaxPk6oJrBR/dP59/uP
H8ilNEKHlOopR7611dj/ER7XtCXlrBCSfKp5cwXYXhMMycgrc0j9udMi+rgzjgqYG6lb94aRj46a
CPsjOb96jV2pFxzf1NjOpvRmEblYTe+xVhZ6xlZEyt9SghFFTJPFA4CniBmis6w5vc5TKEg/8RZA
S3tZDfvQ0J/7P6YeIfvojU7+Awur6JfVieeSFtrwWwftBq5Z+nOnPDpI6H/JkfAMqQgalS46tqkG
TSv17BnB0SWW1Cb+VjMIrRlTp8uc9XapJBg8e6+VUysw+AnL5ImI6lIpxq0ZuJ+A8bkkwZY8/yOT
rbbvLF0bbacPBNlN/esc7cK9ZaI2snoxrBHb1jz3w8AOSYxu6ZliaoFaudlFpTVaeEbcky2qyKbR
/swTgfjCO2hf2Jz/kvZQXyn5JRAginmJ5kzSn52hV6Y8J0tXqWUk5EfHVeKTMWN6i8FI3fBH76Hx
t/i4DUmTkOodKZVgD0ZZJz8X7EUDJ/JGOKvKGL6Ki/lxVZDUC9X/bHiTCZ/i8PXJBYX+QnIuySKI
k5mPis649SjPZPe1wHCs4tIxwOmWDi3KSAfVl5R4/v0+ipf/uUb56+J0o9lu3nUnkSx657n8JByC
aK7nWaaPktQSlxABw8spEfbyX9okDDq7QCqL9Ap7X9D1DoyUb2JwI6pB6sUznAVdfhPL7s6wXEEG
Ap0Xcbf2LX2kesxDjEWss7AJbS91Ci/tNu2OJ4EFWzrlL91JPPw5QJuGqp7jfeITPJZGiHI/2fs+
4dKR8y9FN8teMXsIEnszFdGYwYIGcQ7MBrHrBjtN0AJ5544ICVVJoTONe88upLk4DPqiHCoF1cBb
veRKEc7fDJ0fykOxE/IAs7EyySvFcznsX6vjxiYq/LBrsdZAdmfSh39x+0LQ6vAbKG/f33zm/kRJ
JFgZMXOFSMaBaVASgB7PmmQqX04jbLgaj8pODGH1gj6tmi8+NiGh0rEd0xnSk98bYnntyBM2g2T8
kFdWo6FXXH4jx9BuS3pMekyMBluRRFVpjHHz72mR1bHWLYRmhBoNXeO9qgYBx2SkNKJAweiXa3Ct
E75kGLX2HHzwxVxlXHSzgPnmggP2LJ0t0KmCde3i7BUKw51ge1ptJ35tMAKjY4yhnC3YnrucP7Wu
0l9hsI5bYePBgiue4Xeif8y17czjPq1+f8xvOgPuX8BdjENEua+LTV0T6rhUlVDYme8DHDAsbXu6
QZH8rkFy94PZ89SMfQ8U8f/LgOSlQVOppqE/n7xitquEUYm8VDUAqYx1x1f4RqmSnHXUotJw9asX
YxD6IFSf9JtYTohfIS/s5Zfe0cEhfqxwu+pBmEYttipdwrp/MTTb0Jvbrj2/5TW+W8FcZSc+vsn8
0GMt/GYi/NN6XGwCHKapfmdVF/mrWAhm9f2TTDHlJIRoiv2w9G28M2sDPl6i/BOf/kBxruTVPq5x
6Ytg4Dt2oYq6f8rDbta9tHtL8kSkNfU6NiyBlYIfH1ddZFuonlbDkYNoTGcgLhI2nvsd+0LDM2nc
ns1c7o7jRHe3Hv/i4CrwvjpRgzmY5P+FTS4MGXfmNrAieCytz0nn0wVZaF2iQ5yo722THslm+XiJ
2frHZe6uaYq2l0d+XUlp1lZQVEoDhulNZCRqr09ul1C6BZqOp1fxNJVC2rtM+HG0gNFllsdZ59oE
N7kycG43AqLRRk7T0F989yaxSfSrsr6xcs9BjIliaR/PwWmxavyw9LSCje7Eb3z7AHKkQVO08PJw
srPZ/Hc+3IwjULP3nD82XgVpQGo5HZs7GhGpRoA8/qP3g6O96nWvoi3npA4ndBUIICNCf+Ub3Y/w
LJbYO9lQ1JTL0sCTTzgk/r836/JJW7nDNPXQ1CUISWpsACYkkT/hXNkUwflTAKVU9++wrH+zOmg6
8keupGXei6O+u/+RSvYlv2bL7+AME4RPvKskfOZTPSZNdMFmee1vkOg91aSZEYFSLCo7h6Ral2WI
fCtJVWM1tSpYMyHZpEWdg1oqe2cEoUAC0a8ppfZPe+WtUVV77uLglcHOsGuYEfZyDo/+5ucHF68g
A50GMsNwYAzrAbjQXaCMNvqyvleLrpYzgzLn070kwZTA+jvoZkwcpfch+MmxFnJ8J9yxNeKA4LuW
kzmJ5PLdmOXGQ5wkakXrXXj4PWRFHP2cMt6Tevwt25iGl4Jre60+C7dzlOYc/iakEj0I7H1/03St
T0oBti7T5YedL1E9O6t2JvlryPAOVTLzC8mQ4kETSnfI4eqzcCzZ3N3fyOgicYs3lATvlRGolsEB
/VzJJX+yphn+gSV4x1953IEVyG0uEszYWXKbtzlETZCi4VijVWqYhBP0QFj3cRn8TPE1ePw2E9GN
5iFe5ZM9Su8QFDqD5ehHBZXLObx67gYhn91t7rlPZeLkPF6Z5liYmpQcYvWFMo7hRnCiwUMMxrP9
alvJG/1Yqi87j54OuZ756RFRinH1Yk5RGgV4Zf3VQa/hH61La2clG03CVyfZsmiRAyVgr6aqSJIx
NREnqEyYA8Y35k+6WXWdMAygFNAoUfRO+KcWzbR3lBY9a4y7UYt+oy8dRrjuAHupFoKOuPA+Xhds
Nghy5WVzNE/CjAfweHPQH8coO0sN9yf5uo1E/Ka3zgZ4vIP89THONGHAoNxpFQVn582sGV4OP7PN
E+z+d9LlCjL9A0H/CQiJq2tyHNggYh3ozD2Ha4LUe1EndtqXhRDorP88SW4OIkrBkSjwL46sVxG4
Ej/dfYCczHyFkCir+iUKKybs/yoZD/LUPlzk93jiYvSKXFgPS/zMoR8t2fyq1925/TcRiDU8/DH6
7qHTXoFZm2BHJCZPw/ZGgEH3klOicju5zr0u9yVTw2oJVMpiwvSTAvvWzWUauxbXbm2e3icvK/vD
PyTN9PRAE20VDcUWnliO0Um5W7URyphAu7Om7FRR4jKICyKOdLcm9sjeiUuoiIm3ihizu9INGeuk
E42riGlR6gT1/yV/EiWKe9nXe/lw85YLs/lO09/oDejdguCZINxLpY05gFKAHxPVNYMftpuznfmr
lJysDyJ0qlWNQoWDA7eiNdNuUauzlhFCx45mFpM1boPRyr2UjIteSMcfAWynyi76gIrfccoYnmUk
tOl+BH7wZjm/sJEi5pSa+GeVFgJ+Gy+Noiff/ROJs+wVfC6wYN4dS273TqoFVxUdL1UIsqyQ2GQj
0U+qAgMd6/cBTjJCeLw1vGjYfhUBAxLciZyYPbZfAKTty0uaKmBFqsh8r/RiP5KrMHIecD0B2OEr
46t2c2BCYgTTRzA+/wn32hFTlLQkkiy4RvJIMGY7zou3C19DFjhPQLss6t+IXhRcNFhPcpGSR/o7
e37Dq6ZOvkKo1phk/mfurC9iw1Rv8WZbt/81R54S+ZzW2Iyjazs82TWnLrubjs+mzw+rZVJxpZcn
zVbPfGchhdjIE3CYoZKPHztuPzM6cFic04ifjKIOsvV6P7wmSEAd5fTlieWCK8rB+yM086RVS/e2
kKZGVD1f+fxBswZg9g/6Kqzc8lw5xiievQt3nE/TNVVE9xhECoIWLiZaVMMSJG/EWQ3BlwOBtzog
JWGCRyOreHjBszoxP5DzWxNrKuM+FLyKs3+N1rWWkufJ904KosSASykAcF+rGc5leF5/eekTT7pi
+PdqjVw2dWf4KNhbLMktG3mHSRjzMSx7HqFnEl7gTFn8fmGDJWey1T45nW4GU7WkqIu5Wjx18LA2
DwINffPAOvc6qiwHa/8HNCX++OFOlQmE0J/t7f8BpxwuPPtCHhsoODrnBaM025SzDaGKnTYi/VJC
+fNYGfVAoX9i0AOeufQ9v3htVQnEcIf6CypaR2iMFaqjs7n7dhMRuHUH3OTgor5MrRCv9aAX7PKc
s/5nRyiB3fBqwW/JfH/hp6zB+1kZCmaj5yPhhB3Qv7HIg+Buxy7+alAQlzDlUWAobzDD4Gj81lWj
O7zyIwi2jP5TtrruHFtXY86pQ18TriPqb3UDNAmcGSTxvxH3xZ1ajvgS7aBuT1izyQ05w/rUrwMO
GTnPJAEf9r8x8gFsMcZhe06sCyoW2J1/DW1I7k5p56O4cFOnBCCltsG8EDprgeE0k36EOpT+20mW
RWerQNHTuK3vHNXvCshHymY/eEl4ljeUEG3FpLUuhK7n8/TpYjaiVyMQeAkIZEuCloK+i53Smc6i
rQG8TKEq8+7jZWCmK9c1DMqhZjY1nHFEPJjq/4WZhmd+W0SGAaO7FBrytKqFJvi8yzkAx6Xn/gtq
8ycq4NY8+9yMcwrHr1m1ygC2XAAUJQ9JpLxLMviIw7Ee8zgROvRQIsDn6B4sL9MvTJXH9OulztqG
AlpE89TK3ukuf8xb+tcNxVYThDOAd5yJuV5a4zSxnbs/iIzPdGbXNjfef122wXYOt3dH0V873BTU
ItJvhvthziHbEFiYb4yQT5uxf9Srtp7FsQfpsyrc+0rCFzXK7u6RVGVL+rQW3MWC93WLTYIYmKFR
f0a9j9NUfOtRCWchnD2CAS42bO9AJAX23f13WKylA9sVeX5FcBuMIDnZHoaWJynfcG8xZs+9GDUG
aIhWTE+LDU9TloSXt5Jz3FiKQVEJm6pBWiGayb/Y0QRl2ClkUmVzJZcFeBOOdOS0wsfJBQ2JSdte
pPTwYzZgz4FM2NSl71SYxbO40wPMI4wPf/DN8F0AzktuUey8Vgyk6eQUS/hVO5+FhCWtFvwqXLd7
GiO7ANPFlF5A1T3EZlHgw1JwpsKbrONOCsVNYtRK9RXw4vF+m8/hEt/6q9ACZHikbm3g1U2IGWLm
1eiAJBoCHdFvSqY2vmn4HClGKO0yaqxQ+hcB34r2oz0yIiU/nbVeiI6WUH3FxNng9rATeufEOsU6
VCh/3TZxGKmsp8YKZKIzYsLG5lIuXYsbTzgKk3Yl+GHZj47FgPKmJjwYt8aSfw0HdVtCyqsDvCPa
Xgvxvbjkop/KHhKTKo7org0ZDFujonhxO0ZILDJeW6f+siyV3jbQ+xK+oZPqDEf+kKs1ZQH7HlUm
4HpD4SalOAGeW0EEUCcKB1OLVMpfBYVlBXkbPC2nlx9XZOY6ShLk4//Nd17KyxiWohE/nHK8nJ0u
I8mls6FdjmW11KJJvCOBpoCIcvuUN7Y9ApKt3CHvXYCu3XlvMp5OF8WULIyBMVueq2Z40h+g+OLT
NiqpdEfbe1RL5ouXxpxgY43ZMAecKlccQoGkQysFYJsUTWJIC1lG3uqdejZnykU3HvztiLKnm4id
+27YlJ6JhQvKTT2c+EdpmUHSIumqM5UOzigNU66ZCWCQZF4YLPOpxQoQQ3kp+HJKsOSL7+BQ7DvW
GAjuRxrSzcI1gnRHBa/Ceh4zkIBzSRPdAHkqkM+o7/8F0I65y/otT1/HwmL28RaK2Y82bJVyujnU
hKxKr+eOUTAoyVE3F66CO552Llu4+UEnz1YCQcT12yTYepFVQuGlytxUL0Vz+k/Cb6kL9hBFaOEx
lZ8l0BJOkt4V+kzOKtb3gdlUZicTkyphNWQED4Xq82IU/JTzHhMkarCoSHl4LfQyKUzomJM7mCu5
lO/wsycUvJ+NLYzWIJc6kP+EnEmWwWx73X4itfjLaxi1gpIG2kbX+DAq1Pg2/fWAjWGsFsaOcuHb
Cnt4amOk2fTcJ2Yrqxb0BOqpUAKYtC3UFWL6EPr9urnpAzOUxOVOQ5Nr/6+mvTTla7qeWw32UVHF
haWkHmVpp6Xn6HdJVkqnco4LrVlWZm11/8WikYx98NUAVnuqF3ROC9Fva+H5Qfl3r4VciXrs2mZ8
TgR5pkMJqtD7F2pea34/VsmfzPjYiGr5rTqVomJUptW1+V4EBjPSVln7GSsA5eYekKaOwQpa4aJu
eP8jFuqgB2punoC2CggPibLGTN4us96kNUY0g2CSlA7ti4CWq7U2fyHaMUCfUq+q4hCYkUFL3Kfl
I5juuHmyOGUQR9JNpPuIUzRtlBfAgLOO2fD4KXyR7J8twlCCDeyzWSxTACvVvDxK9IXr3duX5ta5
Lm1AsSBZ1s7omqGFOmUwWegL7el8v4WJY/BxjdDg+LRiXOS2AJcPMBTS9dJqZp2LmReoBK+7F5mD
/tSlZ2tBE3ILZH6+Lk9uOOozk1ydSXVHmyc6jRTlHdQbtKHIq94m3axq1gQdl/VU2FDnOo1810ii
1ha1VoznWqyOMFFDBrrkcb82/emMdTg/ObjBgCAq0RnFviC2f5POh7HZdxuBoQSL1GcPf4uvJGO7
+D3DbmPdUahTc8pA0S5hHqzi9Gg6VCHiC2zcoKHrtMhgjr7iNI63PbXxkIxyg9zjCbUS2s2Fpk9t
zJAKv3hlGsTCM/FT0aiZUTJnSr0sDSJxCfP0r+wPENBCOvMabiYUOp36JU+D2BuKb1HyT83Lz2XA
rEeoimkHtG5fZkZrkkYGos0eI1D82LJg9EtOw38JlHcYFYAjQlt3kS4mkSoj8HInbBXd8CdlE560
UXlXi+hMXHcFickr/yRvz9OJgd53DsBzwg8UJpsYpTSAnJ1uKgr3Wy8dsOSirQynELW37IMzz9zz
gc6VJWPGG3JpTTJwrkd1T4P4BUEK7bTbav6208ubQuLRsLXzie8ArctlnbFqTC/iHZjVp6G2HfYG
JiqfnWyUH8R60yJNm36+vFzZsdi7RrXMeeX5Vei0KAOIldhFPOx+JZKSWjwcQydyfDJy3CRdOGCI
de6VT1fyXO+H8hFMpC6xdyaPidhk5wcjibVQnP4hl40P2PEecl1b6sW5VVKF3jFrndVYMInTVuw0
PaQG1BrZULu7eVpCzi6yvZNT2sRJ9qiUhu3OuFkmKiaLYpA+7unG+KL6lB5WnMZTk+mUGWWlPUN+
3wSjh1AjdIbodAEFnfApB0ivgpwamY+lmtd4bhm6zDusnf/6gjUKuHkEBXq7DK2NxiF5o4vOn6wE
4NzpztPsCM16aewTIYEmqvPkLK4cDB9uCzNQtzfyhO9k0G0bGt59nNL1NUqz6wvHPWgzQ3SWT9yW
S11xJ8ICm6vbYlSqO8Jm6Kuxvmp35Ydm6P7RdDCC3Xt45wx0isK47OapI/HmQ0H6OO/jY9fgOoT4
hea5BS9hGrH/Gx8v40hC5+gDbXJq4/6x/k6Sr4/lo17cRujEHQp0iJIhRQqYXe446/hU3cdLKxcH
AK9cwxhaRUuqsViKm8TS+8b0zq+mtFlqFlyJhgNQNgDDKVzSVNPSa/1BJv7qPLs1b2YaSFXR38Yi
tK0W3w5DMEEtD6VZ68gObMZdg8co3GJlSvauL+Vj1AOLr6+HO9vV5mGHrVFFLH+6bu2PcDkK5t4Y
eS3HRctBbeETbGh8ewxy203iSgzpclSiJIB0Gm+6HlH1n5IDO7SvvShk2S32jbnwAoYR+l7RkKKd
5yDq0kWB94+5JHP19ba9ViIw0IszEbJzmaCL6+qrNp+tzbTSKaMCz2fjvqsn/OWVppu809hiaUrc
ndzC9tVHH2hO+1kwN9YiDRzbjWy7y5HFS7K6/viGR808tKJCtvuWAAR6fGJ5hxXA7n5iMWxtd+v1
1iJxi2l5TF5v/B34MkDO0kqXwXSvsXl7zlYSFqpam0I6zWdMvogfLdN3ej0FieNcSa1FaljymtVr
dtvM5ZDZZeRbpw7nDuEKPunUtPEVebv+gNSilQ3nB3IN86bvvFdxdjNlX2OvU9CgVEOdxBr92+Ew
rXrKeN3Z96RS+n5ca7CbCbvYKw6B8bfQoYAoJvULdq5K6lqWehMTFlQEFfBE5OUMnRwOdooaOimQ
Bgn/BozLTvegBBPtrI79xvaxMPgMgmUw838I5mO8Uw/cvOuzYAwy5up+f35eTv0ZXFws5Zs6xiCp
2851gTH/TiwMhG7sgaZCqAfRKqoVjQLiXfYccAiFkAXxzKiGXke2AgZeu98aywE1o12crCsCkFNS
Bl4IwSlgHimAxYlCkfptaK+zVPzGtyZ9oMwE7I8qwLxmnaO4/ItHKnML4I4AqtS7W1vRTYt6SkJp
CzGWIuYIHcWUV8GliV7xqcCJxyq+eFZ9x/8V398YwmR77VdozI2Vf/0xAuuVwaat+VuGSlrRSkQM
Wq8JdV/i88EqfXkuzvGVYjVVDJEilnoygJZMZI5iHEzFDCpBJVcj0y71YtYk6TuozaaX8QWCNd1R
SWaLSzkpx7cOUQ/FaSvpQHGARNihxT8lVXhBta5IIhd72J5b760VchbbeK5qVUjmrbrFxMS7eGoy
LGK45Z1qZH/eOdzCrbmnpslfxBO7drz/h/DjOKR5ZiYPX/ZSFyYyOhWprOHSppVF4AfnsqnCeYqX
Zinj52dWr3XpeazVLiUxxAz1qxa75AuQXduK4XoUljZMunEmGd8Wv/EKxC464Z6yOeUBKv/K67wo
F+c9n+oQsLg6DQM1Ij2svoam8nMpdAvKRx1dW28rNEWjKX0wCcNjMeUnTrPMpkC9B1fXXNVNWPD4
OQdebovg+Z+cCUu8JZMDzsV/iRLDLSZs1yXrEewCTvMHbBkzBHcxqQcf1+9deXO0NUw9bAgN3eTv
/NlLz6v0OXsygQ3MAHbZ9LSUoyjuizRreNQ/9n7WQFH5lIuA5nlRyFud7ZJszMruGJuiBCZpNahs
Eujs5FoqO/hWWNX/AKMwbIrOGF3HBo9gVP+ycoeLnFljeJImnZx6ch/Vv+8AfUEwf/o6ijSRdIp4
kMxSg6YqWWi1OdyNQJydxIoE4zMt5fqnK5OeP3jyZjfxLrxf196J5zZt/sypnb6w6HPYOJWJzYm9
/tfzFjrKbSgRUdT+bVGMsXcttAwW22STm9baRYAtJGsoQJLm1eqtKkJE4ZWVtERWoKuB2kCBKSUv
uBDQMsPc/oH45po3p1ooNz7MHzJLPHetSiJGbkz8A0k240APBnOvhEBLWmYAloU3YHmSSWztStKc
zPZPkQg1uOLCUINqROkdi1OSyZSOl5BqT6egcvdu1Cm/Ap1lhGbpKdVnBGGMNuGptAYTUVVuCcZD
3vQqR5vpDo+LAy7j6j5k7ToMH+e62sOA6UAAgofyyUokIW3Bdals2hp2Ovwbtm/keF6FjL25+rmM
sjKW0VhSy94yOd6/5fBeynvmlWHxVMo3dJfyK1xLcP6uhxZmH//zRzOdytbZ3AlcaJPtVgq3ftS3
ytRSP7P2CqjbhmSFU3yOVqF0Kl22dTD7Pies7tnMxOoTW+g0++n6c3gDZRBLtxL5fe1ItqvKB3w8
pbi4UjlRNq6RZzwvuC1JNt2HMnsIfTB2ocsCa8bsl0nMPuoCVdWp3rBpLOA+0sfsfBfbcWu3FWJQ
5L8849DVlEISjkiB3FkBNgHvM7snttknyYbnSJFhVBOhIfDwxxraWEiLKDPSw6DcPW+N3wbxZ0Sy
CmG0xXkOcWZsNz6KWIWa0wzKgqI68l82Xn77pDZFx6BKaK1BXD+zLkFTbHpqAz+OkI5tjr+YYaZD
eZhmleCKe9As1OshEgTFjqJL2ER0pGGGmSOZT6S3rS9x94Ieqd9KT7TQAuvKPuDagsF+5MLHmOh3
+ENBJHeDa2Ft3sJk2qVe/LC21KeAChm2jXEQYj4nGYedMPNkGY0AW9HFM8ByHuj19cLum/Jgf623
wjHplzRaV+uXJgSeLJS3wgm1wwU072NdUowTo7yR/LpkbwZZ6/7yORoddNSYYlIhsbh9+dvBUSo8
0s8By42Ok5LfTpp9tYWJwSzWTMpAjl/RKKl12vKD5J1kJkYTLuZXm++F9cN2E7wLKT6Vsa6P8a6R
725HKI2mGTxZ89GW/WdV7gDfNmhdN7mbx+3TJqvfjpzAftN8kTTyR1DyooxF7i8zEkU2lAEKSwPM
bUej1mZSj0oJrzZlerIY4nRlElEaNjFXvE0qSpBGsLvBRzouDLFfvszsKwIdE97ZHd001XqNq259
d7WN6tfCfs4JwPW35u88dNGjZzdNfycVrmiLscu1Z54vjB5KhWHIAAKb+LmG7GIRknzC5VfYeKL7
86rr9B1DzmO2tEfUUvxuDJyPAK/2wewitxVOQC9VVe3bmGyd5eDC8jXUce7L6Jph+TKc7YwvTHDx
KBLVlJpGf7Rmx986wtO1a5wintcR5+8nv+CmArII4yCsYFIu7MMcvZqMwlys1O8ooBbRxgBntx0Z
pvWJzc0t1c8I1WcW7Oj8LQYCgyIt5MzwvFqpqJnx0FHChPi35e1ZDGw8ByMERd5pehzFrnALTH7q
+d8wnRUzMFYpffC31pVrCdfLouFcrX84tHCkf3Yyzn4FJyNwdmIIo+WLPUODGz2HPg5x8qaGyH+r
5JwZfsjOFm4BG/oNdk7MDKkurIVsUmKwAbzplNoOcnASq1XoAfvAi1BBldHBqNRWDqOH/mTttk1r
vxHGCufUSPucV1E1J/nLbuz5agGZJkxaXAHxSkpfpv2vzTbNqZGj9mQNLOaZMoWvRrqZE+ZEBdMW
smFcLVnD/OPzvLcQMhiqQ4QYPNgDUDuXwq62gtd/LY8A6SfR4z2KQDMXaiAPXu2pmWgjDQHyBf0S
po5XtSUA2MSB3+ix8nBkNOfZTllM42kUcVeu6EdPfGEhHqjEnWkpblWB14FXdu8KDBjySpZFaat2
Ah8dJ4MOlftQ92kljCFVzwpXxk5CV7Bg2Np8xdTP/s91IbcIcf6s10fyAsZQ/yXlVkcX6muNONnY
2RWJIIPnShS9NSXaBLvaVgrec4QgNA8wf+NJ+hSdxQrF4/KTLAFmx0gNqcTGQ2+48diJe2yOf96B
Hy0dFOvENZmCJjsl3AIQ7QsPIrbuInuKphzSJUfxxlvDH8666qgoyhqqUsWxJ6ArrtusQeZq5VSn
fslUU8KRoXmc1lLdtYw/QYfHHylg8W+ZCMXAH5GvxkE8igEheI7DaZC0kP97NENUSwczk9Q8VBiF
b+TmvpRG9/TJCZ1FTfxCLZhd1LkOtS535YBhlOuSTsNmJjFz44XU8AvShTRcgZGFySAZwxRQdXCs
RIQd2QgqpmklTMJtS1YUCM8Nrr+stcKVvfbZEslxcyxWR3Np+q8p+Vy/fXudhUUe1IX+BxKz0459
eWh4+EcJ450HopERMRSkgrX3rf5kfH8ffbXYHrkssKJo/5sURgZcVvj+3HAxmGTBlkCNyLQcIEM/
LOm7X55FFVhJZJTWLnUz2hOm1NyFy/p0ofsuo6jLXz8NL/g77fW3ZVreph3rRdDGPLE/6IvMFlul
gxnkdV/sBx4O/ACpHsw+D12+WpYZAJjWrdeottfvIsQ+y56zdyfM4iix30g2pUre9E7TmecmCTu8
MaM7ik8gW6gfrhcs5r4uuS7f/p6LXIiYuCEqb66SpnmVxAgpwEbaLqvEUMFcWTTe2sojTVVrMDxS
uUxNON07ycxzKz4MhihUVCMFZVOLYkmbStUi6B5RSKY5m9aIv7HUiQ8Gs+0BXVv9cO8DXFEdnXTa
ZIIl66y5XxtsyyOauRK3MPZtSqPNzgiCGgrFxFCGLiVtr1tFfwADybw7zd0SK5mWIK9Kc3k0U4LK
pVNMrhM/bSNBMRYIfRMpY9QZ/3YgfSjYxkGDdoXteUj3WtHWYBsxcMzhY2Sv7aD369nW/vI9RVfv
qyyawmGBouyMxPO7xS4XOetc3zo6F6+XhpgR4djYjjhWcb09/Nn70WBx4tjZ5Q82JAk8Q/Vkwg3j
N8jZLgRoRwGBhujmrQAVYCAZRj7FjKVs5+TxJlxkqFvRDGvi6iKYwRdRIVIXO9CdUGCNeE1SFSkF
i4s/W1bEZQ8/cMCivy0ExusSkikkq0jFchgf/xaMlefDESGjwZGtA63ExeU0aoXwAzTmlIn+xH5f
H3zvjrl4MzxDYyYUrQVlfQkL1t9b0rKC5hpXlUugEZTHikLxV5ktWJ4lcjVkXGpi1TdlqqKzAMHE
zcdSX2RQ5iAJVSudaFiluYwHDNRpGpkf25m9nnA56NiGr2toPZaIedvvPBIgpkHz4UVWkk8Tbsbe
r0ZG4Bn/VuVjnI3dcAbM/Mx0XERt8GSvEJ6sxxOlJeNPmdVbkuEic3Q68iDHA6Ns96lS0dE+F2Wr
RX1Hanyu1ZG8X94SmCHvatOSq8IHccFIWYJSUYk4HyoT6jV3pcWs1iMpEwL5nNMvwfjQ6tkKOQ/Y
IKnyL+JtLS9kocp41l/171BUflstjeaOJ1va4YMuiIEzwAvgmitY2gJhbu/CbSXMHNOSitMiRSAU
s596wcilzzdcEBTzcdNQuIWkv39W5jDOx3hOIvGdkWZKwJljY/18OqJzuFTJxAScrwQRCOCABAal
i8CLAmjkeVw0lcz4hHFoQvnQlKlwP0ZZWuatqMSRhr64YlcyJ6QGmtzwhASsieAC529Rl5N3GRa1
hDgrVLWjHgBnfbU3Zd3JYQr1SSEqCaeZL+bEvgBolPO6OH2m0nWKI3MbnSHzhwh5A2GW615NMClK
bbIeT6PoVh8OIG6xxp2Ziqpn+nZGZWrTd5wLDTwOIbN1oAX+TPSpB7wgkmA+9WzrwMFfSr+nNTrT
cjUrWW68ZBX0K5AukieJ0IPmrJS2T94BUXiOblPia9DX/eQT3r3rMC5meh6m+O8jlpPju9661eU9
WGWtILzTTCVx9c9M8jlRi59g49vpLNWHQamBbTyb6smbUWElnm9aCIa2nfR8tYFP6Z8gue1dfMqc
hUqBJ2/eAGrCEJhvBaB1uAmVTR//vFi6iLzffce/Y5bKnBr+8NFwTPQX8qNmqT3fbmkv8HoSe/Q3
1d/kmPWu3+sh03Zj6Gbrrw8uW6bJmI4mgNQIO4Plns/I7ebow+F1IiOOD1I5wiDNsOxiUkpFcdNB
ukctpcDiwNLqkBsS/i03/v6/gK55CZ6AeF1ZDHadygmwlyHjnUUcLZhLMmpE00CctaUQEYEYF7IY
1EQ2UaE4pnYY6C2++8w2obXbK2tVORvluMDyenTmkJhuHJqdZmGcpqRUNZNrSdXCiK+CKGViU7iw
rbVmJ2Qa2UmXYpNuQ1gEs3c4hcqBUD2WyddA52e+Vj5R+/eNqYcKIC7ZVn6W99wTYoMuC2oudrkf
Cis+X8+i7BCH5XTgeCmxZt/PYOFQ/TmpFJ3ei3xzDw3LniuLgDc6MRcgItoMzJaT/J/4HqhafAaB
vjNtaxaaNaP4hITGCBEkJEeDz/kBftYTG2Nm0UMUO6w1x9MxhQ9Gl0szzTp1GqdH2XoSN8xaMumL
HxvQXLgSv8LK7//HKhqt65+vu48/h4ezexlsPe1A4wfmYmlxI4YAOnhSButXyuZz9FDsgMhnsUM1
p+V9AYvGs3o3yZNlnr00ahlWdulChEinaxFREYhD40UFJLq1kTrjcFY6s1hvpTZMKT9GYmH6OlP7
YbL3Jn/XTKmfjEW6xjdypCxycWGooK0rbViMosT9ZtEgZtpE0nP7aaWnz1vbGxuS1MH83MmEdwf9
AlbJ/rK+FQ9+i64blDVU4BQjZpWu1yaxc9kneg2zYDp50ZRAHcNWZXud6ZcHnXt3EAjSCEyzaubm
cmpUQp4PdGPKy/uHytc25buGMp9O0tpy+QFJHFAwaS9H5eeUYonFUGr1Xl27Zw8ylbcP0+lbGatu
Y5sjrMlTkwdsapVr6QlxMyrqRv9lLbeecY7fLRzMvKUIqJCjsZD9Akg9CEiQBGWfqHsehYJVVDs2
GHGNaFRjuu47ZnoghJzT2ZJz6vwHtjNf6Dk+yOSeCxKEFRsfYEygRF+GeUSIVJgxCPIxZjFV/+nt
ioeibV4fsa4IIpUhKtUSbZVXGD/fP1Y5g+dEOW0kg318ol4zpQVhCBL01dAsD4SPCKLMEaAj7vAW
zJlVPEYH6pPmLJyNxQEXyavlXZOJHfsxQkKWlW/Z0/wYg7mR3DuIHd9CrrymXxH5rxtprwINPzRT
c4zAvp1WHi4Gz4VO4lPMYLiImwGHYfiS4y6vTWCWPprR9DjkToioTnli7ssCA3AMlOjOfvsPE22n
5DgUy9flZMamHSxwP7L+57bcTxVORSnjhtiCJ6Go2tggHDrW081F19QW/NbXZqa0ikqWrLMke6c2
3Tad/dkOkJKX+91tz6n+T/4YkBeX91/qAAJXfxCetGxH/E99J0dEom0NYrlLWwJGBrS6MgEJA8hx
Olz+W998vh8mw8BGaAVExJ6jiOnvcEmSmqrupcwr+pUCyUH9qv6dUWUZjq+5Q1JTl+0t3TGuVXec
j13FU0wS4EnXpqQtGYuu/PGDp33vVeZSB+evZX5U+ASaJbbBktrSWLayid/mIqLienhjHtWDJdOV
ikOtYlLoRdZJOj0UIgKvZC6kouMRdeIo4uG8bWMtddmNlWFRnC5CljQFZowWBh+t3HdplfTXo5ul
7OAf8+t8psaWdp9gv2FtEsugy6PeUJ1NzmRJAsoeClygdNAwmaBlwXGfCe6vbFm7988PMSxpipm4
VjKoti+uAc5WRNRa64njtitCf/L07xfljZMds4KqGB67aJKedR81aVHWYJjHRDbL5eHcGs4pcRJh
enHLdXZusG1ng29d2T+psF2vJHPRKtLykdS/J1YqNPTsTJkHi9ktOHw7Ro4wqlA3brYtPtQrobwY
WQNt1xzL92OVquxyNIymtFbxW+1ulbNhX37hjQ3pHz4lYGl88I91WSWdv1373wwjezzgLTbrhQHs
fAu8JGNroE8WF3IjlXzInnDlWtGHGXHTUFybZdfhzFL8ctfL1OpWaZIeJfmT3zLvPWV3t4AS29Lo
JClFbnC9D66S+si4Bk7k6z3mVYQ0d+n4H+oH4X3BI4+PgYC4n7OexdFKOox/s2YR1FSfCOpb/Sy9
WmJZTySTawoV1lcHB55g8UJ7W/1j7ajz1xuPNu904E1tQw3q7HOqWD8SOZyKLhrsxZ14FLc+SF3P
S7fyeamQ9uqNLlZ+fYwRqXQ194c0vRi04ZmTKAi/26rc9nxm+N04zaWglttFRwUrz56OKzsC+Gsn
7tmEdH+tFvNSTPThCkqRPMffn1EvoBQ+3fVfQmnFkr+6R6SLp0gtHFcBl1idfCUBiHBcuesgdlH4
CrwZ3O+zIZ/qdecEdPKjgaNVqRztT06ryq9sAtBC6qCJkIyluvLrKbkW+uiMC3oDdDJCz/sJ9JRO
woGZSBdbZUHOxbSJ+wLcOdBgdG1VLpgpmnd2KBEi1opArvuxny3CIs87hs/ybee3RYLDXWRO/gp7
PPHE6kgU5Grz8ToLb9dHCg2ycOhHzdzhqAdpBjQCN+hOvtnT4lhbpqu3ZwFVMvTZDe1D5FYEnsgt
fJ2D58ATZbrkwQlj8fis8bOauOBcQiZW6pZCPOVtYNPC9nTF4lXX+4xiF0asy9va+3aPuF8VZYE6
diUlh62+xVWPqNahmDgjYxGfYWG92p31ip7GrKkREwpxq0hZkfrTiZ+v24eArYtql2XI/fE66j4A
9gnXPDu49pIxQ4ksHhJROq6aFz2HBVJpq1Fm9YrvQXScTtrOHYwp88P4DlTmhpZOPbBdHxoJUQQJ
YDQtzvwm8nr7cp1KVGh+eqt4gmAX7zxBvJhexd+iHEyhwPXpt+w9MWcqSoIt0nn+yMbLrKlQWRZY
IyLXhesMbqMw+ZPDqJT6/reiBDXL3iZAM0FHaGDhEWwmYSnQN7fQIvfyKDYCwxTVW43Xlx3+8Ugi
LaITGEKtHZJ1Tgw6VdM2Afds85XHwI/QKbUe5+YodKb6mVjWrPI69Zo18jXN61vmy9AtcbYFxUoJ
oOkSNPhRmZUe5XgS3eNf01mDjMzBO6i8Lta0WW2c2cnqGTXbhHw0Wsbf1wyyhrzZVZy4B3t78FoE
i4NSrI2H5NAj3wy1Wr7J1UramQiWPK9AlwS6qiuAH1n/O4QjYDZt6GegX/cCafBP+tk8k4xQKosL
tKDdsprVLO9O0qODCki+XSi+KVuiSfIAFBufYyDp5rkRVCpNUNIoFRcn+l2mBlSXufVdowUbh4G6
tPK+gqpCchQtOcfZ90o7Med+j9409mL/C++5+0GerwSnEe7e77bdb/xSoy6LlaBM14k+U9/4Oh0Q
lxQye2VvRMjD4wkip2YtstTKNrBGDOUphPu708Q51RILLV7wtd4dzNliZoAqybAPp60cwwHiL8yq
kMXiFYAIpPej486p1mMAeQzmO4w9i/5IvM33DyeXpHuSkl2VJZ2DtM+2Xn7mvrqf7IioCku3/E6X
t9rT7G53/nqi3SjuZ3f20TvPy44SMSdP1wufgLh3JnAGpcX3w0mQ/RphRfo9+bzJYyx1re4DvNDp
r/azyLndOtsu1d3oR9Dz6k2tQ8noHbAJkoAJTiy+xFNQ8QLNo1YaN7u6DZxRd9bA4MZAhEcb039y
P8r+o9uedwvZsWF2hB7cG6ZPzKeKqUvNfpvOzMX15wPhvv+ichhlx0bKXCYGHvJuA5pin3PRwnjm
XutUBh/aMcsBZ7zwKSZktwKu6peNulYJ+8vK5l3dDpniKb7dQkQX1Ilna7NJ02ln9FKW701oRgC5
AjfQZ+2rBfYINOnTZWEGeZMIDQ8RCBbgrIs9U7Fw5LdxOuWgT1swQTH/UTcf+23UjGymFXDJ4R8O
62BBnHBUSslz1MFaNvnVemTfg09qCaW8Vr/HAYpZ2djZORWcxqgAhVpas8FT9+Dl8NbY7HAro0m/
UGrSFSTHnc7MCoWg3XpHrjAfUJRwIln10BZnjEanhCSQXUJZuPMMx8AoL1yVQZm4KpNEqxjiVVfq
s6+iW+QJeHLnZgDc27MKRjJMGUQNkDr8wJH2ow/Z8adGMuPS+D9JBiHcPFFBabzDr+SrmJAn4aC1
oqED/X8SJQJhJrCcinXVAw3PzbpMq8QSt4m/atsBFFAen43l3Fo2vcKPHJ3JR8sKmmQAzrhAQWGn
35dLTqrQfyfqQ9iabbJaNK73U7xecMjG14JXq/44zXBfMhN5LJG1yiVMl7Th+7IYC9HNaqQhWagv
1ENs/aswpLEl3HmeqGEhp1/S2wp2u1JHNTgeqnhArBghhFHSw7gD4z+ugtDhS5+rw998J1H/zLyx
TSoD1WC2VmN3NZgsGJ4My9kkbVbaW27sEAWiYA1T94lHifGlU7YNCwDlDdShJjV/H46lR7NUwK1L
zvWtf065LQ7H7KGhStnPjAlXhaaKpMaQiy1TirXEDgNFHlVUxKX8TnvOaFw983HFbZ4HUiSawwWq
siMXIi6Hk4tC71TGSW/6l2ic7gdnvyAHLHwlrkrg7tWjaGbau2N3CA+nuxRUeOadwQ33Ve94+mog
K+feHwCiYw+SKTAG38BckAfaidd+ISS6jhseemPAHybBxWyHuaNRMoITOQENch036vymzJfgsqJC
F0noyuIFbpxyiobNAxuxdy2X0mC7cs8jlwMGv4YG/wXhg/ss8S7wjk9e+fNRHrijxE3lsVmpDr4W
Qg0fVJSLUaiNhAzqGXJT7CRpvBSQZAPTIGBcSgjb+sf8or/n7gsW/plUPwmfe/ZWZt9t+5aT8KW7
RyzmDGK7tYG11AbdCFM+Imtlibik4W5tqpQyBoyQAGm96eSPJVxBh+cRcXPPi+QSlW3ATv/Io/ty
TZ0l6tL8DgiaVJOHwr3//ZAUACyXNH84+MLHNChHrs2qvPXrkAR7VSRBbuFjWylxuJOf5haBt5ZG
o/0Ldh0DypuHbSaykD/CS2Lq0pAruE4PoJsT7DBEhIa1BOafcxEhLUzDDX9r8dgGip/DJ0E0OkWt
bfQLetXpYwx2Dn4WR8eZU0qtCx/Y93QhqTpdeVlSjqv5bfAqHUhBLwPGgOSJI6Mjjon+5Z9yAcxo
/AmVlkW89EkYnOHCG7MREcskfpwRp3/W5z/9DvIkg0h7yTQrf6kQkxeKJQZJIa0CCtm9Ec8Iy6/e
Y8VoBxwxfdzHvQsAEtTfL+nO05m1ONq28UoIzgRE/ruEyStaZUdASZsrUohe3ZTk9zXEe/l0SOi7
eX2fWDFg+FXfV+ERqujozUBEfDBIvF3PfcdoU7izux8ZcTlghca85LBRp/vtiTHt1s6jv2kqRvKb
HrY4k/kU1a8gAd4rIn2F6b2hl9MS/Dy3RUmcWOyuMsDikafn3/w+qqINBgOeVmS0K+ZcSNqKKbvm
yUOYtQ+g0lpH4MQXQidJhtZvaf2Zq25fCcVql01otjN/LEh6ypEn1dnFELBqrGITeXT4ZmMpeF0Z
Ib3/U0u86NyspeDg1zUmdugITh/si14zn2tqIKQk5xMNNdFG5pqLAYDzWD+Z3qM3Dgoo2k2N0P7M
eMX3dE7+3bpVojDUZQZeRmwO8ZfLCFquxnXy/xEr+touPmfsu3q57auAn17e5qyEEAEd2C6aXmdu
YhGCdZdSkUnhUV8fguDUTkUVgyDqDt7cu2Ni2T3i89Khe4/FbE0BN9j9Mjooq02chotkeNkT5dL4
SmclXGKNtPG5pjxZm5XRt7JZP6XXwMgRMk5qCwzl4Fq06knOvzM9cgIogxmb1lZhyC3o/F0YwR26
SyxarO1riX3UuZ8+Ktk2OA1fhot91s+G8WYQHGGdGA0CV3pvq3ijhVZOepkvmawz6zUD+Bpc6bFA
BueNcxeG9NBwfnvqDHu6330GswHnfKyBE9gtDs7LHcRJw+JHa/Ts8OkAeweXN3SYm9lfUIY11fQD
KxCfNtDEA2ggSOMXZnx+rpohpu9O1mighD+yZVV1+1aVug8zZrHeyrvi+0mAOfS5v+4h+/KYrQG7
37PHSwyf+D+/3gQcHeBn0rD1HsJLcYqIXcHhuREjKR8hjmiJv0uVNQgXcvw+HRaQqcoJnDBeC0wV
xyDQrdcrrhXqaazk1Kc3sQTu3G+Vf5dMKMU5q1fK6QaB7XdfiRVQghLDzwpjwHbyoEnn2Bvi4tA9
yzZFOGyzIVy+HlMe38/uuOMa6ZmOtOKMvM7zyCsN/eP6ygYcCgkvJuBr5LwT/50nTZo77PRygWf/
5uNU1WOD54wsN66aRx0w9EGY/wtaN0Ht94DqWBbxJxfEpSZsXGVxrYHsefd5dX5sbCaq8sBucqdw
bXurVJov9+CTE3b6BxxnBcvTWr+6byg/rzGAIvczfkg0jGrCpN1vqIFPxHBqnz0TDfRJECrBJ2ar
52OZpxksmfJul2lSYP+ILPOhAHfxGjh5T46ZvIMmg1M5tB3VQ91mZ5PheN7fK0sNzeee+OL+zI4l
p6csz87EZWrfx7h0nSBBYXKkbADnxRoWhPgmP4aYlYMPWtju0Tq6wRJbKCWjBPMccrWOLatAOwZm
x5/anhqylxcyahqOlUIWjRZ68i6598mPgKNdm0kvjD8iDHFqKxrVbu+SlUo8GIriGNrnbjsHSkXb
pzJ8mB/7DZARoZ5cLMHwZZGYLfIW1k6hG6A3YU9bVoz9v1nUyrN50uR8rcUgTYVGRVQ0TaLRwtV7
HPTLrImKyxC9C45+9+O8+rCan4mfDet25oQwbVtZsiThXD9+no3z9xSv9QF3+ArpWkW1m2MgdTDL
gZTy2bXlbzJwhtLVifsjSulNoqv/bQ6o1/53OJI8fFAhL61v25n13yc6yAwtk7MiplwzRwPlgMRs
BwWLDJmCD9a4SKwbhvinMikTTMhbz0st0B/qTTFFvF6f2BiiFm+JQx0i7fp5Znwzu0vs1miR9cAQ
nMTCcq9gXratbJtK8wOwYu1dKUsyTmPybgryOIU59meCaPe4FSS0VmPiqU3ip3bWC/C6sBy/wawa
em95aOp+92yyaj3doCpAHNt7cesFB6RHWyRULwVPQPkR/gALtejBTJtdDGxc2+bNFjXKUh/iT0c/
4EeFVD8u0jyWL04+EdQD01aipg+oOxge3E7K2irqLaalXJ8/UJPutneeZwEK8InorX7h0/5Jq7Yg
LZYZWNTcYMICdg2GUnjM1e+Vks2itpdvM2Uwrn/1V+vN1Fhr0dLXOb0UaUehLe0drBFCMXOojRfM
340H/tWRFtKNAlvHT+pVo3nnDsOQdCVKtc+hS3ygd4HFI0F3tJwBpcgpu04QiFvknbN+d7MWfFvZ
G/5JgO1C9Y4FwhboGUdAWE9+gmWusr/7kubdUkq8q7KWBbr/+Zsc/HP3nF0Vcgnp3BW+FSV5Vmlc
EU40SQ8B9j5MjfunAvgje6L0kVap9Isb9xVJNvZOAccAorH/aCuvuQY/OlI7fVKn5CkMoJ6apYha
do5h/ifMkD+DFfQIk0AbR1lePE7F/8inHujK5FtFFTfmDu3BRRivfaOI/4J/An6+KwGvs7WQERmI
PT1bFqkPpM6F7gDQHPfJ7sxD94uqWArcWNAG6WN7Ge3LnG613nMX9VhQYREKq+bhmHnFimcWQgF1
jiQ10FLCvYHirQd5Yj2tRWtcxP2mYHd2M+LUz5kvwBayqRI//3fSiPXtGuZMLZKLL6RKTxtDwh9p
EBOxIwa9rEcdlN/5e5jBdTPMlWKHb6EhbUMFQUPxb5GE6noDwwGVqxf79182IuWoAliaGazdDgFA
R9TlZLrknVBNHfljW5oQ3N04bmBTtj/FcvvQTpOae5t6I7YOauSJwlLY1xA+eKwvXR+3wrj6nnPn
RLyCQUN1e3SMM6T4o3FCAl6xSfxz6nFRrsk/z5QIOlMlS7vdF8sFZn6zeLbavXQUH7SAXv/CjKpj
JmewrbLmj9dSbRwcGzMPNwwiElZHgfZtmq2CTsy4u1bwJhba/OdgVWgmFgQWds+5Qqr+i2mF4Z8Z
kh9UwJLlVWFyrTsS+C3Yoqy64kscHZcL3pMXn8L5phtC82vRLJIRg/wCUumzvK2FgcFo6KMBuE/0
z0HH8tYelXeCswn4VE2ipqkAoB8WtJ5QWqlRaZfK/oIpwOs7kMNvvXZ+hLFE3SxQqvEclr1O2x/3
7h10/JEV3UZGuAfnV7Ebax3DXSkPK8CTYvmGdaRht3kktgHju6ULWGC+yIs2wIibp0f4yypqiRg2
/xujT4paE1u3UzfTXteUnSOFti2NkAGx12FQMP6fgPmnf5leJ9+whsBdl/JGkPTkJ9vvo1ZN93mc
ApbzZ3CnqMKvM7AbUyNZMiDCDIRT7eVFNXQkWNU9sdzqTfhoCs6yXLWa0PKiQ2OyZNqpA/AA9khQ
FgWd+29iFW6P0B/nxPvBNCKOyNvFrrXd5oOHxAdv9eJSHb+wbaLNMfyZ+WIFIg2Kd9AUmaN9aDUz
eWdQcuZs5tvFMh1Ch1aLHvqqUXv2/zweIWGqsDQZc5fIT4yYvYeJhZkRrGNy7ac08AaPcM5Esv9i
eA8OJSdftOoMUnqvD5sCXpc+6h0Qh27XaiuOzGgKvq+QjtFo3Ptl2Y8UOqOK/cQ5MjMR81nZJeeY
NGxO1zlR3KPfm1SZa5IW8j5XAjDUeaXU8u96rGfjI+jnAAH8jgJCZt6Ic9roRSjwfL96vLjS7MHh
M6xa3rP4Rh4TcqDuS/dKoxde4LdjJZ92uIiYOvlxNgRTOwuGGr1ZlYerZfXmlcOswXBi1ORc/6s/
CrpJyb77A4hmZQwxn/dO8KFbyymAAvQSqxjaebH6npwiIoiekzzVY3mrF+r5U9ubCG7MtCessHFK
dimyRItcTp3rBSKeV03Og6lib21uW02Oaecsi9ZyANcxJozGkGuKiXBjMuWHvxQaS6b2J3ZLPPFl
zPiYLN4eW/HuwY4fRuSnjCu3JAS5qN+mXzqQuItO+rtjksXAasLcxG7GzGSELhqa6ukjOzPeoDJs
hvCcION3MBOnq0iz8mSKlhnSOBeRtSteCiow49ximDQVcgpSMqnLXMaZhBc71ftCOMDFSsKV7Xrp
E8HQdsSoqDD2m4blxXKMtzJATvjBxf7I4HwW3NUs6pwpIceRtPW4z9QaabyMiJ3UWi+g6kYwWGTI
wRSwlud86JIksg3H3fYq8XcwCQP60AD/Rsf8O7wB0qXFt19NGDVVYieB0KDQeKjorEsVMnq2qZME
ohCC46GkA05D90NxmFuF+G1f//PjRbArr/OG7JWw/+KeZmXAEnsG2TLUZRBG7SOJqm5kdFcxcCP1
njLOAi4Lg+zu2iUEUZfN88QQ29vak0TgCoaSBpO6S9ls7pPk8eCT97I/XR/ymYor4yEDR9ERwwHT
Ly5yBfgwp0nShzKS6RAOBTn5vg4lkIH5EMlD1l5s92j46bHV+dY4eK6Exojn6uMsI2Zl4l8ZAFob
gTuAMZwsyZN3v4p84yctxegiCSFGJRt+6Q6B7eLUHUYTeNiA4AtWCiCvzVdWntXh9zIGJ/rvNNmZ
2hHRuIdl2SqZ8/q06uNGlFz02MGIy89MuEGqWbsCmn6+LJwgwS2+bk+EexOcyQmG2y76uvXwaFwN
fDNqWqzjiMaZ002hR9czADQ/oxL225pghVnNp1NzDVT4r2OoalT0+9uqiZZIGELHFvILv7Ebawhz
4EDpIK6sLAyp6ATGCnfL8Xye+UjHlxoKuq4Sk7mFMwgeFKl95Q9Hq3lbuKOv4yEdN1uJf9MlC0Qx
W/3NVVC96mKmvKnp7+vmz30HAQd4ZUbHM2bjMubODjecGm2fGYHeV1Hr7vx0G/l1aWXWfdrwU10P
6zXJe1LqC+Wdi83YfY0HydXyIg6i2Jh1DPdJlOv9GqlC2/EqH4eUwj6IrB0YmGAsr8qOpEkl+R/l
QB0xUxqezyJgjR3qtDyhskhvtClQrchCpykiuUIh02NnTlcBLW8B9vBpoENWOetufhJHGw1F/wff
zEEYRJrOzvPUo6p+2eOguWF0NYpl6TC+/E6+zdMZeITfR0/1n15Yh2V2MAmBtY4Pzwv770wALkvA
uWhHxMIBIB4Sy8dbpscSv7Jyt3M/HeYkkVdhUu0plOrbbEI26dw9fUoO6K3wMOzEASEFuahdROEh
+7noNBIBEel3x5pTqd8tn8daj0Gmw9cewMdPh9uhl8HsGmEpXb/bzoAgWOYAnptVSM5WfhuJlWb3
0lCknEuaRBrasj07jqAodbW5ETdKJOEtLBkQodMOmK2pez5s+W6eUdrRXkuHp773Y8KvOdKmIYDJ
ZAvOj7lQ5/Jn2RB9rXQy6o6fof7jPgXDr22oXR0g3FFMzV0M+tU6viZj99MHU8NcnCgMKUOa4i/q
rzR903hMawoWEhZD0Oa0491mRsW5ed2ADqi6Qly6+Dxzjhw1pXUX0ad3KRNQ4+iNHtD4N38XBskT
w5Yc4WwAnaWQ7JxaeUJLn0nad2yTzZpaGY/EL7xYjJ+eU+8+ntGMl/Cd82zA0ReY/Uo9ebK/zsMv
LyNY6YTCsBIvLg80ELnFxBN+JcfxNjRjzLq9lLq0fLpV4Co2alc3VdMoXj6tm9rWopT4u1Ee4bRu
cduuxang2NMHm6jYvxDpb5/V6p/48AskwCnCr9b7+wUQ/bj9qgGqiSQhKoSY0SEMQRjnWcensl5C
x8JifhVDUairPGeSCWZZUu8G43HGxo11gFnWG7NRqx0qLh8OtVDwGiGYohtkYYc8hjagZ3BOrxKP
o0vfDdWATaQ4PdVrccJ8Az8yS7gT/Cjbp2mfpB9UEnJtvlxmUMHXNuxhPLgKDKTmgV0e0elEYo4n
CNdKXKo7KN6uonG1gsdDj6UW/9iR0C9chd62ee8MMGu+ARQNuKbe7CUdlKDKE4peSKY3dwJOMXKg
mThAdEdGACr0aluAPxjt/FNx90cGNgcwBK/THzu8wBejSeX+Y5Mm6nQhWgSfb2lbVZGg4X0CmJRD
kxoRVJLjMkV7bHm7zC7IReLfvQkniltQdtIBMaNjKF+bk65tdUm7coswQx6Md1rmTDi1um4PHHtJ
1m6gKxmvDelZub+e9cd7kzfLL+EGP2Fhr/+I0Xl2UfHq9ywfFZCLuZhgGPbjq4OZLuApeXvEkdOv
kjdyJWXe4X08MTNEEIZI9ChatAZbgTWfLuq/Ua8dzArbPn5wcnJmnaOMamK9mYLC77SV6LeiHzSG
gIhMwtOrX4Id2qegKreyXbH4RYn5Hzip0CdJImmv4QBqG791LreVf93DGAskWiTD8TEV5drZRYsH
QTKUAAZF9vHt851/ggPfiG/4pClfgJk+nq5jcwNXYB5c0xiI8FEFzqYUiwcZvlKxAFatiSvZpfOW
32UF3ovbVjli4tjbh+KEvRs682eRTecH0dQ+OBO3qDREHTcUAIpq1xWkbQFlhystdZas6MuRxHdz
LFQqgIYx1lsRL4wdOhOtvoMwCp5W0R7fe6lvEs4jK7uwh4wVpZWpbMgD0N++gYWdAR7NckTp6u/H
h5fuUeDB5qcqUlSoCqveH54pADJ5lRA8Pj81Bq11Sv3PgCdOUr+pDYF/aF6z9IkRGsrvrVRWOf5M
XH5acj9db6GRQExctCshVBHWe65uEdoiBMavTSXOjjXXBuafXZYURt7EsuIV9zIrUDClGMlCXMC5
6OotqCEIBNpFLZWjzm9NNiwu3ULxz2TONvCt8vhZ4g+vlkYjU/xasSDwpFX7Fqwkl9mFJVUei25g
48ghsnm8p1+BvZMgOtcyN8RicHcaHi5feUZadNQfEnBSPCLR4L2aVE/JaZn7SrLvITXRxdgHVloF
SU9aC+hkcvZWMuqzNqdpZPsdEi/xTX8JMII9c+AAUtBwHa0BVZ3yTd16TLSHDIcIyWkp0Zrbhlw/
Yg6tQE1WhSkytrlfnQiREacb74wpTYeW9wyw3PmvidKtI+BgFBMBACZ+o27agpkB64ognPgIT+zw
78cuKw+MJo9atvTVa4JdSq1VjHfE1yxSCo51mKlXRu+wVbwNaibEENGMTPzuFQcE5sLqpIfs52hs
YRUZZJxTSS0DlAwZXenepv7aoIBDLJLH2Jgffpq9ApSnTqsZMGmykt9q0bD3Ix6p5uiRG8ztegX9
XMJ0Io1AnhR6S4tbUd991rGwH6JBfuuNduaKHbtxO4KLk9xHdaCPOlzygwf1pGoNWxACzCJ2LNlQ
iNilayKdpQXknh7zwLZtMgqBJcQEuaLnQTgSsKV94rBXvnppcc7o6dQ/zl6quueOM9nBSeMvNdt+
g6dX51Bp7713utUj3L7MCz6XYfHgSB3fC1QLFfYS3YwHI2Zh4rxd/9329R63K/0HvQYwIqB/YG4T
60b0QnLj+cXVLa+tQbg76L9KJ3b3P9L1rNjBpkRkhw2td8R4nrnqInbe8NitceYcvsYvek+I+Hv5
96kSowwMxdny0HPJy9yfiMrwBJnOrwo8+Brf30tDQpUliHFx9WyO/ke5YytUk90xfpr10Zcz4oCV
ob+TkfFAdZfFWTrBwCGFgcMyrjHc8ST9CxERUJfzEkGBl13AHqCcB+MF48tK9MvhqgZrk8sDgBSf
Bkpxed6CPW7CyZWb+I0f6wcghtl3fjMhvUCLuy1S8cN5Gu+ehgVEa4YeYKty78IqVAjIMqMkOz6e
ZabRhYqUDUkFKW03edhN6MElz+3j+XNmxekQVa5JIRzKyzEtiNKEljajztq4QMIY+03z0hBVsRIx
I92qSh7FW01KLyY1zCQe1yH3pvT21pzQJzm1KxKOH1MHO/xmSoEZKWSZdi+Ugd5LPgL5Xb3V08vz
7x5zN8o/l/ovc78V19QDpd+PzW3I+aJrMl1qKaPEkRTwNkRrld7Untpa6ppOW8U+mXxYl+oFuY30
PUHmoNtFbrogstsS4NtghA4PtLQ9TApj+z9NRjjaxZ4AUiMK1svdOMSag3iK0xe4Ae6sX6W+qVTe
uROCaRl66ylpVZvPuqSnjqY9+lRdWmiIS49C1IZvgWb1JdUO/qI/yWWihAj/KCXyczInCgnO073S
LW7lntiDpYUeD3nPpUA67klUI1Ox675EKK8Y2Al4FIMXOWkmI8tbflKf2v7Yqrx9qjP2nGflkxwI
N4rIg0xs7gDKJ23BJJ+Iv9i2KBfWlH9IBbYUUJgF2O2FEXmnexNaf0TaR8hSOzS/kvd45oBsZh4E
SWXDwaNS69OMu2r21dubbnGDxff/9ZbKpfwMM+h46H3IOz77QiU4nsAZhfN5nCWONFrWkgACxIp5
D18mdz4h5Mq2E5Gc/Vvv5sUJJaC97tlFgyj+N+mFzKFx9te5ZVQMkWXxkgdVtuwYNBmHI/+pJ5GR
SEryEV444iQH4mItRforIUo5lXavVxNGnt9m7lwU0tguZxa19j2uFtyY/OBDr4n6Sa/RCAkS961s
6YtyeelvzBbEg2y6YaJre15PimaL49VnGLzyXcS0EKe4Jj656H64PPnOxRh83fc/lBdDX3NeWdFZ
ta3R4HLOIQjE/e4d//vPDdqV8P5bXnEJ0tGxVPoui+gG7DcEjdYnutRrrcZ4Q0SC6lY7Nn13zyHM
yuv9pWXF6iH/CI0IUhJWFUOLOSAXKoidYNm2NSZbaHxhJiNqMsJjmw4G6PH9MGyd4fQp2JE0+CAP
gp2/9onFBeyDWiSwLMcxw4urjyVOglzWIsbuIRmziD1CPin3/gPnpDvqOVOymz3ggWgMZTZ8pa1u
PaOYWHFXNMlCk+WkGVfeObJOey2DUOq9XqX7EXn19DkjxSdEHdBX/eYsp/8V5trI4vhHafRP1tgv
blL/l/PHUQl+3j+LtGugoO4yyN0jJnZQ2gKbPbEkKhh1jwjYwC85Wf/MfsnsnB80jgrOAtfNb5ft
8iTPRD5EqBltYF00bkMtbO1jPWVOrTfIFrdcM2/V5bcqNi6vbMuDT9+iAsodlV/vCGIuRWTfuC7Z
dOh3sBa2h7lYke1gQ+g19mJtIvgr5EbT6evFbh/cU66uiv5Fp812gK+kc/dPvPOTpLXlYBdkKWWb
KBAvrtbjacD51/IqKNh9G5A8K8UjM6R2WuFkce6xvwiGPmT39+D3ZT6CvwSqMAba9RNLuNTVJcyE
Z9qHAhuUqKd3QMqavDWPG90Sp02M+FHC6EMYlXu6KvQsh+dUBLWJxc4wZyziPFGRKPOzVOV8YQ1x
o6uQLUMAHWxTCBnbNwNVC0463n+aN3RmrXP7bP6nAdtU68mrRGGHSDUdgtHH7iLuJ57620l2cr51
96d/zdxMkUDniaiXpah4bB4wEGioKX9MMWMWeDIkWf2XM1i3HUcmdOxJ5hzS+GrhvcnU4AmMamQQ
nnb+kQmT/9ZtKK3VdeokJh1dZ5Zt0YIX+POTFvrqH1bcsMYT5uuB7ZbxphsfByC1nOYnl2SiO3hV
636UwM0ocXxBavvM/eqxykitt1ZFIvbq02jdpuiM31SqrMK/sYCTa0iI9jux7Ek1MV4gA5otaowp
qisF3dmNe3097st7A9iRvA6Zub9GYLn9Ch4QxgRsRDocKb8w7PtjmtzO/VscbfC3s1tWlIvaGz7H
RGjT0Yhqa0H3wT8D7rsLxTMNIF338H6UQn6Qhcdi8AmclWIy2GlFufeBEezKR9vEqY+TW1n2JLA7
iO54b7UIhdnY8hd/9i47qxyZHNTYb3n6gcX5L/kh0fq+rTOY/TZcUU7s5xHmIx4iPvJaL0sfAbxH
0iiqA4GdCH0OqtdOgK5HZ4E1BM9UsmyroRvxGmR1hjeiB80c0u1agQuGG0ERxcaWzfufzkusUrth
VCmVOiFvVM8YsnPreEB8bFe10+FdzFnUsKBpZ24ZjUcWo0pnkRJd7w44WCQX5Aqeb9UR9KJYmvgB
vy3ZJeWoj4pO+/T8LH+ysTPY6SLS3p3aKy38Lue7ae5iPnN0Wj/eIVnhu2Y192+e4Y/aUE6oTA4y
lflRsvE0DptQsi60N9HELefEZ9EEt7305WrWn3x8o5a5FppEj9SF6hq+6yPTdgS4hsrFFUkRBYhG
FzgTXSlxrhySc0E9KuxrJNH5RFG5wdIhXbiVmq+USawZU1Vmy1yLcX7irDPCkFQGY+GSajw3m1C8
sBmz7/HtDZ1P6hOov9J1XKtaAee7KflF32cwQ5UpT5H3Cv+MtNt5COtPZEhEijUChXlI2Pv3aw8K
M1dw4aqapyFFPmCdXRJJz0DGx9VXYWY6y+UX5OwE6WHTne8+oWCd2y9BzkEnFh/CjpzXHP62xECA
+H6NAJ8sw/KshWVW9ujTj6VwxNIYyOv0Yjy84C9jb4nOUTHauiPw1DtMlwWVp+UaaBO8jnRBe7WP
rwShih38YmUb0C0sHX3MW+ddGNGUoVZ43AL4XFTgiCuMhsmSMXTWJ8W9mafSHGE2+YHK8UEQZbWr
BDJpm0XCEUWeoXivFke8J8Yk+L+Y+wfXPMzjd++yenf2/TNRv2tJIvzz8E3ypktDYRNpV3jGW4pr
8U0TASo2sbFUDmFgTlVpwp0CIXZO12bIidvpa3Gf3GbFma/wtL8Y0u/dU9J3sxhmaDZq5Na4mJqb
fKw7qa1Cj2BbeRXKiEdCrcvbXQH1eRU2vgu1QdR7p741wZ3LtjRM5HXX8Wky/ZVaWHZhS/9p7Dq0
FQ/n5SSd1TRmf3S1/APayEavgdrfGcLNUfsxdtfRDS2al5DJDSFLBN0ckv/zU8t4geHH1SF/X3+6
VRNSK1DMhq/xdaPj/L51/W613XkrfYHwBasYrRZBKSRotl+JiFNTI+0YwMsgdIJbj1EdGIIlqky7
EgCA2/ePnwTgD4DMeZrabC7ExIXVUywBWJwr7trJj46wW2Tyuk3434OirtWLdRIaFQMOZPuPajFq
QaVWmdlhlij9CVx4e7dByK/8VbX8BCtTBpuEDETA4Aik1iTedY25AdbFd6k91yfOekW1F4PepNw0
iHlEB+CUa68FheCBPM/OBGVsVIM80lh+kbatEfoNWSY6HNzbNFA+dBTFfpwv1JADpUYt6NoQ4fqL
2iazjgBDYeb/ya4c2v2vdmzaTYRq3CzEk8BtGhr+heQb4ZFQt4vgiRL/4MgUcY0gKMEOvUGpBeUE
zv+Ql3itBkPSfFJISHgK2E6cBbv3k+kf1CRQKWar6aioaraj7zMSqO1tUz0S2Ig/0MzVuEooS47p
Fwk7HYTX9LvbO0t63O9kYexvDrM4CayUnkMA8CihZNblIKV36cEh0QOZOrjm3uLiHLjVaTEZFXDu
kFrT+k3OrxT6fZBhQjgIGRGlNPDjrXNL5WHv/gtsH86Ivsz6dUtG+8xdBwuQDSwpzal9D4J2K4DY
aJipf84U0uv68HxmgkpdfmnobsyhzYpfwd0u5UwMAiefTaQvUHhJTaxBlCFVE7giWiAOGhmbARim
Ml8jeaowe2YFq5LQYEmfaHOqcGNsbTGQUSTQ4M8WO64ud+Zh47TjrKeq6r2vwFx3jrRTPdcoBhAq
qQkcEWSAjPuXW5s9roS84dipm5q8Izv4Oqq2geTG0XXElSDyLvT+9BTeouiP+4C3uSwprZqDducP
4rJ2PDVRTLWsEPJvvDH9/3DxTFRNpAdz2RPqDgwm5dTkPG0saN3fYVRPo/BG/JDiTnSC7zwkgj8z
8DZ33N067QXtP/7ixtc99q7DjwGSz2OB4bbgYgBRyRGib4f05+mR8NIs8RIspjoH7+Q0J8a5ySCf
zuVO7iIgr8Wgc3iMZTq+u5WwycKbXqeDpjgOQgwk5VOGoqQF3WKpSWWJAuBpy4VQqPh+AmOxjc5H
Hv81aKbOPwLJPz29dvf5oANgtSzbQKaj+2lsI3E7nQClOxEzeHPoU7Has3hXbJmAYpQ7QBA9jNy9
tselpYkUWUwWSAB7eeQ6nGE+VgXQxgHx5rbf0oaQOTcwsgjwu/IhnS44FXrz3BiKZnqfe19Ogvgv
W4Xn0YQzDWdFgCFX5HXobgurp7eTsI8eqByQJ60/l+2xYY70gG8QmuvLRBv/LlGWwPzbrCY2h0aQ
R4PsSWkh0uV5kt0nGrJaoTBy6B0aZPqI5424VP0SHbRJoL0WYOXDiI0g1rLdSoF1qTDAN4GWn896
RL8Zag4gBJqFz1jIyz9UsQpEV1usTmiXX7PS3RRCji8jP7O7kp5lZ+htchxtjorUYqy+i/L3Dcfj
0b48x78ef3gKV/mBS1bC4fPYi2B4W1VS6MQZMJqaTs06JEtMEXUi1cA9y+yVyzZjuBoKMiD3V+L3
Y3hyoMwRYhx7w6ZkEjZVbsdD8wlqwOh0qolPEJTHwzQfR/YG/wc8U7YxBeOjBr93YD0LT+2rpU36
6po7sOr7alP75e9vvL7+vYQdBnN9OY7+MNkgo7OtY1QYKyaphBWDyibkLNbHaPfapChLB8KzVICu
Kbw7jJTnC7kkQzbWMQllV35eMBm65vdpAX+wA4gCtWWOrr1Hu3qQ7aNK0To4c+LoBMJ5J9beqJtC
oU6SGmhAc2iUuiEVooqBygeflaujiE2mSe0ByE2ZLO5lWdztHcCcFB2C/5SCcJXVOyXCi+bsoXAe
4mkdiP2PpE29me+jWQJyFGKh0807GKBdGQP+gWvIzXBf+YL9wVAmMhom7AFdCxc2HZ4npFK8dUR3
pmsp467vKSpKkBtpuFW8Xj25ULByTNtVm3fR66KVheOnmrw4Y+frgfeP2XfzCDHLwUUwFKPdGwKo
x5C6T/qU5J/thtG10JPJV/e/RWrnZQnODZVTAqeB4uVRqZnHwK4ZbwQ/SceIYl6+Ee02ea7lzYyC
gonekw1d55q7/X2SSFy3w2j1ZsxWTOfo1yRpSLzkWoPn54YYY3hQ/8IfIDpgvaUTwb859YhNiNL+
6QffCCd7V9SdVrxxXcXGeOBjoyZ6gf99yApHKUdgMi8yz+NBJn7tw06a1Xabw72y0Ax5JSw2PI4X
iNH1CipVz7WRZbAOmm31047R90QupSAqC8C7u5jPHBv9pZV0nPc73cLrZKVnuEFw91nWBTpNytHi
sqhvCbAC168eL9rl7oaU7rKqkZ3cJOkj/9ThQfMXY7+EcwAgSeLTRq8NLIR1XfXWie3xcVLxdO7S
crxxIwwnd1L4t7lloDF/QpEUIedKIyW8b6KCiwbjppb808XZ4J8px/surnZvmS023NV7T6F9XszJ
FrOS+ZUL9vNAQp9JzgKD6Xh/XlsIQqi7zlLd+DU3XDQs3QdXWjxHDnpkqIAC+Wt7aRGgcLh2uVBZ
kt7SDU3h/LNzYcMa54s0Ep1jofRzedIbs4CxEJxa3+ZlqT+o1BDq5S63iHIA/TgY9LYRh9zplqdU
ueIu7xywrKAMAoyXsSE2ijUnpk8UGWxzS+bZjLJT80oiIbGGHLALpVKpL9FsQlUYVuIZiXfBJkHc
bMxOIsP0Wo7aaC4eDABXMas7wNXlBVMp5eFgCWmd6YlQn5nvipZv1/2L8KprN8phAKQ8yxVRBnHb
ckbf2X0xtX4zLekA/UM+c0xtWgEOyj4bpdxFSHZCshHLf5UVlH1O2RzMZJvVSGlnVQuYxbdZDZXa
ifBZi9o4OuvWTS//hh3yXm/CpglESEAZzYM9vbLOj95KR06MYuqp03uyzfRkVM26RpQ1vsdmIgXy
35CZEfByEc+hcZE3HfcWSvAgNip9YjjVEZ8LWuyoFJr+EQ+2y2DJ7Z0IYOCZM7cl7X8JqjJOxGX3
m7w1cc2O2IJdvpKvQFcUWEVoCML44SQ+SU8+el954JbGVcivLjOQtLlAh0ABbysZGK1ymWbD2Z3X
vTzWvC/tDVeyOoMIsm6ZBQEn6UFwESHCkMoj0+aWwyNo1TtcpfacvU0HIbS0QQ94YgoQVSWSzW5I
lMvclezy3sG6//GMhct4PjTTxZVamLXNOjWCGIIVkMRcEkxVa/CARifweLcAI4c9l9aoqQE5S7q1
SSzera+6iiOUKBAfGGz4ncH+mVWtPct5VKH3XR+EnT3UZwKiKhPiFlW1OcG8lnKbMjL1U/uMZ9Zo
Ep6K+m3DPACquUm7A1YOzH+zp3ppNNWWzKSQMybyKNNRkTJyoDkmwSlm33rnJln811LcDYXFpkG0
RfAMrLVvIS4SPAYWBdpauKQBIloSaPfe3uvIuQw01QfNmbRmb3mxlPTCD6ZNYMp7O9ZVPVlKCFSe
qZCdyZVR3AZxv0mC/JsxGcVr+vIXH275vmYFqTQROmJF/fhnmKhuDcnfXdpD7IYCZ1SEfJBIkJWZ
ApEWSVAwK30QGFyRTd10Ii+2aj46IX1lfdejVxL1/KflyuZLgTcJVwhnX9xkdmvvIecdcJ1d0jz6
9Ozj9FDOL0DUFY5srJLex5MafOzQqOdfkvdMjy4VX604jTDCpo1NUZpLbKZMaT2alTZw06MrtqYp
eRDmZRZ/tjAoXDqwPtuAG/mRoPFXhDMlY3lud+1xKatfwiiE0GhvR7Fov0nsM/J/Fw86r2SI4T50
IUk7qaLzMSaUNM5qo0Fp12Im00tTlSlXyjF99MlAO4IAHB1vLbdFuvS4IbGBe7sB3+i92quhR1tM
4moukUW4LAn3ScRHYg28RTME2iGlg9xtazw0GBgK3Eg4d6Ek54CcEZ/8IdVPWBVrSzTBVilQGeyg
YPgw285wET1bymt1H0UWbjiLcSE7XsnXq+WM3D6Gy6iLoPOgXVGvT4zp36/xQT0+ZCFYQosD6ySf
cvh+e4U+jPeVFAUTmHLs9jTZ6ydPeK1zYwrQtd4KCDmTtfWv9uIsi84L38S5+BdSeziNqFo/MQps
e2YzxjDTjszEUBHRcupUhFOO+uanTSlEa+tk2AtBmMR4ZA430/QNh9p7XIZq21l/GGo/LFVilpWt
DLlmh0UeDzNaEnCkoE4vabngx5QKDB9yos+CIU4JQHhT4xli1Tnpa+7mzYnnwz6GhYq8b9QBx/rH
9NBHrBlt9eB7bX1dyZAMx6fgcMWHybXp3KnJMqwDCNxvhT9/oNbKgggVQX+emwq+9ipgdiRslXRv
olkkKrIrwv9SDLGZ+u3GUYZZSPQ7ZDDpUzDo6Esr5HW1Ns6kuFPxMCO2CCRaWLUYVq8j4g8eTB0k
ACXvHDsURXIhUVlB8onoriTSMI7pHmxbBPlCkYQBXUdcf757vEpvjd8jPmoDv4EZKBKfBvPA/3KL
a5qrAiWQK48QINsk1DnI0YDkdSdnIaIV7IK6ffUIAN4rm5oTqjzrlDyrF+Z8ESXKjqVaUB4CQbBZ
gBkEr0rnEsivgjOWsYLE1PVGV1toCMox3Y0weXV8BdeazqLk3/RuBNG+VOR1tRJ932H6EE6s+ZH9
lR+nIU/YV7LI7BNUJ3sL0aKCvG77Fi0J2ZYkh63ZAGUgiDGq6HIOdKDk+iEMjiATvi47KiqMPhr9
lyiaDBtHPVvey/yu3A3iAXhR4zCUduL8T/VCG+YNBl2qTDeq1HpFkWfntFHwbtJ8c6asqFfLmfG1
usvU5UZaLqfuhyoYR6pSqfvcCWchRgDZdfi6TdRWSl5pZm5Th4/lGaVdfy1tjLgX13ex1HwggMDB
k8jJs3NllIxwcyDU9SkYyd07QlFaQ2kI8L0DEHQwzPJ9iklytWmo72H2Zx/EaW+bQgQ7IH7cUguB
wrkrRTo6kYXWslQPo6kcTEr89kKXvBNaZyE6t2kIF2eiKwySKHQ9TIuuGXmedmkqZyNYnXdYDIRU
e4w+VMfHXgVaNnpgS+fFYqsu+cNFYsbWNkgHgoeTekWUtPpK0b3SMhcVz+L6MmrmpjUJdNE9KlEd
Zdd6M9sb+Ev5lzRruzqpnw8R06sXmLGSE4jTzed43AIPKkMW3MUIOdrssA0qA0qAfvSTqyE+LYPd
+vqnGOADj6/buyujWbaE2inM2+Ad1QdyhzYtNnIDCTuHtBLmPi84pAd45D4Njy1wOgWaL70f1rli
yZvvVQ89lUt1sjHIIC4t0cJ5SCrTvjIm9TxtrI2T8D7ejwtMJjf0KOsywtdSbDnSf4Vub4v6+0LP
JWh6bbsRcdKAgJ7TD7l9aUH9XNbXHtQtAl+HZ3mfHmJIecR0c1G0suVh+w7x2/IZYz6vtQybFOau
JZO5aMRyfZ7qSyqt1Yrkuv9AMhxUkGeW/aaIF4zzXCV3FUKCmfypnMzZbghJWhnYh53aXLu9fX6x
ejfw9fq5PRpPlIy67gc6fy3yfChJRpTItpP60gaWgZeNoUu4VF/wqnH+kSb0N3JIUVs97EpLoFaj
baLAATQUfspzjXDjDLNJmhgzAn/Xz2B8HiUKFX7gJ1aSYaU52ekkG3oOLreN5XSd35CoSBiC3GDU
g9mS8tcESuxVSX336r1RmHZzZ50tFnwZJDhGfp5eYif7xzYZYmuQldHBEWLAYdh5K87kwIk4omiD
sBE8iZFejJDsla3lUJa6KhqYIACvFRh1v8nnom5KLB9jGfz0Gi2aqd0FdZXgmg64814vS3wDzbaA
FafVG7bHxXsLY5dwB17D7OW5BAEAehT4Xyyt1o01mv02yUr+eBG/Nnfrq50W4PJxugicj4A/BnAj
CvLkq8vdbXuEMWngZZn2/EDQeCL/gY9lBDFbX3V+fBptp8wjvoEntDvla7lQPINrsJzzkQCgMdos
kX2EcH53Cj7znXayTYG2QcJqlct4YwYM/jcud0+IHnZZ0pnyN/Bmas7Gn7fM6aCHieaKaJLJmNJz
8wJtYveGNmwfGEisKvwjDWTtThK1hCaw0ix2PjNH7e0r0lSql/FNHH3UHiF9cYq1MTGizK9Hu5xt
OJtzCevGGG4IHR0KbFN9xfHKcGIHPVhoyNd+E7LyH5sVRL2prnoJApRxnlSjTchGu77b/2yxRm02
xWvz1zARt2bvRXIT2TQFDRbhP/V/VxBP/bB/cjAqhWKrvBTCbsqO6fMpft8XIFZu1iBIzlhXZCfB
g/T3W79ejcZk5WY/yAzpm6joWgcdHTgyP74ruDPH3L6IICh63SL1X7olR7iOIid6bQCtUeCHtsYn
LT9kT7Po394DRIZug/0zRQ7XhbhHe5rnkhJlba/c2x4fnXS41Ent2TnMMGTPbOUEEQRB7r4ql5ru
9Q0dzp3myFMRTZSwkjw1okgIxsSiu1pvEEVuP76hpRBs20v1R6g1P6zR5EP3p+SD7g1gG+RJB2v5
DO/hh568WrhDv7PF/bRUxj90ZRmrXYu1aTO0bBAZlmdrWliBDFY9s5GDZ23+rtBvJhXxHs9v+XBE
oBaTKAzuvMtQoTtGZ+KYd2LuG3re8u1wq4JblEt/e3PnN2OpT5QRuUKEOKwxCtcJcHQNpRnjdxNk
UCyDTvTuITuSJvTCZQHOFt7p6t5GibwgXR+WVS/MfCxfzCoFNByfhk74PGg1p1tuRS8fC6A7smc0
7muju3uuvpO64Ri3m1kxfuB1sOnAw/sOuLaEpz/hStlDnlle6EFnaljxhMDJHAmmWUNFDq1byfqC
ennfT3p6zyvEAEamwA3cl8eezv/zDgBVgkq7Qsqwv22JGaDsQmhPKaV11yj8V99Q+tPulJ1rFsqx
WR5fhLIuGOmTCS6NUf7k+ckHh0xxdOzg8uagau3gvDwzIUNW2b0EAeNhshJLZPADfK0mkm+mgm4g
Z+KP1/c10B0GNPcoOIR3CWPq93h5hJNXao6MakCZf2jWOB5fAvV56JIx+NHMvx2K8E9kVqD6aeeL
9RGn++qMWcppFByXEv038nvNM21pu4OlWZljMT7htQt4S2J3gP6mFPNyKp4TL7YvwNpFmLSRyk3j
W/X4QqPnuxJ5hhPvC4VeD5uI+DU42E6PsMCD3QcNtvx8QyOk9T1sNlooATmNQwyDIEQKXcWMU3hX
sNEYzhLxkXWcTNaiMrCL3YNuRtSBYt1Qczbw0Gw6ENzTbczRBfKzktc8Z86GXNikF/gRKSnvHCCt
EQVlX49JDs3VkhqYIX0lHtGORYOqzJkpWqoDAG0am5Xln1Y42tRFKC5HO8qP2LNMr6hmDvtgUFN2
Fyq4yY21kohdYwbPvrwnEp7EcNHAbOnVZbU7/vKFFhunkjmGOlnCYm21v1xor3J0fdUPmnavkTpP
ZwQRzx9oprz+dIq1JdCaqth0hMYVdxZeNFNf5jmjiFhQIP91Mgxnt1MqAaY9K6YJkJxdxxZEvtsr
58z+GEhH1jgPHcH7zn/qBqXA1K/kvcRngUs1vp3wNaS/mTHPFvhfF99ZSKh8r+9g6ZxFiLiN+5Ft
/mkuihwuWda/bSiEtZIilWd5aM394Z/AwTzWaZShILtSHeIyMpFgaIEFyL8uqDXsJYqOPbdjHueX
ftPsOvF3CA44bqKZcmM+kT4Q/+NHtLHlYOjTfZH6XQe/BsMVby9KeYBn+fQGsFBpEsoEuI7H+ltr
pscsZ+4UvE2DKTGMPxjHK4NaPvOjp9Tl91Hd46vwm2QqArMnhz2CV1+CRrFsc6Tlrc+YTdp63y8C
c/QDD/G3BK1DUtIryLrMSZy6+M0UUuXK5F53tyQMp+H5NupKSq9az1lK44PGt6Pajobg8PMsjJBd
GGM4j6ioxeQuSmlT+K5zJCpvD7tXpoLKJ2wrXtUsKO9lAFh5SjoT/37Vn3/iH815MTiVMoIMFudK
tBPUsh3Km3Uhx3WIHdj7JJpA5FGngfNQ8In0E0slzYGGwfBQsZc9RkAsy962qH/vCzRdLy8/qFOG
OJpFTTohDgPUrEs0jK1p2GGqKizW1NsEkjIUwJtU/rgefUD0zENFG3APwUfmQytvWj5xcBXQJl3h
RbYAuWDl61FrIDFU7c0+sRR6yOp92ins4mpO3Hg09csont2955ZMq+PdJrci9ZOZqiObQVP9Mp/y
zScWO1xoPbs0FYQL58fhpTxLsUQyvv0px6rdyP3V+/Vey34VxJG8vPNI7u6her9AnNQ+H9sI1wco
Uj6zLyGD/bl7sgbrh6PdKqRPWwTIyFiJZFuxa9a8YHEKRyPlMLfHWvXLBSYMBdt+Pu1Bm5uuelIV
wFizmfS5udGsotk0LUsfHBYKa5NT7dmLKY6hbOTA+vQnCrHvQ5pskF+G7uLUuAqYOpn11kIwc1eR
o6ljAiZ8NRQYf4PpSvi4cP9jNWBXTGTqWgwEX1uwWDsD6SkyUdPH8hZdJFlmNQPSHZcFuVvV13p5
rNnzKRQAEQq0NaHJOf4731/MKAq/63/cYtAinb/Ehj1gDuSKSucrKlilI306NNZ114VTkiRe+75v
N0p3FUubEIQf/CZyJh8iM+0eRnfWoZP4q6kLwNyKAcGRmwM68wCDJDPq3WfwD6BPnmxwKxb2iKnS
QDgVCMBncy6m2s7wlMtE1XZGmX4VAakQuhEf41BZ1rPDpDE/VX7SNhnkRiCl6sTaFbzacmcIQnCJ
ZOrTkozpZ2VQRD6M8W/OCbxzQ7K+5/LjAwXvt0yWNIW3W0feTyqg4+Pj7+JhjB8S6ACzZ/CiKGQt
FfsRc1pvPqveS65Zf1c6Po6wku1fBhfEYtxCFC5yrPtuIoadDXnoo6vTN58v/4vUj2Rk7l7EoOHc
7P7XrvifKMO7ffHnRLZ6Tip1YTR94lze3YEcb0njJ92u95cgE5PF6uabr2rPLK9699ec0pnafMv3
Dkf/qefsfgXuSit6eZnaVmz+/l+3miiMFjcgZanUxTrxFcolhTkA/+tISwCQJpcpjt0JBKNBgIQw
9OigXw7dCa7puXhLmBHJYe8xxiv0sEhxayTEjfYF4gIjaxOwKLkgUZl3cRr+L0McunaCWZBIornA
S+BMy/i8iDecVGkLksukIXfiOZwD7Pro7fJsZ1WQx/iUwFP2IKVIs3xck9Eaw5M/wai9PrMUyr/Z
XTSCmQBTCpb3R5TiXtTtv/RpFiSza8EAsGFeni1eAc5CzBdxbcMJ0KPlmfrHR8fXuAf0LCgTK2i3
32zDHCMpec8vziIRLxvQq1G5r6PVtiT+Q3TecscEL+znGGpZ6F0IsO5E1bWo14lzr6qGGOVCDyTS
HuH+BKuSi5xNMw28i+3QN/c3Uv17Eu2CxsDnSSfxRX0f2ls86QAvDoCVL+7Q2/V4ng1n3ueQJrC0
V9t/bLXshJ2FokWZRO6r72xTBS10rY+Nfd07ewALDxSIr6WnrvMd2yXgQvHNyWtqWBZ9zgzwZj+G
U8yFG0YOU84xJQJWfd/PoQykKm9tObFdOSCWd4f51TtRkAlbFO7r5LDmllMK6KllBBsYHaBsHzKR
QtkJKTeA9tMdD46XRVJK2HDANBEyKRVPhJTCHlm9MrTPCBzQlvcg2GPn6EsUjjDph+RjpJKPoNm3
KIztAbix+C4j9rOz9Kr6M6bBmIIQx90I6PA91h85XB4Lerxn95HTRQ3DUEfXoeHax6aNJB/oD0cx
UHoTjltEJXESHqOuLJkXXXaNsgV9Klmb1jToPr0dv1mEdxh0l7GtcxLIsOGvS36KLrPaDYmwZL3n
4OU2b86pJUTnQaJ8hu/8uullClFNSNeO0y33lqWjh/k6vAKNNvn2NU9n7o9+ytpsUSGH/Ca3uqlH
vZLySLEOirquIkbeLCVaTRIZ9/FO8k9uQ+goga0uY31FJX4c2Fh1vzNZ3XDhU8qmSu7WOL8qaL3T
Hdvf1S4c0wUCHe/9I3e0vcwCGv9G2A5Inx70nDQnBBxIAAzYWLgUU4GczeuopIPuS6I1Pu2AXbhq
EUmtYL4Bb85mAR5yuUobhqo0iTOe8IpLPA4buU3kHEQiEQtnOQ==
`protect end_protected
