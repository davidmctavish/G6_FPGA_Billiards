`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QtEdBvxo0AJmZWlM8Pyu692KA85vDyKkSiNiwKutaDqpg6Fl6Rkf0p+DVS/iCXR2e0Yw8oorKl1x
HioSTExJmg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
M/rSH4ws6Qvl4e6Xcgplc1YOepzhryGNdxTcGXd2VDTg+MXeCfFK9R6UaxxzE23Am/qi9j/rH6qY
ycRdjHGUWHElwvOPyEQiRzLcwfn4JTOwZbrbNGXk9FOYGJYwrGWNNG5HRyV++t+kxTFoysh51MBW
KII1WZ7QFPxlmb/oUYA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Gf9zc2yd53XpujNrvaA+55+xgM0ZtbmnQAVskCR86IZ98IpZK3KqhOnzFpItzYwofXQtrJ70C+gh
sBlSTb9AwtvWOszE53K4Ty/ceBLGy/HY3BPymdkszGBECTeEEOSoo76zuTrtrPpdsKQETi0ywa85
uj4MxVHz1k9WS4qja2fH7yzDjhKFM01zNNFf3Jm8yg9vEeGWdEuPimv549MaiQp0Hf4H2wffR1h5
lPHZzFlrJ/lWHwHaugNLDKKzVe25ixZIlKxBlXdgd16QfMPl4/SKTuev5ZADxIAPj5Y/RrL2I9x7
UQSEkPl1f8DVpZ1g+494E36h1cJNYVGeKhhL6w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ekNzu2garNE3vM/EyYYHSHRt45uAdUHwyH8Y6Ji0dE07fvU358ul9WEpRLxFprSGq2+j1KnpJt5f
CPsz6U6COLaJY0vm9Lr99baYsgpjV3vwqVCotgHAd5VO9QdzvyhXbpiiZOkXXOiUykIKCJiwmUFF
AbYog7l5WWUqeQeAJLE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RMWzMni3qLJCKQtaL6U72jxVjYFAM1fmnx086iBcboH2DHhNVA+sfb37BxDWRT4leTKwBJ8HtYe4
xwAKVLGmbdo5PYlm9J+EHH6E46jpmOF9HsNxMHiU7fECZSc5NZv7xjJ0ATqgYg6b46b8IpeJl5QI
GYRShiuaujoYTievp4c1ygT8jENpDjEGxNeA++MuRLUqK/QSZctEO3ghEAdOX5xN696qAgLjW2xc
gI4FMngTT5PpkQWiSAzUMVaxApt968mSGxG9wnhWIFIKOlzhs18A+9K+993BBr+eOlp+mwVYFkuv
2mD74ytGrh+nxtvZhiWOC7hrP3NVEPt1cWmVGQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18432)
`protect data_block
EENVSZcfsLG5BWNn1aqlrdDSK8vf5ahCntHS82RMpli5GGm9u+tJGp/7nLW0wlCxJ2tdwpq2kVwg
0f76Za0Biy3/x9+d7IJ1d/YlieaWU6BckOts46ra696zQn/OFAuBxqqNF4JYdamG65JXnzHcJJ1M
h2BpdLzpO3ZklLdAyRH+IZRanX64mKDJLHUM96lOZ5xhpTbrtl32FN9YTlXqXDuBQ8F+cHfPH7JR
XE/2wXflwhCbEHq+1brdj2mL3fuq+Wad7VsclC1bHcv0vAj9Jz7PHTadCum5gPLhw4c53qLR9TJv
RRc4HokBEofXqzFDhB59aNRw6/1pnz/h6vBHu/ZTIgSLUBJamWRDwZfNPfIrE9UNqQxn9XswxPuT
vOo7006wbZ+2VDvfz7gsSTZuGupQTJm9QotFhKd15qV0VZly5LKseI8GOAVoYmPNeJE+6/pgd59J
KDZ7ZcAnFOd+OZD25b/VLApduhqjvznJeiogiphC08G8Yr+LrA1fA/cAo/f6sRwblBs9UW5FbApL
QpjVy1of87ZRmeBbfS+hpvKw09WDExHMXNx3UD5qBv7gyLV/D3R/o4WqFsr7jziQFMGv/dVw6CPv
/EFqFPKEu9wpLAjH2T3fWGxq0bkF9DhdaVAo8Hr5GhgvbSSrBxOkM8CodJ3YYTUZaouEUiB3ZsXJ
o8/D8+XHvumhY2RtY2r4oRRhkBX+6Ga2S02+p3NOrqTLeD7PzLyir3cdrykOkKfW/VTX0kugnAqr
Fahtk6IQ4ZdTYV2KPj+r6TH8AdzB7dNo4bzUEv6IhQwAtNHhHEjIuF2cSBP6qA6ii1EN9o5O7qUa
wplLm4ZE+Fvj58JW/sQhZlAZQ9Y0sIw/mxPDWUXSqw28L/miAADLqLgelRksfoyJ8McEN3EYkDNC
Fa2jUtrducRkbISXDLIvdNvymjzY0dscwUZN/Ug2Zf8M1yxjHxOTLrACJvGhwVLnjFprOptL7QPn
6pPErvXFncs+fySg8Cahxy3y+6vBPE6oOqb0RvggcYtAgRbyOm3rNTDGtSh6G5pvZLb/GBVv/As1
BuRG31WrVVNVssRQG2dvYr/s9xb1c7IE4MVYKOnvIVmBvotH6GFku8jsrWHhNoJ5HsxfiK0wXsaZ
29mxxYZYORxJgp0kON5qkakd3JdTGFw1aWk9ORUnTh/wtsR/W/sxCCEia2H06zwVHym963V5ImU3
bFsxP8OCS3sCHIv8e52i7dpKV2ajq3gmZ0OqaFnSwIUqpJ3gK7M2knefHbCbH0P/2pYZZOY+7v+U
6uFbzDBwr0cMdHxEQSWuRwSclKwaVHuQ+XexztKqb5zxRUjdvUOO1dK6FftkFZWfOOj+4gpqaGj7
cWG9q4n5U88o6M9ELLxQVfqmmMzr/mF0zW51XmpocOB8YRP7hJiSqYxBa77f6y2d9obaVUoyoTny
870j8NjxhIkK6fTlgi6+DMg1idaKbUPNsreI26MUi4odhCA7KWK4VcY4cC8BqEra/Ffte//jAQyu
WJdSw2KF8B752f7un1TzXKlQkAhfJyAFqfsCcLdEV2KggHlSaiZ6RSaKyTb9e+yBrxsOMMLvyx6T
jgB0CQ/rGNW3IOU2RT7HeGcPs+FJl5OnHf7YjUlPn0PUEb+I/+iS5q0l9wWC73PG47X7Q0XEDqaj
SbQHV3ZPl5fFTTZDPHF5fIIuoInbu1lbdKZWT/miVHDzNsRm05hSjWJ90Mo9tpucL46VkDKpobux
Fyq9OcE4TSM5nzDFxn38D+uZoDwq8cGiM73j8P93z2WSHoFnHDEkLKY/Hkt2aV3XRIH09kV+R1/X
J4K4TH51knputPJfKx5TZODvia6K5yDbc4rzeKhVehxl2VRaBc9lT5S3YjNTVV7mjEdSdDfWckNF
k8ARk2KYnTkGwMvDv5FCXse+D0cSUIpJ2NT4NrEa2LkHewsYRD1/HqglEGh05BGHQq2q4V28Aity
w4htueI0bjFbwJz/pyBNEVO+oq0IKEjIyAFHXE/VD4NEHqKHRKss+jqFo2ZPDizbMfuc1x8sMIMl
7JLuzpKFGClyIwekX89OtyVcNORrnHZtHIZzWTXOpTjPl2h1GRhrvRwPssR2hJxM9+7Seg1CnQmg
4nMCYVzvwpsqfGCVtud/OL62eIH4PX7qpQGKBcYTW0h+J3jfVdNoidowfXM5GZyveDq01HqYOnhd
M4U+V5fz/Rd8RNHZdMTJs12TuVYNI18EYV1m5pD5XmKzNIrLlhZqs/MxKc8LvSgrzXks/zKVF8JH
8CropNPMzqmnH9eBKSWXRp8jzIzeJrzWKvOyp7VYwF49th76qrZEdKPG19bq+ob7V+/pedEPyvaL
sbc2KB+uUBDJtMOiDUBG0MKMIYUnqRr78e7+2sYy6TBH/DYvrYlyKtXUh/zo0sOSqHVzXmlNBvZC
3uIdHCk5WFoZ+DFUWHIha0Jdmy1A4WZCWcyENFuVGW8NinnxEzxS797pTlMbp0AfBu4IG/6ceia6
5qaiDHskHPrGH/cR8/lyuDIQvwf+k8qhJDFZAtpBqGQfPaWaGO0bLAxngQ6DivBpj3fC1qJ9Xnqf
XNu7kgBUPghCOv25oLTg+Q2XnZ9hvvGXsbdz8dfkdLYn3B2+ump7Wb4vcwJfjPp+I4KaszCNla7R
wlAuRCnPxv6V773J+hwaYU5QM9hHJjO8wEzNYTF6gHpA0cm9CnxlZTAiT1yK2inow5IPkqXw2PYw
TzgRJ2sQ2Oa94izSGJTK5fIqEJDBEH/ySxFy/hGLjYJvqT4z9bHzXXgvne4gafINxSNKUiMX9hM0
J3kA/6Fdxt/1oQuMtdKQFVGm0yaZYohs8zLCkgc4BdA8dGLuAXBDp5KPQPQPnQH7k/yr3MTCkGzM
fisnAyuLjhT40DTxMQV4AcCOlOzsj0uxt72KeLyfdZxHOEFljMOnRvWGWdzTwqK1sN1fuPQl+I3e
bu5gQ65mzcXxFVyroE12njH7CMLQZELMlHmHp7iS/6xkGOpRYOuAUknwN6azmlvjlHvrMN2qCE9h
VbWpZKRf2cqVLjZNRNdZYvJLlWZvBFu/CBjP3P0b+ghMxeZpPXEWhIGtk+zhWhyYqIRs0bhpm3uX
bvX8SbAunllT+ymKVhMJcLA9r2iUs5MuWHQKjzdBnTQQEBhZy0ydfmWBJNniua9n6QxmT9Xao/dl
vIZcp2pwLehK8fcn4JNvX/kVcABOhB4R1dznp7/aBSYTe7nid7uw2bmcDn5JfrwZaPk71BBsJ9c5
v5KTP83pL9EIm+Kd/0OV4nwsiVLO2Z6CgxZYKrhIInAWEJSrOMddvCfwKUhzC4bKk0JuDKR9WidX
+Z6ms6tieKLxaMT2hA5r3i2gWQFipTg/FvdGG1E1SvNGHBIK7ou5MO+xZMa0tNYrjZFgF3hnbzbE
lmXd5YD31ho0W08+qN6V4nfndKv+x88TsR6tXkX83sNxC0ioFSvdQsYXgI2GVYMG2Q37pt30zb02
ZS69hUfiYffAQMR8tj2lHsW9OHXjBtj0Z8TNBJsIaB5Q4xCoB4mAqGnW1CsLv4rraSA2j58CXdTG
KFE+pdajs9FkrBW4cT0S/Fnyl83GYefoOXu5FEDiuiIbK/TtUato/IxDCNq7DY44S7Tb3YThzDo2
D6z14f4FoDtMnDuc5zIaOfGESClQqkLwYwtmsFlpRhFxc3opOEI4I1mCJRQV0hhAB1xT5UBryOCT
UtNLee6IgaG9to90JbIj5UzetklMQb3QPGxlFy8S+R7rYGx3tCcPzdIFNDnQKOe7G4mdcYm3LyRF
gPrmir9pW44YwsJCCkBWp2eYyQTr4e6gONQEKn7+jt1JnWCYsq4gOUqMARsilfBsC9OOVRC/QcPG
eUg5Z2at0QOeNpE5mfHccHDa/QWjhj4Tb1uN+Ky0l6dS3Cv/xzgGdSuFf1/4aItvNBTCrRU9IQtp
xfe/MBXagpd3pRkujDtmpcjkcLzC1w+RYce4HjLaz9Bf9k30BVVL7RO/9NgHqk02l/sjXQvLmgGi
CIJJ3DkBVgTWNfRCHSmAoVbVOavnQsCvRC51KuPNh3szxQ2vBqmWCTVvo2dtzw+XHDUiCavf+UuW
1OmapR+P/xujlSEWAtMi2JFPi2NslnA+/9/bv4rS39i+KYds6EMtIR7slERXNCctnxfM1PMtdaYi
lj56m5BVl6n52+uNvKZFLN4u4L3SxEO2vvitQImAF9XEN9dPbDR1ektk6tbJvYI3ZkSlcRR1rhDM
o/os04bO9yKTT/a3Fs5zpwXIAEUfqJESz+4Wg0bxJzudk4W9MDhcWxXlF2kvjBOEX/sASiGfn1D1
y9lCIjMQqCQbzgUmWQWgiXMM0J/q56xe0QtZhZbZ8cCeUVduqtUeTjqPojrPJWcu1li2RswXJskD
36hSvVjGp0mE6z+qh87fTIOdxGF1A1fLycLsWLIMa94dVd1gN2rDCXBQQVuqHMfaY/sp4klExZBr
+jcwIbctQKza8+Wvgr8qAeSrlNgWPXv8WyL+fRPKA6Ts4blKitoBlmGXkMPqAt50k5PUjFRpHKAV
zcrtQ6GM/3v2XnROmUgWpQK6wvtQIiVnLSuTQ3lf1IJXByYdYUaFVm4i7B3ubLK26XeNE6cJfBNs
29PT3QuGdRX+ripz4f5ZuKkdLXw4MzjEkZb/KwMsnN+4+CunwOuGM/zTGb+iYKsbh0j3bp/ZkFXo
YGcSyjzWJWtyBBl9W7cU7K3kzCJINADlqjXO9w9x9PvfMBBRQVzNnsersYBJKVe1iaDd4wkyDi9C
EJu5YvSEQcxJ1OERZRRmUrLKFBEvhxpcugvWydMHp0JAAVqdRJQGY173l7pvAiRqJTfLeD0d3mOh
szCM8e5TPPWM9V25zzRmHIcdzj/WTvmrPehgd4Hg27zFu3xnVUYi3uh4jUIxq7nJTpOD0fQa+8u2
WlLcD4T1jf1XUIlnMW9mpsuKyNuiduSlCYJFr6gR5kR1lSZKnrddyP//7Hd/cMV6LbdRT8MaDXTC
Gf8X87ccxdUzCo8JDtkfXBnTTffPjeJ3qOwAEgDeD+qVlqL4NR9P3GnMsue38VF0kC3CUklwVom1
30AJ6wJNkiG4mslxWp1Y5QbE/z8dNfR4o01F5kLDq9rADrn75s4GVjkrdTB5qRSTLjVXC325FNn8
cVc9SIOyMexR74w0dJ5yLyRlC/OES+xasddPanDusOW5KFmp9ZxGInipLkyiP6UfK4gqb14g3W2H
DbTjYypR2eCBy+T5AW/IwEbsftVmg/mf05iL85JPeo2Wl5jp4KUZNrgyuOQevwiUWK0bpyn3JmMl
l3ojaIBJmIvCmxjgiGSJRh6eZ6qpNZ3SeRMxEEL+Jl7pFkaD8U/IfGuX7bee/Ph85qBT7Gstjnkj
CpS3dfupJG2JE4jhj2rRs0FjYLitE43ju8wIk+kX3vRz7xzm63M/eNC+rVwy87EF12mQ3CMjzaMM
XENNjSvxL12CE//Pal0O2It0n1AtPVVUR0YnUpullbvtTfZxjoEfKQuwhKCg51pRRCX+7SlzqopB
8xa/lmLNMXQytROUQiO0taGcy80XHtaZqzH+cLFs7B9jlgyf6r4tlTEW49uAtmM/CRJWGtIDspDV
wXnfQWUR1snZg2eEol6kFzzA6DPE/gOXkMb8mm/g6aLNESzwrU0ZdT1pjvpKQVEvVtEuRvpaCrc4
gtOgfp3b1VYxJ9PlHWUh+u3TixUSLMdw4NDv9Qyels4h/k8P9WEWm/KKjWq/NW2FuH4YDVWfsRaf
Q+VB5Is8hJfOEX4bDHxrBLz0e9Zjs2Sl/zkhWL+RpLpuJGGDdUdBAPCCRjEYcxbn6g5BXv7BeLar
JpbJ0Fq1g+0f0TelJ/WsC5n1c63hCvnbugMqZDrSTZ9vQp5rjbeqthmHiyy62oKX0Ehn0eie/drW
nmxuBa1lPEo/SUCv10yovghE8v+8wYwdhp60KuOPpOd3ZBpzAGfhbTOogYU+nMRH7J47WSijwDnA
zQnlDGf4Pb95LULZp4Hh5Nbq8YR6f3vxDLaKlUaev/if5WF67QNq7AKHcyVbKJ1CcevHem1Ki2ZV
1b3oKGLgJo4VqkLgrbJ3V20pKzaiipev25KypCwUrqTKPcdm6pU6k1ShNXhSgs8EHEMJTX7m9lBO
m62r5O7jd0DoWXn9LE4tpQQwOKtfxNTLt12eqhBeb/oWafdqNbCFhkxDN+eACCTaomCRPwmXWJfF
V3kd9Opyjzf6Gv3DCchXE+d6SFe8y8fx2kJ4eScVDmIH5fqvoDRJPbFJRNzIkTMGSJYq+l4PP27e
46hocu/YXaV3wCHnvlsiq4rxeQjO/bwIHpjJNSbzIFkcUazAyLqjZGEMWgx4kBTTJUhbIg8tGfdw
wozeM2/7nnkDQISW5IvlIuY85EfnRtm/dFXkQ+btdTuBJuCZ8ik4ji2HOF1JR5MPtXAKNcyK4s9k
aTV1Ey81gHfcUzpYTlUMGPKt/YM0D+ospI5119JPfK65Bg3UElXSd6RyjYkCRheOgJjlwUsLrevl
OAktFSRmAqQ/B1TPYCZ+bWjaZNcl16rSMr2ClFMvWOQYv7VScC9ZNLxgOUCC0ho3h7e8NSWEcQxD
FSd3qQW6axit00naLaNHp85dVbgAXh4Tgh8dNodhakBlCbKvWaNJDeVPzT1ZG8JVAiYcGki9Rkdb
L/690WeBoCepGf4OHDElTBaaDVtyrHJYMcw19T7aeP+Ttgj7i1BSqV2eweF+cKa5lY8GXbkU5rvx
1IvvxC6Cav7IaL/8yTI/mjjW15R2tcHWUiI74oR2rcp8xIcGmP6XtNhptxH9HWEQQRkqvc7TQOXS
at+SrKw0ZaatkdXm5o+MKrbSO7Qp30FDed1CqTHOSQxIk6keAwozuMBHWzSXY1C3aiiYWRikJjBm
Y3Dwkux/7mVeZU4w01kZsxWqr2vUO5gwyrGFYAshXlTD3MsEcHT3Wvam5d+vGIknwtm7UzQIyrOn
dlsOwGdDb/F7lpwn/WysX23PESYVCt2dzfXmbIGONXesjTub6QQdx36T40Q4i5rtWIR/1105LpeS
jltpC1lBo8GSVdziQg1wYrXGBvYtvrP6iymkWMiWaqTecpmtZP2mZVlEykst4h65Hbqvr2v/A4WS
kWEi5QRMRrNb358UG2EgVOHGPrtSqqy+wyWNhyKL6mcmgcgipsw7QIYVH18olMQ4mkd8iVVkIigC
xvtI4S8RMRX2urWXn1JMcxVqe0y/1FA5RCPvIrXRYUf6cmt5EgCgnhwrHBMpN8Yigp5SijGNZVc5
C1oYnfGCzwHsMnC/Osh4FN+nD5//aTuf/A2pKRMXe2hH8Wh1DRcNaDrD4ltUN9Owiz1SRFdT78NQ
KL8TSrH3+ng6rwIRWOkbTgYtCwDCDbTVaJKKfwnUOBCLASyi28SrLT/W7sKCNjlVS67y/F3uQEvj
I0VSA9O6Uh5jwQVtIgKD/gr82H/1EaOGwE62sLqPrVm8tIrJ/SGgOyIKo5pKqANL4ZT7Ys6rFVxu
Wmq++UlGwBhMFKv0aA/LHUgjhz0Ers/cbzI3ViDcWXSM2pwE+7htPY36fba9TbUeZPCqRELtzp1F
vFL2RMadE1HcUoeXi/4iU1hWSlBhSpIU3rAYgEVz2uRQCxGh2VlXBDybiWAUcVFSIT3GBmkR1adE
vVBHSMPcMp81UlHHVU55C/A/hBWKBkgF+ZeBxSAqIGcV/uvlmkS1Bd+S8PTln8SHrspvKU3u4ord
0+eqTvgH/6g6ONUZ58NW2rNmmN3hMa9b8m9x4E9v3oN7jkUzSRo5vq2zCKUxbaYyp3yL6/7MhdOi
nUJshRjpRLVAFeIAJ5qeyDYHX/0svDQrw3QmXAEBUjyCc0JoXwg50s/jQ0/nQE1Sn0QnGOKHLZ5Y
j6dxxJtcB1orzvc6rCB9nqQN6+VtOkCj7sM8l9RnqVmQcPew8rs2awMA+ueiR3Wa8+bStoNOjn/e
oS+iB4gWrL6OjfUmBl+/iWPzP6gdpGXbbg6FrHIt83RFd9AscIommm8DjxVNe1cCmqHUbqP+25Pr
zmZNwOO33XooQgTG2Nutg0FMcCOtD4q7wWllLA/oYcZOq7IiwAGHcK2QhnhPunLA++Xm8xdjVB+b
hApZW5SVyPw9RDn5QctvREeKwDP5jLQFaVvMUhoRF6qpTQd63wXng5fNr3Vefp6ewmgu+x/9oel6
A72o9LjNIe0QV88Cp5sYMNm46eIpbIL2EHE0CnXz4TTWzKqk0jgFqSFaJh+tjorH4HyzSlzJiB08
zAY+hEa4uCXZh7vtNrJUp8kar6nIDvzDobBXul5OItZhL1jIcGbjSOVHJGrQFJG25h4MJZkypzAD
0tg6QVc46pnTdCC0lddLM14Pt0SEcld1sidCuySCDEkK+CUxucFOpXDK71f71r47kZKF1//ZsRE2
Y7/4yUUo6cfTtizLKoIS22t8CearV5dQNqWq4TOTg/rVsyudeq9yYy0/z+xiVTdOsSMn6Ih7vj7J
n9h7sdiW4eUxE2SG810hzatqB6+4IGYDkZtx/meqIclpTfeB0VD+gb2XGYP1gcTEn/sWLNwR07hB
lvu8Q0cNs//dqpzylk7L6qfUZMUyyk1ET6z/uzNlkX+b7LJZlRmzh0AIRp8yRJ9BqIRDSjH4D1Dh
ff/ZBJhTHUxuYbddEuk/pnx2hVZF2zHB8kTfeBtTLusnU5qsDn3OXOtzwa7HJosl3pi+7sNfQQ+P
993dz7upJrwwFZpnG2X+HMSTPFPQGht8WlGk32BKoNo6bVbcWJPWwesDe64UxpGGT0kpWI5/qIq4
/6K1XznExWB5JNuYkXo9OWy+yx9GTd44X4ZjzYO9YiFkyarTS5loR2uXFnMN64UoOwvsHW2GdJtE
OcT7MaCQwTMPlOcuRJ/xRQ1NPrd1OeH+97hDeGhg8KQ9kMkUfI3uoWmw2smaVif7OkS4L/rEVt2M
W12jeE6Iolf6k1XQ/VBDIp/GIvGcr5dRYvvDX4MZgpKEHXQIdGrP1vQKur2imk/nbmoumwoUBytE
cbad9WaUjy3qY8Bj/Z3nYERUO9dpSVv+66ecIo/Gua/CpxisFIzRavdqClmUvPUvvD40mwagMEyv
/K3MvPznfSbihVKLVwOV7iswFO7recPJ9y7Q/5ilkw+3bkrfuztFY12PHhNOFF4TY1suKxxHAhp5
vW1HJV3HC9tN1piyH+1qgGshWbx744nNi2MgVP0C27JNlt7dz9nEiQyoSIDx2nhhJr0QsZt7zHRZ
RXyXu26fVwq9ZPBaaud2i7NVrfCfj+U2RZYpqHuUh7jIwRuydPtx4Krxs+zRULCL3FwtNHeNsLw+
foRRyKtW5R1LrRSdrYCuf4tQAOXk6634szkXzUtDsdr/E7W7FqSOIBDT47de6MZgDKObcOBoaS4g
exV3mU6UzkqSaleICl2m2GU+HbC4eqT/DUXK0J1523AkWFegoGMtB4w9mzSEcm1HUHFquqLTIA2Y
LgbJNaLyj1HVUMsbIykyJhyZ2ZDoVDYSLfOJTNn9XXZyQz6UneCKOpCZfzK/4qUKke753RyzIpHL
0+7XTj/Ba9VlwjE2o7gblDw+vmaANvwEwDXhFDUNGxtJUQr8OrhllhHre/tUdnaf0x6L4DtVb0SB
Zlq+fesc//c0SNTzs/KWaFoT61oJ6IvScEyJa4rQdDKwesYuVPyIWOD6Dh/NWqhW9nMKG836ZcVy
L+vtb67dWB3REIgdHAeZlg+MmRZ2v0lzj21RJMkuEKzf24w+5EtxukFvJI/mtoAsogeSUQguyw5m
WCJjj87BQ3O90sNLLq0Kz5fAFbn90lINBeSyIeMRTrJeIx27Bo447osqFAIpBn+ZBHaMlZ4MIYip
hmMjpTePcuFpNIWqB0oym57dmWfroMcVOWeqIdvrOxbbRGzjq20bAke5bMZPd7zttBnU0Q1Z40B+
Yo8ZEF8xEJleWL0J7p41KJ+KPInB2tO8tdjAMSeEpKBi2E2TVzm/pdADKhNIAnCn/4SUf2fGff0h
YseC04hvfLubBUzUVSc/7FkkSzqCO77xvLnCWeZrOeD6+908iw4zn0dGza2KSoUQq1GHk0xw//Mq
j7HzjyYUn2/qb1yOVgnnHtZ2LB1RkO9AR3hUVcRNXPSHmhZ8tjIzdyJIBIg20pNZYi/F/YDFhNuU
0pXXHcbKZGiQJBbgHkMWBnmk95d598T/9j2P9WKE6PgjuZXDCAL02u89XwIx6U0NZ1dCVGoLg1BN
tgedhLuy4dfZfRi/oLpln0ilw6SLdZ8VYNgv9kPoTd6LpEtkjB2N+WI3k5ZD2biGJf7ebcx8pX8V
hSoTU7cH51Cq8/azFtuNs2PzvF+0J4Smzlc02XEMyfzQ07J9UgAGAM3eJi5eksYd/0jv5O9tpU0m
dmjBd0v8KSqKU3rDQdduBkTbBvoNwZ9CBSIYydFbzrdnUAUW6+9YWG9WPfb6JtOcwqqIMRreS3NE
cT/PKiR4MUS6tMeieuyyvS0l8wnO3Z2j3PJlP39zHrb7FdsY51fasGOIoqi7lIGVP0nSydL9HDaa
AhHE7Kv3G4SF26BZNGpiOd/ArSUYw0LyBhoG7YZc/44NLfYXe1BNAUSICLNhnFZQ4brT4CO+WMwK
4mhqX+ZcI3jZjs52nFGoG/gypvZ/vjVkjVspFYk987sO4lhzu0ZBc8MwFytLM5hjoNQxrPJfFDeN
wzJKpo8835Q1X1xhILR2GDywUgZoeQYjd8/7nWBnWKtEb0V0H/8ahjvHMrvQvKSwrF8iVoB/gFVV
FkZ5YP0GJr5gFIzVm3PBX23OAIhdlSv/Yw8J8wEPW8JdfmNqxS7hrfQnNTb/1RVZlMgmHwVOjRWl
0CUnfYFdBVm9SP1Uv4i1k3aKxIopvKd/NaP5Qu2jCBL1H8c4YZskUzpRYjhAFsITaCW5ewIlpsbm
esiUoakkNVoOwKnb1z0ebLWQV7XlWQR2VnGr6TVoxgOiUb9/dT1C3RjA+/wWssxQiNhlo8bg/6+4
ufV25/76JiOgNUMAIjzVNWL0I4PuqFNyewqlH+wbCthuUxzaAsyhekDisnkP7k4zHavtWTsxHNwP
5UmUemuKv3IxQIOCkff3IdpPZTkEgJJyndC7+OXqgD8SIQYVBp0RiPG5rs8bkdUBOSkf0a920ysG
j2mevs0f7nptIaJwCCEh8diNE4PDTSDj8PoCO4IU5VALyzp0PQ6lWf8tgzh0qW8gRa3HcHKm9+wp
o7Zj1h4kVxMnlQ817jcvuYUMAQtKb5g1NTp4Xf8Lm9AOFw87KuyF3hZuYXhX1dD+NVwFPaSmvQhV
14GZQ3Y3ovzZWk2bbonedq+hVp4oJGIvVLucRwtKS+A2UQXTj28y4OviMIVLLx1grdISEBPqCqD/
2rosOGKmpuDOjS5wWNmBya/la9V/OtKL/RsxSEh9OlrV17NuN1NsKyJ8DIhB06toioYKUUDgAuUN
4DhCllyCOhczRpV+pmsHCALEdOZhuXCTL4Cg1Va++cFIY2vfN3+iEXtfMjgfFFNO0uIjXZxQqbAq
2ktuc5Fvh5P9/dUsmsPfXfUCvcpILSb5yi3nWSAu1j1fHTGty2ZvijTuZKZsRCZEjo9eqBLRmrDO
j1rc8v/dBaz42UhVykGYtqNROtu5vDTBlX3NG5162QDL3I2YPAFYDmKC9MQd/bjEf02y/3txSFgD
cAvwPbIdhNuFZXlYeGBo/3DhOzCyg8NGVLALumnTA2xoVPqznc84xZ2sBDDZwbEJ4KPdTHR3afRJ
xl2zGWfmcZ7TjhPmxWTfzZ+eggIF0l4arOfur8W7/gyEa8RpskuVmKI6ef4U94xkdfI/ADtj0Uaa
RBXC5decSeMvG9ah3yY9CE9xm9/ratx8+0fKTJNxK6wDcTElmSvNUy2BSStlWQdcmFo90cB7C4Ac
9dBQvS96bLJHyBW8ikEikcjX7p3JYue3+HVjP9u9ZMt9TwP7JWXrO6/KhP+XboxoaH9NU6yazScR
95DH7vNj2I+TS2lTAD1OIjs81FoUtnLfe24QcelNGHMwSF6YQtcSE53Ywf1MxUSVGYLiGhSpU7Za
+sCw8l75qAK5Idp0DyZYQ/OMkbC4QSbq5OZOKcDPGlh41U23VkT6yBViZx7SAY8Ajj6CAYnao2oj
fb/cFc73WY5qc6tNAzwe/RMq82GON/vbMleAc9UL2dHoFYigv9SBSCd5YWDM+qtSXPRRAnnNXakp
PYnyWA+lJtNZXivt5S56NP+Oi1a4VBZsENnuJjo2ctK8A1sbJ8BEzgllCQWbF8Jq72swe/MdGy6k
q+6wvHKr6p3aP2huoGCZoDQCZObpu5yOQDVlrTnpymfqJk+RzMvctoqnGmz5DoTN4NQd897QaOiI
ESl9C6EurD4RuClxuhjJZMt7f5hQmJeayoy208XtYxXA3Cjg0aEIaIlHr5jV8hS6I2++CYIl0lLp
OJ6arhuQO8/vr0J0KGeM6LV5hl+IjjBQ1+L67zo62vUN0bzGOf90WPukhXwMdV3SWzLONNDdSjFG
WOXz+g0mzQFXjofl14thn4tYlAxctsZtiqdNaAX8PZ5Dw2U3sOpwFR8lKWWLXBYhqN+nrNt7k+jq
tjWw7kHBVZ9+r2d03DWe+oq6rj7VcUAog1e6h4xIqPkmjKn5D2Sl4W5n2jFLX4tv0bIpk3DEUuTu
6vtssJq0X0L6oEPpy9dYVx5Wi2hMJawQTGAzwG62bE+YNm2N3Fx4PvhcTFaLn4vLes4GRXK697Mu
ikfCY5EB3TzmK7++eotHKkM+ZI5+dSbmjqUh9hToNIG3ACNe7UNQ48qWJR11Iwsqb/Offf+yTBD3
/1fh1BOYPSnnbiEqT4ztAQzpDVkR1046nICzHga6mifghXjiX3T4Y1ryT8CC4/7ggWkOi2M4N3Z0
L1H/SJDQcXY3WqV7zcFef/C/TqS7hiyXAXv+GghnSSxTr4RNEpOBD6dLbA7swy6206JxzKEj1gNt
L3e0WF5pfwxVUUztUBNXBjFgVyFVmu7JccJqfuYfh7TPApL0SKmsI43h8v9ShTZDzPO02w2Ewq6j
0R2nxitxTw2umF1STd43srpg+Px2q746KkDWuCwhChMQT4a4Ik+lzG55jjm5ddGEb8O4MFCPizAo
Xe8fPUid9fB8QHjAkV9X3gQobtYiyTSlC39j6efynZIlOd7Jtr3DZw7biR3KjlEj52Yi2t6wCyH/
MCfkA9d9ttHLWDqjCvHa/NCxqUi90rGvuy/fg948zcBXt+HrgDASOihp5t2sUlF2P7SpjJQqZ9q2
daG1WJDREqJrpbqzmYWxQyzR++asWtC74EfTM8DIFcxX18WzQmAplc14pXRZxHr8bZMGcyZ32JD/
dS0IH4J3xA2KhcXV9KWRifNeWEXeZjxPHwE9w/QLe9bHIan+lf7pT0bOFHdGjMK93eHZqN0j7Nqn
fBWqYT51fVbMZMN6VadP0Be7qm8yOHEeW8GjD+S72OrSetvV7XefRGhY1+sqRvpOCZZOLVD67ILn
kIpBashoZv8WicziMPY4Xf1G/hsyx67TadVEXEZ8phTAfoVEy+tTZKISJGveLuyJ2rmF9Vyjy3CZ
+YK3zAJXo5QXUoCBKG1dGNtdlMmoFqMh+Bpmc4jPUHSMAAlw0m+D0aADB11rv/WkQGeu06/UeZl0
inuRVK1yP+hYAMLcIjLayk5zUkk6lPzcNq3xM0xX8MznZIdCnfYUwV3Seo1ANuHKb9GJWlHbWnFT
r6osrUXVbWTJu9k/MlP8KM8hhcOnI9tiXQ7iR3YKo6Ps20E6E9YWxNfyvL+jcq4yyp2ECDOcOeFG
ljbZViQSzYqHQNqu8dJvmumq5i+3rzz3B6QYefoE18DlG998Xv0NZkonroQYcWIdsn4z86bSjTWN
V3UUIuHqyPQzJkk+cquQRLerlnHV5e04ml/9PZqK3N1i/nK053zBTtyvu+jtoeU5hl0lyoUpg/4K
NgGhno1Eqm9MzSxmBLXR+hukHHeGFjNpUm35GZS2GqLb3TvPsxU74q3ItPn2bghYwlyeL3hMEK43
Tf0kL80ENYl+iq6pTUOUodm0pcxfE5DLoNtglV4NsNar1UOIYvpJ8/qv4TLxFdmEAx5VCC5e8KGg
SY/OGDB8oVlD35kUAqcnHOH1hrW+uYzsSqu93oTLKmIzSraNKMisRMYIcInVNgzDgX6XDMp7vzhM
3Eap+/VnN3EAyiQg2k13l6Dyu7CeM6BHvAPykHQA2MUAszsSDGLCS/Hdu7eu0RhpKT2WLhY/501w
skjUAsynAVbiLl6Z8yIjKveY/FzmpgkuT8m1/5KwA8Ozs47eULQcayM14nKIjcbPGq9NRwQeKwXW
LdfP92WR3znWm3RhUQrNe3YMRXzcrKGHNxBl05iqK7SZA2Fi6pFQXF8Lhp6U98JgeQtsLPoligAS
dfav5c/B+7XRLWF0WJtBImBHWjugvUDNi/H7FP69prFqjCbxIehyLP947OJ2bwPgAiEhanTV1Mzn
vDlVwXp360qolZun4vLQxbuNJDKlZgyA/1gvobiMLfqWAk4SWSG3hzEidR4f3X3WIJE3DbiPMulZ
CEnpTbTmRrdjYRRcpesjRhTIWP5ZqZ/wKjpwLr/HuDKaRijzBYlIUMctNPTjSPp7cmxLiQe0XSrB
1mQVecozWw7KJaBUKeNdY1lgm5KOvFZr7lTQRJEOAmvMFmzgZh8BIqntOp8+/EYKTP2k0DCObiy3
OUqzqbrxh3qgTLuaSgBfmSK3oaxr2HjagGid/NA5VT2VSvRA1aWwjCU+I/7SjPUyuAqyUrAs4Rkt
CrE25nUpAXqLpvOL4N/DgoVfaQnXi8dx2sNk52Am6mCUEF9cXvUQc5n6XsmQAudHKOruXMPa6swi
oMXJaFVJ+++cm5n3QrxBAuUAUAT/rnv2v6tj8/7lJ6KikkHi9r4gQcr65CwYHUaIBqAvnG1Lxk04
6DPc2nUAzJwwO/KoWlfTWSFDOs05O2lGdmSJ2K2SClvdRSWbdRQomTsDLvKdmLi90jCKgDRWISCK
sG1MOawAsoPmJlDIom2bKxpQZE3Ku/9vb8lnjcNU4GJRd/YglcCpSt7tH8elgtSl4LK7barguzCq
1W1K8lomYOIB0FHKveL4NwAojbPbjXXRM/AX7nbG3cnSjdr4+E1NlJdiatVjWz2opl15c5GgVcNu
vovu9D/BxEwi4mh19nxQ85AnIckilUBjpgMOtxGQKI7ZcGR75GElBuM2Uo8FPfRRPZhcz4UgtVP1
fsNp6xRqVUEKB2UFzyhOHlu8H3PmG+DTQmPRkTZUX5ROBKhcXqQPmym6sIxH4UJOT550Hms5skDT
AVFpLYD/gKU1QpB7akoaBadDgkO9kR2kdLwe8E1OTvXYJNFN9IjWYjAoAYkb8aV3X2N4IRF7+48N
awpupjmF3GiuOwEJuzlXNmzP/d2Iuey+/0hPvMPRJoFIL+dfED4zugoK/Grkcei/5vc4X4rucayX
hwzO05owLh2Ur4LuilMmfoP0GKSNeoYr5+qr5AaEMMlL8vnPUR5C8Lxr61sb3l/qZHDtlegu2nfq
9VYtiP972k0g4qY5ueAS1Jyggnse1VP5vV7stWXkPtXCNeuv3QrwztbsWOxtXc9+a0nEgO9fJ2H3
hH321yo2rcBElfF0cEV/hWhdfQ2Fh+7UY4ZvCQjJP0TuaEQCOzEtfnVlTrKyibi+SRRTaClsQ6U3
8E1ixyPDWUPxCjM5/33Hg6OjUuWIGuRIJLYtd9pJqX9tGgGZBh4ch+wzBmaNpoBbLlWFpfQo1OLO
TE5HdnIF9AfTLuccnG8I3vjem9AiWbvPDjoo9mR0NcYO3OVDJiwlqvBHVx4umYeXMej2LWgDRt8A
wV8QYq/d7d2XsNKmbitlHxBh1g6I+bLJhVS4dtlLmW77bOMiLwlI9rVC2+j3HZURfDqS744GJQIR
J5E8P4N/cYT/maKU6cGFlCS0jSUauqx/1wSMeqea0C3m4zBNSNwgPeoDwAqJ+dIM+kD+y5oGFiAi
IoOKZ7AVq6UPHMkSHzQOA33XvagIOtgy6LuoZpnHmNyysP/Y/G1ijxW5CY+0+fuQO0KzJ8oRNF0P
zsOiTYuAERByxHpjq8tUqit8uHe9NG8J0e5x7sSYaSEJEzH7l3LUkLbpLgXPwTLCp3rt2BDZHTck
tEKIVnS51NrYjhpkSlxMLT/xM1qPyIDgw+r/LrYrED5z+DMJCk4ITbG2AygkrGi1BFjWD4qPV+EZ
2u3BcmwryU9wQoZo16skBgFzeh7Rh/gJ9u0pQit8Lw19sxIJv22neVb9CxvtsqVteCwsTVQVJint
IRBrIR8HNy7eLK6eszno3ki+kuqr8lCF2LkKSmJaasUj/uLOuF7/yTocjBwMsolyUUC5jpMUgNx8
/l8ZUm/0yFA4Ts835Clf+0KWQ3lcVLdLbCX+tuuo00hzwt9L+CFVlNeW06vi0eP7hzUbcGUkAwqJ
VuH1HwKOddurhS5AeuQLiuwk+FfgmRRTEermUGVfHFbJb6qsrq2RRNEIV7zIHcRsUsOCjGgHg46c
KLLJo4xiPjJR1hui7y9jf07zNSeM/k20snI883kncL3tR4ckS7kbbPHeMGfnyAKQtzIsPUrqNEp0
CKfkED7jlos9bU1evLyxZLaj8piPVxbA3TcCILuxcOzdQlLfk7cRE0X+npyz5VJ/mRxX6AuQxWxw
HfdR0gcFoUwYHa3LbEW8qrWk9SBysSXES8pA1xur5cXwljl/LO07afgGNLbSe/lonq4B7jxPI/0R
3s3n6hV24O8CGzlR5yOh5xYACekwcJK/2oRy3ZfLirHj/UJVBpL9u4dTDL+K4CwmztYe3UsE6zBZ
Gfh/mI5fVNtBd99ZltP6yJfcf/fbcSKwtnDF9d6n9HOyNWNyO+FUkJ8WZTGrvRaW6l9JJZ6hnnCb
xh2XEFxQ8/KQY4/L/lbfyTYGi2ePjmwGXnuipA4rLNejCo6w/3qiS3rlR7dz4L3F42r8ER5wrJgi
Z2g61J24R0LU9FMTbJW5bfJcTVi/uOCYhE+q+7/KUXm/ggdI6MPsfFmokvbaytEpsI2GqOeysCms
9u2QHIW3izbOr4lTJmFmILg45xn3f8RhUYpf8HWN7l8lV7xCjHeDMCvPRIH39QHSDU8VNXbcgRrR
OjTL7zJ1FW7ByOS57t5FOoyfzJ8E+0WJUCuZM5TTRLRQlIEuwbD6meFcU+GRk0e2QVSMEVebsfHU
ydOQjaaWgyiJ5AGVy1B3VDyhZ5csmi00R3L6CRTdZwFOh23SlvixRP29/OPLc1fB5XKfpiCeqZdH
tUPwOwFE3TYZu6SsbjWpPQuzjbGv0J5zAzBWET2mXaieu19yZZfEFjv6SgovWxl+uezJsGFe1q4q
1/2Ht9d2Bf4AIukLERlekSbIDZZhIsC5kzlhf+y7NWz/ciZxMqdzjLNImstGHXZjM9cRsgALr8oN
B9Ej4td+PNJJoi33KNQ6E8/37wJnYOeBXwXrTS2za0Q478mQ6wSFCNwZ3gDHqda5ExFUJY/r4paf
0W5SnrVJ8O5aOtev4jhamELlGPn1C9tf9ft7jRy++BUX7UkWdCIy1pi19Jr89mFRR06j2KrtIIQ8
SoTWx/kSVx+nxN5MBZQ6wdVl2v4NCl5lkLWFFw6R5/hK89IMuPDKQ/7sQt05bIwOVoBptgDvd7y/
5HfJ6er93Kte+/7M8FgGMjNS1EEmaN0OIvgcnzkES0fyR5/mZX2VlxRMVnLu3MrsbfhoKKK7WBZw
nVgXF5mOvA0HUUXtBhnMvho4pQKT8s9FR6deWy6JxE82yfXExsN1+tnclWr//rPElo0lLIULjAOt
3dz4J8HGeVHl6+IFLLh+bEpZqkeLpibf0XZqdbHfcFaG9ouKw+DY8Fj/BpWJqIUmX8ujLtjT5oAC
XAkgu8NoOQpu9hq4A1a7rmsG8+GpVTDOlacXJy/ofqd565Qw7AR0kPQPwPowQXMhm/KjcPQvzywD
bnItjN1dh4VqWQq9RBYLTAy7Yu+6Iqu98yLMrTTLgh4yoe9DazQ65r+CdbL3Y2TW3u0nVP59+4if
Vhr8NogASgqh7Mof7AGIEpm2sT5YWKPaAuDzlp8j0JzuCWsGdXx1/DIM95wp21CdR04y6d2Xu9tf
B4p/VpjTeQXgXcUuNh90wRfKPbTnG2BVSHGvD3PXo/oWWbZCOZnNYPMpeK2+j7F3y4CPE5kPAZXV
A7c3v922Z63Ldtf/DuA/dKZ1xlHj+v+JuBXWFuYy/+Tp7HS+uxPqi51dyPPzGHUaewlxwWD9AXP+
BlfAuXzCaS3pvCMZHYd/M+QMPzdR7MQH1VmJV7wut7juGoPxBd9QfbUxPa7rM2b/jd2u/+VuYu+K
PKGUAL8wEMi6DTi9Fi4K3SgFOulXeZiN68VJYaNMsVUD/joAs57Tj/ivq03mwdcE4i2bkEsNAR1O
ovwRZvQNMAaW47txUxXmG5CoZHQyMa4eL6e1ncPVPwNSvzjUcG6+XaAgJnkvvU/B0Xb0DOhHmf0g
CJOrD7mmMSozO9jsSEkXAimve42JeH6EjA527QGvwjpBOj5Ucqenb8pB0GaRu3Yh50Rk2vSnnIr7
QXLIqKJX1UVVTIycsY5Um9xHT2TR90xQ9qFnEOx/9Nsk2S1grQP2jtwtw3p+B/U3o3BeK4vXThiu
DGaKMx0u/W1n1sq5KiXxQYuwSoX3b6XsUPz6TnRfMxDIKqNhHk2mwOVeFLPDZa1YluWXTB7ZUGwK
g1zt6hCDoi3K0SLpqpVOuN5ldtP2I4wrkRpefm/7eOv6F5kBvgLWWlfBYG3TkkNz8WMAFdV9w+OR
mkpo5RZePKDAmbdb7I8qZoXk3vA0QrrSxaM4RRQWZhbglEBLkjKEGsq6FLfqor6VnkCKm0qlzt8c
mVJsIiXiGnzWix6VuxjpjATGDaU44jkFG1qYAnyeArUVg5v/BQygzUy/2q3Di2RXgAoOQKOsg/rc
2svLwCkiDEmmgwyIvVC4Vstag+xSatpgrLiyR0tC5Bkz4ghGHGeV2pt34ZExSiEJr6I/SIEqPTAD
f5uXAxt4ewireEBeHY45borrqgGd3pxIzpK0MfVMm0HiyZVXpoSVWajxCXTLDScTRtBya3Tq6K2e
+aRO6S51zIlpCPkrA/4uoL2V/9W5DUKaEbb1SxCOo1kE6+V6bd5/Ku0Yxjx6Mzu8rZMO1GsnwHww
XjJHGcwrD5H1W9d7/YVAGNK4M4DsiI7EZ5BrmttLULSEN51uBbMgXI8/SEMzV4BgqXbE8OyhW7BP
jE+spXhInOKHmNUgRCqWe0ulErYIF9LunWp7+M4zzaWVGyriiZXDt9XsGCmxRiu7hccduT8wC8TH
LgB4XRi3z63iwbNGh7fyrhyswZ6OVTPprWzQa5Sa92U4ReWprG0z+6OacdUnjUgzm4MtlSG3u9n5
ajpNczG5Mkvocj9Pgw0dHca4Q671L4BpCO6dbXl6rg5564kdLup/iVaRvn8cMp4qDrkpQ8QJCGUI
dzYcPonfniXVeksadOh/f9jLNKi5HMxCu96Swk99hPmGdL0Y5sRBwyZL2DUCia0klwmB6nMrZcFF
a08aDAALJZuzxV/wKFLyTavuJ4B0kVNvY0aDoxVYKNXxiR/lLmh8psrKqJBn4f/bdl4zgpxVvbPG
lzFDaCYMpjDOBJj4XJImBc119ok9Dsop8Uz7FdTrsWbnjBRYGqw1k21NMrmq7QQqn0GVDq4G/zag
Yv+gpbyjK5iZeTsAPYd7xZb1DvINqZOVzUFf00fFMRE361j7+kbN8Jlb79c0KtK7+2FV0Ns+NVos
8euyLvtC2u0MLxSyTwVftudsHNerL2s/3+RLPNCG+82bg+3gouiVmAvngsgdOJBPn3P+LnIS5mF6
8s4SGoYxJySU2J4nPgbzG4s8r54BlbpBzdvC7IcvP+Ju/bSnCzIjxcUg06re89hHp13mxFBajber
LUjUe+VjQbJnJgOysYGqnRIMDQJewGQNLX0VYOyIF+Z3ZLcwJUgY3aGUdrv/20T1Wag5ANBoCbrZ
5fiP4W6uPkCW2GbX1P4cWOVhlm5wxJ7OXaydXPgI2Txm1LfjDlhnDeMmh/Q8AN3k8C7I5VC0/bw8
EsiAR/uLcqKH8P2RXsKmsbw/ysD/BhSfziZeXI+Tleuebu7jDKvI1r5BWJFfVf0FOi8wLAA5Ss2M
B0OQb5Os682QGFDjNeNJXsxZ7ixf0kCBGaWFKSuPjawFyKVtcYY7dnrUyVMx4EOlhrLD9N/L12rP
uUcIliLc8dS5fhz4jF8TxxRZsOKw3RIScccecsEHBsXno1OAuOe6uxzs5OOrNJvE5ghQPC/7MyXJ
uWkBBrYkvN4Dni5+C5jZTFOdWFOW0lkiCQhgvozLFsljgZ+xd/pNh2rt4Q2bjMGPXEb6vnbjHGFD
Ru2FG4ua3R7O7IS5yehnJ4Rb0MbbMtmEKD0IUCLsEMjPo4L/VeuDOfDS0K/EUJuPmVCWaJoyqhg6
RD+FqtB49h3TOc99Wy472xjyw1ScvNSp2snSgL0a5T4iXMgYytqH6uPMFG632tMoiPEexya6UOg5
RwkSYAp/6kINA4Trva0GvIfw1TIqHpUp8C+K6ZCJgO5cHXP/4C5DN0W+aDleJWjySxMZZE+RWPLK
2hycIkRcUpfltIx2ZbWwTBrTYv5qm80TOdU9Xy3RNm4DZDnif+gtxwiwrleOXhhb8pv9N7wF2ASZ
QRlL4XbzzgOoQzdiw8rap6UY2ZxMsr2Pc2MRhI2gGtyNmDn+/67g9pMbeDvIAnnk6qDLiKVDl1kU
ba103lylfsdNnYwRlD2daD5XYDlJmuPuFh53hFo2Lhsf6zNACvDTKmqL2shcYtAqsudWGNbt1js0
RykF+Bxqucj+YKbzhbihI5fXTjVP7FXvZ2ZZ6EAWoReri4yPfgws0BZuX0L/gFhSWHc+SGGLLwGi
qn2FYsLSNMmmBC68W4dsiZz/qRCjbNNxm+2IMirWspHdxeHleo4XNeWLmCcKxINDwIwSx14bWaOo
tld8gseZ0w38t76eGXcSkgYXyHKjOL/d1CNeZ8vEt/fVPvTyCBQc947ei1MlbZY4yTu4VVANuhDg
KO/1h0ehMg++azXHybhyzOi/tzgf5mZppB8Oa2jQoDzdz+cGujswy9LrV4rz5aJ4ruiV5w6Wh0FG
ZqVBLL9Q6tINUCCk591+fBf2QFSNzPin9rl+ktiy6nSNbZ2kRmxjrkGYueAQMk/6vYTxmFXd21tQ
GN4yP4DkWsLgvQa9cUiiiOZchtLp7NOnAVNGloeHCvZij5Tiy82mNJiJTP2yiHolt5L6T3caRAlb
MkrUkUVuj0TRbLqJzshGnyjzvGfkH74caPaoFDrxmPQ+Mz3iQPz7VJD3jWBdxNWDFle8Qu13deV3
doaKbsJT2wVjAAX5JqUCnOLLUVfWYihGHCzITkw6yVd7ZM+GqPNVeuC3XKSUkdKmxP8k9ZtNxGWl
2JKliWXhpTjtpptPFLEF8LYDdW8QPmOlAmrpUzVKcEIufMUxjFEKcjA9M7uJ6QEeJ4MtEDDByxrH
j6AFz0TdADs9YwiblvuxdfWCQEYOVhlmJmvjkL8nRkqg54CeLHShvUmHnht/NSvD0JN89ZpBjgX8
iVYM7cFqy/mjyFujr7S/Qf33RIzijUmA6xzgm20OWyApTMiFyFFm6cWga2Wd7zsH0/yO+D4Yi9w7
Gzz8N5eC2W/icC39+aHVNruXsJEmFIwZXSJYen1wRXtUVGZDCeornY0jtn3hQeu64gXoA2Ydc3zd
CdGygUh6gTBRq1SzWTQze2OO+j2WRWpj3bHIOjxSkiqPgkAoAwICrXA3612OMlpWEzAZPI9gw5eG
fUpetxiVd/JvLcysf32sjNH5P6AQLeZdDcA4O3AKvmgpL88LZrGkJL8vLIqrMMg7QrDV51fZ9r0Q
vZu5m/8K61gDsu1C7MBwNkWmmHVcqI0HGgb+Jhabgu+zHny20pYX3hXKaArtwQlPkktZBMX8HnFq
unNulHC66MKvA1xYuDShmdPQHO35jyq9X7h57h6BfDBbfYGVn/LnR7LE8sjhQije7nVf7o1BJbvZ
r0u1x1A9JGVGO/wQ0q8t/xeeNkvzNDNbM/gZom/0DjAh6p2hoZLCUobeajv8lgIx6RKx7r7bNe5W
E+geHtgoY1b8+TgopRkqJqvDClyzungTxBVcSIPJ3Q789VN+jggBfMjWIymmIdAqurItAlhOCEf0
Uxbeixb/PinA7FayJMj2sQqlmLoK9CpaQ9JGRMdXlJQoy6K+uhpMs+dg/JmWj99gpIyp1IOH02i5
ei5BxcdfhyicIUMAp/ZAKK3ytlqtCAZo4jvdjQ7uA2TTmdl8q02XQrcDjmnSghGBKTBkQ9mtIHRr
3w1FFAM9V69b9Rq7WGdzueCKtHX9luqLwFBZRY7ZjswfI0OI9H3TtPvzE5rWmfHwAWFCXAhIK6Fv
9adLmyv893fXESWXOMrrC8dHpk4bF1i4Eo0uWW8nxjymjgtywoiOEuqvjKvWcVsKQuWBBQdjNRRu
4e1HdMqpTFmkz+tSECnCf/wXzmFNgZFHcjgotZEm6uQABLaiwrdcXEci+HEtGDyiFfYPtYc2O1Zw
pX2jWNNfbvnFpd+JPs+C23rLFm+acnHA/IFM4pCZGgCuTkxGD4STB2apgYBsuKCnUxx1vUNSXp6w
mH4zVh5oh8w+jNrOn0x5PpgyCMpNc9uG6QJJT6eQgtpMfjQCOmiisNjznBdMq/Rtk0xGms8MRDl6
qMRDkH6GDKzdDjy53mGbgnMnghG4SLZ3JFfSsoiuEbPPD0yfYX62k0vmDu9Db1bbqUaiBRlzoc20
2yruWKCD79VqxP+TQDqDEEpB0x51WcnJc/EUcslRkniFRFPDF/SPk29Fa5MoJ7+TP98OveXq8D7H
5aintx4dftiotJs1zdf/MnHYOHKFvWqKm0ST0Ge9Dgu3/Zq6pUvXf3DC9MajJQzfr3XhU5pkpbap
9Dd8E6UT44hnNx7lxz3ABOh+NXTW6JuECCqhdTrIJjAGRtEvxrgN4tbHDaexDs2yoVvI32JOzpLu
ylbEwaqpsEfPRdgKI52bt6rmXs9KksjjI0mIMUpaJ1pfNUox+e9nPqRCL0PrjcSn4wl/v+5yrCD1
aMn9v1y9MfdPXEjnLxtmX9PXocFiO6Wdc+vjxtHA73OorEXz2drT/SaTYdhL9hWt2fFQmCVEByIB
HCk5fmvcaeeSVzNYzP5oiVCrHBt3tKc2bHQA+OHMeRwHxx1c3ChaqSIikh75WhnR/GP8oWNWAf39
EjC66RrojAQFFaZxhYI0pkhXrUk0nVTeFLcFbfeSG3wPM9jpEHMktsJdMwZoG81kz/ZDuQ9U0m5s
ujtAg4tDA/gEGlSSv0cLqpYq4xWseBjeoBRlh6lC5wzKyadnmICGIM3KJxGwNHBp7mRvXB/RLskR
Zu/Fko0bQkYfIzc6qW51aLyAlO2n11gCqMNJGhck86JIemhdCpuQv5GpsZW4rYIGJox+WZnAYjWb
giUgEE/AKou2mlrolspj/bY5Nnf7QCUAVRAyxtedKNOfaYYRq7oqU9ltSXUwrMRczHjqYR352vL0
nLTw0KWwoC7davgYMeG7/bMO4666jkUj8ZiQ/R3zVOsLjhPOpDwEN7xOEPCLxctocNRtTilKojYP
IXZd/RHKhaRW97G66BTAVTh76fO+Y1wl0NkiVgfSR4T3fQ9XLUaHACc3tt5eqQxes+YthTsUH/YJ
e9O+bz8HPYLYVY+k1+MciDSiSbpUjKO8H6r02apdOLDeQ2qpeSYpZEmBpaKuNZZScL8Ts26grm6n
Yun8BQE6MxZAXnjV9aPswqVZvZOkBLlgiQlVbewPQRj4FOVZpRIVNlaassBiH/VZheK+QdiUmdwX
bE1gx67iEpab/HKDyj6/JjTrRCEP2YdTRiK2sXQul6jMjKMl+luIwUfqHOfxElPWkY30LzRjwXO0
LjD409HZzTWOWoY2Ag0B4uKYZU3yU5IWfD2OlMyijDbbg0KcajDIXnswvl59DO5O2pnfBcmtvqeJ
xmD2c4Khf9h/29JsCfTLH989OSvIJeyArorboA756HbeJmlxrWhVh6WylQT5HrOhq2ib+mFOMoVd
Yzwr6w9W+c7cJJ46CXzml2KTnnDbQinOMdpFi74gQX1J5X2rVBWM3JNgARZRJ1CWgfqI19To/F0/
aYBco4AhLaMspXGwWPXT9+cLadWKZosYCatjaQs+jidq4IfGnx0g8z+27K9jR0aPZTQYCeYJTSr8
rf6cydCwKFiaiVR3y6jtrRQFQguFYpN0CJT2pGusdLQv72AhdNhMZCl4Z1bgiCqwJhvo6eTx4DJB
DK180MLwj4PPDQBFVMTBmcyU4LvXeX2ZKT+hRhwL82LFSXJt6BWC4CgbFBos2f7r4ZV43ffJfzV5
+LnxJ6JYPyE9Dr0tRN4i3SEbV7Oj/trZCP6is2/1nN+Pf6qh+GbM+lkjxJYFItLF+KH9Lu6Gxq6h
NZdM300SpBBkk+Q4LRYkHY4gkmt+
`protect end_protected
