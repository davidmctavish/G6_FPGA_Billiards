`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AaugILxRlzpaYcDC3tUPKT91eCwq1E9um2PL7KEPKsyhd5b398ij8R2DlG8bHJVXN+pXZtOCd8MF
76t7tVBR5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AfPnD7PDy2nDn6cvdV3YMMwK5nuNGSdY3Z7+HraRnPcddyaAD38YI4mEo7B8jpNOIh+p0BbHGi7u
OU69fkx9qHCP1ophqa/IXnRU073OiilX5nCL1iTN2sTifv1WIa2p4+KvZYqWYbQbVZhsvTnJIVor
qjJm9GGdPtMsW65zXMU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hv8vzsDEMIZyraFe+1Q8gcANU1YFXfP9KNMJTxN0KuDm3qnH5AKKYT1qMEBuUp28G5lEEr0SciSc
aHk93bIM2Anx0MoIsquySOPWl2UvSzpaUiR+n9aF6q32AbJoQYWArIfSpgoQkMZEvBNjIaBPFsBj
y4VuPCUv/mQr4hzoIm1dPRkyoEIe+lcV5gCO8kpZtHVJj2TNA/35Lh2tb3UwzlqzcORHidYLl1wN
5TkKwPbW085smE4DRb9GZq9TjdjwJEDXnkHuEzWwWw2HyG7fyoeFOtq7AsBFc/qdKxyWygpODab9
J3pQkk6NVeYjSaCJ1LXto39ZXlfw8zY/Xi4d8g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N2P3v1FDg+LNP8fd2G8Lo7K2iBaCNQXdGoSUYoxnfhhERVikF4Sj3/T3HxAHKzQx4TXmxd30syxE
Yz9kR9TJUPsTh2sEbDXOorg4Ie/vyNJudrkTmhLA4ff8tPG54IGhuMehMWhQBdu11FQUgmrrw0ZN
vMivM7Ljz5rCvYYLdzo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ASx6IsJb9r4OKrhHxNE0jJl4zOvNuTDh3c80qBlgjT0cOLt0XVVVe7QA+Fbk6ffN/7/1xoBX9Nqc
htdowt82vSE2ck8mulVLxfesX/ImhDMOsezsCWPfypmnhnhBcz+WZiue0Yd7szyC+6sOOgA0KDII
rY9JKcJBZyzBV0QS1DXpGbfI5z+7qT87LQNvYG2mME+EmEhryMgz6XxYfxqzNz98S7jyZ01IaVMM
s5SfzOTc3BClKL7PTv+TL/K1Yvr6r5SiHQpAqjKSdi0Fl5hpTvLVTvnsKu8W5lx3CwH4AptoJekX
eLhsu3SebcFH4Gur2Oq/qQKH09gkNEnTT32JGg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24800)
`protect data_block
RuS/BXJG0mIiaDXrb8f5lQ5nDX8aMuPjlcvLCvPLf9NjU/0f8GX1OFme661905G3s87Q+TDScxfh
RyzMNK/ANIQUoeaFw+1Shw9kryruAjlBp/wNW5U1HcjQYApO87hahgr4Sjv1aKzd8c27iBNlSHHY
aCu7J+eR3jHGMSjMSZ8ebK1MgOP3hKmXse7a/8ogIJz7sIH0AA/Rz9KR07HRYoCFMCn3CjWX6m3k
ZNsHUxbhQT6LYmm4u3vdo5FYxDWjrOYvYIizkiltISqugOj86yL+JCjsSi6BFFi0JWl8eK0+28GS
dvQXaMnTHSlY7EIZbdwU2QlbYnmRCaiDy113ADMTlEjHWkrBVswpcER1CsXBNGIi589OHl1/Th0s
1CqRuc2Vd0rl3g2DhutmUK3MQCVMZJQWDvnYQrwq4gn3/wQh+SQeNPbhi1q+C3fcMFbMY6oOeCYv
dgpVSkuEJdvfqNqKqvj61SVXNIyUV6heYhpoxgkDJwtcaJvn2g9hJR5Zq7BW59GdnBT+W4HadC4P
BMY8dSEyarrMuMRtrt1Jk7UfDTy7pSk/jXzGZhLcsubcIQ81zH7MheMI7FdY+BaFUiHW4fj6VFQN
du1hSILUHz1cpdVd0pGqJU1Rbehuozl426xNJv9l4lvucQAZdGBVr64Y9Fu+9c8XsUYqYHdFAi24
5Ns/V1ROiTtTMClSphNxZnJKjss899Wcfx8GAph7ByxEioUp6w2H/sdSYeEmGCY13zC4yuG3D8bk
3N0M4L6IJRfj5bZkZLbUOTHbaVGofpXOkZGB2bbWC+SByl0dB8FmLwuigh4goFlSUC5LxUTRFDx0
VTPrDJVra+zpYDJClSaj+qHcq8ajTLleZEb/SXfzJvJEnP1vc81Qcp5hlVmJmmAHH1XzGUbTT7I5
hEirp6DPdXDugw0dlxyuEcdkbVZRDno3U/IoeFNpPqBZpo9MND35KtUNtZhdf9UvI1yXIu2cjm2E
d1vua3qsDfWlE/EvJVqFkPPYZH8wx2lfSDFz2TyQdMqvoRPbNUkh/QGCLaNxF1WO1Ezae8l2NC+V
MS5RR9gITOHFozVFKcoXQCTRBF8b5v5fpSlcJdVn2gS1LRXFfPvwwwtzt3e2Q4opD0NJWUnHI0ox
QTq/AZ6CRB4Glyb5HH2pi3w6VDJcu/QwJkA0FCQcd+bHrpfz+9y2alph4mS3sERz405Z030rAbre
AbEvSJtqODDEqdWmOHe0aQdBC5ZotsHBH9QNnSnP2t/hb6wjELi1V9FWpLrnl+ro6Nb4l+9pOpRm
yIibdh9lmWXwzslFeJTXB8rFB5iR0OaQh1S7W71SvEIPPFnyWcNvnEL+FAMJvjmO02CJOvIJfFku
Z1WR/x5qQb2xS1XmzyIOOE92nvskQNCx94rfJN/kx03O1jvRmYn0K1efK8hA4zq7S4nQSSMC9YbS
qquosk59sRPOgsRO1jqtzH3l0rnzgafgcrJHK+ffq8E3PG+AD72bJAIUOWsjJiVC6yFRhEgTL0Q7
0Xo9q6LrmjOEvME9ZIRUy/qRBsMrhHbfBI91vpwwWsgC+gQagFD5FH7Kjk2/Z/SZsMIyDvYqw0CT
I+iKUUwX06UFIX3YywFk0SMaYqo0v5cS+VsEMSHvYYyq9rtsCwJo3HOuGo0rGXCrCn79ZjoVyQg+
4u5NOmnCqOtgRb+ZFS3kexo+SAgX0fOukXAXxmnRgXTZk1Xtry6d82vqZsk/dJI3cPlQCsyweQao
nNADtkX9CAdu7yfD0xrcbhWhW9tOWCK1eMBbOzg313Qbw3XylnFDCCbdIhXdpIC589mwZCJBDViO
T7rxBd18ul8Aw6f0+RYIio+o5KWeyDxneah2SjWypCTj2cvCYkkTLUxUrfPrdGimvyvJBke4fQl7
8BruVHFQG3R+TcPSD7g7+WJJz6P5TJG34coiF6WXuZ8hrRpII2snv6bwzHjR5YreyqckPAgLwLiW
7n52KQtcUa3p2WItHkDoxD/8jkD1mbWf+ds34CS1YRD2HnzSa0vaW/OibyfzjSn6oyQDV4zEPV2o
Ix61258DJTiNH6YpSYzPlX5Qol7Nac8jiauuN3c/RbFs0LIbLfu+rNT6V/LJCYQ8CBEMoqDXmK8z
jw+pIG9nxR4VnoP0/YL5bvCjRFZMgpd+3Pn1p4ToWI5GluQ8L3i20Q9qTPFn6p3zePF6Q2cduO0L
kt9TG74KwdpSgEA3TPKB2YbZ/xUn3lZ5HppDOr5jsD3vag4sBfep3mEmNBOBBAgSpoGsoy/wTdkg
XtZOAvxBDU0Y2G80WYIVuEprG4khVNHBbi86KDnAacT+fXfZx4pX+Lt4wWNksk0Okf9Zy6cR+H+4
idqqLzcfiTzOJY/3PCMHSME3Ph6eTXsk/0wjfTxyU8+Zkt8TOIzcmJIbyj5biEMK8xQLsA3CE/Mo
Vg2kz79vzwRf+xjArMIF35jP3I9a9lql18MSWnyEQ2ZAdQOSFpCYo/J1JjsEuBbNVw7ONrXNXj8X
Kwwz6aQ3Du66ob4RIW8ROvvH9YTvZz8HaP3Ob1tPzyQBhd3ynTiGy7GsSeRk4i8AcKXns1uL+UqM
eebtYSjkRAwAW5qVwAkVDevVhsXCULDq5SERkpu8fCrDh6OAARiOJPy+GTpO613FqhqVTEFEbBz1
Ox1PrTUDUw/Axf5I/tJZ0jNgNfs9mQMu6j+JKtNVo5AiKhUS0VG5yIStDoobYDtD2pyfIZTAKA6v
GzEXu2uR/JXj/LkyLSCaLzyWg39U8a7DR34z2jUePdJT6qDZ5Gl0NuWrpVWre8mtF56LbEIU0UjC
0tUnILCSdDsESrasbE8URW7cbDkbxtq3dpOmgzdP9xyClDIpb6G+Uz73uXjMFVWRgpjUYgCCQ8Yb
KPW8XAZegimMqtGNbsO2kEv/8rfbN3loF6JWq8ESwJ+t20SQpcfSlaa3E+7YZbQgeO1/2Wsz4x04
Bk6k0xYOIc8llzz3CN5a33B3kXcqE2jmJ7UlBz+D1xGzZ6TFIlMm8XtLDQUA6WFtnu7ZPDUzyH0z
BcNLKv3U2ho9F01NNk47nTkBydqlqNiJj3XhrheAOihydM3gfzD6rQ0h44tEKdlTF4gANB/XAKSR
nklHFo3ARuexbjM4x1E6q4j8W3id1FfORaBx3+9T20gyRNmrAM2oLZDwzBmCodbJDdloLVftMUfe
fVMvdBZhJBFkxqnvs6ILDm0I9m3OPe5BUXgYy/gr2fAcw219U7ODRM5BHj0bPhGHN6l9zatAoYYp
qOaPohH4hwAsFEakF9xIASqASjob51n8mX7LOmglqHawpZ71t1rWry4hotDfP2+JqHqUyr1wqv8j
hn+3Uc7zjBw9kUN0JiA6Ew9yzorCidPo1SG11Vpa1Y4Gu1p9yEa1TfH49cdU5aUO8OverdkYU2ft
AmuHiBiQmeUUjdle0qb7ylMDZu6a4/v4ekoP3suVmWKxER5SPsfmbFiYm6DHKwljbOhimy4vcsNW
1lmx5DuqFXJC6TWE5mrcTvwwfpBWIDVJ/LRvrri7cAhfVk+tasGx6izT4rrQCqbH9MYEcxAG6CjE
Cij7QRxRCsCDrddVaPNzPVJDP06hc9L+7ALOaZdJBvRmMEpAHb47tj8c+UrMEA35vNOPjpJ2jI7a
MGKnX3RoeXkoieZbNCJIeK6H3YWHP+8X0xscUw/QfNdP0pe4ikL+nkqnvJ3ocoT+aNVx5LMH/c+i
7WQq95n/xntw3hdQvKcMLW9PbkZRLzpQzahNOVuX6ek4rjx2KeEu5N7pscgZvTkwF7rgOnYt+TE8
7/DQtHkprdu9X9a8lQXJAvP08bbhoEfv1LftUaCHKpU2JUaMVZQ24YuIHQPKicSCdtgqVHhC20yE
K7FWpNFhcOmbvsbQG1zekQDHKvNleI+43v3TY71k9JM/gOc9VZ8Hx9BrCVdvV4YBtvRLbWuIKoYI
DJu3G7cHnriqPPPqtpbhrN0en+72gXNMz1GkGbXVxqLe5dlYMryc7BPT/6BgBgW954xpcHNrl1yL
6FgeVabwSXF9euFEkGbo8ffXrcKyVNGnV1RZsBcfkK9xPxOgvxTCsK9oE0otPPydVDxx1t+p7kZm
wIVzDKnEEmi6Rj2V9bBy2oDrtoQXf70RNdzRWl1pKMLn/hKbZZYO4IrWyMk1/6lS3NVmeEmaKrcc
w5/dVMT8fdibOen6BLsHQQMxBZ1jA8v2H2fmWyBzYF1MiDcix9Svcxdep+VF4BrWh2Coo+kiiLPJ
ugG+/SfQyUpCiUv8BDLrBZ4qzMxGfcSzcgeSBSMyLQpphS5OQFdeWbiMBYAlzc3R348EEufCwZr8
oGaQKrYdoKyBKB6q6hsWmtiQDLLCc8VK+1J12Lp0vi5lI5N0/YmbGBE8CbOHcNrRsMjkS6xrGstn
urW7cEj6T7XI0OB12kcN1c2ie2lq4Hp/rbKYsxSB0Ms8wmISYTrszD1kOMOJI9NeWPNlSoY3TJB3
EUnPKZOJww3c7lj/2DsVXrGbARMq0AZGiJMpkaqVXBNQ8do+1mD5V6gB7vYtd+Z88BqWSVF92pxr
YuTWYl94SRKbc0BGDYCfWp75gzAFKkgOVWoCS5PYNKEDIINSBPZAPqSjCDu224mr3B4oRc0DwBl7
Vf/598xEICtNSWgDYUAS/n2snsFzKviJ4Yb7ftK3gMrMxch/VZMX3a9jsxe5Vdp2cdI1s74o5Ls0
Jw82seC+tP4zwfBQNeFk+MhVMlpAxeA/ULj47o235/G7B5nI4ZhfLKCOhg10aXZr0ywSdHS+ZCis
Bi/cNGnaqH+Exz4mz+FCIMQ6/hdC7wNqHn5XNLkzY57bUB6wkwVylf3k2ATNH08R0Zu2JVLJspPf
mKAM3tDTZ/4AhECroXGCvMuj7YzgckJ2+OgbWy6n5lOceaPQwKm8GZRY2nemEbxrIXC1zJ0CYZs1
8rciMT9rKe4Ao2R5cxcaKxa0QpX4ZF+QcjedqZUJzUI/ddKX0RuwbRmy5Jchzsu+m4SmxXBKZlPI
PtnwA9u1CtyfA9E+a28kAi3OAWFgWyQSUGffpD4NyBBMgBCBTcr4kATOiRrTqpljwACb19TrxLkC
g7yR8S0u/Q1gfkfnOK+U9SC97a4l0hl/MZwTbIhvAuyZ7RUqcTREOJCs87sGIDU4UaOriEyrQh4A
1teiuc0ScGgaL0FvuiVfI5Qbc2ux0Oi0uyUgTSiwUYu+SHjcG6wARxBJZCrnefRIXEgr2VmlJsLd
PZI/opSHjXusZZrL5Btq5wtRaQ8P5455P+E+MbEW96vSQhPqZXN6t/ZnBBkax6uAUhQQLtQ/GY1y
pt+LAmzlQANp1IoaYBUc9fmr2nxArDXYSO6fDaSaPGfsJ0OGisarhH9xfANrZYZn5zdAk7QX0DQy
x9TLf/035AB7jgLHhyBeKn2AG/zCsscNffjMbtlm3dyRfbEX3xtBxD1I1LSTdxClw2TdSPqS4Jbe
y2wr9774BMah+OQPLbSBKLVddWSLh7XEal8XbDJTt4eOtPYw5K1fOvJPf0e+FRrAQo32wxeZg1QI
fxxQrvbLS9IhVZEyuq2LgYu68f6QRXPjP5YzhLlp+LyBdNVCZ6v334cpblXZnchjaBLG6k9K+pHE
hcQiAVY+pifj3qWIW7RsJPA95Cl5n3rhPQDzUPYNICYXL+DUggKugnq8ZTZCnH5vJVMVJby300cA
CGoFETw7g09J6BfT5As2xCYVwJH0U367Rd5v7Mf67MqZ3sFLpZc06lJgEcKP5DeTY42f9KhZgvHq
rYql92+AMnmFpL2zbWlSdDqqFnebcuVOAhksEJ2W5IFoVzgxCOKJh5CoDhvpJsFo/q0mC9di2qUz
2kpmQMe9A6ERPfkeY1sVjtIQSTj6Ea6pLP/c3sslfX8u8YE1VphpdlJtZCyzvkw6/BWRILvleiUi
Hp1QJcD6cZRdwz24AUfPnVu8oIvpgNlbY6aVzLBXmdYFb68+3hM19QZlz3Ay2QezsVlwg4NFSgUA
5/lg00tUBY3D0JieALO76brpfP2VzUc7togWTmgrE1O9eOzPw5KYd010/Ofw6wIb8cXdGNQr42sC
9+wtOcs0L+pBW29kxUWCyeMhlnJvfflIWCJLitFNxwSBT5WeuAqPHExwDA+GIhyq4E5T6zMnEsnA
7eDCEfR1YarcWMKcAcEe+Yw+UEBb4J01oQOfkqJClCXa6nXOUXbG+rtrw782Dt3fiCkSluwl1YiF
JHfWm5dWQyac3fFAucFYqemtYqj/3atxwCq/yxGcZBE42CNyELkC3k0AO6xZ5kg6DBmz65DnIxZ7
UNDAUqjYpKCnUX1nGgEh6ion9PmkPqWtCXdxgDjJLed1WQaNGyZH2UXtyy9okHVJQQ6gzlFuZx++
eD38A5TBah6Jvc/IcMgWkso8IrwuwtNse5slAyKruQQ5X4eoCkwaNB7dVmQnNPfgpmrhU3536Mgb
DblOKgbqHNt6KzMez8F3/WAyH9RCwm69i2DduLONGPoFAL5Iqk/SiOylLDXVVnCAG8aN0Bs2rtxh
d+v0L28eu4lHJ4OXIOXtEEsS4Ch7MDrkaVdomC3mZDBB3LL7b0gH+erg0u5poRqzxmZpFeqWDpeT
I9vVDPAgBGJki0IKdCtme0lBRgMyv6jPbpI8uDA1ZPoaQ2sSkEzt1QyOAcuRdP2CK5A0NCZ41EL7
KUvShVur9y7BKm5733ftxDIf2YAI/nm5Y+IDcl3ERJFNIndaIfWCDFav19952KGgNzMQMpH9h5+b
yG7KYnGWCTDgDtOqTtfgR+M5DnzgWBkgVqRyCF2RN5xTJUxJUHWlwtgE4dK2DHhhKNGEbnPCEDvr
PQWhUoXVoV56CC4jUs38UYvpknoyAudSwruLosyXZpnK/UsgT0n8IIDVeAkthzyF7Dge5WDw3BgQ
09ICOGFazR6XhNrcrRKKGfHKp0u/u6GP7u18rUCd1CAtegpHbvNSS5zABzEkA5hK6RdNs646/LN2
mGfpqvakagYjPS+8vBW7RjQQ4DrN3axLG3XoYjryVX24TwHmbPaBceWwB/MKfmN/QkGO5kwtQbou
Z+IhhiVkfywmR9JsfxJAqOMMK1P5RPHCHNCxnyUpGllw3Tjz+wmBfsv0hVhq/TeMmXpui/x8Kr3X
OI74mBEwItL4gNxUzBaG/x8ZUM4dHYona6AbFQDY8JYXCenlp1vR9hA0KW7DhS3qxztts/09W88e
dvl6/zI1mD675tIMNsrsmo6sf6Fy1t4wTk6NnZyzRJBjjkEKyneLy62Mme5XtyaFmbkgVU5jvZAj
bHIRnxCa/ht28LDqGxDSiCLAqkOx14D0SLqzVD9eN/yLIfIpsU8z8MOwcChb80YvBWgDWA2jICXY
R3y8RpHX8EZAJRiU8TBmYq1URdZjeR7ZvEJnmRl+ANmuTIJCf+qVN1iE7q+wtcm3opSLMuNgDRWb
Xzwyr7bc6TRQX/5aZsVRvEf/i5NN2GLklZtk1k9qfsUmOvOk5uj8PKrITVzTeYBfyX12zgbXEKdS
3Us7nhhbtpEbXkTo5/PvpbIfVzUNqyICAfNSoGi/PG6E7L78uQTT+zqPbYv3Psuk+ARO35B1bmUc
MlfBX0MstwTmh49dhhXWzJLk38B35H0RwZ7aUy5jZ1BQ4dm1PuSR7bB6szLsLlxF40cy20I3FDEK
ZM+ddXNbRm7P8dBjUInm5VSfK9alr+Mt8J649YixbZd7vpwj2KYP0piULik7ADsG/EM2UKb9aIKa
EHG2tGgZyrG8EVaZ4OMh9xkIarSA0VH6AFZ0PsPZyeyt9pMasaMU8ZdZocUdj8xSXmcPLrw5V13F
PBRy0WrVHtRZyd4DphxRFAkUybmWMoWfby71u/iPgiYOfHqodt7pkcZPWuHDOPVKWPBpr/lDg3EQ
uLnjZ1Qdk0AYJpTJOa45c9IeNEyYi17uc73nlTC2glDz2ORj6h7g9KU6peWDcJ3N/2e/tLaUd0hu
OgKx/b0FafKPZwroZ18eAQ27AZHLOeNctdMkixLWNmrepBLYVCOod+noOqQoHppWUaax+LQiD572
U+cwOtTjziRl5aeX7DJxWmbVmtVZ8Qlg7m9+EXy03N12XRfkykWGeH4r7zK/n/1I3LRtGVz+vVll
DQ3Dg7lPgNJ8aKr6ss8vaJymSyLXtQBiKpMnNOPVmgXl/cJK4dQa0aPzhyihTNMeX5sqnNbOO5GR
oWOF3CLggwtzcKz2NufeyXfkKp5Nzkm+TjdpsiLKIiky4f5CYdzgvH24TOmsSxpA4SaQq1gwfot/
lj0o+zxrjWT5hlhkQVaeqRcpERmtQ0pfN8roGxzuHfynNqmrFDHAjNY7tDXedBHf9FMeHpT29SLk
gTpcS5LAtQ16cKuwdf1KbTqAq/GUcp9oZdD7zg/yZBhoMYaRh6Rpyjp6PhggqF0SZLCnAHNH21W/
kGEbpNPLrADO2mqHOfdILSEFEPrPg0a0yro1oxRpPeeDke33kZa6hvpBXcZmwVLUxTHPIGf4p7jZ
iFtpgFoVuGHtHFshklkKxVU8P2NGJfGekadsJtzQ9gO4twoRF8TP9/1zftqXZi3PcJ2u6hoxtwTY
RVVgIEyGKZ4ha0XY0InDamnWWQhyzc1uOtYBG74YN+MuhKhAjT65l4BbjjOWH9KNPAYrPN74l23b
FRrmliyEvgicjvmWG7SnaCQmz8LWK0Ru6JBn9F7ZJvroSx2UqVZMdLQbPAEuRODsMk7dInPnCiYV
tfmvltlcwfWJCvPU4c4habnSKLv2raNl4Z3Y91xeT0hr6u3GpcbdESHw5w1/EWYKPqPkbNkJqO+0
EFFS4kbt/xkvKKK2Yo8avZiyXTXjTYr4gEX0Rn2qXDKPtUN7KM4CcsfqYfzWYta8KnrLesTRa1Ov
cQ5iuBq64z/D4hWBEN6uP3G4W/7JkI/VvxRo9FSfXSsaIJo2hR8/0vhHvZqdeoKYUkwfx8iYOFPc
GnC5mDV+OXm7ZHQGOt9If50j/UiHZPC7VLnuhu2QQojS/yaLn1INL1sGeKrxHaa9b1LC7ZMPXFvf
6xa6uXSNvFIzvNhZKnw3ElfnhVb8Fyn7U9HqbL8cWgnSyfxB/0vOma4Hx7L8vCVsRimJiJzaoTDw
n9MkA4u5guBfsLzZw41tNONi+u50/wQR+FmGZg6+Qyo1++3iV7DPE0r1x1oHF6mITV6TaRKUA/6y
PUNUftQzNI2snjxtfHs2p7CT/aNjOZLadjthqd34HtJp1TPMfLqjqwOVerKjDQaMCvpYOE9lXWfn
6+q0aA179B7/Ow3epBiry0fKaHydtD/vtNfRxgTiKkGqTVKK7CHiEtMkeHCZPKoBK3OHHKsoCXPh
ou41omLF8QpmfWp8lKeJS4Z/K8GRJ14TNe8kPYh/YzUrzzU5pQ2DD3yVAZPByr6fyIK8ShqenctV
29yxgLMD95WRRTN1krueadOnXgFnyx8OWG2nXNWS5KEp/rzVSyqHLLMLODQWd1leCZLrEZag9ITc
etEoH6C1jzOLbOhfBAHuUSmSIAT6etxspubkLlv8dvW9mZwd/zG9JZn4xuO6IF76zuH/XyRvtamO
Hq6NLNnRmHtdg93SnvpBhG0vWyEA8VDkPxtrVmt7OXHEXdEpEkPu/YvUWK2TDLrieNWZyv2rMU5C
rrxqV7TTjUiTEfmHoXUaz8l7w0O/RxWTldlcBXt8JHICcASnkaq09utEk8pHNyu7Ym4rKhMXl+v3
VcmyHKKzkNsG2jv30lume/4gQdv+5KuXkDodhfipXmJGmTx2avcvfJ98lmb18hSgNdGTF7tylzLQ
DmKBrEXLpdB7Kr1hyzCDFVmggUBUPdk9t1Vkv8xdXCFTq1ZO4xslzvUvagfUPLW58Wep1Xv0KzLt
AnKnlUHfl5FgSDF8Ye0CDHjYTjQjwPY1l5aKKlSAWBzO7h5KNQOkLiIwQ6d5e3ZUSWIhr6zVuG0B
VXhzOqSVphWM3TN1zZ9K16aNBh5HuCSTas3CLCGgYc7Bn9qCJfAvgmCIa2uH07oWZ8/JcEOGaANu
KXULW8J3QY4lpu+0HTjYRdMzZa4BTYg9kkpDPfvtefvtw2gVgVKd9boZ1LUd3cmB9TOWfUWpYE48
n1X98AswkVY/RS7HGxEMxTaaFgqW3v4vgLJOZ0LUspwcsOYf6dJN8ICa5qYeRjRVQHsVwHy19Dff
kQbqJeERLUpZu9SfSyPx8mkjDJ+7A5HMiRct44VfaPDuTpPga73Y2nS8lXKN/E31Xgzt7mE8A0BK
+aQTQiksmRqrVwEPOvIGjdo7f6GN8WsJma5xK2VLhGUaXTFpbm2n5OBI3qrc/n82GyfTbvpZvE26
eEk27zRdIhAaNiug9sSmM2gb38GpyURQUPSjOXOL1EeQOmAF2pk8znFswE9268+s7M5g0byudPWx
aCSpdYUkBhnSMQRa98HUSi5YbX4YQHPTxZ0spSr679kBlCPaHfUHq/luZbgIlUBvOIAIz8cCAD71
1cLqRW+ZxOAD9MeDljueZT4IcGzgJ8VZUGQSrEh7ptHNqQee7eHcLfVZguK9/qvZAYYWJ67t27wQ
Fi1RQFQ9d6wtpjzbnitO7iXk5hLc60QT0CLe0VjmnY0RjEQ2i3A8tn2upA97aw7+c6dGBjJ7UDne
cB5P3UethVNt+iD3LMxAN98SFTaVfWROSMRdPsy7XxDtgxF+pldHtQmB1ERrK+q3T2v4z2GaXtw8
BccKIoekSz8ne+QjVsLof+Uhxmv2BKmXbDIRjZfuApUUytvrKyZhz/OD7+QGnndA8CObeKg75RiP
myjl2gdj2XUvstrtWbSl2UXjFeNSUaU5h9gKtaAIdwWHRbZJV3+6iPX7B7KtdHtyS/kPPzQguvgR
bIBDs3GR21Z8+P6jRnphe3ACXuGCny3nd6JZAkQcVTdAYxPMLNd2cyltAymZD2JRPWgs0gr0UjXi
GnOdrYYYeV6tg96wCVFZ2UZ6wcSS8Ova+pUVaPV/tOn+aVqZO0r2296/AiUsIL43Ml006OeaZDQR
1PJZJHFljIj6f5HZ3nzQVSNZ0m7kih9BhcSYDywSMfntNzMFsCL19Bkp0H+a+jO1TC0tRxG9CwzW
ZB6zTXihqh886289Q88+KtfwsFLFWx1CZrH+aBE1IuoIIGV8zbY3ARU0yAIk4RqqXPEDv38C1xXR
tH8ADKTbQ8X5joeAeTEKFbQTJbeuXB1bvUnL/eZghHL2AgRi/cfdVLQBnjdvUdrNKuUbufmTr4j5
cM/duvZv0g0d4GXQFGsJY6amRbZXKvlQ0RGKNab0GRnr6kooXqUygrsIJNIQp8H6/QQcMqQI4lzP
rj9M1Ipl+DIK4RZG8GGGKndDNxgDUGCqAEQf3sPpsliBDs8KbiGUpW11eIZN83dgW+rhZ6oqpmYF
2OW8tGTWPMuDi2fEnK3UcIWUrx6oKHCaGD+MMqfj4uVl2TrukIolAFlsRmmahhjxAZ3/pfX/sznS
1Kf7hGookRn1QwGDHkf1Al28/7HYCsCjzzVzwrk38KFwShBOrzpNoVNu1iVTnuIrLGBFK4fxDgAW
Ootd+3OT7sgXf8uF8h48/eySzpoqrKUYEtIBcWqkijVBtRm0jSfgDBX83sem8n8PXimNRe2Vkdyn
ZsJx133TfoRLZmD5W++ukT5b4C60U2+0RcGZZpdVrpgwl/OMLIVZpt76KHphfEugwHiJJ5iYNMjR
C0KSGO7mcP6fhvOaTSXAF/6MnpAAmCrT3TxbYwGH694Aqy4a0bQoK8X0d7NDCVk0R8uqbUopUdVo
AibEtnREE3cKbIlXblh4ocuF39/mkpnVMpZxY0F0athGRCBPibNb17hzdVjVG28IBpLyxs7TTOjQ
0hdFfJq+i+7VXAVWleXwqJrMYrfwAp4ZYwb+uTAmEdAxZhJgM/b3zhJuMX5CmWeja4GOSB9IDQ8n
vcVtmh+jIxtfrKqrj7hBDv/7YFlqT9a8ElMENTonZ13PybIjPmYXP8EW2NtA7BFPbzj97vTZSYau
4vbQGkw5bTs4H0lDP1ohfVdqSYVL1xyZlv+X7M23+ykRHgTpGOQHZMT78ZiRUFaZA5FFV7dPYUkD
IHXqvIWEm8bIiiGOAILMWdXn0F9w2QdGNj12KzEzm2hi2WUzsMdnoPh3JwRndYfw3WXretfrXNY1
0PuA2+6cPNnKDNrtboWoEpEiwzjVkzDqnjsxzCK6lh3Zf55Ioq04uZemYI5SHMG0I0Krdyi+TFGL
k5lVKTcQ6UTrfPmXttI4KfpsDS2YtJkID1P5jn5LVzh3hZlIXPpy+rNoID928libLa1AL54DHc6a
W97F61lfCGRA1o1M9/e/G2edB70iBVdayLUHQPh+c61CJQdgiCxLVhJHmaggoZb5+KEmxybAJwYQ
IS1/+/D2vpB5pkdJy5TPSt8dtS9dbY6fbUbwq8IaDyGCicnWxsCWaLFVKdtfHXvkFO0cA+geXdPp
j9iudY4lIHBpw9cG/kTgY79aWOviWLh/JIbsAnHGSmNAkopxcaHR8XkuOMVIJWzYthhmeZAWHKRv
fqil/bc5FxrwX5oMUlMxTWA1QeU5hbSU81n9iH/Y4x6fn994u3iQrSaFKXjd5IRl3y+jWbfrgdZh
XcP+dANmQdNq9oTYGYAsBnIz0bkzWdvFrOQp1HaDl1NjiM2od+tc+CoYj4adHdMA0hMtA5Z4uU/D
QgPWRuvS9SBwbrk4Z5BV6dKdlYP2llkt4VJED/Om0LHiNw6QMMZ/Tf00hEUEMZSRM3AwcGh5JL3N
98bArwKOuPw3gOY7fGZ8YKv4EDu4qCO2PY3K3DKquyGFOjofx33VhnjbtXNBup+tNG3eitNt+mBH
QBXCqBGpJ/68x61zx5j+s5rGkDQni87xpBQOXzJCg6AjASMopFTnTBGpws/zaZ6yLh66EzaXMWHh
xwkFI/CJatT4+AXqawbfJLJTZMFBVX+8eCUR5EykgW/4nwlzY83f4KTWdLoRJ+JOzXo5fEh5X/53
E5A6QPOInFum2OI0lK29FYkTa+MCIBztx/c/DhukMri6kUgN1D9GW7IOXVfi67tOlVuhmkdmVI7/
ZPkxYR5kmjQ4Uq4E51Oe3kqp2CJeSNnbekDx1ogtFgUjWBn+f9Rt4Z9wnMLOZ/IsOOfvX93kGNrZ
E4ibtIgv5vVou0q3vA7aYYy0yF4/sB30QC3g2E8flzrP4pehQ3Gt8ZtX14GZNq14ZAK3pUIGe2zE
lNumJDgoh0fopB3NRsLZACjPKpFMoF6A9eB6AN7PZm9ud9s+4fNodGUoT0b/3lQy98kQH5iiFy/E
rmXOGsmFuksgPNrEijNX+6AfJxbNDbX+sXyrxG4v1Se9YgL2E5yYmMH0xzVcVpHHWnSIRKTWQZTP
iir+UcX0QR1yGNxQLymQipSBZFrNmDI3asMAfjPS3mzz625mAFD+ECfwqirURa13zJ8xNBrkK/xy
pDfIrnOUszLPWcxBVcN5kXarqlCueG4MOVV32HOLxfuUqM0vglNtGVeMhNPOwtb1U5OLYAGza/G2
+GgPA5OizgZbCXXBS6aBCYgf+knIYrTW7zaLI/XWxPSUvSfPywFNkFNRi1yZAJuenGCvY/aEBX3k
HZJktZrIo87eEapWY0seY5i4e/NEGUJGclyr8MhA+HoWRtyNxY4gWjfjLDv17EezRPK60yPet7dm
OeCOjpoeARO9CROzxQ8+evt0wNhXIvoBNGypwiWaJeXXlV8REzOL3PehXbVLB8qJ9l4BlAi+InKz
agKScdsdDyaBiQX7qQNdohM6TFaMrbE2M1hloWqreLKvvesv8vxePDyu3JFag59why+e1K3mRY0p
2xSifVeP1958UGNFMpABosqPzUH8EI2N2qPvX33az8/wdUEYwvUgckQO+6hl6hgIPOwOo1Fe5bqF
LwV+fBKkzz7p0NL4qgfsz7A4H5riLv0H9AzCk06ip88b2F1fERHihG7o1WDY7V1GV/MZBEW4mn/N
+j+a+pCVw3EKMQbUoYVwIU0zyBaGNUKNmYmCMiMBRhn041URIJSQxnAw3wByMHFyittcw6QyMwlb
i3TiefEDKa3Gvc4SAk9fzEQYYpGq5EtUv0Hc084tEGFK62Mj+zaAvqV/jn5yiDsKvS/M28EA/is+
v4rU3G1wnu/sp7fiuaf/iWOQ3SYF5nBGve2DC594kdzPebZO1ho/m8kwE1+sQsmyF05djugOOdTE
hdq59JsRE2nCti3KiFJLgKD+mmuTV66fI333cMowC6tgFo9cnGQtCtFVdC0MEnzLLpVIgw6OpnWD
10WXNa4FiuwH/OmFFW7klkclaCCPr1V8sM0kZLK8EZurnBkpgFvEuu5xBqF+nzJM63lvkjYeadQ5
AQ+3TVJvzpaPfG6H4FaF4r79V6hmkGOyNIozjS+aCSMLoL5VkQ8cFx7rTVfOhGnva94VfHxeUGs9
KFPItlPXKSUX6S5PdRmxVfzTH42h0JZ47gFJLUPtQKTyJlDB6ne9g/0wIBN7JsVM9G4AYZdFB/3W
24nOaPMNdTUKU5EI6P5tQ20BzQ7v+CJsBZrTDwtf9/yM96DCKyBPXEvy0u5XW7RuyBTshGn/4TrC
wLsiNBUG1uWwRCW4srrtvGPYVhRbDuB4RctXo6/qTS+S91ySO2/REjPAbEFNIS1ii/OmuFZO0w0d
s7sil5x6972oZzJAvtHngfr5voHAHwKjw/Fak454ws2p79iDrSij7a7wDp3UkiJnFm3lad1pWfWN
qCoz0o4h9K5OK6Av/zjOFCLP71aYt/6ytUS8u0pg6qP6HLqIuShoMqRXi0SsvrAHhmCqjR17DWTA
sbe1NKkSBarHuefsyiV/JV/Dlr+dFoHb3ttNMBLRQx/EfwhYzSj9//dM9hK5jL65RYZkes3C3EpF
4irFck9+PDFAEw5DIjasDAEE2FfWItZv+9bPDhF+1lxUZBdNTppDkM5d9OzHI+XEAEV1nOXXtIO/
Bns1TtGP+H7TTUWebj8AZSD2k9q0HePYU70Aes9xDqHs47wVjUAkTHXJJeKq9YKBjEDvGxuiJ6BO
j6qE/Klu7u/uN31cS8yJlu6QTqr6t1zAQBwx911xmONFbzGVj++UVHlk1RBcjfPW9SY6ynfS6xZ3
JZVIt8Vm1mkcp1w7upnv39vU8Fgfthvt9foqQWr24h12ulw7QR5hfm1zxBYHmiK5TrIUcGiyR1+6
yYtocpHi/M6l1/KWANu1DtXRqJyftmXMJ76Pf36pTkuWP/gMuY8ZlrcXdw1rF1uOsog8Lm7MSwSB
df1sCaROWO/7+mnM5vLeq4I9FMD9ToXYRMXrRH7PgLDuSRFNxCDr7wziyyh8D2YKghiSFAquhp2l
xfnJ7hGRgpgS2YalS93Txw14Aq5IN26vDYRt6lRFtIMGC59eHxah72FzOr/4SuH0bV+uWXJ6phFZ
FlEzU6OI7WCU4XzhJaFL5nNi+zxCXHTEsPJKbcZ066A4Y0O43iavG+pxhfkr9TJJXUMgosWxXom5
tqH0Lw9z/R8irRIdQxkv/T/fhC3e13QVh1vmmifKRkGq8PskLhkMc8vm4HjXI8BmDZxf27BH5ChJ
WBP3zh8DX6zt8i7GODHcz0vrNzh1p01iyPIiPz+dhihfTEp3UqQaTUDlfXGO8MIZVy9fThkbwAi8
DobdAjoSYTgcGKSMigAbAlE2UonLaEXVpyC/6jP0xFX0Xwvnt91DkhBP1irIsRCv1Ez1wsCrFTF4
rdDdPpPo00GflX3YW2UhvTV7UOq8Ok1dy2DEXDlIIUnsCZvFFS1r/jgyZlYnLXIHnmW9jgILfcNz
2Xkv7/W/o8fKBeLIrxWyd5bx91rz7gfsNSKefh3BgFC1cUn8/eK/PGK4bq8oMkvwPnkvpAdc2ESh
hW03GZ5FtCpsJQMdjMmx9hBK+rgebuAXbv7fLZ+0VAwRsn9bhzO8NwQDVt9LNWZUQJhaUBPIuDDQ
u/bcywtI17PA9QzXloweb7abA93NinjPM3EQ0V7dDn49NL7UHJhA1mqgQOGveYJgrZWdR2UWEcXe
Zi27cB9uDQIb8uNVnssgv3/A48GvBTeC/irH/+FqXyTd5nARugd3363XN99fyJY1LbYoGzVfKTfO
7bClYut0FeAPMBOZO/CHv1+ky8fq6CjVAzDsmBL1ahHmANT50OJjYBZY5zQmO7VP/nrhMBAP1EUC
1AFzObkjPI0rMPlsrIYt3famPlmcrlnC/nDZi/Q7K6MAFHDS6pS/aYVK1pLagoT8qwQLzyvcJvm/
lTI6R5aAHSyvItV+cl1+XC1+7wnbNhq4h6QcrQY3kqX3rjHFrmnEtb3Xd4+z+yPG/+025FBeYnqM
GY46DxEoq8PrjSaCjHp+g+R69bpRvhjEBWp0HFdTtF7mDeBc/iIq9nD33Wlf+XWgj5DeO9mbxcZz
sFzXRm3xr/jnPN/vNb5AO/poHDoaz2OjQlopNKnHSSwPNAlRoN/v7l+8TPAQcCTgTFeqtc12STIF
BBJTjGKgg+cf6ol0uT2K1ixYoE+2mVGewzqITKItkEJ97TiGms+bYpGbrfewNg8c8fN+NUX3QOlu
Dz3TgKU3M8miqBE4FZA51JYFbOrK9FapXD71A5jQTvmtE9/+nLTuei31QxfHukNfj9euNoJ4+NIX
pwLIvkqSBuGpyWHV2aTV5LiELDkUOrkl4yWC3HNaihfn9eogIkpF/w3p+fbUulhuH/3xWiFps8Z4
W2syLrOFZvs4uLOdSG2R7dtPgSw00CVVAVg3jzN9y7LU1YyW8npQHCIVAgfKe6gVHnvjrJj5BmF1
TCqNtdvTen5PkHCIoL1f024cfFP3liJQbyZ+ANeB9TYC9XTnnmGOgzbyCuQdtxhBOr0pfZVjex8m
9Dy1NwZuvCqdK+fuuh8aP+dSrYF0K2/yvR1ZG7olyzpofaCVYSENdCWU1ieuMbvq5ZCezAqDqrTZ
gUIMrQF9NxgT62/kR3DVIUth9PvpaCRhUx4GcupP4Zib+RmL0aKG79x3FD9bqleT9kuHbrpFE+E0
rSOAM7jsQ2qU/+hN/BGKQZhBIdWQ0SJk7MQPml0mRM7BpUOCv//SorBpNvNRIKIJqSyhRmdROxsR
VSov92VbUHGGBZSCcIUnJR6hWVfWOQm4hkmbn2pDQa8Jsl8NwOwcArEKIMjmZ7ky8zezNvw5ocD3
AbV8ePwidSM9En5vmp/SHUj/RtnS2Zn4FkDCr1x6tDQGQMqN0aBbwXC4tQJ2YmVns4Y3atd+HEAI
eJKFOFF9ljVanldldWsf7k4abnHQPjwPTArh1QaRcmsuCuVRxmCaF5TqO3OdJGcvuOI8GUyAl5pE
R1FtwpKz8czaqgByNd/t1aPpeDrhwB6drv099ZBNZv+nghDcapArk6j8ED5KT6oEwM4zlfKa+Tzo
/KqLqiE4ZFxZhwujIYaK3zX5Cyv+SuSCnluhbgjvCWipe0qpGzztAo8NbylSySJ39KQbhpQtlTlu
XjC0HLiLplvq4AxBxqSGtcmwk5kFtaK6K+A4FsGejiqhGgLwAJMmvNt7wfSdZt/2dPp1BN3AC4Ms
VvzT94RcxhVSrxUm2AH1FkQ1d9lWXimO0cJvOAkzv/y98VTYr2ZcFr9lQMmVZdxcqHm0/S7jfsJd
Yq+NDRk31NZ9JshpIqwKaofN5DN55jbvAYXC8INX1Z4KmeC3eIprS5zpG864aOsVDikGTibSxKwR
sLTVXNw/Ki0e0r+8Vs00IBxZ19seMmDs/sna7wTnCKfSJzsmRaFo94KWi0XaVV0SzWDJpJfFvLmn
fnuvSCbiqFUoOcKuuW16v4VgKSO3XI9MXBkwLLXghdamsVA3o9clJTTix4sN/DDLjyYAPlaMWq44
ciE7DyVoIhjIsTziCLUTdqZ/m/pVo+jfRHaVHlCJeyInChtnsJh/qQh2M1p8a6UguL45zFg/H8J9
maVeNVwPyDXAAwnTpSGR+4DRHRQl8/32R1M0L/7R5+Q6shwggt7CMFM8ppxVwxd1Sw/6fpF4VrsL
Sct0G7lJPR7zKeZbL8ZY8/ngOu3HM4vAaCYUT1XOGQzOdqbORC8ZDR10TGD/irxg4+eZj1yfu6ST
fMdcyVHvwaZrx+vpvWq6h8xNYG/uDZZOacS9Ps8ZBlrzixl2BQxUYyQUq/USbit71RVBhCBL0d3q
ONslrReoIvpwc/lzzyCIM9uy4NFlBezB47sN0NTX+tfLg8mJRMjEs5YCkuRccuYCqkr7cWM44ynZ
5KWlergn96YLc84Ywa+NgjH8a5SPEAB9r8RSoNnYZrYoakuqKpo6TMOVC15BtjTPenvS7i8blaFy
B+ROo8/4AeByuoXTA1/pI6+NQsXv8/0U+O585/fmGQ7XPcBqDw3erCG5A1iRVxXbNVaZHVYTaU69
3bSZMIHD/vGwVXx/QNMv7DZ6vhFx+GQYlwgYnHat1l+KI3hr5T0FfyOI2O2VzlGJe88Qbud3xWEM
8wuW2QPiSg7kAgofcLsg2HqLrh9mzR3F24VqR/6w49L+9/RP3zpVgUMLDr8eFVB3Z4h3w9EFZAEf
5+WCdBh4KQW35NNEmhWnzc9AyxHLFYcBagTKNu4Czb3Fs5Dr2eq55f3XeIiJMAENuMatBhJe+NBp
mhAO0YEt/IA9EHDfg/NHD86vgyghf9F9rhpWIe5YrDNyflq7Qys2jkDFYnPs4ofYBMzg1bskYtpc
yZn+3ykBVntutAyMICkpGsgRcI14JovFmuBrOVoh04RwkNTWPGFfMEVe5a/+VlXc7DJ1wTDD0Srd
9VouoDotZ2EAnV3hacIDB6qDQ01/2RUjPiCMxWt42rftQpH3t9YOuIvJKrMJ0TOrzRTZZqdCnRk7
xadcoP+iqgegNlIhg4gQKheGEDdCiFJLLbE9cghN9pD/ziQVoGbVzmNtPsLMbHoyltJs3ssU8Ssy
bDCqToxbPa+17paiU7uj7PWFwnh5YHpboggpyEPQzZCL21j+rcAPUtidSz8nThsT1Bf7KbP2ZQXE
6H8jBdu6r9vUmxyvpIRj1DBOKcJPITLyEHM5JwPsvZPjLsaEIu5IS3AlkF37D6gScn1U8Njn5T5z
L1tq7tG6Loh3TMXUI5zNq/OFME4GNNAShhOW2zf3xucK2qJ3N7G3byUQcauKo5J1XFo5Ha9+PZ68
lH8wL8/pAbECznjCJbl2CYcCPD5Z152LSooOwJ3EABWSbnSi55X1pcjqieZRGEKIRoMwTFZ/fEgg
zV4gKEacwcoh9H0c5D5vNnOhQ2ERHVupX8aKvlMk2A9yhraqq8QQaWJydCrX+IA6JNwzzoWajDe9
JWiZHioNpziw/9sAbPr3grT8jsPA5kSP1AW2YJW5Z781NC/dNQSRu7ggUYkCppDrjTFPt5h4hN4f
CJKExI+JmEA4wPM8N9ee2N4v6QOXY5BCdv3Fu6vo8U6+DyfGOCc5wOutxtR6YH0y/plKQRPqElBR
QBa7+71nWDysfDTX8HJXtH5WfJnJNN/mRfm6lWD3yMu0UM9oOcpCrH7ZHIgXHFXfCoUyfjo1YYRM
7fyXRPLwa1TSNkGbxq2z7CrOqf4QvoKFH857bFMT8ik0XB93NO4ecYn/+jlPItHHfUmJXhbecYoS
6OuKr5kjjWsCYj2IRfrCu/Qxy+t31nH7+FFhi+OlEMZspUans8pYNB5D7Tvd4U5kzNoG7UwELjHh
o17YIO9UvAujogiw6aseTNW0o9PTdf7R0JopJFDboamgaWfa6oXXgxQ2zChvAwvZBjCohT/Q6LQB
1dBUzUL8X6Mp/UPiYEs5FE0beWvl/udWlvQMBDDAne4K4PSASscDdFNjNzG3sMhEwGFJJuQUK/w2
weCR6kp94zvjsnuf5kNAFeJOg/G984KH4fz4ilkCUOVMgs2/+eYJUTgKDcEz0zsxovp4zOzs7hBH
7AAnuOOPfi0r5NYcHm5ZolsFfYIbRSGTafmCR5ziKdXdUqiEcxGRevEAJK0o8Dfrbh+LFaywP3OA
sj5jFdnup2DAk7JO1EdEYrHcxB2rs2c946/X73bOkKtOFtwO1ju8vc7jQbevHxHX13u8sP2/4poH
jHYkwVFIjpy8iEO3hDaYO2qZKRtyMVDXjOXDOfDijOWZy6NZXtGL4SMvHjWcaGCZ90tvI5OirjIS
U9k5U2oLGNqldrDlpPt8v4r3Zay0SyAQNLlq1acnimT4RAuV+EDb+5rUl3GQFpFHsY9c0C6/SOYF
h5zBvpLtzuaa1e+LbyI8kAY/Rp/WEarkznaZEXt3wjePw+v9e474NaJfe3ssbVQIWoiEDVlHV3PX
sIFAtcy+q2Hv931+EN+vjyvokYzfQYIsjlgf9/R6wTnV47M0Q9BpYlqT4rY8cJbDOzHyMroEWWBF
fH8+ll5ymfiKGmwGRNgI5JTAH5wVTbsut9w12CU8Z51ja6ktytTkCY4mT0TZeN6nOgk/ZtG2lVvi
D1FpmVg6yDjFjsLjFXXzoWp09/tUQa03Pw7x4mauP1PX2KO2TuEelnWL2lWdrHslmIWo0YptVjM1
hMIuEEbpZ4bVTjFo9RoSeIIg8KugR8SWszVVXPX52ImoFeu+C1C7is5KVlBlutQtqIeh7KKH0OOv
pG/PSWeCVvf94KC3YPMStPY/Xqw4Dni63KMci9/Zxj3Frj2O0kkDP0hoDmn9BG/q21VhWftnUZwS
SvrrEeUSig/d+lp1WmZI09peoRWrlT0uwYRpbV3IG+RJS2PyCLP8Ifh7wKSZXsVFOgcctXOCoTTU
T6WUL+N0QGAtbgmFPAzj5cKCFkmbEGJ+RDridjlCgIozH3RDIIc3RF4wv07hqcJ4kShyoPNMOThg
RHKSMzYLwv11Pon+jwW7jkY7zWgbUN4yvyw+tWzsf8rx8IrzFMd/RSkN0ySCH8+UL+OsbcoEz7gB
GfhUwgp+BGHjFxwuEHp/nwjuk16z68Wx+7hYSaDWPjrSvyUpMqUFrQFr2Cm0AySqe+0YYJ7mX9I5
CBVg9gOazRZYKaX6+Y46g2KSmgLy1sfa1NZqOqL8p/bsWqNn4xr+Mm3AKXEKzrnW7meSVL16VxUk
1QPTjBs+bU9+X2MiHKsC/ymWXWLdHCsC0MXlgv0KNSSwCzMrTAl0NXAeJ23VBwwJ1Q2e/rfvUsJ3
14vA8TBi1zxM1QH8r+ga3mOkazxg99nAX/P9vsAMeuQYjJ/N10rE17JyCU3zqvNHHo23gSvE8X5f
veDutxINRx/M50NeGugjvXN5avmfX0sSuc2hJKmt9pPDOoDL+LvGVj5ipIfwsh479GoIdpIr+/wy
geZHmqe7bqqeJom/GXYoapJ0LEdlY0p6cioGqBWuQc/T5egRnkYKL7CdM1sOkUJfiT7Wt6zZgGUC
oQjyG0CPLdhKvr+vL5984tFE9LNPt2k7voPlDmHlV69WpPNqBXJct5A9rdevgLkTSIZKPVu3qUv3
mBjl4pK9qjpnUaFqSTld3gH7kHuyFf5kyr3+Iz/fsVvQyJTsNEZzYmexBx96nwJ2ByExCV1AYyQT
IQ2d/4sb4ejy4fcuHPt1OeKzAbOB9tfIBQVAZTD3WSp2sR8S1tExTap/rlRhuwY1/FDwLoz3b/yQ
UpxTDj6DW69EdILetJT/BHn0ImAyf75Xr1JyhJS/4nVw+i7gybGKo8zdh/CviVfPWHlA46dJPK1Y
RKLBXJxzSHIP6q3HY4BsI3wcVUud/xhxGFSNzMTQewFpDM2qhWreRhU0pJcycer1B2DNHxCOIWVz
+Bk6jAFPSFsI8dX6TrustJ4N8YkoqaF9FZFyWfKvav7O70acT40SuLuILCQ214fwvnshk9hdt70U
gV0uy+DfLKxnp79BgEGUFpK/jo2JJUy6Tqv/3XILrjQNPGaN4zI+Lc+QDml33iVwfm3QeU7Efzrj
CJ1/IMGtZlcdPEWho9kVJ/H91jJ84kaoyjypADFbJCzhQlbHGXu9P/P+GNKmvgZZGUPaumaheEnR
qF3pDDoUSwI6QbNNjzu/R7uIamMZ2Yk3RnXthG20PIo+rZgRL5iaVQaMMSo9FAyToy5QayFEv+eo
poAOsSspOc9DTcr3byAbLauqm51+ynPujwDF5by1X+vDoJYc0CAw8nJX3JO04QELQBNE+7W7CgKp
rwThwyqaWsdOXNWyzmP7lRUI5avxk/o+KqPL6gzYhOuDeTC0Q0pI7As5oqeGWOFWKdP2NzwxPhrW
LBTWytiP0zLHJKrd9cpp9ckR6yDAbhcj+s4/4ZrLMggY5sVojVg20w8WqKGQ/1/ttWRGsQFBD4Ry
A5oRxUR6O/PjHzMf81Kdx8M7WwfNhKdTcnXzchAB/LT34Odo0NOINfChNKO20wM6fbDUo119z2Dh
Gjc/ebclw7wPmCC1KoRFdQxIkbN3r3xhZuN9wg+m2MAlr/Q6hpKcpGzVOeMRNitLiwJye/cPnO/1
JKDC/on5tfl6XWQafWfy5lt/NFCdgNvzUj2Qtaz1M0PRPuceg3O9wiCoJSakWc5VLbFvEmPRckcO
koWc6cz2YYGnYtd8J1q22bp4Uw34lVlKg+C39kSXsAZGb18ccLq1yrBDawWzVkBB4Hx9nv0wyHt7
Nezc+QlNDsR4ND8w3LyFzFRXz/fd64NyNFbY5VBuleqwo3Dvu+QJCcXlg5l8T1hqne/8Kyt8/gZS
TK+phnkcxOJo5UihNyI67CIzK2MfEZEtl9h4H9MH+vwE3IaVTe0LRW4qQ2uby2NX6uCkNGqcb5e+
XkRVhxlECLp79Dy2eC3cpjbG7hPRDdEARDE1nAPiw9NMEU7G454R5oCq4axgZ3Gp+dQ2hQ3wS3yp
xfKdFPE6axXQ5vIxHN/tbSWdybzjZbcTFihzi+QBogNQEAlCLVb1kgmFnJwey3B5nLJq08WO7Pvf
XYLFP3WwyeGrh1nT1efu1gIe3GhgFi8T47iVsnveIxODIA9mtsYghn5wiCsM1EDzmJgPiJOIex+0
o4Dx0+3J3rEQn61gKW6OOD1SrzcZsIxib3xlRIuBLCdZdgAPJ9YvbXb/wc7Oy3YN1IJnAWK8mD9f
QS+YxdX//ytR5g5hAOS2X7P66qKith67uki7Ms/4rjL3X8iJkp9dgdC5eyuZBV7VZXm+dkm0M2My
Zh4v0shlBR5fCjifrn96s9l4hnVF1vMczS2dLV0pkPtqGJlZrBzD7k1ZGMOAVMkO9NuObb+u6zJ4
a55PPv2KFqYvCjhZhOf3AKn6kvhMPvPmbAawtrG6wdo7+ZDBqukizs2ld1Yta4RYh3Co8GMu0JoL
WXcu7KH76WdpXXz6VwbxoxzCmCk3oQmn3o9JlR6z+ta7XNSN97SrdU7E/4D2iQFKq4oat/HIs++B
yBpIqglrBOu0c6fnKBUyBZ6zlTS7Ciy940+grVeJUN4esg9EljkPIeKg7jq8y1ZIPlmtiAp56aCf
IeCD4fOLPzjlfT0wCiCZ1QSnGNvI0VghpM23tUNpyaFypao+xhNqxBrumflfA/WZVpccEYv2SBTB
EMk98SzErlE8EgbKdSwHZH7YI6uJ5JuKz9LoeukSSAm1CnkZG5THBcW8lI0V7JjO/ZF8bmz/F8YS
eRgJrxSIWixshTWPRmGLvCkRF5XyQBqptTEmGdEH2ztBI1OvWk5g2EliPK4bzJa4/a+uM89y3IQG
jwbss1mHOfl0p41d91syUDF3xD1gIPNzuGtF1ih5vRCZ5PLQZq6eK0e8LaeAtC6u9T1kvUL+09xx
FsokHdguwLSdFXXs43F0PywWmjDvAKrKeTC0u5MS6SOthneHTmmmL6nhEwS7RLUONNxzziyPB/T+
AWDV41JF4d8xCe8n+1ujHK6Yr/NgVSIDo8DwOFqgmfeTFSWNYj3fsV0MjuHEukqsiTSPgsKeCRB2
5b0N/hvYeVGfuPS06GozLKGorVFjFJpbFERrwAcohbO1gkHfx+kWa9gVBWXOSJgNn7NxghwuNQQe
SkFjiM+cN9zbrHD5kpZfeIv9hCMDyUs1BYtgIoyYTN2Y4Z8vf6DS+NVKmlmB4YObRQK2VK9AMfIN
45OH46bjCJ5fta01KYfqUzrjd+T9QDYuhJ2HAUnBHMLnKrZB1p7OrRMLmxWwTE9SUFXcNzzrR+dg
7uL0r1ryLwpZA6xWdzBX96Uzn8D7wLkXCMztK/KN/ov6P5RgZNdl++za8RutHBzlPx8OWYWEWonc
fhEExSUvsG2KbaMf8DiSI9CN+vVP/yrjpaz7Na+JxUUpTONB7xUnWEZobO492n9wYtaYSIYlHegw
z+OQiQZGmhzD9rVJqoWvrhKCRsjRUmNUQsJVijydKnwabBdZ+XOa2nagGw/BB4HqR5ezfhNmxqB6
Syux9rgF2j/zncInlFP8ThIeOY39NAZsEjx9p44yGy9PfFMp/Wfe5+sL6+8hmNfwGxsO9eDNvD7T
SqPYIG9i/weBjVhGgzDqtejYUOo6mXMzo8HFInn2CZkvS9BT2vyY2FP8BRR07gpVdrWclvZdrjHW
bVctajiozSTEhldNelcTYiZRIXCtfR8DsNIF6oi4wdqs6FSxeb7GzGW+TvH6QJtrLzAPMUpC+4NU
PFBCWk96HtMrnf0pbH1Rbziuo8mAJldnmC5vSaK1QjTOPJ3BL9uONqH57W+eHijkgUL9fUXGM9m7
1z7sGy+VVaniTgtYoHsUO5SMVAD19xX1iudOkwOpICUiXW8bjnV5MpvfbAw4AiAB6HDD4jiH4aKY
jab3tqIp4XZ6dAzWg+ttm7jsc7S9OcNZYGzyq2WsEceFIvb2MXQSUnoN/EzKooBHrPRl0nPTqXhW
VB1V/4w49DFdkS7jwa0dOGOkpHVAmR+GKUvYZ3bx2okk6fYEsH27ojq7i0SYb6wOCc9/OOa1oK/B
vQfevs9lcQj2PdMaaYDxfTS78g+ujiZ6eM3Z4z8/hDTT00FQyessfhQFqX5AblWFtSFFcm5B/Qyk
JfaREAaOQ01k+OgJAoXgHUdtw/eXOmsifaJ+ntk9Wk45irOaeqgGiaTReHNSr8ufOIy85TRlp73Q
gsYWG2N3tsHkCE7IS2VI/TE2uxIcyrTXXV1Csx6Pz+j9jWdc6cfSDzYdTLUZKaZfXb9LpkUEFVHK
rwOvC4pYWyNqKbDOCuarYXkrSRHAbQvgbTOkj8ZYhDBF/ud7yvGCzNC76MbRDWjuF0qdV1EbQx9v
zZ81B46EH8ysV3Cx3PHzbJFZ8RyR9iN/bHtuzbL/FRQJNL0sSxoe24VHFfVr/U/776FWUPdVDbIo
goBhOVM3HUtu2uX2V94FDk1YB1dZEN9NV9yt7reEu+plOd2vlQ48GWObwFiBkRzmrvsLVJcaHkxv
bILf12gTAmJUkl1eYFPOXXtuslU9NKAxlPOTEsCoazN0Ot8qsP2LtLy85WMdKnpSoDvRNCFhcyTl
LYdtOF7t/oS494VwDJpJ1+phWyb5DFB5gIFOJnX92gKb7Gdc2b9fX+kMWaJGCJUAIrFnhwHHVZPF
FwvnEZ0PWR/pLHOHfr0NtqPz16n+fTUAvqb3g81EQLleXBF43e3J1NcS6L/9aIzIBpVptUYYokIf
aDnV+rsk+mACuMYw2CVTVSLjakb50N6eF6DevDzOm6pr0Yaq3H+ZUwE/h6+v47cY1w54VQORSzS6
nQVj6z10z3RdXhU/A8ddffzYS+3eoswYcwUT6nawkbhfOsGqk9RK2Z1eqV/F6xzOG7p6ks7wE/j8
Z4AnZJcj6JIUVwqWPK4S/6c9BDEMyjl1tnHJs3MYvTkAeHZmaIE3VWOM76UkNvkmJjm/LALGnocA
nVHIOKKu0U0zPUvyfAXdqcxla31DFeYaYyDxng85+7vor81gZ5rRBw6sdvT5nQwwtiaILmY8s8HV
Cn0k2kakwI6y7jzpM0PfWcme+CA9kZW8XFbFngcucSKeanyJx6e2G1ozrUGzCd/G0/mbnkweIor7
KDw2QFJBYtOCxVPnjtLDT6F01Sv3eSfN3F3KZXM/2nzADnw8DWgjEZJBM71a446ZzQimy8LFgbbY
eJbVZs8i6mG/Wes7mERXBRzM8o1gGz6y4si5TDS5opo9Uo/Jaq2YJUcPsywDmltSL/oit2+3j2EA
oXyo+61AMT/88BkVdV3u33xIEPOOCOo66EdVAxCxkj+515fo9YvXKEGZWG6u6ph94XF6VZv7Hva2
/jaIYtXtuGBp+peLN2hZOqBKQuXYmIV13/Om10HEJfjrAXlG079uF1HqXRymHDKawwTB8ydA+QIh
LQrZw4Go+IDNy7SMwNu4netQetYGQMVUc1CcNIOmNCFzmlwpbjhHNYeqGR35hq5m6fr+2X+6YjXz
SElZ49255S8lMSQCAS4Ne4eajtKTFNgRYQuMAiR3z3V2wfMlBbCyrXYGEcmheA8FhbZnHrShjCHC
Dts1M/wY4Kc0+TtoWJGH9J+U7V2NCP/+Bb2SfZiKewa6lClS+sZDQVkvT/VO2NGWVkTC0Oq831TH
y7ybWM9lU3cPq3jhE1XuT/GhNySQJncxAMQQt6qwyHV6WHaiEADE/sbvVCxCFRnGjMo6PP6WR2OM
B6q7UkcbWuZIT1vqo2xB5H2lbmFDOR6C57DxdCpLrVodXpzJ1AIc1L1cjaQprYstAPgm2YCSjVsV
3F8kIsHXtrUgFwNylAhcHYF2Yug2HZyGJrMShA0R7oyR8tIS5eY98HrLe+ikx363BUaiP/WPWXuj
jgijY+1awmbl386/zYRysfesGd5GTKh1nUNlLpGyrr02StwO5pkFa2YQocTaE53woJtR0O/Vhp+U
9oTyxHNWPedth2JVCLsdZvCWcbBAw/jNpSJTWWWf40Qm6uKnqbDWIZmgYfJ/WEcN8teZ6uaePsCh
gq2NPeEpEGKJDOd9L9F5wbh7QkgcKwZaXJOMy2c1QMvv0qf5p3OU8scba1GptgQebcF9DVGplBZv
+wkXExc8zKWnr4py0xTYUusBK6qZRfk7fdkOfY0nCzsjXMsE0hBytx0U890Q6pWnDuWKnZ9KOL5H
SXhZMEYtncx95nvZUMHhpXNlneljfkRPHyPcmOARxdrvDJpfsNFx502WUXWBvU8FtxibubQr2fFr
9Us2TCaDnnhGz5WalGeisJZfkpHPRRRZcjwjQPZlJHvGAQVO0Y6acEip7BpN15pAWTZhWBBfwhQP
9FGLsM70/R1QEzxY7FoxfhNpKtcPj2eWOuXvNuv0+2lgGWpF+9q0jHJvsJGESzG7T1AWT5AXdnKk
uar2LE9M3Hu6sLv6M+QtrpA7g1+1GRP5/P4VnFXS0JlErUSym7JwmElFf0BUHp0NVJg0+Io121I+
IdaKvhJTSoWT1CDPMMxwLSpJD6UmVnW5tvhPE2y5+NKKn0+Map+7crWQimKxxHhHQjFV7bWYlYCR
rDssq/B3qaevHVbUYdSAWofFf9UZ382hGG4Ey38JOVJ+BItfuo69zjFGE7aj9ysuBAbnr3FS0iMV
Ab8YMJfo0vLGrqtz/+nJIjwfzcdSsGWD5Hc1GOmUGIHjX4HHZRuLezg4rFwvCuzdyEKRXhhXdpl9
O7yjz5FEVgb0Kkb+l3YRVdN8nA14FGSNlurOXriab+M1A64D60F1B5ftZyFf0t5uGYQml0xJuwEx
t2AdgarT0alEX6yjJUuj7eUmaS5YDU+C+pJDehTczlEwkBcRwoupKowt7Xne4B06tgrB6uTuhePj
lY6oy2LTcn5k+EMCqB+zn5CSXKYY65trKpgBtPqIAOEPqi302MKk/rSnB+bTB1zVIarwDjG5SvyE
4Mg7bcZZGiDhfnW/0LbvzOW+d5KsaCO5sxgE1JWnMxNP92yb9MXrG8IO9VqziukGy/70q7Nzd6EO
wlGB9wzbjpuN89FjvAvlg79GQKqNVe7qZgeS5Sj0Zyl3mYD7ccj7h/g8qzisgrM74eizVDDylzkJ
nzcCCim734pVOk3GSWYLOheOR2qsmY6wE8wi7v+3e3do2lJtEbO/A/8IF8AuhMlvxJBq7iTa8+dO
KgmD9cQmr3RZVZHHoJxV9xUj0OorInIwYAhjkc4JQlHDh6uj280jY9BkNKxplyIg2+pNwQmuC4El
Bac/rjNVQN9Xuj+1gAdFfN/uvBZmleJEFfy6M3o2oqpiDCRQINdNRgrmq7QxDbERfOHGpfiAjzVC
HQEsCm0f1MpbRvUCrtw7KSCXOgsA75JAxb41VKkSMzpE1/SS2558L4piRG24MIX+OGD9FkYFAUQW
OMFtaFLEWHj7vWEMuLLIBKlqMf5UMkcI+9QP824lg8XmTMVFLWYfb37YYCALkpMtPY6h6JiZ/Lmt
pChv1LLu9k61F/R8vuVzSqvKDzhQJNHqV5N/RMG4GkEJry7oQ6biEFRna3mzLGh3y9naT32ObjJW
WPYcHfPM2bdqGR0PBfSxqoefEVVUMKjVApgCu8D8amKg9wFngk8APSbGbsk1zuVo/qpi4DlmKtsG
Y1Xh/85igFqOh3e0iSzdvQrJez42/r3/4xBYi5/JjgPZXlHoxtpR8XIIQ3o1BPMTtPcqqEmjWXTT
xJ71JaYcW1+z1RU6XuoD3eIDexskLpP1oHxJHB4q/PESbdYww6UUAFUjOTgSpNxTAa3WkTpDFczo
tjBzjxviXghDH+sH5djW4HBHkwbK2aKbo/v2u+d2OEfsxyN7gYBjsFYEvKqjsKEST3ybKyVWSuks
41QlxwRrCq0ZyIZwb9RMii4dpDvh8fU1W2vMuqrbtuVIR8R0eRUQ6kNF45Jqttae3eV5dbfmeMsM
dS+Z9zTWrjXDBGSqOT9hb3YK9oWZ+T4bdBb4JCVuwS8esBDQDKlnYLiz7IXcQV+iqWoZiawv4MWx
u333hMPFqgkk+x63QJtJUyds0xmc/ig5KvZkSMPBaxghoH0LHLOXWsZ/eEA0ll3+59Sj755VamXL
ycB+1aEqQC8POZOMyxwIU21G3rsesj7SyNj4WPsNxCnJOLauPD+7smyBCwX0fxlrt26zw3+7lRCJ
H4ZST1DVI08/HxU9OqHCvVT/OoWHE++BTPPU48gaVN/gtsMtNYlV5YYVUaCq6xzb+btPLuTZdEBm
dVG8i2/0zuJap2aKHhWX/IsGCVasyMgfNPa4kDELosBbcSPql9tY9TcWw6s5L/2ltw0WoqxGrBGd
ZqMAGkzKRl9DDU1kQwaY8AyrHP7z3y3ZW8cSyAWsuZkodiAy2dVQrOVQoFF7BSYyHIZx+EIbGuf0
0xW+nuwc+WJqg+9hy9NfOnL9BkM69TO7fKwXWYiuv41UJKVA8TKLU34mJNXf9En6jSpAI5f/urd9
pQzVdhenjsfGU9eJN0DjrJmJ1qn5CdoqsQMeqlpIJ+6YT260QG67+CO2fDuKhhKDXb/nlZ4GHPya
+W9omqLHLBocJbMAcA3ogOfRMdG9oJ0ctEtpyo+gqsI0FHsHbBVY/cfKhYWwzn4uMaE5M7+pexcR
wL6H6rDmGBCGCWNcRmT3JY+WKZwNDXBO99MmxlSud4HarqEusN5t0ha23ePM8rnf4OXQjlKVzQyZ
ctEmvFrA8iosFIcjDBSGLyaBEEoJPEgOnonnumwLaJ01MeOhwqCjNmcrfCbsUSyYOg0GaD06gsYa
Lw6bNpLOAaxa0gmNibq5bJTkuQ0JIgeYZT3EBQ+oN/z+HKZS+bzqalIAc3SKmtSwm26h+4KshWee
+c+LDksLTT0ibZG+FdB2Jal+yj6Cd5hQT2a+wfBLHqrdAVCA9DBfIA533gyoirVK4fevJ4csfnY2
uQfATQXjCAjiiELNwgCZMPToksQZRgKDUmMGGNxHeNny6nXvQM1jCmRzGt645gVDonO9mjMv00pK
MeTIoDR8AV8eiqZOtFdTbJp8ZKyUGy0BqHKdP4qndvnMWlDwbhcrcDFWMuHwlNDojmEy73EN/ZzY
SnNANPf42zqooysOVXqBBituuX1EnnOUkkP/LTkK66sYeuNvdmYmS1IzIhGtB0YWh8OuyWMMGGUa
zAkslJbnq7ATei2e6R2LlmEeblMQdKdScASmSbbmeA9yefAUA12I5X10VpJYdmbdOEi24VlSM9Yf
UR0atP57uwThUrLM3VzOr1ydiSwpUSbyF68Ds6mK1316BR8+psmVfmmPEftib513T/pPbttdOB97
dXBQsfYx12jn15SeZ3m7xAiazP/JR+UOViNWG3xilLTey9Dn49nyMO65lInthftJHUqsBM85ifjU
1IxOc7gZq1RIweHhqSYc9aS73akQvFtXo5W/ZaWXIEwQFXSI+PTzf+XgyFjX3pugVrXgQmrKlJuN
54BztLILUw8W7//HEoHnk2UAA8PK7+x2M09urR5Wv9Et6PXvGAqrEJnPJcilnruFXpxMPsIjde0/
ShAabFQluAx+VTzXVpnd+IXEgUDE+awo6AL7VxNv7hiwdGrVkw8xsAwVxnEqFVsrsf1XtyQ1/05X
sfjjlEAfAyB84V2T8V2i8+anX6pfFZxX2NIIk++EJS7CzJ2Dv/QtjRjiLrEibbilwniX2H1XNu0g
BGPVPn9lTZxpzXMjxSFkf3bIvcmh2R5VxtvvA6zThDnTan62e/Pnm/tTRwo+Yk1e6tQXMRNF7Zna
UqiMeIvup7OjF3uos7wKhDIsH0tgM+xHEqPnhAFxbnkSYJrObEQ8i3dGX4644x1jJ9nseyf+4qy5
ReK7LuV7gQ6Qnn/RcX2s8zQFHmxHEwC1eG7cXh3jLPzpADD2h+VA1n+ibW5D6T8k9pv7GGqcihop
kMNneZGVQEScvSOc3+VJ0Sme//7nFtYTWyv4DUmsrvuAfeKDiOIYO0DwhsnEklg5+WAVab64Ehlk
hKQqX1Gwu2/ep0Qwn/zd622PI/VWQWMb2BZ8NJHkrn53YHYCVq6jnZrrdXtRPDwR1n6OUSuO+8jA
PIEiYxts2/CUpvRaIXszLt2cMpxjYtCbhnrEQuBQqLg/iT2w+BZN7FwzUq67EVkZNuDPpLfnB7Ww
2hyMBCLO/7+a5qDxNaBJbOKpvDLqUPxnuM+K2d3Hs1/VX4VvytmjMtuadq2Ks8aJYd0OX82eWh9h
IgStEg75kr60yv5Zl10zxUqgpXQt76c5kZtajjh1AgXaexiGS1qmeDVlrDQZKYoo8BwIgE7Fm0BK
8kTrls55gcEM+PToZnXEBK8lC1pLpWeSSdmgWIS62vBdj7R8lB+sA/x7jSchH6VpvEvsjYTZPxHH
9t62kxYb3KSSRr3KhXmYbLzPQ7oCTrjeGfAi3VCC5ya/GA2KSzeP94FnBbPlXqoaGb2JKz8JJPEQ
PmnVG1qiexDYM/3z/eH9Ts1Q41rfwv6E4VLR1wwDd4Whe4rjMMMV98VOo/4DU69WHXifHWrYQwiA
CqLmZg58rpvHes4Uhc3uro+D3X2n/FX511aM9zll+5zVMZY7cOtDaAGlz53rwslcgkwOHt9vp/Ni
LdCs5vFOFSNNMY/81XyvySf1L9xE15HTsV7Pw77RbruKXTNn3Pr+QzUIBKRDpz7Qta76zYuZJdUb
ZPvLTSoIlUPbndWteoKuaPUnKkcHaCvAwwccS4KMq3ovhhfOMxaGZ6Bltef9/5zZt74QufemB9AX
nqjJEJFTyRi5d0rqpwr8UR+cnyYNCxMOoqiYFY2GTidkFw9mPmUyOmiUyhbORLTpGijMrDV3SKyg
Gz7okAiKiuZZdMZhyQlnkchigThQ2GlAqb2t2Kjgjp5OR3UJAlMcQJ8eq6n4qBJgVL71gXTP0ccD
bSeZmS9+1F8mj1M1mbIhZPRx/8pY+2iu+/SI34tjyEZRLEs85TR5w/nlvq7RMWUd4jfVyb32zkPf
4/G4Y4M5Wpm3pRGDOCP/6SJUsglr8hJ7LQ6KZC9uRF38bF9JoT/U+daw1qqIaeMuQZ8qfkOfBfBH
dUGshuM7gjTPiU7+LDkAljGnH20rXjCp7sSXqONAD1cd3/2J7isoCecQ6ayk4vN7TN+grmNEnwyS
aD+W67FVkoHW9sfUbkezye+cqxG7AkrRlPPEY6JP1aFlL6M8FBRJ7x5v+l9Em15q6wlqMsLeJvcA
pXx3Sg+m6lzYi5/yd8Nj2boBTHlS0WbVxlGsx55aRfADUEHRXonWCVf9OxhQrNN3YXdw/oAV4EsR
nibJB1TxjqV33Zgj8d3cJlbQWeQLwwwotcT+nZNdVZMbnxyW0OEC/fcu5A3dHvVN7iOifbWNFpHF
o2MTKuXsd7iYrw+2ARz4BLC6T5XnyeuOJn/ULNNQDOT5f4j6G6YJsriql3KOjxtok7n3HKH0nqNl
N/Cfl2THs52AdDDkrEQxbBWm25QPC84/2hMB8toKpM77/2UX5qDcX0RiC+bGt3HNwuoXdVnTgtgh
Gu64AgkFk5EmYa640Udw16uKmf1+WP+4RR2VlohIxFqcQdgW8ksy8xFiB+aYkilT5TjXPWakaIdP
0wNEJXreh9t6Sp4E+dypH5QW0J0i04HXcHMUpm+ui8hmk+4DGAjsjJS5VHjz7cgweFGMz+pqpF4q
lYSb6X+z1k9rpZtmjYUe+Q67O6cvHneO8CAgYOzgyMfCOlXUTc1ItRPYDfWuHdHlUqwd70UHXFzn
MxKZNGbMMZjwhM79zS/9XdSrCzIXds5Tkr2gQU8WMSxtZLYXCuoX8s1vwzPxGW/a1qYrG9XLcjZT
SJ7FXo8GUgnWv7Ep6AYREPhMR64EeP754VPOH+zDOd3ulRFnzfodBaXrPeoRJsJTWDuZAVMIeebU
/YJFPMV16HaIH1b1sC7zo554t0vuGgmcelfsaUODnb5+eAmWiHF/FJ11NM8+v7OIdl25Q7WqhXwQ
d7jfy2XuTMowr6XYNHUOqyXZd36IW6Ej+DPh89B7PkAZDWRUfzx6abPa6dbupCGTJoTdlJ0/sLLc
K0o2BFPz9OBxIl3ejkqpDQ/7A9RhEW/GvO+HxI72YuzIBsEhACyb4/U5s73mE3Vb0RC30IT3IO3X
a5h1ZLNoWwLzrnFqrULw4AytJTFQy6uQ7lV/vOENcaFZ3fSRNriLFIE9v1ZE3GPJufJb3P4jKZT/
9YCu2mN9vAV+hQPAko5/vPr3AA/wQQ/ZSoER4ZLQQBbtw0xog24/cxjz+QZvC8bM8gIO6oP7HhEy
FV6oYKk=
`protect end_protected
