`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i5SV0FoM+ny7290xjjscMpVS6+OrLADrk620H98azSSK4SOhZ/DvQE8YtSbgHjfcrwWJFF7APVxB
651wrIypAg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b4s5HznKkBfPLK2+4/TK32fG0186IhLrz524hcAJx2T54TwhZGbpQnfYA+DEkCvT6qRfvnM2ldqw
L9tv1KXC80D88HFwk9q+MgEXZEZOx7mKw/VdGbbF7v7IQvvfRv6f6Rgj7eXDEqlAGYbjHOl26SWt
+lp+yp5gJ2bAVVaD19c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
glL+d6Bw2sM/WjeeBr3tF974Hg9tcP8Jbe/Op1F4OolBgZdN8jHnsFFPHdnrOC91tsz60S9rzCUS
MwOfdql+NFNIfKjogQR6q1EkA2PMo8Sly++25gNStx22TNWDmcZxj+8k+PERP+H9jzfRAuvmp2NV
/CEN/2MJ11M6pBMhd9pB2nwbvm0wX5biflQAMLSf2UGU0xbiIuVyHS7CRP1iTZDEeWDdS1PW1APL
fUxVvHc3VZN3jGRAlByw0pxbA9hPxQZ/tSrgrdvfZ2t7o/6KcRwHpsca2XTezAnaOou/hlbCegOr
cLk12DjsbOi2/b+fsIFcyb6cpocm6XzIk2pHeA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f/McBdlzSrQvVfq7JiJ7oDVli4RYWipBSWzNozk1gMFrYbygHTQSPM7xbNXdgnuK6bazOa76gdcD
W48D45txtxCR9j4OVdOQXCteaE3nO4a8ckQc9I0tnP9E+R9HK5dYij1a3iDrnRXSyE5jcIhTzF4J
ykAtOhqxvVuFA3wg8uk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pdd2C8u/6Tj60rZNNQIdWAYEOHlkDvRzvxzPmOHZpy9CuB035I2/jQ8vJ44gH0kRETThh59REAWd
6Hrn0OLhJyYhpYC/RhcnoAaKp4IyDXsoEhomV1eXN13ffkwSYVp/WAB4b7ZuSrUbObyKwriQS+ip
rggwgOsh8p0l/+mPLAoeFAlUM+tZY34bZ4vZZbo8b/I1pwogqu23z+hFHl0s0yMy9qaewT6QhAP7
30RBqNy6EeWQUE+4XipGYkkVmm47boe0of2h/AKzpPhNf6quDlyVDDK9L8q2qGf9jAo0AK3y+On1
DZjTfenaoumwVXtqvfoCx6bFnWWmF1a8sYdhAw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13824)
`protect data_block
eTIKjn6ZEyzoSQr1nAKky5Rrn8zpv8n517BplOST6/BqZotqpqJLV2tf5l9CA/4qCqkDSfNg2PYh
vrt/uaW/vffalyT44vrJWcRPXl1A2bVmjKxDEYHdpnlnJZzC7oLtOAQTpLHrCK14h/jNOtWHZO4B
TgMrMhb6RZVoMoN7svR9a9x59S2iGp6HFhEEuUIA1sf5uYBMEeMNFfhJd/UZ1NuX+ddPC+yQRZIV
dY8Nvw472GCv2I9GUCnd55KnKPW2mqPGuXN/6BqFqaE3DiPQkNMPpp2rhx5o3iAgreAp3hWRr5Tl
DI9wTu/P2GP3a5qaKd/EXdJo0X6oQFWVfZpPOsHyCbc5otFH70XttAXO1K23CZRNA35FjyQZBYdu
S4MfdLgJszAHRwzORG1UC52ZT2fway6Od3YzwDvqkCSZ8msvurm6zE6Ai+KUdKUtwAk70ixBpd5C
B1IQ318KGJTCxTMcgSBZS1Huo+5h6kDe1VOboVWX1N6ZW5Fkja/7VPd4Exljbdpn9cOrm9sWIuEz
P5bFkO70NDfiMgsuG5j72LiZU6kdr3QRgPoTHgCIX/+GLRY02EnA9hJDR0ZtdeqVui4ccvFv5J2T
9uZdFrTjrdcffKPLKYuZkiZVjAXNcs+WQ/kvXL+Z5EoD6xDJtNNWLdLh7lJS/YcZItTzroYeMIRw
y7uQTjSXkKAbBdPSORQin6JfmuUUkbGuh6dJaZ3PaK2p0TmXn5yjdcjGA49Ipz5Ddu6qTz0ogKnb
Y3LMQROs4aV/+o9Pox4AxP2EyZy2yitJKj6Lz057Uvly8iMR//iD6luo4H2iFAyZayxX+DR11jNG
88kR1/2mKwW4E8y0Mthyr5d52pxI+fOU9ZEJefDV02WUFE9ar1u7o7sVOrapRxzzZJUC9Tj4VBgQ
WmDC8wp2LVlNi1KlzkXmb3VMK6uqM83lCRctSTGdq7FYi0BQohMfSf7aYBZj6QZZoZlOxPP4zDrg
+2W5Sirr7lGIuIjltLI2GAlCDRvkSZTRE8PkxE7blPhOkdElXWpBtMZkEO1rZNcw1d3+bjaB1XwG
6CtPtS81Px9NxbugXJwzNS8vVzDIQ/j75lDIey2DNksTCLE24GCzzkOVZlFHxI9K8c16b1LN+sYi
G2jyVOX2Fx0vrV6iYM9/kOfBz8DF5288G5hWKaAFS1pw2FcggVMtNtiq7h6azPkCduWjO67wxSTv
x+bS1x2ptPieNSMOMuEVP89pTNsM6hOpFIoH68rW7/GYPuxN2c7/90zmds6X4XF7RjfVDv2Y6aoV
EEUMMv3tdGv0tD9+c7IgKepYp+/RD+gRomwWPSo5z7Cqk2MIshZzGmKennlRaOt3ZlQzC+Y8RSmO
59uF9EYsfqQYeGI60z+IOCiB5znXThe3GBRzqhziGG+8LXz6bGU20jfSNrradUFmwqzFxx1yRX63
dd8BS7I1rxd+wUx34U6sS3zEqXz+CI3/tCZAEYbMIAks4uQS7EcyVu1zUcN5FUIOcKWGpcan6XQ4
7M6F+B+QC+tZLMWoR0pFFpAKN7jYLxbTDDP9Gkgnjo0lhMOLB6XPxiy7UFQqtvMlrVTW/X9n5qtf
RDhRWbFeOYgEtxwUfkp6vOytW4Fi+aClfBxsgVdS/yleIdgIe4p80duR8mSbpEh/lDrvUISgW+q1
ceHIUTDTfBh9kn8aqls6rFvC3NUsTeZfj13LEhJcsmnZQKs3+iEFplADCpfNiI/5stNYDGPWT4Ap
pggzG2gAv+Jmljr9E/NFMENt0Q9DWOznp6YdBwFm5g3SqC/mMX2pC19Dhqec/mHZoDGqfb0sva4p
NFesX9Sws+UmPhI3BApl4XcN4txwW1y7x7eEHeecMCbn5W2joHWEzTQjI2Xo4pHKtggU/y02gss2
qO+vyZvERr4/4yo/6rrvjX3mpD+6/WtDCTE+v6SUrqGLyFhp2njtOmUc30LauNE3pHpowXZXV5GE
hKbl+aLVv1Nq7jNizDjs8muTzBL8ZP67go2dBn0YThcEMGIK3Tyi1OxzUECMVIkt75HaxzFeopvx
RCXBlVixsy4jNYF3Q2nA24a8C8oUvQkoeviAGEPWRn3Mmpm5irQVXV14DMsz9O6ybLf26GNEczya
30ypsTm3cusNRzjRUvxK0mTAZuuTwkby0sliWCcthckIP6GktpP2JAjiHkFcK0aRa5oqT1GXikFK
YrP2IPWG0cCj07wzCWhpJanyEzfr5KAPlgsvDen6gb3UiITTmZ5had3OM5j6gAMrc9qYE6lv56mm
x+f/HNkgvf9JT5/8udsa78Dzw1TWBUPqAJXsNNXgU8njj9Gngq6lG0AorwQnS6fqPVb+3ILXQHIV
3xzlcgqlhAc1PSzmeWgAArx/ZGqrOjiAr84KrYPC3hbBg9Hgxu1yn93ROlpu+A7cDUuKkeHZKIgV
YnVNCWWvi9SBOhyr8KE6fLjUFE6p/wgfxdKEceLa9xV6+B95uf6ncjgGeON0mJ0bEL0AB6MJeBz7
UBRzz0aHD4KNJBJATBukUhUP4QVbT2Rzro7mVVAALPBdJK16C6HmS4LFiOeFKe+CKmP6dGWrcd7/
ncUTu9Q9WsPbkaWLUaCJilkTxAmdfePXKARW2rPI5KrmKnB+gSr7+0fG3XSythC+MHPVzxzkZmLv
f/6PZqxLOHaoTvXoJw3cTOriXdb/2i094P00F/GbDv7EWbCOwgZiuBoyfnshocerTJ8SlsiM+0O+
sK4HNB5SQnhGNWeN3U5y1lIQcgOQQzvB2Fgu8HMrxspacEXiXpZAdpcKDM5rjY4Fhn90yXFLKK6k
8XVrHd6rPE7zciciEgLPuThRuW+a//8KNxp8zvaIbkPGbhgJiK5a88XfKHEPqHo6Q9YE7tRtk6Sp
Fm/62fhj+zDjn8fB7J9kEFw1A7Cx80ZFMaIKkTtD4mjQNSOB5lwABIQK51bX4Z9GphGz9cMF5vTp
7t52tCSvKbma26R14eY8ZX3BlL3s/l45UZ7QOEt0dYtiLZnj4xnfEy8lxtAwWf7zZZpwbcZEsxyo
5MxhOdwk9AJ7Bd3nDPobcuATmXxC84UcFDXN3SkLemGPHlUtvlc9TbTXTnPDJgW9oNdKMk7BgvcO
5L5qYEvxPeED6W+GfR6kDejtXeLLOEOr1BQ6cwqKg/BhHuEomQ6CGus8hLtml4MY2nnXwUns2gGi
bkdbpwz4YoG8thqudKC2O+ftjX01X5o1D84VE9FQ22rTXxH9cQSv6Y7eqlNeY4l/oAZY27TJE/39
KHRJi1YM4oS0tZQoeddRnk4uWJYOF5v8Ki/fxPmr//ZohRQy84i8EUx/aGJsUsL5baejLtxFdCIM
+r9Xppkobr6e12Y/gzK0ZqMTSQxvmM2SXuNPZz1Nih6FmayFH9S/H9gSXTdKNnE50UueWY21EMyW
lyKwDxWzmLGdDhr3fM9kWSC62NO8bRoFLcrQ5YfZlT3Hs7t8uBy9aExMQnmCjJDepxAM+YITNO1+
nqYFQpbB9yypciEv8Qf5Sm2qo44mPx5PbAiuKs8VJqD3OfJlzGxLJYOib5bkPZSklLtRFpSai2vI
7n7G3NNUPzdO32rceLJ3MzzyfNLVkX5QoJtWGsyBBgSRj3xy88IdkdI0PAiAOnskc2a+Y0oofOri
1+Z2ai1M27cDVMvnz3kS/ssCbTDo7iNifvl2NDALE/J03tWrWmF+QSn1H2IKaqTeQBdRC2HtYqq8
WXd7pVko0WlXOxQuNGpwjTZitfiBY1WPF2sEMoboDueStrccw3Gf17lVwDWYbr1V36MnP1lDbBP1
up450fdY44B9RPtoJ0r2alMsotFUKryT0RLbj2UIM9rys8K32glM+EDA37bbOkVpEZeSH2fuFVzc
ivkrbD7BtX27a1+KZMEyO9Gww8DgF0WoJ8EPVP5uJKebslXPUVhzUa4VU1fGc16HxmAkzfj6MERs
xiNHsfm1A8X4ulhPbNuAVU2zA9K6uzLz0TtPYh9lhH0I3dB63thGx/efvJy8WfZRJgWgigXkWw2M
ck1/YcX4tjKgHrnGQbelSREgbwZ8Nd9jt+zknyPG4JH3RxxSkiLCbfhukILg2O602NZdrGCWEJfe
puKyNMRW5TGMAIsGdFLeqC7kNPauBYB+2xsntPMhvx/kbq0ltwpeuJ2eeEObA8GahRxBFptAkNv0
lDjxVfO2TEllzNowPSkItpA+bdt5j8HuSXt4ApRkHsrq+q6csRtdUze2erdCvzbPUJKp90+O8bwq
sQaVwS9VVPx94FQdBJTaKqVMsj6ltmbelE9y/S8KgcV2YTndcoFAvA+RWrn1Brz2hcabJ58+3tbk
1WJXM2xVBtXDIF8Q8XikFodJeFZ+OaAllL6NblLIZb19spoPGTYbE7fUqYiYnhq/Fx0ttmHjoStV
nphSeO6DwZ/OuyA18aLhpMTqkVJiEvuSAUIPRUYcp6+rVmyZ6f1LGXB2zUMQeJwSE9XW6kRiZ0uJ
Ay4OqnfItt9xMGMXAw45Qp+QyIfu6GELNyfyJY3AAZ+vE6WmBNJYuDS9qqt1XPtUSG+Xe6COJ0oV
WXb23r2Gb7OSZFtShgZvXOtquHpQB3tZw9kHlSrukkmNLD7lnbo5OLLylChsxt1ws+Gp/bPkX/E1
zROUBOfGOPlEUBl38O0WqnTuczsvjoB3xCY8RzeX4A1mMBjvdJaWYBw2/8lfKMbtHksRK9Zg5rfJ
89GMo3dI29GRJeuHaqx/ZXvp09q9HT+mBqShN/URL7MjWTsO5OF4jrTfMC9oENF9usnKt5t8TUO3
utfswCqoocl94P528ygSXlaWVimtFTfio8Qop0DTCF6Tx//SyMva9vE5Z0LyXAZGR/J5rZY36ayt
DEFyAIYyba8ff23LPrZXk5eLwtJZaDzvgibNBC0Hn0xlFXkp23hZtI/zYJXxam0LhAYU+SMLZPPu
Rq51kwOJ0Y+IaJuPKoDqbjNZYJLDBOXfYCedqt03W80GMByX3h1Vc3Lp45FnCxNFud+2sW27jaiO
YA8+aIcAMBbzwNpmWfq68gWxz10beVfqF/nDtT+cMoS03SxULyFlAYcxK+ffAwmylxoCZfaXTddY
vTw/3yw4ETn80/LyLwf+y5yKLLjLcbV7UkF+m5fjzJ2zMGv3JWwdJusDWQM3aibNVwoRTc0Brr+x
cqbyi8hLW89I/T6uADzl36UKb2xdMzNBIqD3pPmzxGWotzVFW/Ej4go+DZ7Nckl6gHfdBltkUR0V
ojKaJ4U3c6Ww24C+UpKLVP8866gacJ3vQNZi6dBlBqXSLqUU1/R4QJv98UOGJdb4rpCLZhZ0SsxV
OR2A2jcd7mqWzk5EH58guIU/uSOG5DblBfo3HkhJgo3Njvf1SySHTjRU2AbHvwUAOuCnybRDX7cH
yk7O6jPoqUi1qnaZa92fDZLmf36Yqs7zcshH1MxqUHUetZySt0a7beEbzG6qjcIVAgX/yOaklx3P
fKpMJ/ODTNC3QK8scbsHjtLNP+lYleVWF0g8vgjooP3jJlqYklKd2Is6SLpzdjsauUD7PmSyqRWJ
wUIIEaMe4QP0eNmykH/t8fF9qjRvfWNT8lLJ761zWBwTJPfusAodVA9crkLvyDlmp9FL0P7inDZE
3pFTcrrb1HUxUWoZq1kwi/4l3AhwiHB4oDXMJfB4V3pE5DvtA++r/5gynQYhc+O3zOxF/b4AXUd4
Ju6M79dkGIbkvSXxrhojyJvgdrtK2nl9HcqDKZYybNayayvbyCoFQ55ORpmv9qfPZbQEvFb9ZwcY
SPVhFAm4g+JDCfGbBo67l7G7GE90gPk0Queesf+Uk1T/XBd6oSjsdm9NPs+TvsPfvwopWq6ERZ7y
BnG/GjMguONs62rLZtI5xYTyYXk3WF9o/cA4c/sijXNAiYcTp8tEElEjG6j2K3g5PFfQFio9YHQ0
g72FKOtBtBqqKrUpQ87cnoFgagKcSo8w+bZwOaw6r5maqG4ODr97jz7ysXYZQjPlUx0jBlUlcjgV
zzbO3NTjSyEeODrefdWB4o+zUmWIi0yKk+lgCYG5dxrveLEvX3QnVrgHiwQcwhjIrwpzo88e85ra
H5jIoNUfXCT6wf+22HoSA1l68l19BWHY4sLqjsgERFfL0SI42+LCJ621xZvNPsCmzyBdRPUfLdpZ
ZT002yxFNmVB6RdwtWOWj5DnUxqimnOemQZ+7I0KbTHadvvCPPSZSSmvcK+eTE5Q6h3c+QZ9nc5n
yu3GH0LpWgGnNXzhRFMhzKDWymVi6QNMt4LSVxSGh+HCCruE9KKM6N/YfcZ6YC9H1H592D86KWdV
djD/5AhONbD7Vh0FTQd/WItkkXBcb4gGX2RGn5Y9xcmBgwMQ38HhXS2aRBBfrhx9SabffIWNbf4r
4CBii4ZxaOh0bR5bJsk8bYr2IDASVaGgi3qUoQEdyO6C/83uQX5T+KmBXguSajrXf5ugJG+oXRJ3
cGrMl8Xor3aNdA6ZRFdh5gjqZN0PQHFlnUksjDEOczc5yUiJHgvE6KX+Mv3cQcSLndUSoJox7gKo
QqP4Y+t92esF+UQwbEGn43IWPfQLsTWyzBzrkiZcpZ8Yh6LO1Ne2UuO7uBhHSXDajuwnYt/2F3NF
iOGTziCoFcn0Nz8/6AdoUAxU02MhHdAEKdfqAMFDNlifFu3LQ3eCekUqmhmR0RLrRGe3aTwexDeu
/sgavsMz9fUafq5XkN4PeGWX++586G53Cwp5wiXffcM13vdNh0DH1V1E4UXWs9oLpUSIxK3/PvNo
IEJn+6cUhoLaVm3+vZSKpVLiLIgPLssM4llJdI6EB2wzPZSqMlmU3ubWfhiCzX9WVYbBxGPdtfpA
33AEc6zF/fn7ilqFERhxWY6TcAyBbvI5Cm/TxiGTrAxR4TJ5i5O7DoIroqIDMsJPOjm7fJ4N4SAm
tXzcurBZ862/43LbwmwEQopK0U5lbliG44dp8HY+mjd39kJsfRL4udFGnXLIsHtKYFS3tHRKRCPR
jf58YNt9GBnL4mF7T7Bx5v4aff4nvUxcG0Qkj+xvRRQiAnk6j0dW4ONTcbBB2uNF4KtDZuBOsPb4
SS/vaWl7WlWVYqrcVsboA/ogY6QwJ9IUoREAwiV3mAKb+Y7MSJwJOAgDmTVIYJec2OtwQxfnpybY
xjfP9h+oXruW94FqmzbQgts0o5Ewl7IeNw6nqLGbJ76TvYyz0TZgI4OT61MZeGNNoVKBAVzlS1Yj
WjvbauD6Ex2ZqufXcja5Ikaa6f3WX6GSaLOhaBU8xJNe63NKu+fHUHDlU4CMc8iax45QPN7p8ueA
lmLKaPpBDsZ02+tZfq0ia9OVxz8MPAEYgniXVjVUL4W15l3Q7sV7KP67DiQLilSZ1oXSDkDigKGO
o7jpZZMfkBWKOwJQe+CPGCVVRrXMw1YYVYQidBYEb++mr4vQ6UOFpqmCGgd7lSr0Gnb96/k4AKhS
1W8ohuIeW6UKyvZkteqg71k6oeTqhi75FZZnpqqIO2B3nOqDhivx10LW0i8dFirtaSdr2xIlnryo
9yXUCn7OR3tePXeCeierGWNlU9FITGqMB+kZGgSPsYkd8FhqhZTGc7shqi5NcgtZZ+oRTCgsghwn
2A23aJoUc3pc8gE3XcxaiV0BsMHk95KpJGt8P56AdyBIwmpcnr7Nml7xOniS5RjQbVM9ul7kxPpZ
Z9zCuCuWZK+wo2FgIeADeOT0ORovgkwoh1j0IbOViouTwrFm5MsrrcflpkEQNvZTZZnC5EjnYcxv
6zE+HSrHovChP2KKT1qfqFKBvYdKdZtW1qsiGMG/eVkKRfOzw2DsKkbqOHDAsNq2rYQPrMyfG9DH
15PJ6pwk0wUEJKxsAyX/wOwxQW3itjcqWZCaWEIq7JlyHrnag72Edlf2TCH9/fKUFwGv6vxm0JYe
Jj5z9b5+++Ct6jDQXbn+rGg1yuNZ77rDV0fVG87/0v5kamxe3elIBSD3ctuwGWYBEjeTdhiC26On
mHT2zSplMvotoyxI7bUZQ/JxSNKI4dcFGF/zH8rGZOTx1rFPiN/jsHrPHgWxNavUd0SSFTInUkHz
egDrzX9B5S0P5Mmqba50Fe7TbrCJ/c0CCbNGm6fHWthvwOFt8sn5FDsD0RydVBQI+iWOZvIv1mGt
r/ub07jZQElk/DizrDKaql5yFHuaTMuG264/a5ehe1drHVWKllHpcvEo5d4VIqhovSXNV2fBDKVA
xgNzix+TNv4R3owJ/I3aj3/dUW4lFBS5GENpk2vXRW0eVwzf1npST83xrUmf473Mbh65pPp1IpZF
lbJ6p1USsCeWKdMAxB+pMlnAp4nXqoexAuySTksuX9hrsqRkR2DvEPnkqgctdMgicF8sKXcW+Crr
hVj0CU3gcJ8ypNwjWnpkxj1vNzBPCQ+m0gpP7yYczn7K7mJ7nPVidMXaeOkC2eRDHDCgZR6HmQ3v
0Pwkljk5/fqmK4M5Y8K89F6ct7jLDHTowE9qHi5lNEEbfxwC65W3Yawy1yw4tZblAqRrDhw1+QGj
BONoTkrlaWNU+AnoKpSRb6jfJQ3yLFYZFQvSKjQNtpqu4rHyhOxJnZBZkFK7sLJMTnHmuSOG2LQU
CLt+AsP8AeoCkvCyj8xufJczoANvRNchgDWMeOdMXexGjUjdscSEwedIyxR1VcyalNLeOn0D5FID
RZRRiN3UHQ3XjXoKwmnUFqnVLOpJubnQu+qERFMtBaGqVJAOLPe77s+We6K6LtS12wD3mT2XJ6mS
aFafCfZMDN6C/2BsEkT82SAh0QLJheTvtgj0aZgt7n2DY8RAnbGESBCDEhL8khB12mbGJ41Dlmjc
ARCFJ7ZC7vZZrFgtZW8fQtz6r1/14lcJJbiuWFZIyrmh9Gznb0wqV2XCwPKISg+BCWGtVqGafVAE
GBvtr8lfY2WTP5TN/5q3zJah1y/6xUod60H0H8IGdun4aBFTUFLHVF5uNZpKICaoEfdG1x89kp2A
+EYOzWLswPM8EHzFU4c8pnu59RMw7MJQl2Cki03KMv+FCs9116UIhmWQ7rDx2g9U0bbUFn9IjakZ
dS4XHps13xe+tIHrP43YmUEfBjE7/Kzp9qSWQbKs7tJySkRk/Q6BmPx/mmxFNaN9w5UJzpp4FL6L
PL5WcRwIgjcQdPnY8i9Yl1B8gc4r6Yt4/FzbVTi1FBDEntj75sCMzG3eVH2c2Okq+Y3TO5ZwITCC
++g9PNZHewNVn596FB6nnUQQ0J5rFeXd7WM5p3kHGWx97OLd/STN+Xs+PuQX3xFuA2rWfKGU2DOa
jV2xPXitu/tMY+TfvyIyWXu5BK+o3LahnnPS8sk7amEzSqSveIK76nR3kF4Cnj3vnkUR3L3xE5Gs
av0M9iAPGtABIBjdMJG77KpT5ZsSmtBRc9r+HR0OXr289wkCcLPamjhtzzT41cEYdx7MX0kLoUXd
K13W/bf53s8fRNsOajP3u+W1aRH4dliUio0LOmDucCLZ3UpxE2WB+AgdPIP/BzlVs2mYia3LyrZd
fj6oLXKDqIaBMUr4OHSM5ZKNez60SxIg/wpRiLbpqCkxgyCmRkaF0y0XOQmIMK419q7jl12XwOse
fY5KbkbF0abcgx53pF9eMbtVXYFR1NV2l6hqjN/wK9H6exGgAt/7S+n302nrEas9oCVQXo2QWDxE
U3XPIO81EhmC4AtsATjihLNgvXqzaaHS3RWPUzqITqBqJadH4K+2uw1T3xhZ84/AAFnfA/uwPY/6
AKmczgRWbiHIOqONWbngAmH/FsTLuCqtY2wAQaBenT+MsjSoXnQy8D3kQrtmnATgDol5By7csUdz
/unEChtwBWpIFdATg1QF4Ujva3CYkyx33ZSloeOvT886RS7kUSZzXkTWItCCFgPqbE/O8A3gmFF0
vnO4oUJyON1aiUTaIgvXhcmfXcqqH5ly0UUpsFd0Gl2KWEsyKN/hCvfPZRDy19fLnw9HcUjC05dj
h7R9jhtev++kSZe2Noi91GMchO8+akLp7Hs1IMjwhm0c58uEktfrkIcO5PuLyf/6zC3yK/WTxMlc
cfvreHVA2tsLIDakzkM9EPoKw6I0bSen3Yf7+KrycXxVZzCSN8OV8m92vXKHgzDJ9PsKskOz8m9l
PYKGfxTz44Fpb0FiP/mUEeFE7I/+51aBuErUqBtNjvQF2qKh0CNhOeAheS4h3jEEwiuhQKV+IqA7
ygKyhmKR5uZOuCs7Gu8Hu3f0eILxxfr0vcrsw3SXcWY0+fCRPefc0whj+8z4QgGIzHnrxB/AVUuj
etJehqPkN4AdWTDHQZkTrbC/ms2Yte00WHPei2WDaPZyv6lgIdy9kymoPD332sqo6tc7aYiAbR10
bt9/WwZXaWMYI2SpIc+1mR8qZoyPeR9Lcra4rrXJXEXTsIZ/UE2HUHW4oEPR2Z9dUkquI37DaXy3
/QQAeOGHPRngCumBR5mMxTI+Ga10oGpJ7HPPXjmzXwgHQ3jTorC+phoYrlUmUtGd5yOFp4KOwqaN
mYWCM8aolX+emajTsSz+b5EuSgyfFAEfuHwCMhQDrp/YMErhjdbV878fdThQT7z7p25ZC6LFFEJL
DugneXTxNYzXtaH3JFMGa4Mb3lIGeOY01sJxs4HimFboRydUr8t/nHC/ZwgXS2peV+I8Znrwam1G
687jm7B5y+/cizJJAiwiI1T07kQWA5JRZo6kLnPdblcSj0kYy6EZ2YaJy4aoWiMOlWrRvVvHYuMQ
003sSsZSm0FfuaGv8G7/QWkf50oH+DEHihgAcWKQIGVDCRd1N72oWQKssiGQdNjRHbqgc1ePAchZ
++GdnYxoXuwTSTAraYvC5nuOrYeVnqIeKZTZccb6UcM0+JWNKfQeI78n7wlaRtUmM8Ktz84LCzap
OEETHEz/PgaTO5db08wq8xuIMLDGI4MFhuWHyWxzj1jrWjV7qzp4rsUNpFRIKSlZUYx2SaO37GS/
iBRY7GeTSJBVeHEuu63OqWRRs9EVOmzIT1B83PLicv1DPd4cYzwr/fHRkruAU6RXHGLjW+G9hJ2b
g97bj0/DHnwse0XK6a0KsRT4i/6pgqqD52JfilqtU22BM8+ZuEWICM12tJNuN96UvAwDhGyH7VQ1
Z5H/4OEA7FCTVpItJ1ir26GCdMGQhzloOcsLZr5Ir9mtBceDopBUT7JK1NSd2Pr+1Gv6CorILjnH
/JcN4euhGAUl9qeIetowUr6eErcOelv00NlFK9goPTS4hiqFM+5fwmv1iZ0Yo7ygAofQI+ZtqJly
goD98NOC4z2kvdfvDRGuQCdXBNtOVM+yDkYKwo5Vyfn5lP3oCfneWzEiQxZi3ZCy+jc7ebFEcmCQ
RAnPY0MhYAKeN13G0CKbLmiaNmKZ3lTtXxC5EupSe0c8mWyvgfvTLtDKQmnEfKVm6sNV5fy8s7w0
2Hh9svnxQPphoBI+v4IUFOungXxHq48HEwF3uAWFyzyPn+3eC05Cze6WfdWsSRU0pFNNDsnayL6r
spXwirgNYAu0qfZrUSw1BmsltZRviec59QYM+p01Gs1cEyeD1NpBLju9id5d50193gZtm1MKxc5I
IyWMPu85dVf3RnH9yt1hQueK7ZDp+Ls5TJfRfDkGbSIo+mN/0JaMGm2lz8unI5yfqkEdI/dbH1lZ
3YDi6srkASwb/jDO5nCcj1l7QG4qBpz1GSnlEiX4qXV2iVxg4p0nzu/gUXf9bQnMIyKHmrPVA9+t
aswWxMEni1+ePdb+zMBYSsCRNZGHwIT3RqLulBNTAkoWezuZ6vDqqncGUkxRMci1YybmcUmfpWJa
V1kg2S1SyED80COekhbE4BUDHN14EGJaCVtSgCyRKVpMVfBP9ixkFWTbmfcAfY7qVXx4SPPo6wgx
L3xRqZk7Z8HLLOaHN1J+BAgiOufnq9d/c5jOE6gQpWzuQ1bki/5NuwBqWrjzfhR5xapo12VFKaE1
4WnxjhEYeNzeeg2VFBcRgUJaucBXitNCsLVLFLK/tSY/eQ4DU7lfeuC1+dptwyIQp1iUrQL6nTks
d+dgVdEJzkFM9XuwirGq9Aloz75M2Rrd6+J8o+itlp0h7/tvCZKK47xUmWGJK+dQaqRH9Wms4rji
gMl6UXAYtuxtQ36bEm0Fbf0TV6zJ2Jlpxgk5+UMiRhrL/7rtEc7TclS73RHdOvrkQKFfSbI8BDZG
bXA4Xb7XW096UnVOZR/uuu15f6yHkgGxTlIoejnNwdb81HDTljcmw4zDyk4UHL5agVbkiuo8mRg8
paOUb0rZcGYssq0VawuS6W5qfJVTyRtVxFTEPbYbUSDkQHRgadhirD27RnVmbeeFtjI4wtELRv+C
2SEj1LIN3uaOxwoipNHcrk4ayemFeW/U+sam/gJVt38Tr8UBGbwVfLrCTVNlaQtM+vqcSz666YNE
k2QY4SGImlI7QqL9kefYCt0Z2CvzMYCsB1sUqi55/w1FhjF97U0yCkTiFU+nVV3K/pWx8gyC2p7J
xn5CVEXiUQummqTIiGL1URcY9KbEUdA+b15OdmfiXmydpWqeHfEfjg6tqIVnNaCIQUu5tGESoWNb
P8GcYtGp7me7FhIyuPC1EDkWL0sB4nsFQ6Rj/DMpTD/C8QmVyp2NUx+Ldd80QFVrIhrmJwFraMar
QdTDzkp6IgeFK8lrtVqK8NifMhF5HfProb9JyFHJOwTgrMorOKSz11lvKnyQx0D3TZ3MID+4ZTis
OrL7iqMSKd3Ms1lysRiyAfd0jJu4+8VAIBMWEMRoLzfs26C0oRevfakCjtcLaDftlx+0fiIP9QGY
nRiDRn1T6dcugwxHjuWnEoyJsGfD8PluvroUR6obmRwjTn4V6SsmuUQFO2gvUE1LfpXaHlzpt9Ty
w8iXyNbMRq1WZOOEC3ZqeanjDKSuIMf6MjDFnVXgZDrChkXKMODp6W991vfqoFg3y2+mOcf6ofFv
4JkMmFcCvXIIjrrP7lrPySjGTyJ+ZubTtDB1pY8HiFAZnM+ChehEEX8KfkQTBitj5TVbHPxk9gIr
hDZtOYpO/6BAdsW5c09pD0RvznI41lIhkduu6chEuJh7aMM0Fnpaje26+IldrMrNYYr0Q1ABEMPB
O/UWboriiH5OtwiNCRRMyeGm5HUcFyaQJHa2+WFOZJFXHnh9QVaOmr3eFjAyoi9Ti7xsRsZMiLMU
8VLkXcAtf8qkQ3lwL1D+YHpYDraN4Z0veUyQZvNRYfXvE8ZbFwLKT6h+XUDmYgrDJ8quqRaM3JWQ
CvZDfMUhq8WloIXHypiKDDYzz3ToJXKwKQx64WU1sgVEumLtJhNFiVQ2yrR7U9ArA//zNyfnO0xv
gz96fyusmKT7/EPdBN1TtXcCCQDt+10SEC8dWgVh5Sx2F9yezWk4+WGH2ZZqaSTDW2xMxNWTQqNR
E098emhB/kOK1KNJhWpCvDveHm7C5N/XYADFYvZP1R3wsbB7zlImtGiTJuNSy2Q/f7p1KV7hAZ0n
GogQK1TtQjsn/3IwbVrz5khD2dsqVlzleTUX88kRZcuoNJl2b3XKcIrR+nJLnocQGVYF+CKS+t5q
2Vd72nL/JNcJAGLGKuklVqgMLlJOOGiv4S5hueWcD0ttZ4LzAN4w8pkuoJCpWJyE5XqS6vvSI8xN
+FdEbWxM7f9AsSC7mTad/5fiT1lImXcLK5bBz4c1W4OLtV1J2noOSdBfBfpG+lcNGe9k8rZmiryk
DhW2kJi2+vBPmw/O9fpwOwcdl2HjGS4x6BavGwkTLX6qxL3oTEAIrrHpy+iXyNb+Op2dvGdZSKR4
Gx+4MwMFFTMXf4ii9WvcB8DGmm412uZfbtMncGo9ooErutZvJC37Lf414F9YVIZlBPh9RBLxhwL9
2TRdY1v0e+va8nPcBZAW91FJVZBxKdXyqkkhaxPObUQJcxg/f90cQd7cdZllUFH55iiOLK3WE1nu
PMDE/gkAaTVG3Aly3v7QFHpWl+OLcfgbPisTO3WOyQ4baY+Fu7qn7BGqd2EafN8wagWZF0iUqMQj
fCxRYnBApkuX+K561UURRufchTb21sZwYOy7xu+UUcR/YnONRt7AAI1pxqXljHYLFKiqHQYR06gc
+voDHwSfqkCJga55AVH0ZzHwrKKkagHfbZU942YgLgu0R4Seo99FYtycvgnqxN9qsQIxKkB1Orq1
p35/Hv2eBxQhE/0Xep1AGjXWf6vU6c2OA2mrzt0x3cb4SFkJshpZ1JGD0m+8uloSiKtG+1waVmV6
2kWSilJVo64EWuNh3BvvxHYS9KNDhnpulFk2o71WlAtRB4Ro2w09SywDHCzBk1Dtt6HRci5pm50X
fao3ZK8X49Jak33onclvcrEEHY44XEelVWRPqdwzrBVv0UVLTZU/gB0z+k+ibI2AKw5M0wk/B5Kv
Yr0CfP3IxraQ89FOmPYXS6AaDRatnQpIiRdtA6WdrUQ0MBxffvdthaE44t8qq6fAytP1hTuggCDr
r/yD1hEymcKX6QdPY3MtsA1K+ixq/PUPc3aZwW64ue99aE0rAN5kgNpdu9n2cGt/KaGNk1uyQhVT
oTUwqpZ5j5N7aW4hxGiAMqvFKNV71Cb+eS+BIK7jyxAslr4M+irhIksWp4wXCxo0zYmgG/mHWDH/
Z+qrpbMPkf+1APUmCjoc1GqWxO1UJ+Q98NZr5heClHN/+BHAVhWLjp08pjkG15WbIzPZURblxlF5
7s8y/rggAwKdWEbbUG7QWIJeHxf6Gkco7pC2tiBOIOTQGW83zOtWCqd+04bqnvdQW11F3jKx9DnY
pQnLiSXVzDc7GjuAmxfDDOm962yrgaIqqam4wiHy0eMH7wpzJ6lq4/l3kVHpehqtEpHeqzNjjqX6
fenZzV52N1rugz5p4imx/VKvZ4pp0h892NrvJ/BRNc5w8Y91RLTAzVqlb+NcejrQc2GWBd4gLz5R
Rs8ozNgUsf7IBQkvrz7pIE1zOQYtpzPbY1iJbThvWs23PmKe2rTVyVNl4DvPpe9ZXfGt5vO/eWHz
5mBcfCD6zqbggBHQNjuwDtP/LY2KeycRd6qONpjTjNUWbxPIOcbSyBWYYailecWZ/hIXEtdvCxwv
d3fArrRxPpXCGz20Twgmb+j3UEP9GX448icTjh85/z1hGlYKvR/N91oZFWX3ZCdEmaSu/hLv3d5f
sWQRM1itrRm4XnWDuveumlUy5qauVulIaXnern3zMAhj8BvIItO4NSdXlod1GmH/lqulBKsZ7OoW
vaDax3JGDjxwCTJ6Udv+Prkh2vDcXnh05l7i3m5T8z+UKf0T/23mrIYYku2ZNrhrp3PuYf4LwzJV
A6W8Dm+aNkbGzhktER0i3XRVujmAa+PSHCFdhzAMw7rME6Wqc19Uo771dMrOtLE93eKlJ9f83X83
k77LSM6xWtMqpeJDf3CFHqXC2/a0HgQxfaqUzW4Hdm2UI60gsgIyG/NggjBp/LPmFQhZ/yrRf+BI
A7CY1lkCu2Q9vSucqPUYU7c4CXyctDsTHpqPU9FPrGyqCyGO/97Y1zWkBmCd/68MBtRilUlhJZHf
ltmkaFdkcSD/W/I4eLYfIp3CTqLB0QrRvp1HuKaeCjLWjSL3hliuCnj3OvQehz5q97ajlZFHJFA2
NBpfe0tXmAgmIarU1rmnKhDza2imp+SdpIno66DGfjat/bMkPFoFhJsPy5q5fbUoOGN0ky6S/0rP
7TnHzZ/QhuVSJp37gdHttSHQV7ROOuXZc25cpTloVDS2556BaGCLZwKOZGh2nH6pdesXjM7OMEZQ
casWULsLurz7uRyi9vs/ecI/b+GU1Z/TXofcVjoAIQT5K1djYoJnivOfs71nxnJbfzsWoO0JtTNs
P7hfsbpbXs726WR9WnRFQdISVmr9X+bp3T0JZMKi7xheEiNYV8Wd1heWZkJNsjU7fgb3DjRLgCnc
67BVVPS6Q094mJxIAC2eA0Ux+kQTkhRE6F8poC8KgeOD8nC4cT2ry6dBU94dOcjuJNlDt8reUXkP
xrQGDdJqhurwRdet4ZUFNI7QMAgWdYoRKAgsgky76zEr7TtfwDN8a7rNxPZUbdMPSQxkT597IBH7
8QJ099ZEA/NV/pEQYgu6ry+hsuHwvAT+/Zw0KNkqIRBZhVWrNDNeNfaKjBG28JrsgMZFCIaExLEW
lITCam/8DlfDW0/QaKxYk6UgWib4+OP6dXzBFgEyhWxUMw/0HmRepV8veU6mZUhcdVoKHRy31rX5
3egPrYBKNMJE0BILS01fwnz1USBaaK5FjIWuOTO2d7y86m9mFK1DXfcrdtQTX6VqmxhZgnq1VDD/
GRPYkqsvUNw90bCH4QrUOcYcj5YBSTCBY4/RzV4YPbSmbOMuwt4ldN+nd4eZaGnIGJz8/nL0KySH
JRhzFcXgKrqlbh7pj0ocergTXLUtcMwCy3Y1ewd5361XIloz+hqOJbKNhBkvp7HVp2iMcjaIx6PK
jSVHPU9t1wT8988xpU1qzeZMhUA9Om5m0XV32a0+t7cSvrBpfjLePLZ1ucBsL7KYNjy1P+EUwgd8
Cb6E43ixvOV63KWKCQpWJKXHIkOrNdcqcbSUFLeTt87rN1n6Nbp+8DXrum/clHv12t0aSOpAIYQj
74F+MeJdOY1erOSeEXbywmdStC/vPtkC3wvnROkR7bL6KUg0Aw6kbVFJmoanWD4JlGMHwGmW2sG3
BYBZ1C34njrC6SboPs4r3/c1Ttm+K33OVqqTDZ4kGAqpmpMiZoW/EJysXUMrIDGAz0vACLjjSAAF
rsJrYkA7LgDcnaI/Ox8/tRiepahfqIxFgoh8EHMUWiOTb3G1NehhV2O8L28CEvzdnJvWQ4dTaiqk
0v8Wo5ea2psq6k1EkY3HdG+mw1h4oa8DlDt2Ir66RVcoH1qpT2DQZjKClJxPoqLPQIrWZqdjpSH3
6nenAjH43tRuXPUZl+U086zlDjW5Ny2baQsuhrp96Z03OFToHsMQpWg8F06Ue28PJRqwhRLRwhy6
r2JF1BaPY+HsURUz9LT3jf1Q0lZlf4i6bYsn2vZyXcTfoZM5z7ew8AHUm/r7HduJ/7Hg5NOBeuZp
hgKpEMnPjPb2vbr0cgSVrO8GQevaUE8mmnDULjf4VDVjpX3PeVhEj8k7v/d8E4PXhnNqOLWKMq+u
fTIm9xU3QYyTdd70zQxHsm4puA3vwdwvWUl2MM7D1e2sFDxNva4xL9qxgywMHrQfv7t4+ZV3NKr/
gtrxtu5A1qJaAkh2b3cBEiBLmN7t0vyNoKhvf//kxZuoPzSnypyfJ2Mfq9Uka9pkrBi2A95eKXsD
67ztH8kNUzNgNZmGQVoOo786vcNd+9khYwQZhIa5MCbBOdXrIBt9y/HARUW+Gs+A2/7CzeWy5W/I
uvEOkE7geEnPpAwTwoFqD4Zdn6/tPPZ8n3yYTBhpfoSVwKy5oNOESn0HVg/D4odUG+geENaX4Jk/
R60hZPhAzg7P63WvN3C3cXyU2/F1Bu9XPDKNJ1mfYWmePF/0PYmowMwHUhGyECvW+pxb9mmighcm
AtIX/7DqZAlywaHhoVrm2YXOpAaFRbOg3+nIaNaWkMtnMqNqza9kAp6q9ALArFLy4w0pDWtNmeVd
vhCY8bDxvr9OWuH9oZb3RU8B9+6dMGGvHKLQFGEQlBTCNgAqeUagOy2ra9K+Qg3awpsoPen0UW4s
WygFnj0ZS6BzpSoC0X1D+oVjOyn88wXcQjgJkcHU+YSoKucYH+oNO4fUxLBp41tRj/pq3XfSCSqX
QzYORarJQ597mmSwHEssZyurjW0lRPX2hrgHwSL5RfrJ/EAG3PVR2kHTW0HwhhJ6XQ61L7qJS+CQ
ITzxq2DiXdvSNOpvpBw9lJgRu1GOc/s74jvYtKmKV2S7SBMXcsupY9+Qy+Cd8Vl/7TWMXSSgeGJA
ZY6fBrZHMKwgB1en0RgoEW56BiY1Vcu8BaWzx2fuGs4I8R4wYYahqHXBQ3dAV7Dj1zV+eW/b/LTT
F+OO+3Dq40ontxxHhkBEEdgVO0tIjCrI7XWB11giAVuSIdq7qJDw/6yaXTPmglGEtc4Yjpzsnovi
GdYT9MH17eCzJ1KpKPq+KsXuVRU1gcctfpJk4eHZopi9/+mm9E1VJE/Lu4gkuy+PATKBr048XF56
NYrPgaRDur8mfGE2XVuGZ4r5a13/qbhK6o1HaeRwcc148XkbgSwXll3ckRUsWcXP1w4vbOscp2ie
y5KObJsEfrAo+ALioFgCOYixnak16hzc2glBzhWnZFlXCA/LhYu90BgAxXTAj2znJjr+jwsODhSH
/fNz5jYsImnjJXyTi5pSHjWWE9zoQIeP8znxedFr0SHxLztAlM3lnWmwAqxrNn30aSaqkW5dpD6k
usWT7f3M9TQMcEg5hTu8GrVS259h1jwF7k1MakTzJI+mnONUDBlr6HOUxftmIZyY2RdMiqm9XRq5
tImQuk9Swn7+fsC9Q/mtRx0qCNy5uxJliNDiDyIh
`protect end_protected
