`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LNVz1rea9NzMbeuB/wYxpWpB5zAC8+id+gCCi6npX04jbHGHheRT0ts+7F4dt0v1u15Gzh9+3BJI
WLNBbjUxMQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nX1ESc+52czLSuKKdtdwDeq0tNp+aF6jgwtNFJ6eql2pu7o2lDJrTJqRrK3O7GGOCQNv4SbAQjjA
JQR1kZAWKBACedP/a1vcmdxDCsdQef8JX85jCfpXg/G7O0esTj46nPk1MaEuMjFRifI8jJGbnlHl
aY9qGePmFcudnqrwPtg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dZIwWFGIPMpuhut1oh3Dn8pfai4hZPkaIZb3RSIhhXE7XmNEvXoWOKSkEhOadoPPPQcj1UkQSYcL
AkHFiviziXxdjaNmwztrdKcSri3jCsGwK7cbTqvNqEakdVSNzVw3c/zRgDmMJNBDtvsxyMlOYFgO
UY/2LztXmpnIP8jDis2BRELrHLWbYBPjbwueLGpj/15EwDl0UeKvDGohMsmtwy16h0yWH/e5YAb7
NrsyHfLRc6I61W6eg2+BghY97xqguiqdXlTuuaUal9z/3A/ejZl924h1yljfI+Mp8PpdZN3XRpyh
8IPomwrEZPtCCFSu4PHCDITJnE3+VjHda2MPXQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sB8ly0+ZP6ribbYUBr+jzZ6Fk4c2RStpcoJFRHS81HusO5yXvWhiX6TwKt4tvPW4Cdbf0Qg6VmCk
Y6t+ZkEWp+3gv+OdaCi98z9Z+uzVhRUHAdI0EdFqb4MMaDwg5o58O16uYDhKA+QjGAUZnfmTOFqp
93DMHN0QpVrgbUhtna8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
phubltgmQ8rHKwqYtpd4LryV05/SkHoyA/5XSEe4D60Vd43NL2RYPpMT26mniOl5TVLnZ1/TQVfg
cr67rEZ+H5MPHQxBAPqiCaCDAq1PbmKkLWaSRxVlMCNRGc9xp/BLwEC4CTEDwRVuQMuOiVjaov2P
3fN2qkJz1Tas64O1ndRyzOn3kFgY2EYfZ7t136DrDbpER5AE99sTNqXfWbkwuafjC1V/hy0CI/oQ
5slO/3Le94w4dIynBuzIYGZurUJAOAPaJAUtICQ2shPvOLunrJd+DO+33Ur1ECCLZFV/8HoB5Z5x
2iKLzy3DzTV1llJFLiYQMi3H91svcnVTK/m2rA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11792)
`protect data_block
UQzAvF5ALBk9fqQJ0QUJbXewcPqeEGBMsu6l0VXNC5YDTZQjhGOIQxErbNTYThoG8n27zhqzwmxf
0ls6DIeOWMwsde0ZznMSOefZtVM5yno3Sm2+RLBsDo88qYcU+0hJ8nI/UPeyLKdIIzH/6wuWEXyo
Md/R8UqGp5H1tbay2/oL4QQWlySLCBGuIiMmRWB/CZ+urpkp2Fj2pba3DzKwCsaBK7BybASvHhO8
7qxvDrvKPTIU8qKJ4fcKWU4tdUKLJV4EROVAU6KZJGh6EGqAxtOmi57JJ+SuxI+4xYQuEnBiIqWi
A5IbWpohMES1GQfppFKVYbYKpW5SWBRwJkkc+cdnZiBUmyYjmvkFKcsXXHc68JqwEzLLqG+bIwGG
ss7w4qggZnBmVPDiDO3lD1zjkUIP7CP+UCk0Ecrhw5pe73yut6DcwmUtOApzrypiz4yR97xzon2j
iRCOutSGkgp2q9AEU82xES10gGcvzlJSMBWK6SoN6gC+SfflFe0E82RkkdbzLLDW0z0hOvd+2BrP
XClrmOrZ5Qdn8kiYvJJ4IrsPCDJVu9afXqkep7opiE1lMh8t6EBO0IHXgRxjzP+qxNaiLOJx4tzL
CasMkknIVhnnkzvqM+YlH9JenaiElpKUZDIU2374SAQ9dvcs+Vdnp006h409cvZEj6/FMMF1Hoo7
CaBhzqfXKwYcGq+8NoItVNj7yspbGJQxJNV18hqjQ5khkEWjGZDABFYuRxG8UpVTFy+GNqnOL0Pz
RBsqidwRneyQx+wLrDlr5RQGOpqpE+x/DhWTeGsYy2kjyd4PJ+9t6my0PcrJn+vLIj7UX9jvCWBZ
Tnv1YQUAhjPOR+lsazFg0lwiEk5wDRpOAGdJKG29SeJo/SxZMHG3V4iwLicBnwn0KX6wiR0zJmMF
xtH5RkESzdH6N+zsqBkLCCSCo0HXpCK4Kskl4xsLEaZ1P7STClcxL6NYGSHzoMd9SoURhewzC0+M
OL83cwmk+UHtY26lAgEM7u1XV/+z3BuNyfY7uOuD1yVw+Crl25A3z2vChNfeJGryq0ATEyK4JXjc
61E52Z5zRbIeTpE0ab4Y+RnELDZXtVjIowSIlnhV2fWtzOeG8WCrADYoorxdQ97wWLa4L7/dvLse
c5QSPB5dM43V2R4EtNJJU+qGNYaDBbghNaLNhHKQ/ZozC8hGsI1bssiMC1/96KitwBMZ/CBFOCY/
OUe+ws+xhUa7HGAVO8dw888XGtFwuXdO0uXlMsWvspMXqo9T7rK4aTgk6z/lXlHeYtmtbBVbFoPp
RCHmKa6roEWaxamXew8+WghZCM03UTcXNt1PCtkHMv/5jTmLHTDD2z2woej+MmybMuIivSluv+/Q
b1DbtXVYJZCdxnpVUdchEhgeTYS6Okzja0ZjMFwAqiKRLkBOzCkdUzTNcIb05npiCBEbHPERgmdv
tXPMR46b571ZRjNoPZ0/b7vPrlo4t6kXVXttLfyKlD7gChwBnAjvO7vnoJVdgDhcaI8shKcOaLhk
GzksabNZp9IINgq09UHe19npZ3Y1754bstvSbWQERwEJo9+CuPVO+GikR6oHBnB/2Q7mfbltQ+Qx
ivyKUrcDEsoD7OhcpdTu4+HSLnMRvzm9jOszuxkhgDhMzKnUmRA1HIDmOzqL5OBT2x8pYy1Y2yBC
tmXOadE8QTOjTpt1HwNCE3KsOTdqliJ/hDnVqX2rNYgG/uRkWy8oTgNy6eedkehhzZkDlFS/3xcO
T656ztbfQqpWfpp1I4ch6PfQ+KF19Qghfo5Di7NAIGly6oo1bSqUEDrvEw8qeI4mR6X9flv4UIFf
QQMvjVGr5YmoAg+/CF1D2Nlh4L6XmxJLPMFUUVJOq8uAzYG55BtWaFSgOZCTdu1+OMCOwW3AOlhx
bgGB+t7lkRg5uAsabog9j8epzpQ4OwPVEIrJdaVpx/nAuBK+fDyFvAbICfws2/M+PBkerGIoE65O
HjDKYMF9PyasbzOuGuXxFuvbbQU4xnbTY0EguqIrJi3asGbq8sv98bAU3hcKUSU3ygyy+4qP/IsF
bHuAbG/viaPeBxlhpG355TNO+FRt2t3RS/HCqeJSvh+fzlvgXwG7mMy0ES0HKNvUZl5fd0kPLxmQ
x64jeZQDXpZG+fKwzAAE11dPJOUMPJ5kTKYwf7m1KLMQDBovFLiwIsVjNMdgyRTuovnYA0E3FyB0
G+0aXxN3ZqX7hOQdl1znJt/MZOhXPQUTerV0JstLFC4LM/lh+HLRxBxtj75L1PSZbNNIFamFHRC4
r3HEtB1ucazVEgw8ZC+2ydzYztg2LYwun/LZ02UayDAuouEx1hoApdoSyP/s4xlU01utubEgTrGa
5v5e4P/DRuu5zlvqvMN7/I8nIQWT1xigFptIyarWto6+lzcmlolQ3oF4dNWzftgTKlL3UTcI8tbS
c2DNsQNs6SRcP+DucMnY0EM8ud1wf/Y+EhkhrR+Pfu/WVZ5TppXiWiaQHKX6+ateP7KeMzHHeAe2
bz/g6SChd+NJNykJTR+0vVlvKcdnEYWPDvy/WKPE5wIKEkLZdkcQfQUhQAbmSLq8l8pv+rQelIi5
FDb3Od+o5AMP8+5Tc0d3svukDRYx2pYn2a6Q0FlFgYBHL1nGP4HoqLkZfwmGqgs0TbWbpJGmOZs2
5c/bsRe2xpALsBEr4JDbf1HpWIkTL3YKk/EZYOiIcOTRfbnMgTo3ylpX9QZhXUN50JZyEMe4jOtm
7PWlCGUJxWA5wbxGEs+b9WcwJN4BNPQHkNGByY3STW00rgurOxXzNxPATRuBEGH/bm7L8iSHPh3F
wKR5FUzUNDWZxyCMtaqFzb6A7JSMUoVUZ621StVhFmoClwCPpAlFWJy1BCwkFbXDfibmScPf9x1V
s8F8/MQgwqJAuuSF8/raa8Id/ccNwvnr1Ll0FKMyyypHUlTpPtR6ozHqW3dDeNcuZcwije1H+aTz
gH6Dw6RsjKbrCHLyYnBbtnyjXe+0nVi1IkF+/KlJVDDzjeqGHG0Y4HmagXel481w7arosNOtB3Fh
V29zh8fssBWFC5seZefaWhbKAFjtOcBM44+/AmfVaGKFh+eSgoWICZ+6eQLTlUhN0LA1BkoWNxxf
gckPGsIhhE4a1jsz5CqPpzv6/XVqKmNVt029OZL77r5LZE70KqMqgpV2K5grNtTpswt6rbXVEhif
KRj9aeh8KxaAZSj7GZfHXh1va6ZJReYWnQNv3DDPGu6GFgnb06e5YING9ecAFk5izmvPsb67013M
cDcb5W5886KU8pjx7ruat/bydnbQiMpnBGvkZfLA7U9K6+xmdsZvmBqfltO3IgI5LHrREzIDfYSD
mPwnafilbtHjSXDwedT+9VytuPf8axzfVsq+RHcaReY3iCcWeWld//uvolv5b4g0ZaxodOvVwd1I
LsoZAf2SPVq39qYbktPGrXiiptJO3XygyBSfH8mKtYtZMoXVnk4lWXj/I8EfM7+gx7UzdsfmVeN6
CD6xdy4VRn8y1MIzGb07n5B04sGQrnorBc3gZPAT9dp/Ya/m4lhy9WnEBYtNVQ1hZQ5te7Wp4ZZu
R04InNDnb7JdWPIppa1KVk+1bWzSAq6+0c+NRvYn/Ji+t6AS8qYW4966PMrasOZgeQoIIMSBF875
hhTlnQB8lUEPuFO9dDyH0SIP3soO4j167RwnGXlgrJLJr4eGqQKK4jChyE5Tq7BpOtC75MzLM0MG
tBaB8ImUYdiOlutWDrqO5OkQKs2LTz76Y6V4MC0PhigHNaFDUD8e55QWv3kME5ikNpkrX8QixRO5
cZmaQFM8RuE1xinN0iRuAcvLkwRyFVpL5drenGvMK9Tf/8vAGqEv9yxCnJ3/iDGzU9ISUkbCsa+z
m2cEh5Ot7+R7e61TBxk56w2fqK2lcMwwxnZmRmsOQ5mIva7+VPzSxAbO6nd2ND9PISkYoEPUT1u9
XnMuiPiPN+s/XUO0ByfzdIhNE82nlqB4V0nUY6ZrwWP0qY+bouEXKafZoxZCLvMgtQn3++h03AH+
hCiM7nfmmqu3toYxVuogibcRsXWoNi8rqWHsQ/ARu69SxPNT6stjW6F6gIXUoLhdJYTP1FR9AzaO
boY98L0q+gCt5XGGaZ+H/cEXYQmIprZOeYQaNhuI4alK4q50bZhHyNXwyjPnB1VJPtKXR+h4ZOHZ
GpX73Pi/glQj+nAdccXUxnTgIxtumYwwLo8sch5vOdKLcfaAOlsNH9qEzSlTp3uXRef8YDfycQCd
Ik7bZhdhEpjoZgMEefai0AO0XBOdLsg8b4pO2fxE3EPyFyZOr08P0szMnrKrlK/OW0xzWFPF1awA
XvTr6D+NRdnj982HFMJe+4U/T38/pMEq40sHcYAIuws4lwEQ2c8qnihiY2wyoDBCwFpYCZqlHodL
OTELGXM/OdaiMau2OKWtyR4VeGJhUZ9+qyp6sn0dz6DmkqGlOqtx9Y+EFMf0xoSoDyAjpqqY7u2A
+MZwFbOfUF/lHa5l+RRbLfcfaI8OftZgvVDTuumkdypkp13iSvxfcvuybgC41uwkAa4vZ9L92o9m
WV4zj9bpwsa9g43CxuRr3Jd0q101Xj1FtONm8qZJhX0P5qecdZdiBQHkps5sLcQj+LBV4xX77ynP
ZYrfFPSpWySqbn6npe9UOX4WaSVClehWjqznrIv2ysUGAUDxO1YdudCVR1YdFCQgm2sWxBTlxREH
eq3y7oM9ygM8Gp8jc2C8SkyrTr5IcdQmWHqmxESmWtCFkKFZAQ8PoWih6AB5aI31ySh/qIzWc01a
Eq+Ogqud8d/oaII/a9Sx8aoxCJ61+X3heQqXAxLqIztJ6c6yzHTGaEFKHw6qqz7RsVA2HvW6vM7g
EvOHn4S/yomudfsmcN+2LqPmB/qtYVEhVgNXkGekKrJ4BRYjK2o7W2APmVcxxV79ulJpF+P52+3a
pwFQxXwUdh6OSoO/F2cnuBItzoUMaK2GafIHb46rBYT0N57echRDQhmklFpvehAuloD2OMyaNiXs
zkl63dQ4LTy5lrnTlMQ/suvC7dAtLzNZ1DYbWNaVLld24skN/7z3Jyc4XgYBtOrTB6r2eZyH2DZz
QJT5F+bRkQ2nO6mPJIoJUzOWOs5tx8CE7xflS4ACMwY5b4F+aBRkfvGeiRBBmyIWgtZCpn6acifi
M9yKCnF0dYBLy+OsHJKhhVgkQkFUM/Njh8qIPHnh5pzfaB3F1px+fLdhFZiKjU+lbumUCDxobB6R
HA0xZMQQ3Mot8prm8lO6VsM/f2+OKlt6S76psa0YmGW3J9TzD0T5FEeccwF9WQa8L3zU4wb5s3tH
DHDkLZslgtc+rnBZTORMpIJyGvej3EG1AXtSUHjQtjA5FXhnqY/zg8BwxjBd1PYk5IbPaMPuVp4U
R3ICkL16GZhDL8PpZUGFOfgTmJT2tv+KakbwbRK6y/t8eHOL/Lb8lbHgAnQlTq+fOgJlDa6e6sG9
jpoEaIQxRnmUFOkAfLFfqdz8z9aYsBr+zujUuRMMS7I+iypNxU9Z+Y0QaiF9en79BZVFRv5KAtKr
kNssZarX41zAaovTFt1+4dX+9Rs+zBK2FL5h+W6YKSmpvG0CvLmLm7Au2N+KbhZH91q3ThgUQljG
dg7iO6HnM/f7oSD533AOvtmjTSAlLKYn7JCWUD/d1xhYBZMjm2TL69W89LG01vD/fXlco4Pp0Hw9
ST42Z9Fb0h0gVwxk8HcgddiBIaZktPax5ObWJbVqKramSJ/cs8vbeWpBfXbCKS3HnLZ2G/Ev4Kvt
KcM8Zal8EzR1K2AYu+GFoEOhgsB9PLjfx5tH+7hLsh3vcKnEl4OvdSFwRGep1rLZdWs62oVvWk32
88hntSxfXTs0VS2D8nkWmrpo3HF6b28NqbUqruuHbA4Y6nzefB+vp4QKE5gnNIkyDzgfl2yShiZq
zJkhICKbA+X39p0m7DiIlErYbIADqYKXvEYso+OTYOjMP8y/sU+wUlJnwrn1+CD1GbPjKOjSK0Oz
8bp30Ul0MW/Q5pareb6tOcDrCnEgR+w5EYM3kmuLU+dL9ULgH75nOzMsY8VSzU14Aht472u2TYVT
2GhFM8VFR6mMu5C0U99Mzurs7h901HDb20htOZTzglVPZDSpVSSSCr3miaeRh+QjLJr7pQcKqBNf
0qE6T2WISdM0adq1u/nQBZQoEq8T7i8lgyQXyA8+owTBb66EFXiNnemUSfq2I9AU+2/uIN/s3kZ8
yyx+bYAomQ5E+J9kUtuNJMcdfKKx8m1WgMq0uYmrn9ebBtLumU13dtdOuqNqHP3jFig3n5spVPXs
/YJ1ktrTyycysHGcLE9v5pjb34itLgQK8SkX2jGpnx15yC5PefU5ZA44mUOcDHpjaKmFb8kGqr4l
yOh24CZ+YuNPZhaWeBHmX8yNtRA+235aNwD2v0TVHUwZf5ohrhTskHAqj4+gVYcGatv1QuGpTQI1
8pD48yBeYznIktg+t3Mgx32BG+Gls7dKtp1Ojak4ffHXMIWuD7T5J+ftfTWERB8V1Y5EuuPf+Ibc
cWZ62eOglxiPW6ZEkjN9Jmxed7qC9PliytUPZrz5xI+abTYBQVAO6bJtqAp85aDKWi6fj33SMB+f
Ebtq3bNaOOxW3ZP7/9rOWvxA6oRGIaL68wz+iWsgCN77c8a7HZV/tVtkqbjkmaSC9yzylF8l3rHy
tk7+fPg4vGA2je0ts/IQ0rwN25fvscnDBfhOHUFN3KQ53ZPdW6jfu4rlgvt+I9r7uQHyWrN1YG8Z
ZLj82dorBozN+4RTXumyYf9U6Ya8pJHW6iGPc523Qm2hr6WmDB6pp+/C6VCFNh1DQ2fWDpb4ttKE
2RAY4WeR1yPBAakuGYbKp2lhKs4ReIrkU4pfdA+Qyx9704NZRH1+U0s+CAaq1apO9Hn/7dCUi0Re
x7AOk8pnN/tG3cynxZbPVYI03vdBeqk5Mx9l5+MZqJOy8uTLhrDSg7lYuEreSd3RKxafwF0QVyOT
/x2oly+VhSII1UG7VT4NoksEsagdsm5bg2nVR3oEGXgcnXS8cWvtw+hhSLoTaiSoxx2/+wZuo3Wc
wUn+SbV/SixY8MKW88MY8WNLHx7tapBSphktLQq91UKkWbsYbMvbWOCEE2+KyaaZZP6D1FZwGBpR
09JyifXcv3XqyqJKIWR0Fz6EYSaiKneZHmqs7ZDtWckI1OI+cQB0LZ4KhAlEJljy86fbhUNGd0Y4
kYH0X366eNeSazufYoIKqhAVTsd8ryGOFzxDR0NXNIoHNBxnqBhfiH/xsMOPJ4K80hlGLhX7Hy2c
bwEQwp+j25ojbA7RgKfypPrUUP5amc+Igk8UEKjLqyEJP2e+j7xBoA1b50OQlSffYtxXl1DxfY5E
HZ3Pcy7wdw+5A2WrYwxQTQcCy1ypvnMugf7pGEMA5PACsmdMU0puKWOHtRaf56p+PNPiNL4oHn5i
KoawCqWcsgvgJ/rNOKi75N2JcQvUdCJBd8P+LyvQN98hUHUD2oLUlq5wP89Ee2+Erct4t6drO70V
zeuh7nKRLvIi/NzjPYF/WIMGZE/+gt+O29Fp/2/53Wr+Y2PJU5SdQlzArBYZkT7DuhOKdw9eHY32
zE6oxeuZMKJ15dtv6tQdQ+E8GGJHEsnzuLtV4jvA9cNlpOX0Gauw47bvVjTQMvfSO2LHkFN4oSLS
6SBLQT7PW0NXn/d6I6CcQitC8fEyJ4icfhy2FHMYuyYtqn+7u7GoAh76aSEwQKFmw7gBsTCZlme+
MCYdU8cwWwp+ytVQ2gBCTd5l08U9irIz4ouaqWDfaKjcKzbcSlf9YeHWgL5MB63TNDSviQn4yy/8
s2bucw0mpjE72jcB7RENuzW/lsVleXew8RpPyWUgSiWFwxmLIEYJn/oUnRFuUbDF9y8cn9PS4EXc
8tGUYZPWGgfaq/9QwKvc0QbmKq2CpbxJrYOQhYKudQG6plWxhdoHodQmR12j1SJet/ufvEcimVOk
hjytEN5lglo3ixmzZLXcGrnQfx8ICStbMzVRe+xkvyoszVFJmAak0QjtpIIFrISaxOGr7q/xG3vA
rt3w4/G9EvhMlFhLYrlADg2lo50cyWJGvgRuBtlGHnENvjKs56Hrbry4OmbQppFSTDJ+R3qvI2sr
edsuhwwedOHVjxjHDAqm5mGs5hTDQjSogEDfSW+oVd5PDkk7vezzQ2gCg7nEgpKUc9e5Zl6NdLG8
N5Ig9n2Z4iftxWBFtgq+W1hFo9qhTOusBojnd8mg90HJE9r6wOdxBjydIrUepoqEA0wWkDNDxAeC
sGRfh9Obxnu/qvIMuYf1n7pO0Dx48rX1B0f9Ke9Sn4NhRZssX+PU4sniEtg/6WHDdkF3yldkN9bZ
I4E8FjETIXhK4DCkgGzXQA/q7JkinTRgCcNoRuJbIL5cePY19AUd2AjW8jIoujdFWBpJLHn+F3Qt
7jRrDCA+IVliotGDkrhXZuPx3pPtPsHg9i2imLjXloI9rS2Iz/ZXhyHofeYItf4+McgsGIz5bBds
c8+GAkBQWhXJOJUkMF0zksAJVbfjZyzbD2GhXOeVzp2wdA4z/vwuc9XXgGqp3IyMd3Lm4c93T4Tf
ltEVDUE2d70Rilbtx8P9OCkoeoPq5cBbRw30hhHm+wne1yoLGUc+OQwwwVFAGyWoqLOp/28yHRsh
EpnTTZa6AiDlTwaICNojcHo+HNBk9iY7BYQLmZvqcnv0owTA5TfCJGMNc75S/hcNOZ1PwIQew10a
mbzJDZ3nndKXdSY8PGIOkuAelugi6wTnWI8esRRKZLOTWKzW2kFTIbS3pyj7/vZAgdGXbTFOqEyv
uaF4O7hXQdB9a9S26W7labfoxC3jFNIBh/XR5iBiPyocQvMTyHXh+ksr2+KvA+b7MhXXVF2YZL4x
j5LaA1vM7keFQfFPmVkdkLExUAxQ2GMlurBXnXhkUb1B5vckbhQCRfiyH7aQgOIqsZHGFSO8Rbv2
Ej57mhj0+gTOdPjJZohehSeCsnnlsHzbiaOJJ74c2NhrXuI9SZzy0tGDKI4qIZm04WxWrh82NLWU
VqCpopb7za1PLcJOzSsMf2grdlFnSBq744837CP523+8GFFqTLZAAwv2CbRfrQypL/02vULkFXcn
U83/9I2IjoJaRANaC5HBJFp1z/2rfTaxTv52RRUH7DlExkzlf5Xu08l7yWxXekEFqCuROjAxAjgy
6r2qfPPHUEyP5mSVNxL4WFUz/hSDikZEidnvHFLKDw5MPpOhf0ghz2rcqDHk+2jMsaRYjsoqjnM/
HS8fqQrZSfEJyTUAfxdCTAXh2x6zT8RpFcKd0KoaTORiwurBGuifvvS2x8AItkM7rDRdKDN6bbEn
TH6AhATwS9PvSQPQmJRVIyWVmzTvxF8KSp4xFEHw3CshZIVKurCo1K3NlSPQtU5i1yYXuGPrMFmC
FYTCgktKm78yQOVUeZAbPtsJEpRgz3pUb8rDgZ2okdJVljCNf2cxZcjPTD0Ywr/g26WXDXC3urpu
JuyWNrwfkoPSESQuK0epve34YQXfp/XTT2IvxTiA5SSPBvZFH9HEnzfU6h+lWmZPlyD/la1c1Ec1
jgDtOYODQSv0rMW9D30Lj+9VUEcTJ9bvKe7TU+Oz2a419WshUun3TNkuBVzSlz3u5NlpPbWs3dBB
zk/967YVme7HWNOzE1LE8UAlaEHxtDTp3k2MXI7AcsE2Msm3YGBbMcpDsZpvhmOVdD6pklZp9A3G
7DdwI4t/2NrApkxC5BU9IJhnRMkuxkQvGEc1/J8IyQ/C3aLvH/lWDAmxZwHB553TKjANZqzhTDyT
R+TMJiF6fI89SOP93sM9CLpIyIkfm1GUGQ7iaZlxeS0FjV13NrNKDwM0DjQuX4lvLGfyHLg1ZwKi
UiRm7NHEQcWgazNGAJcuEXDdyrzKuqFQLBXsvtzjvn2eCRJnPcbPCjRv3d3XQ5GWpGsiNeVR8vnv
cCG3GUWPV9gA72QkQtVuzWLU4yZrXHlDOkOeM2deAqSHjS9UDE+DjzcYs9jSPUsRzaZUiKekSosk
tby7jjzuwXskugqGGb8Rk+KG9FjjUnHhE7SXy5KJ2LYLZDCDLf1wENY0bonbb+Iwp05V9Xvv3+0G
8qibYAedX1R7i1gWFZWqCa10WuEz9AB8/rZfxE3XVI2X8kdiTd2wJnvFFOJxwwHbMbeHIdmZsS2r
yimtoTDEcOc98TV7NvK0usZvzhFEV8jyOQEGupgGoyVUdllPzXJc9NWQpXB5tkqmTkjmSRr0j8S/
SxgrgmTLZg1yqPUSsxm1fGl8JkvNVTWPQy7STKCBU0jWR33K4yq6kuh9xtcU7TGeilXI/Ld6f0cT
QmALogb1WoOC3nSmXh0ANILqV6aa6VpRPD0Mj5eE95SmaqEtAoZ3rgytee7iBYEVnlr0B7HTdZd+
sVTFasQWcuakkOAErOjv93jURA2QOFyCZqDawfs4DvWNxCVPS8DWv7oo8jfzcYIzuRA5dMNag0tR
9U2OvgbyPlnvJSmH54dKcRkFTRIugESW5RpR44bdzpGu+etMhSiOMfjjtd/Urm44QeAlgbJ2nr+F
3B60pTXvdPAT4orGscEF4cQfUji9xfxFcJDzoEo0mUwnF47pFBpkRDydffI4cRNa8gr+HrCO1ZC0
OUAh2JZhLZtgEGe8kWuJqTraZpFdIgY/dl4vAKgREhKfIjbFKb0CSnAri9UL/UPc/NpUo8HN/aap
goFOgrQpXnhEtIhWmM9vt87QRW3E8BwB8/r+OzUPnOYpNpvTJA4FvHtGdCBHPuj49EubWnyo7MpI
dfAj57kUEQCdTNL08SWpSbYk8U0FtuaDiu/iR8Va4uwwhjvk7jNOW6xX4VORp7tTGRJoN5XEatYN
BfJHVKj1jX8U+aeiqOBGPz463bfuaiJcT+wmkfC3yyG/vMFeNatzM1lCX9aq1mKCqDS4ban1t0Vp
31Gk6JrKQ3gyK2s4AGTMmBIm4mtVXnNfiWmjCjQcgLlDXuIWVVFXDb7TDLpK22g4KjUy6s+rv+d3
LQtApIM8gdWtJKvgPl0Lux89s8VIp/DIBf94X+CLSwMiqv60peSq1PTQu9a3Re78oFsAEI8l7cIM
Jcsgwxf/66ZSVZDl27Br5x+LBtA8fAPR5TlfYjYTbVtU5qphF1WIxwlD1cb0pb5g8czvwYTB21vY
6ZUlStap9LNg3Y1iqKbSqm/WW86T0xvkE5PZKdMiN0UM9TeOPMg2TlhngMB1U7sGbqHcI2+A4jTX
9BaXtb54UVVXr4Di4RRYkgMONCTLQfhyt/nTevGZy6cx4YWVL/FpM/SkmXqaDHXG3bPmAvnhcGwa
5VjvXp6uBTotx+hw6ZwRMIZ2u3lQ4QfYpmEyN7E0bYTsNZHoCVeqVKjA77aIUZUX5inkju6hTcPk
s3x6XSdIWgcJqBq7z048IV2QoCS508T6oYDKmqyjUxSPBPg2rKOvdl4wxg7TnFc+l2LXbZ3fUaNI
lYcWzizVGa+Hw4DuBslSGWo0hg+A1VHxLkMZIr1A/tZqKzqDP7j8MGr04bavVc+e7Z/+S1UyvElT
nLlTskVmaoKP2SLS2q2kiuzM4O/5YOKPXZMRO9Q7uUdqVvbUS/He7+ehk+9svfotypNOZ0FT3umm
uUBeKYvz9FxEikyI2Jvf60GI2lfVP6vRPPF59MPs1oyNCDZYD53dSzbH5HQXUw7Y9kSfMFTOp3gx
9pCYICDcQJqXHafj9WIXMgbgdG75l3IsXJ8fhLTAZjvCcB9lVSlcJRqcKv1Y1fWUjZh3BMTsqYyb
PcrmElVBgsTqEEHK5OlIRQIW+J8XSYnjGAx0nmTSN7/7OgUk8xXkbr/dPnt2I0kXl/Qln9JrOu11
TmqZBdng9ADU6deHreXkCAcNAcTUbTXAuGidnsT1rctNWgiiwPeRWTVHn91NopjK10Liytrrm6vd
vdlSd0p3rCfrXPaynpJamSMl0qNsivOSUVfpSXuyQ044XaVskru6pQ2ryWYzp9gZ3/HWtuqpDa19
Hw7VIdulWtF6DmsMbXo3hDnCzzBHj7TGTJh3t5v+8d2PrY7m/sFcb4Wu43RlmzLLvb1UNH5prup+
lk+1yUJXRSmXzgaawxuYRHf5Ng5RXa5i/WBiVCY2ISD7ir4IAGrvd/MJZMDQc3kQrI+f+L4TNkXz
Ke0qVGZiWz7Nirzl+m5uaANFyPjRSKMRt9rixwe5nwoeDDURZmKxB2qq61JG2j+kICxQuItOG5VX
2dSLeZC5d4+Ee5EfBXmnb+vFjWyoemciNBfQ+mpDialRnl1XHBHm9HHsxy4OPSNbrJdZ1R3YNCAA
rv8Yk5GNnGz3bu3SaUCM8BwCwsTaaR6MJMDQJ4u5HTkN3dZyLEiF4aVk2uiOz3S6VVOUCSd369db
HKKiNE3HzWqrqp8s92fQyf8gQGwBXK8XqxW69Fndj9X1BMjOwjemY4XPkCbkVKAnM7zSWDlVdPUO
AO9EI+kzm6wo3zAtQdLT1oxh0BNG+E9bGa4QY2WgQS7htpiSWXoh3tTOMTofZoOCEENwUhwnfq8N
5foI8ueK5trN+q7qHydXgF3rafnYJvTXnvrhE+bUMFznsVqATG81Uzfl8s99j9Y9lvrovDLGbAWI
HLJfgV6uxx3/moNjMRfjViSBEIkHUY1yVEYPEcBJjaVsJJqRMcGhhFXm7/xuFXOyy416f0eLXPRP
h7uIxPV9SQoPcZkB/klhQsc/eVqsfzPORLw7tMi+swSwvd3iiqo6FfUT+r6b3Q7htEtq1pR475dS
P5FnlCp94iR5fwjXHpCBAqnB7mO29VSvc3LhsAffNg3wFM96t6U/j6qYqnAh1WDkgsWVeK1K0mig
1Lt7+7mhcxEi6Dj/xRR86WfB71OOtCMgtZVeqAldJvbU8p9whipelV+/MVDYgJJ/34pmYjuy1h1p
o9YXSZhKNcoxer2NASSnwtMmFI6qb6TCY8DCJ3QtRRLyuOvbbezsST0eGHMzO4p147XqVqKw6MLl
APIdrMncku8sq31sNzn6Fegz3aF9deJdnb2G5Gg+g6EvOGPAYzjWkqw4HkB36LBYKBMyoc0ObBYM
yte4zjYtLYuWj9RIMt/SzwiSsBOEFp2zvmD9rrBakPxbdLn/ByZ2/TYKbfvNOGTL1yYZcqjiUCam
JnwJnB3bX3+NbUIZX0gSsSGOJyUdDesr2DNN4Q6iw52dfZxG3f0OMPp9zJuzSGCbx99lbJ/x7g4i
orzyOv6cRw5OV2FgPCEOkB9zoF8tyFDtf2rvuk9nGSNjzpxElONbOw07mMn8JkvPetXNsBoJH6s+
xV+95AmzUiojNn/3RQieSe4VSnFBAkYIg9m50Ynn3Qdg+8I2wgdhWH+yLAKsFxZGbMtQXBsikCE5
ikybHieO9nDYRnY98XsYWugROH3m6VDkkl32mXcUz8BMNN3poTjBhfaRYz82RFDQAbuCHuW9NjZP
9os+BFNczItncRgV4Ccds9DXsfsSBbibqmlpf2yk/CZa42VqcEy2aiV59Sf/c0zNDx6aiekma1AK
R/qgxNhAUPNP3LTJkfyCTX/w20axf7ovGIjw72kdt1Ilnp7VKT0QeXVw4scJWpNgeSU8uuy70dyK
8I06Gpw6vZHFXix/YXXOk3mEwTaJmdW1j5YzsRXsB6jXHcCvfH+Aqy7ptPs5HDJwakfC34AG1I0H
rJOnVBg33R0nnTbCWShULcloVPCA5Uyk+H5ZL6ZjlElVmCHGQDn++kfKae466doLzvWuGALA0MJV
dE8pley5mudec+uEsKdAvLTRzge2RhV5tFl8Dx+r+eCyUuds/pNamf2yHuP3EpNg1zBhY8mAihqG
DpRL3AGNmDcsi6QZWFTmIXXGPOYu3Ohg/8cK318gQvh3ZbAg1Da6UjiJgQfgLA7oWcWUjwzdYmKn
iCNVcbTnFezFS15yQ9/Dc1UIUw8mLBPuTBYR/vkaRFpa1dMi50SeQkqDn00Cpr0UHzhsLKr03Cxy
4a8fHAlThkOxAFyLtsoYVl+4HyBsCcI8VcIoJ/sxSjiKs24vFKutgkxSHVqzrACtZ07hHwqgy5M0
SOPv/5VGQUDgHMvrJZBPLe+BkFbM9nDsjoscd3bo3lKmckd6Nv9ejlC/TKgkmbf076PqcU2v2Irk
I8H/W8OPorETjD2eEgBBD1LnL3VhQebqFXT1DekYqOeJWuKxE28fbIvJsTCgd2b2em0stqYBwI0y
mBb8umKZFgTjC9lAci1AyqMd0i2tn6nsR6moFuUG2xwBggVVEq3ouH+ir9R/R5uWsBtFm0Z73rd6
LG/C0dN6pAusrz8Y0jc28a0TgBehPHXtLdU1EBm6WQaG1oeEGY3TViimq/uvy+zLCi8VGMryo5fw
HxelH+dPG95ojrw2w/GzldJBqXOdnHD8oMweBH8NQ9JqOjgxHcon90qynx0SuvPzhQ+v5RbO1cuj
BGfJu/4NlnhOrKquVohT4T2Cjkdga2x2dNw7HLJRaTqbdgp2kUUs5aRkZEu4Nq/D9rIlQlOdVgAC
jCAGViLFBbmgAqwm/Te+Pjdm6LOztUWIhpGC+QNioKn+cQzjHPqOAg9RMFwd+jU9yOtNpKEV05y5
b8vswJ4kbJgq7mjFbN1mNfjUfFwtqQN5itD2ShokMB2cw5xUwtedZBxDCXtJmeSNv/qO0bVid0AY
F5xuxVDRuPgcQGBi/70gqS3dwyUoNA/ohZVutYiYH9CJ7WwwG5nH9XL7t5q1vvaMA81CpYxk/HWk
oF8mueg5DvgCANUBnYmT8UxIpSGcvynRVi0YjcNas2mxOahfckyNel+TbFGltSEN7mErjMYs14DT
PjtGXQPly4YALSIFKm1FJGEFURnnsuUq+++PvwlfxensEGUAkhhD072aeea7aBhjqm3Y+edyVc4x
JX5gHf247YsHlx3LnBuKRwbuMwbHSO8/RvTe2BwEVaHBhfXNcTm3oiuQ9GADdFraSRc8cRR8QRbR
BduaDXgJd9yvWdVTwpi4nSXWin7EKMcfziZRLkR1EXbwGrADJsUNln9q40Xy3X5OuDEz1qMBSSPS
HNDtroO51NOA0Y5WV8J67TdCXqVXEEAU0uHAk3N1ancCF0Nrg4z6gKRPRtd+zN9QFoZcKtIpj35U
bCtIMfYomD2mvlg53bR0+K7mHNOOWtsuI/ibtNyTGygZefeVtCJGZiBDSTo1L90vo+EQvKs8A9fj
FbEqfmJH1MwPKeaMIB5x8sm3DhVBAqv96w3+V/7jg+DMDQwgOE/iGeBn8ZMU6y1lmwijxN0SZz2l
fa1qdi6owSgWPQGs/12aOt2d/h8Yet4YRKSQCmKHFHeXqHcXs5HSaCXMrCYFfFOjehVQkZN/H0Es
HPSSRW4y+IJfNaJAkYr8OIGmjfdMGP9B4tlE4WNH1Z9NwsPdTErwS4vHHbN01HFUYbZBRjvj0JwX
13HrfJnpxQuuOm4jILB2k4/VG5mxx9fhtdH5zGv8tOE8CBBg9go73RCGT2OzyFo9pY7QauNco6+I
eykMuUSzWLxlcob9aljmignqxbvWA+PjyCDEAFbQTMmXBSfJxh3ZWRtBu2c+5FVPnppKH9w9BwRc
lxYHddUap/2pPNyK1nqTmeYFtEHjM6kEpg/KjfvkEMkGQBIawu79iFzW+v3gxMUM+8ySV1ohvZDx
GEcKfwlsUi0RQj9palFpz4LPoeniqIln5e0KkNfy6uoYb+Oh/9M9Kzhl0uWVm31ot7U=
`protect end_protected
