`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g86+w1EDqkH55h3Phg1cBsd/30gpVAefjnMZrkQOt8wkL0JSclp78L+cxzo2VUagK4qLQ/M4oeSg
72/Z7wkgLA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ya9gadlpf6wN/RVrEx3XLHKOR9to24rxJWV0IbMFp94MiSKpGcLHh+RuDJ6Ickp+nzXWuki4YYFO
6KKIpsA1ubLEEWDGV6sUQbRXLWYd4JxATnwaVtcMY5GKwT2kKEU7a2tN8IR+f4n+b02tqsGfob11
b9yGDFUo81Few/+BR2A=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRyUHZWmhO+6Dc+bqT5sXgQZ3pNikgfxj1Sb7hWUlsjmi2qNoiSE7/EL2/gbouT4mn4Arb42khaE
whKfowzhqFMh5xANyAvK0XU+C/qihy/56debHx9BLMECPriSKFuY7637e/O/TE+I2wNUoAFRTrh4
G8BIvMicuGWmBhSZZ07959LInqIdE+YRVUyNzt0GTABFUfuw7/rwfqHPsMZUVayhnRRYfJ+piV+3
Ne2xQsPvl5ytI7bBr6sDsfBXYwYlH8GEfFUzBAlADdLP0L41O4Rrzps+Uuhjw14AQo/44WWGJGav
+EGJ7Kpsn1uWxQ34Gvp5yzs6QajHpK40vbk55g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E/bdDJeXibOIrZCRxpN3N6R8ckd2Oukno7jCQpmC2R6DgUvsyRs4B+3s94zm+MFeyrpjwykVuWml
rdjV2rNQMUrLAfyc3OW5FMJDIQ1XsUUTXCHgUpLS7KV01LTle03SBC5aGKE8SU7ZwYXBQf6rBmzi
/wJcIyM9N20xRfezJRc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FLLP3KSxgwbORoyJqLL9l0mGzVYvVTwBPy4HbRo3DSxd6WAjh1peIBGjCt8WX2J7iWh1uc+7LaZk
lmzrxMkZ0VBpeBbpUAxcBQ8SefccV/tXQf0rP8W1QhnrdlbCtkxRMDDjwdRJ4bM+4hS/iF5MsqcA
k03H8SBLVvAay1YBSO4rueftsBvatFTLweFU5kp+Ag9Uk8sl/fcZ4zIIp2s/Xz+lv+o852gdQKOi
5adg0VqtvxxOIk4/Q/8kkqTwxam5BC1PI8CGiIGWCGBU5bZU+ENhSYtQYvkPd84pUVjCGf9fK/wG
fXncNhZAXgYim4Aa0LVpjWTrJSjnJqsGTJ73oQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14112)
`protect data_block
wabjrnzCU5R/Q92SNEVe9UY7r6f1dUYFZA/RIncwwUJ75kEldZdWsX2CYQ1TJ5gsFQkobqNr4Jn6
lnPI5ET6MXtYkUeB96tamZ4kglbxQxWpmzdz4Se0E7r3QZbERnoEYBcYJxrjKHgMx8WMCYQzHwEA
UDSyr9RL/kuPdEJqd6j9O58SpYhZHQzVpE7Mc41k62ZZIQpTNSQc3Ad2f2/7cZNt+wB/MnA89bdI
fUgGIpBKW0fMPWc3XkpubIygKRKDpA7aRa1ctubr5I72EZZhTFaPWeZlROdX4zzUfZXztfrScOF+
/ZJdifOa8q7KXT68gTF7Fdaag+MBhN/YEAYuEsIPSx7S8EvXqbr61BOxplZwoFsV8fKgl/s7FRoU
ayqfFZgDy36RbpZ0af/ZBIz/Z5dXnMaxDmG7r9ZUQj2ysABdDvjG67Bp8/+QoJ0EnpBFsfMLiXPV
FPtlNH5VvnOTCs57IRmWCFJxQyE6j1gkWwKQHHhrCY56gnX5dOKk5JYZNJRlU/5puQ43EKOtFSAI
aMWWCpqqt7BNl/758OqLWFy36LiHt//ee95Cgtx8/e3uzWbaapmwVi8kds5fkryi9buWkp/5oaKg
vNBJgdO7u9e2xwHi3Ugv2W6pQS59YN8nOmym9OIB3/e4PDxowUPjv+3xBK3NEaZKZ3Ls/Qlh7j+y
mzEeHJDj5WIPQyqiwVU+EnMjoCZzlQewlfhmQdKxIOl3TznpgQIg8OdkjbvPfpoUjz460ePZXtvz
DutZZDosh08z2bNTuT+B8UHAARk2K+n4gIawMZumb49h9W/xi5Ch5s0KRAOU3c2NZ9RG0UY2z3rj
bBSlktfz/n59NL8z3iEKz8knxFTCAHh5Ef3Ic0xNeEm98KF1DxhsFFjKYJ1Fgy8FIo4zQ3tkWDjq
Cui8K/u6+UGxBHMiC1YIfeBVufqUBEGK0i2WeRVkVLgmXwoaPRIPN+82M6HA2JxKsn9l3mB6AXcO
Tbt/CVAwsx94AA1WZkFGiDdCJ0z4+uJyqyTSm0twZ4NoFl1ocLhPRVQ7pqTU5MSPp9U29JL4EyIT
94Q+i2B5VMiNbyu98LUDYoxy20ios1SjSlU9v1pngTy1+DqwdvBYZb21LY2Bh2R8pGaqN1t4oTTz
pRaXmvPbafXtx87CZ+o/y8tVa4X5hN80ha6tw6X5wFxk+/6di3LW9IhXB5H96lpuU383vGIcIs5Q
O3bxGOfovqXhRlPTNSovXGUW0CJ1G8+XZXKwxWOxSbjobnvCb2cpeyzFpnNxWcvHQOu/ArPQGRCs
MadmPQfjG1dt7jVKtZhMCOHMzS5gESCdbbZnWG/ICXkf5A44e2mqDF8BUXz6squzc9d8v5bX0m2y
tfFLV0M94ZeR1/U0thEgVAlccqgOjpV9RZKjyzu7Ak9utaCPg1X0AO4SHzNZ+dS7Vc5MynZ+hImq
fAd8pBc8zn/cASf5cSPaX1yG7iN9daTX8hpDC9Ygktv8od8OHzYyHUV9NAhxnqYtP2zku37ptxx6
lYwt3/xH2TaD8B/8SMuDFOJf67DnnDwIfPkPe2crsbKVOQuaqC5BsalQb1KGZE1op+ZipqI8gbis
VZRHTSg/h9v02B25TDCW4n4LEo8beo7LGVvQ094UvU4v73bP/jbIbfougFmvDuy8WvjHC9xpkpxX
eEiQ1i8EbS0pMir8wVZOAy5NTPIxcTRoT9KlHR6YwN5PUobTr/aDDGPg1joN54uOVOfWiVqDvW2E
K0lJNoJpph5kPZys2Cya2hI6gRXfn2GfDOVhehfJQq0bRU8sJUivTmX5gU3dLaKqOWqFrNVWy3DS
HKMTSUPrZzaYfBBQwFkexsGy4XX3n9s5yIgR57btZJ3MytHUg1sSagky6sZXMFDCLC6XC7JBDF+Q
oxKcu4H480HQo/XNThywPvWEe+HVEl6HT7buLNI++YZpCBVGAFu8zj22L+pDtbZ2ohWPHO85V3dJ
PXSyupXvE+h+fz1+/Uf3D4DCZqAcdRST9xuQ0zmRun7ZAD9Qp1h2d3K2AHnHpxADrplP7mSfYZ6A
cMzePQJsNp6Ua4M5hoFRhDWTTfuQrIkBOZOeYUgVSazj1qkvtqUw2OxJW1sa5WLPf4ijUrb2PvLw
qZ3WtjtiOayQoJgRAv122ES9phHFRgi1Xu9vlj7+M1WWNIcS0b6+7cySu6tJqEfZ092wy3rGZG3k
EsfFdeMLwe0eGsh+lIYaW8y64r+gJhFnk+HQODEHWcOOcGNXeI+e5HMGcUVY5VpENxyBHPurMW+n
BvASUoSzStqplRY5V69ZOSQsMTGPsDtIZqcmg4XsB7HkL8gOFUxQxff2LAaPJRXCqxDdkCUaGNyS
e4cBMxE/gfDh1FQiX+UdJDm+IAYcZlJhke9zHJm7TEgZZAgf3+oBIzyCeuGeKhqt+3ONr9V1te4k
Z04hfUwXeInOLdMS3OdyCTW7Ez2ajNKfPCtXf0itofX5KpqSWKObCb6zgOFxp9p49bBofGjKGz6b
6OzA2MINRugk9HG+/Wdnm2GBAczL4UO4SvPGrh6URdFVeqrEGOI+DNI5/y/TOrUE2gTbBIHPFhSe
4MC8It60uZBFlO0OqeHlRg6HlsoKR2jrfNo5NQM4c7r564qza1raqLbs2otBnTYL3xey337KnAoN
ClJHR7m0U6y0MecVn1oRIXeGr1OSVBEAK8bho23LN7FyKLM+gJjrdCWrdFD+m0ptHsQmWIWb8QxA
5MqAWqtlqdjbqDTRp9sLGtwBus+0l9ihRXQDEMQcSt66+KvM9n6ohIS+5uSatdGAR/6h/aMAaMGc
aaE7aQW18+eyLqvFqV88wP05koWrARpq5+2X4cpglAPgQzwc5dcG4u0tv2K24lPgq7axli0Gop2f
FQuuUUcMYkbqhDQ36C4dFHriOt6WAdbz2su6DXWNwGbVFADiD2/NsZlwlT1jzvJ6wwh+iIpJzDqt
ySf9p4jDlYH8RXbkOO1I7iB2Mj9wKSfsIPWNIEK9fsyNjQCssmmuvoFz6HAlkJxdK7kpqH/sqOPN
WKAS0uEEipJjq2MNg2PZHN10XYkZhFbd3i6VsqLQ3Max6wVuRL8Gvrm6m+gXBySx7rIt3Vfb3xnK
1RbV7UIlZHpBKe4ufm9qbcKSn3Rm+rh4atlB14tyuu+603rnx4+6oRRNWJh/bU2+WhIs9PFZKjey
dxKPvuscmiPUlU2Dm6b68IlTfoI+R2g49XznlJXNfd5LxsmXt5f3jK/YsnOGJ35Mj2b0OnMOwmHn
hae4/DraTvoMG4Scb5yyDLW6sY/uVbcLsXKqfxK+2ThmCsZ00bzXMtj8Hx/mAA13EvHWggPsdQv0
VS3Nc7XC80xVJbghH+237k8UkY3wFhElF0e7O8a+IaEkPFj/OeG+yR0iKDW9MGoMgQGdpnkiHswC
uMKfIVu3NBc1wyYmmhAvV5Klw0pVcaZ9pCv1pbzzOVM07ix4VYPHt9QgrqnWyq84uXl9pzHkhn2K
iK3Q2gnufr8At5IZICPtLzr5v7u35Vlq6Mx0U9XhKkQ10lSVeFk1nlJ6DbgLwgEITe/ZYTNUegSJ
3ISOilmopKVqPFugLSYrivZTaCTENS6dixU7yJ5f71tASOSk8g4RSCftkvhdfp0gUgEtt4gS98Sg
YRo7/dpBmp4+4ho1FNeLViiaD+ACzByAy6X48llX7LEknR3iVbTZO7SUCKhOScPIGWfkBlkwBQWg
W4/hMwmJtim6l8FqOsZEPH3vMV2Hdqm0vD6FFOCF3Q87l0ioJbHiro6jNemHvq9mMV+U9mnkTBQI
CAajtk4DBBQXI/RY+GUzlTc4qTzcnSfSWjpi3RcGMxnHiBOalDVxNa8UugdtLBjh7mLaV8vwJdat
bBuHppUd5F7IPzXIPCJykJdfbql+cwYF1gNRgmAegkZb6+hniUqG1kLhDeQGpl8M+I9RA/yoDqqz
nbDgL/edzhqVI5WLHE+dsms7+3b2pxi7XfNaVNOBsb0n+janP2qNJpVWBIEVtTb73xlrSeDJJGTf
nEOENDmGK3Zt0+sIfEikGnwK2kDWReELcGTckDkI2xzRDz3mm8einsvtDCZUEJePX4a5jjZLjR+k
XhOP6EwQf2vlOuyVICNDHdztsCJCNELZm2G024v40cnnnyeune6zfDHw1l6INxj+h0p4N24RGQPu
S9QLJulhGxDHMsx6bROEkUgThXFiH8BhMUG5Jclw07kI+QrvIVaAI6bo+L2fp7W/A9icul4w8pvK
gFNNv5XiVr0mukzx5Lkcoy1nCeCi5cffmdVuoXcyJi4Ky3llkUrPiKWehmcFrRjwBebVaimCZpx5
EQUDJ0qds9tMRlI8bbOmmiKFkR6AVfFggqB8UDl0MXZ+8pAVo1paq5+pjxZYwaiXockbJHNz53lP
O2Zxlb708dmgpHLCqVetqEMt4HL42VmdOOI1p5F/k8Z8kO3YN7EPf55Abqm7reQiKIdI7uHINSI8
Uf6rwSSzjwg8nIvyy4WingYRzeAkXlfJkgrO0w6H3QI9YmAK+MXeFQgLvg56uda7wheE12HdvnU+
9lQ4AEg4AuaGwQHeGRHCeezoDj+93YfwjSUNo8s4eXIP2AFUhmSx4wqjm967zbDoulV7ILg7aSY8
JiqWz53RWnkSu/0Gt0NOwkH0V7R8rtvChVNHKj7MyzFbz7jphPun0Oo84pH41NvxGzBMHsnRRmpK
UggjdsRenzm7u1kPMCAiX1+qZlhHPd4Jc3McNNxil8VOykAyFjXeEPzVaq9j3sAP171ZN25ez0dq
BeUq9EKHErGiIykiiNUTTny3L+k2fUa5W3E0l9PBo4OD2e6l1+4JamPmZzwdcRtlht6Q7mvW83YB
b6IUyhT5YzxfykinSUrKAT40snTXK4rQgC7uhoMcMjP1jB1n0LGsW4HQ5yTUj9BJmJ2D8y6SJWil
7qTs7Y216GLxq4GqdjsZQ5OMO0cUp1cskpAnV1UGzQXzyMLon76B/vYOo7eNgWNdj/42BCcA55lt
S82d+/w3mMWau0b/+P+cH+J5LbZ+exQM4s4YKGBGHGxSQ1C8ooKxX4hk2AxQJSBODesfh82NZIMJ
DHqhNbpYIklPY2Pcu4IIUcfWMQSbi0wukjPEl0iuCyuPuHw4P0uh2YxWOyKSCuyxkv7BkJhFtgZi
e4nVeeWMHxASvlWpE4r3pJ1Xxk4AxAKT/28omzvRTOgVZuGZvGdsOaRswH2/6sHVq7ggw5izOIFb
YHz+7pizGvpOuWdF5Q3gUfbmSjBPA7akFlenU72oGGKaaqVdaq4vPZNElWIqTEod4LjKlau+eX0m
POP4CHjNSnOTt2xQupVGVbVrYNy8gKsl5B/UHNf3JvIytkMJsHG0z9i39ci9K8gfEJuWDTwpy3AC
SUffCDVkIEu0MfWhTqINRFUU+4xAGtK2bEy3rodtl1F2LHX//uVAFxO5GkOT8a+ufknaC7G/X4S3
2+2c6uR4GCCB1IF+VP+lAR9Q1Sl/6LR13x6iDf9a9JPkxs1jwswIeiiNHnvvTx9tP1wVMQH3vQP2
+kNOFo9cJ5U1dNMw728AtSQexUYFHmZ4iyXz7GvxJID8+vIIYEWH2Tei0kVnumUkLgodVWFzFHEs
V9pkj7U/p2JtQIJhjIjKBvwDTP/ysTHlf7WKlmRE4LdZUNegCnr9qr148dVxjF+oic1mU+vneYTK
pZ9GGW1Hz57ZqbGuNV5BN0RIfQ+xcTjCd5skpj4aCeF7NFu4jYbxpc9c871ydwS/ufrQkWs/a9k/
8vSCy4BiL6CYnyU0Q+jtB+xjehR5CjuYdSXKA1C6/g/6Xh/n2JgZpRk5VD9ZrIyj5aIOjk6SkLsw
DVUf48vjz5kPrLI7jIW5n9yqsvt8aB/YtfOEZpGqTupOuOWJ6pXbjIHrSZtjZ89L+os4Znv+givH
Ig23Xr/vvpZyP7Cyc1l3vqpp4a0F2GO5/G+8rUnkymy2hiEhMIYoCaIGEJouu3CzG19CJv6CHrL4
uZ2dZ/vJ2ZYBfLb94WD6M6c3F7aAe9rcxVwIjgFde4nNRzsDw+N3bjbr3h7/XaK4HDURAfLivYZ9
aTqKtdX5KmflQkPBZyliqqH8sFlaOAJKAAEaQut/Re3CMSUY3W7+IR19t+tsfx5Ri9nh9zD525YS
l/7iIRAkU77PTxt2PYpWTaHdh8lhdlPitWBP4Psllrl/V0QH0fiG/YnfVSuNpIrWVgGDA2J2z/gv
b8rA1iu2dtV03DzW/eigz6CCknKzffq1z0nKI98x+sEB8TSvRu8xgByWAQ5MIfBoii2/+n07eJYf
GR7Fhx+VbEf1gxCSlf7I5Wj6zpZLBXswdrzhTbo81qWwzSVNGPgdB9w++t5AZdla7/jHVHr8Fiy3
Meb1CmwpEAzdFbopZ3GspzTqkhrCuji+9+iRGIh63EOFRB+zBf48OVAtC5t0F3ORt7v4di9lXXCs
WpMI/5k2Vf0tmzEhT+6QCC0/owrT2mr8WSHfvSdPRkJb4we2tHDrdF4CKE/eoV9xMTmkw5bgOeW1
bcsFMaQv2dbkFLg2UHq0UmqwATDcJZ+1rh5AuE5ZSKMPHbb6zYvZ+0SZZfDmXN7suFJ0GClZN71v
bodkEPdWEYnMwekjV3Jy574xNb4PaIGiEiDc07mqS+Bg/wkhox08gstBQbZf/Ukl/2H1pxHgp+4O
znuXpnRy5ubg8KePPk3WxuYQzPG+0W6OGJYYO0MxPgGbhzRGxopg+9XdPSdG8bPgfA4y4MQE4Rvy
9tOcLD7KwRekV+ZTde0J8owaKRNV8/ThmT0YNT7hgL00k7jARGBdt8CxWGyNSkYY46Q92blNy187
27CBslxX+9BfQwEuszpH7j8bIVIy5TgsG6YewhWE7j9W0M6nIcnfltOhanKvpzlgiD/RGBEkxnlQ
alacAavLALqgAmnb8t7tFsC/J+yyYwwYHr9u47pyxPpF/d+pFnDcmxK/0cbTtjWiQOns0tJagz2U
FqM1v+sSTcL5AtCmu34/f280P5vhKnRx3++J3RcB8VnaMXX6kzHtV5LSx+FDLHdQOmpswoKvVLhK
r/HpXAkAN/eT7Wu/QmnaU9nUelh44gx88ej9lN4T4UrVX04BR/1fScUyEtD11gBBoVnotHPt8p3T
RzQ68bStPMJj2KB1IKHldWOgX0RgI1pRtwjJLmEBdsUuTnrOKiDIIO+8rJSUrCusmxi389psoI7V
bLaNpDW5oeiLdXHrH5T0whp1ShplnmwAVE8T5p13VjULrK43EvPWVQo3J3q1kmz0NkbBCm6+Ozi4
5UjTmZTuR7PXfXXOU/OuXds43DzvN96DBCk4WVCigDZ4QR8FYrYo3ccbh7A5Nc+cPlqe/b1GrX5+
4mRAtonbjw+TrObxcsUdchJPieGpXZGeIPclDiw2m/Bg8lPB72w7G7Wjif56Ariocl8d2wSPT7Xw
dLhrsZcm3IFNlJ5n7KzaTeaNEZnATG1sYsCtwo+ZC5oeqekcOPzAm69tZ46yFBAwq/OV6mVoDTYe
9IuDDcNJKgkFLOSGtSLVKxOEf6XUcXZ1RXS6ps/xdLTrRcr8aXgamKv2hu2b6nPVutvWdF7z/rSw
/gIerhn7IhvpOnVtkllTzcATlpzDecozJn43RMXgR+qKEoimrorVNy7a6U/PSWuNgsOuUgm95X77
INT9h+E9WUl+CaRP/tNck2h6HhV7eD2pzqUe5N08b/s6Pb8iMfLIOQnP0kG+3ZC/wbraC1jKagUR
LGpy7dc83gwzbGZDCeArpAT+U1BVs0RAW+xMX/zkvGBYlykUX8jHk6ZxuO1ZzMew+zpYc76waIQO
CxTCfY1ngw1vYlyIyJ+7nDwwQaHiy2cd02dLnoLD/2rF61QBJDxozyrN0aXTnib/oKKNm6QgsHNF
3ysPBjJf3S8qTc6Tpj8oC+kXr4DUjFEoSpJ8TuUxooFnV2sVngSr/ptdO3cJONy1Bg5JD/e00wDe
WgtQCQ8fT95vWwDQsVlP7sVcrtRClWbW83BmEqhx/F8CVa3BYc0bfpHHYmnprffa0hw5nN7vRotJ
funcg6ZyTGXF8X75fke7CaGrvEye7Gjmsz2sqWPQUeXCdQa8+fePAQ0z1I4cM7KRii3gLL26vSXt
on1vP9T4T10c56TYZ7DsCyS1Y8r+GHYBfhMXlhHq/bKVM9WbcqQ3d75rTO9VwPxN93NHkV5uwjA7
ABrY3ul+c4oAG2z+PKSuBlVQJlzstJyRkaHqraB/4+uuR0Zdc4Z8BZHNFgNtryUPhvdyGYo1VyVW
0Y58e0ZjSO2AGib8TcTHpjCaKA7meKO33W4a2j2aGKWB0tZ/Leo8TiGbZNgTOV0bKwLTIz1OBY8V
UvG1wzT5fa2RmkkZ2Vd19S9SjApc09CHmSebZ4YRaPTyJGXp6Wrnn8hQksvOTtJkZbvL4qm/RZIP
lTnArRF1IZUejg9IFo7qW4lVnAjqgZjI/NSwWWjlKG/T7VrqlM3G0qBeYMTrf2u5aAVh/hGPWP6E
ptqy7GPJfzLxOmswJD6FXLhhy3D3wQooT84+05IRj6qkKOHRk3+ksItHrAuWCCGGQcH8N0ZVyI2k
r0szRGt3p6s4eqzhCpO/ZajoF43lAAqesaSvN4B8OEuPhssy/9pzW9Rc+VmlTDm4hd3Vwdy8g9gE
NrlrfPc/7v6yOtLeFwiQDBN83YkKx29cZQvzDT5Azp63XptdT7aBcTYh3ReYvT9trel/wpoP4Djy
0CUyysllmZmspB61z3W4dWbrwgLWeKTKme9fZkzBOrev1jPGwJWQfGX7tgYLw+I4OZEnJkFHZMeL
bebPuMeJcA49qV8GS77NTV302dKZlMXNPuBOeu6v31i/G7d/RyHyDSSCz1+GWK3Rh0zx4YGPg98w
PaV0jLaJ5taNDqyem/jd1B5gYTsSnNnvXELWmErZ/MBGNCHHxUAe8RgrqokZ84j2nWZVlzf+eogP
lQb11QqSsOk4DexGP6DIxry5i1Vw8OyQRIqWokhKK7v1QXGbvGhJOJBwyReGWd9Nol068JX3yQ+c
90sAcr+1eJCd4AQcMZTA/NHfD1J+i6whbuQmQdrPtJV0ESslJawPy3DV2T3gE2j2wGPxddnIx1BS
2emg1caGu5JDpoBp7l6iRnexvi7JiJjU9ESFkzaTEwN6i4QjdeQHopS8zbGFWWGTOQXdWvM/oa1l
hgdreWlZmVOQMBLEOSZ/b6ce99HcOO85qw53EbsLknzojS3CeBolgkjIfTqv6LdG9LXSE9H40XA5
VMZoX9C1D9fIU2LjFc2NXFxMfAcrvnsxGZfUZ7g3OHLWhhNOFVkuW9J4oDrxXZAa6TxpOd09R/zz
UYlJ8L+yzSSLUkCV4ssTIC7lOZA/xmyX3hFk3YkqQf6OMwqxR6nE+HXEldHFw8bAwWY8rwIEpxqo
Xd5ud0VZYXrG6qwhJzF0YvcnrifUyVGcgaqPdapWaF0OGl/J5SNQjOEeN4iaOrm3QzMuGbqTj41/
ZLOgOpH0mXgPZjUrNSAmAz6/4ukgD1WJtdWEoWX/pS5cgt/AY8zfjrFYfxg4ZFGCXuu/TDYnXvzS
hYxEWLN/4PvxZFaj8IUdVCBbX9FrWjHfx2j/PSzfdVUAIUmWlRpc0yPlXMD5wZVVYQ8SevIjIbbE
Wr1vxoRwwCX/b/2cOxpNp3C6UPILfrOlhm+rfF9GbFqO0E+v+1JRSPrRve4/vDLgAdZL31MlwKR9
SN2jnygTuxYI+FuIfWba/vfxY+V0JlmKN77OaLENTsTORdeklFx47CT0i/2ztt1dlEe3aPkUjBqc
MTDQTm1kvwQlU1NP1HvlJC6uHL7oVNBw71BF1X11Voi0OOizBbCTim1zoe4Brh4yjWJWzScv122k
CyrFOv0pJCO4nCbW+qUOhEm3wLta9XWdRtgSJODHToci4pywO7fY2MmmJ2MhXugBqC3ciQBumO87
IoY2m1mwbcyflvOhzSFibzgvVy2g+lWHX1muSY6F74hLIkRWQVFJ8a5EHVko2h69ycBNVa891no0
LEzUr+4Koz+0/a2l+2vyypUiPpkLI1U/46GC/emCTNB8Wido2Y3jxuMQeqL2DIuQPb1FoCVG6ear
bbL2zorey6GBAm1c8+3aTf6hq04mtgrN/ycQ6bvYeVQvdIvJFrrXJ6gflrIqLe7CgsTBdpEkFpTe
tFVJt4rvv0KwkzL91Zm+s4xgzo2RkJHac/UKuoI/THyGjEZFhV4VIsYbDm0lPGGZpub4Ijne9crd
uWCdW3cxR8WodBfWamWYwenUsgmoQ3KgTpniWQkzkUstgBalqpwRlW/L7Rt46l/A/sj4WUOjXwUi
AY/NWDEJoeU3MoGHR5OABxN8wcjzznhwp5vzmHjcdanrCsFk0ZZ1nH13AIRjwtg1jVo1833XCzDA
WA6gTF7yu3dqfymuWYclAd/q1cgtmOqq6o4oOPWT99nbUME4dvKZ5PZENIcybvjOZJ6c/nSjLNU+
Lr6hfwCzDbLDU/Dv8vPZJMlhgMccqeBqVdYxzZSi9UzW2cbiOmaAi9YnVt49CTgjIqjdgq8r23Eh
xohffUtF5ILRAtXf+UUlVRz3k2OiMAd5kX3AAivkiEvOmTkljd55gITNrNxxIfVBRDBPy/GZCI9d
kwoH8GcuinVvanbHa+uzjTfH9YIUhkcyBlCUNX7LIjODkyAXG4NCCLc3oRQQHOiFVj47q6AeEc45
pWxAJYsAllyAAvcWFyGA+kR846ui/n8mckQd54GZ/wl0gEmXOJICnCVCVbMOdKlaHRimOxjA4NJO
cNm2zVdSP1UHcpg20BsP0w15Se3OYnWx1m2aiwDBZH7vEHgEU04jBuKQ1MwAxpylUc+vPj7u8S48
YEGoM70KVm85Y1OqvPQJwax+Qo9r87+7UWkKvB8yuoHLib1vPeVZRWQ7+Sg5RqkbltbQ0QEbjxP8
GAa9jsF2Hn2uVJLxHcQ17GvBPeIYYkmajlaSISQOwa2768L9hodNIX8Q1FtLRIEOpvk1H6819ZAS
Glkax2Su6vJBOIcSZV/W/NAf551Z/TYlaZc7k4J8sk9H41yeZLOuJsw6ESzIDA6wmTMkrpTfWIvh
tZUzch8EKBsRLVJffUArrT3e9s+8ZiUNOCO3dcdcWUeAOBWBwoqf032VQkwAIaDGbmjV39gYqQ/H
RDWq5Sj3huq+s77CMYPii/JUXij2JIb8FlOiZVT/nZgj7nV62TPvZ6KhiQcMvDcUIu/McL6A21DZ
7FVNQjqxPAlLuTmMjWNQUnXrc4QRYAb8wmVGu5V27XXdj3pwPHijTUgxWpqYyFMnWl+5YQzd4Rds
199sftzyX6rl+/IdIJo8hAMqScWeYTfgMkjnMe9ckR+JxxYlyraQGwLbGzN/gM6RFyxkUHVACZlK
w3x93JyonPeQBoxFDojppk/MJvMUstuqrVbouG7MtT5QSh+Cw6sY7zadR6v7aVGANAhmqEJ96Dgo
rSRdk32ugT+SDte9gW3YOYqojS2mWgNSZtAjPxE7JPLpXaE4t/hS4G5mRnIwq8AW5FU+yN9TyVN5
Hwi4hDZ4RwWDjlRjR9+l/SvEdFjNBR1xcUYMGoP9XSj7/KaSF7QH+W+L+XZmOeTX7mIQXv3cprIp
MOl5lT5qP/mTeqjLNfWbEKkscKDdB30TrSOYit1VJ8kGsGur0snB9pvMPz/sZcivl2U3j+OhruSV
364jqUqcZohgRSeSJYz2lN/KqGKbw5i6uYjaCR5DPPhwmEr1bUqV4fapB4QFWrl9WeUZepdFxwcj
DlUTsdK7bNGVMiqkQ/+qUgr1Ncuf9V945o9epUSeFv5YZxpFfNoYuMkQV6+21HFkPQ5pJ+a6bMbG
aEgIGH1zFMbsT+zuC4Wx1WrtmNHC0BEo6JMCFu50YCjhnLWGjX9YV0ZiIspCWiOU/dJnerh/AmPv
5tOM08Islis+kd57EPUC0U89dc/DWvJ/aMyqiztPgjz3y/9abZHTUoCFUf7c4Or1EfClkayUT/Lp
YN1BVV8RbCMdy9aWL3iHNrP7ROlB/T+lc61g0CAxcZ6jcVcwbavepV5TW+n+5rkAoSQQA6gsRXrB
w4vxxhqBfTer7cgGaskuUfgCbioQZE+wBuMgR6lwLg/NQcXSM1aVgCeOXngblFlFUhEAnEZh57sG
8wYDVhkTy7y+JW6/pG3LatjLNBLYiIfrLLTw5WZ5cSGtBYQSIC/88542f57XVRDImFapG1b1WmMT
AwDEw53fQWHMIzuEKD2vjcC49iWWGYdsEeLJIspXIrqF/Unn2U5CUqR8eaiUO4Bgvk1zP/94MAtm
VBhTxP0u7cDnShCducwcazBl+6OoSyvpH12yKMuSRIqjdiREcPoDXhXN5obTzL3C7S2TKuIvO4Z6
T/jkd3zeWgGS1lDrj44TAiNW5q9vscjjgUlr0oEiv2taXAx06l7CyyRDdNi7Wpk316rzt0aBo8Pj
aHJP0FQ6m/ltgduCq3HoFa7jfz7uuN1UnxVTbm7+4FdinhlHB92/fDY4xFwSqYjnNYt6aGz90MnT
vhnhaAX2O+e0lyw6SWLMUo2YYq2IZJ8nRWmtgroOSXXbR6Awor/N4s7sEf6u8IUsKlQqzt5C8Sfm
++pB6f1m4/FCJn7itGQjAB85/DWr1jYu3zt8DWgQMoSMLqaMFRKpLkTlesusvrlwZ3mEmDRe1IS3
wzHBUBWljuW9xO0r7Iheto/rCeEIvsj00KN/ef5ZSpcQprEnxAjeNtawgs9ZqfctSBY/S39yEykZ
noFsJoE9lDK6qagqw9pfHLtC8Fb1kYnRh0hA9v/eBRkjgUibr56FtMiQnOS0S/xsCTmRoJefSzwD
srQGqxeljFSb4mqF1oHLXW5hpNlB7D0oSqya5HALAH6xWroRYXcWvqW8YflCuFWlLv5AjyxpPwB9
DXhiX73cTQW+aQn0VTnf3N7Kr0Ventf/DJgpKo5JvkvSbIf46jDsxKiIgX/7WOKwvEh4uPZsAmki
j8uHN+BJGvO9/Lx6G7CVEe8Q77HD9JvR6Nkw2joyRDQiAOST1fvar6jFp+6D5ihCX7wmSXqxL/3T
u+CZbt17AUu+R1675FPvXSrOjXQAZ+Z5Gjl7b+q+1JOuBFGoxIU8Ianm6TLbRl01El3286AvuMf4
1F9PXEjghZfzLObF0FvQ60/tnpBwEAuulZxp8vU046mnpS807EcQqTa2orpkVs33Q/s8HD9ym8KC
RYBQer6vh+iYiT3Z+kr8C0oNkFGWvpv/jh3nEyU4CFI7xPKE1i0oahsJXsqpeci0S95wnDCQwXHe
pyXlxToRvgRu+UX2eaW7HRCVtzYgj/fgHJwgO8Sc4uYeZNlBFTgboSqC92wr8QCzTMJ42werTmKx
CGLdG+522fBjIOWyPBIFp2wtyWxCGyEKPh/iRpkx24j0O+bmWPEvOtJm7v4YvNT+ehauSIwAGZ1L
R/c9CFSivivL+AlyQZ9SeTYT3WA7CCTT1pZRvlevcqmcejmSqrLNscljh7uUg+oaZam7KA5Gpoue
w+zXoLkX5/g+l7C8y2iTL2F59xasXjItTBuCFCIHEiJSTZar1np6wBb273c2tpQgUybdxiz/uaxZ
yezcq4kTXT/kLFVS/CdgkUqb5/oMgnfbNn+Kg5g4owMABJJY0M8kYArC47LjtvlHRCxoWYH7tU53
JzgAE2H0IpC4D6/lhIcMyNic4mf3wnkKj+OyY5hJ2pen6TFxv5n3ULNKGO5aU21MX6n1+LYIGEKc
HVTUiLF+lCXHvNAoctMwhmpyFZ1gS08zqOVk2kJ/R5Nwuhq8p+K3aFKfKMJVL/c9CyIn5pOU7ltp
fIydF6ihUMqag7BG0ixSNyN3EkqYwzemEVFqE/xuwcBpMcJWtLQJ7fpF0RazjojhX3t4oWPYQCqy
obT9F2I2Uw/0DyLJsNZXgiOx46w1zLxhj5LKHFkvHi2Qx+5E0lnHP2fPUbYz7b4o67YIQMgoR9nE
jmCA77ly+TqILUcXfaCzYmVYtd8kP0cs9GT/xSMCL1tAelTqlp+vcXhML95SDWjoQPSkRhN7kUPq
NcuHg5kgg1tJl+AG7a0ZwNeODISXdH6+cGqlAkEC2THTIibF4GWjm4jrRm659O+mF8nkIDhUDv7L
DXN7/UDISG9efIcJmfrS4fJceTopKUdpUCMa7bMtaVQSYPJh9t+qxMKygCneF0dKUyL8BuRPL7MF
M87EHHJ2y3noZfsuKKUc0VJXJThx9mX/gFEZfkvefSwAKVR5DIFmrdajng1hLxC3KyOVw4fle6Ue
GxNtJy1huQHVAAMI3SMwrtWPrwg+iiwjpp7oivoeY5hYjpTyGMq10uMaeloKZsiRYlwljZCwBhgs
hbyYOFr97C7hMhYvEMXXocAByrKMSQrciWV649zW0DPoG/pN0MZw3pOQjT+nwwHEecxwLk4J/r8v
TSyFLQr+OxDnYM+ESKcemJrzeH8UqmAzdYDxOmOXAULGU8QXTt82iPWSlODcvy7aI79KfPgnTOMT
fAYS3Omr3bHB0N68Ycs/L+nT2eg2nzsiWwDRlN8Jk/gQIB6uiBIo15IQn+4/n/8meilQ8t+VbBY4
sbO68c8KDyxiGNH3IgfF+UBKmsLp+p9HVABZ2gHYQHpKXzkDP+FYZO/SvpfjGHafDi4trKMGgenz
YxcaVi8NxUAioyYiDW0Swfhyb3r0beVOpKp3SHzb3RcRHPILyZdX1/ZdeChr6/bQ7w1oK/G8jD7v
XQNHSuldxeLc1xQY6nhBYE6bVlWd+uvbgimzpeoaIa2rZTQ0Gw3gn3+Q0vbu1omBOGwOjSUSV2ot
HZwEUQmD2pcbdyKMxy+/PBLWYn+wAQZBrEu9NwtcGzLtHwjPRbsaVtkB7AbrvLuYy15K2IWbNV0m
/4+0xlPfS6/s8C3glXoyHUgwHWVcYrGP9GI8wzh7TFgAbwcf310gH10IPVp7rjuF2/xoRbmxxqqy
f6qRQuy1M6uH+CS4siIxKZQdY4122gqGZ8JYALpUr4lwT7gfB+2SMSUh+KHYaPT02eSrl0iNZNlw
+udhb1jO+W73gs6G5GXukj1TibugITpJ68uPsBgxdqelszczYVa9dvz2OAD1BUlOaYKbwSQkBD6h
lSFtyyd4iHGgCe7+t8zB20mQnQ8HiXCOiQyzhjLAAyUu4zzPJxQ69tPS5d0qtuUBw+MsAYvvXn0o
WF3zZRHE5J36jkMyt7ydhen5JFnaEd0XroD5bHrrkRDNpauX4tRijF5m0gSZz67YvCeXFVx+1Me8
RzjPZq212KhGBkGD3gJo1FoKQRlh2osQgoUkCPFL1BjBbf8XJHJHBA1RG4NRcuoEjdwZd7KTPf2v
ybnuXpRQTM09wdIRkPBbkWGd3FM7FBEdXJVDqhPoHb7xMET6F38RNLRZgJIT/N2iG5+GRzW8JuSx
9d4+VMhbbzA0uQcXEMpOvZzyRWtvih6jsTLsLrfItcpeZaTu1bgMowVk8DxuFbyx5N0fOgUA6eXa
au3UwpIjKwMTpq74GxJ0ThAVF6u7iqP+cRwpwiPOrlSwVl1xXXmhHH0308tKA79dEyqrFSPZSDR4
WRNuaCfhmax0iqnsUlGDYZsKYL3Jp0lTFupsQWeGxAIe2sEmDnOdMY4626ebu6v3wM4IAuW/Th09
o9HvhzWtx4Umll+9ad/SVw0IWOwZWm/InLjepK8ZWRW5Hf1ZkfSkjhIHTbs2E7/JTvR4aZ5/HX5Y
JGiqTN++AYzXPRrMB7qNhPjbn2qMnzl0tYMw7ovmllawdEewigjWjslUAHn/GAdm7uNqfnW754Wf
RWFUzxg0JMuL+hc6wHRutC0WlM4vd5fA7YrjTWKv/vYsBIUrnDk+eEBguCvh73j6O3invaW06Cuj
erwazI8Kg8szUGR3hCR7OUB5/FdctxkHrBSgCPRvaCJcjaar7GzFSpKMv+yj+SAz/wgIJ6/ZgO+Q
wCKuazO1nXWxP5fBe/Qptxb6/R9HJypADVb7HTn5Xou9hhk9goFtxqAxQg8sAxDQ0BTRoSYYIKKE
z6LdVlr5tqxMV7tRit9FnaaOOlttAbaHnOXr2sRdq2SJdSPUyFzYiuFNIBQwq7d6WirihvzXazcw
15Z9rrQgdSZ4WRk+ChwffHJThUPgJ6/4znS4w35K0bkG8aiPmsOXiQyJuar59oXcLQ4fPqMVIbKG
PbFPrVLzRZesdufSDgc32YZJlbxTfaG8QdDsDlOYXRXAYpnXeF6DGg+6ZGIUlxmWxt0OElp4clyU
Fb3cwSZTbF13jxPi0cNqnI6tRSDIc0OSOHxBDAlXExBrulIucuPW0ehYU5ow6aXVQ7D+fbbNjHgt
IBXw4JWOoGjExDJwGXkpUMUrk6f0aTA4YvnlgsobpQFQx80OIw1KlOW31YQRjy8OubzL6q49/Kuu
GFnbr732uVNsqJr9zltmjd3BPE19n4NB4qYWDfHltIVIAlXKqpu5Ar92SVVzjES+QfmY0rVyNNjf
GDPqILNxMpd13i+0WAmyJ8JGGGdjzKZyMeLEPcnpTGTEaC3UfbZW+HmrD5qUuwQT5A7omzWMgErV
UxcVSn3S6+prUqpmalKmP9NILWQGgSJydtVWgnEyF6IO7E7iFzpCNYBbNKr/ur/XHN2lkfenxo3s
h5H9aqBr4/wQzAqqDBTaonCNjsimmYYH8G8AbdMA+vovImEkXCmDsSZ7RMSoSzdvB1iuW10Sn1OJ
YCZ/YnzHP5tOyl96Y3mtttACY7w6640ngHVRvhqVI7C30QaIPC2jhIz+G+Hd5b9SUzCctdkJ3W58
n3AphemqU8d6YClTMzWvpJC96BSjVA3o0DBwG7elZz0RHhKgIfk/4aIS7z6sCZ8SC0Eq5V6fCVaN
4NLSw1Z1A5XN8GjAyLZQEYbVsilb/Dxa/UpmfA1ai7A1re7j1nWJo1WrNQ08VXVezkL0WqxTF+cZ
e4j5btO90oXSbKcednpKjDqRHEMG0apDzoToHL2D55ztWhYjSiq2UPFYU0Q/ECqQx0zp48Q5MmaY
3UR06EKg6u6oAoqt2gxvWSTE1GcbpYDxzNfnlEQV/08C9L9A/vkZ3kMK61DCDFN0XU9HCRa16TsA
h+nSMLl26Gdw3ywkD4ONvkyt4Zu3cewhmZ9B2dLOgshtARDbCELTXT5TT1yPm+kL1wzpCtxF8owe
C4wp/5KkXN24Cc9QR7svRiiEv9/LCxT2HZqgWYtdfS7MyVZ7hsKqZ1uQBC6dq7Z+al1SWfd6Pn3d
2CdSckeCu56/wHATKvPp+2ZJgZjO7nSMYKfMMFaRuvOAt0g0Yz6N+8nxuDQq/Sm58+IQG27SqQVc
3rcqrO59rlvFcs26KNJQmgHgZrejHFBm1CE0QWKDBvW7BC9WmCTL23bPxbPBRJNMWYmJkpxw4X8Z
/Qlgf6GkYrJLW6yGo8zA3jmxCsTtqzvifWNsctYEsI+HQqMu/2OEHKeV8of4O8Vf2PzB+oP3Dc3k
gAkZpPPFtqeh+wc+IF2RXbYTWlT5GADF+LmS2ktYaIFVkoTtl8uHjCqMuSNBOTIVNfnhGPTpbFlq
atsI4KZu8bVApgdqZxz60W5U3yx916brvXc2NQqMLUhY4lCT9LNkWrDygUlaI+IqOheLuyISjYnM
EDB+UW03T3PpeX+qQgWi8y1VOkDsdOVszT1Nmp+zj7BKdEbPZnqdpa/ULjnZOgUwaeQUWxr9D8h2
RYb3HxK/rFfNN11kwD1/ScV6AxwQDrb50smjozGuCDXG9qfLzra/8+OKD+tvKKH8FHMZuGgzOgis
wdSYGhrmtc7nHHXwmUsoBbkQZKZ+vruouYFFM2Z+WG+Fo6/m+u0oJljtltO0+AfYdxnXgCVza6Ct
NmtlNsq7FpCMhbAgtFiS5jgyxcuim8Eu/y4p/RDLWGn9NNPZAbzgELwDFsdWhVM6J3JuoYpYuIp0
LivUr0hbiTy2DhB9LbU2R7pmUpkIhldkoKwKZmvdYrzAbai1jvQIo9R4wFGqIEDtlt2+FZwALuRi
HGIWRPWxUYgxznyrsxu4l0YsZzBeSkoucdOi3EtSW0dpVH7b/axIpWQFZqJN/mHMV49GW0DE3A2z
/RghpbtZJ4y/REK+ePjxZnXMxmO7fITfsxSlGijPvtMlsd14R6WJjq7u5HI7KKXZRy+7UIne/dVQ
9lbjWLYKZLt6ltaZuRAFC12PkHnV+mCK6HNpdK5CLJI66ZZY9vDOUdxkwL4BCTvo94gD6h/hJ4sh
ndZN0VwuRQWRaIuaZTICnSJaXP4Ranv2xXimbOUjxAgoSGKClfkdlcvbSg8skAKxyvoqK+qxZPtU
48IByzMA2ySPC0tHPReoXFK237/YcR4unfsSBl3EVjMRbh+3BZuGNgmlaB1OvhpD7GtM2/smhVeU
W2Q9dgPqhqUlC6JZzrWtJxQE49R/BeSC1Ol2MlfBtp/8Y6Yk+e5aeCNi3cl4jTqitNplM+7KXueS
oo42+q72EZDxmiTiQxRVFOC3sY4aNsBp09j2Qk40Q4P36cfnJ32xRRF4uB2S64XrVgjvvNIBcRP9
KiFeiRUceXq7KaF5AYEIWNK6V7tDD5EbeYBVCCJYH8nG4IPfhAg85OZOlYI/gZH10FteAJnN8wef
o0uuul6cjM0xRz0luMK3K4kX+Kphxjxk1pGiaWUePqVfET03IexRIWn6UVEOsxDUNoiOvK1Ex05J
/I9cJ8t0vr0UMwsfg5IZzZmoQ+nlkmDmtDah1j5x3hwMQ7Eqp3Hu1gwb2Ff3mHrSuiI+CzXrnA+m
sRC2WEHnGh3+z08vrTREVuhqdQSDWRwbGw0AVLCYDkL5
`protect end_protected
