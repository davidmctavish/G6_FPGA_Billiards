`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
h/0OcFzs5jomMn1+7BRybJ05ZCk25BtVaYDllF6RHTqh2rIQ/jWwCseJOtgmLOxGBX1k5mlgnBHx
Kunug4Vw1Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nIq7qPYLjiL3iR7XYRtQduFLRTKHfUQcPLX/kVdSO9tziYivE4ml4Q1wjdKQrdYvTUMIjJ+S7JX4
9yfyUfKWzu7zp/Z+rayYJk6/OQmVIw8nqSjg+7cfeoNSKq5T2MVfIC5JrJ5H8ZhVjE/7cuGfyoM6
7SYV4+sjUe+LEv4wcEI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
g293fy/pSp53ZPe5szWBxiVuZzJa9O2LSjLHYbfagjMSFSU8MetCjA97zIHCP/i4PC2saQaOO3zw
GtR8KXV54V6dq6qXiWsb3rDoUKT1hm9TZ8cICcsLi8f5zo/3TC9hsMOGzo4ot9LAflL0aAETfgW3
ksrhTLgRkOmz25Urb9PwHEORfn6sqmb1hw8ves7CpSud50KhBUTfa9eBjBOr8M3XehKgzb82oJiM
63kkZpkTpuHOW/6FF/IOeTy1mYd9TNwhYllMS4SsZEgBpvUSjbSQKCYLJ0FIZvWSjLBVz8nDDMmC
njJZtQ4T2djm9izhItloJ8n+0H+x1ezk7n9rfw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WLcBA29ILP963syrd2+3CQFcQNx+hLd8Y1eM7lwM49rNqWX5mN5RovD1SG5MLK1steIbBh0Lu+Zw
2l18R/HMuu66vER/A4xaM8kph8/L8e/Pi6XKtLxFiCj541eJqCqdFQ4nQBjzN8DYtg6IN84a7N21
/uXQ21F161k2xB60id4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IfJigQ7bi9U0dOe6+t2QLNghmTcLsB8KBMQVciZUlGOtDxp+vX6dWKEXv3PGYgcDYxpryoSr3sUr
4TiVf+7zQ6hOINcs4ZRPHlhq+Sl1+DZU1rI+rcfXI67HlaFH6fpe2HWrGUynTDOxFeSX4s95Ajiu
PXidxQDi2REC4o1WSrCX383I0e/dVQC1KMGb3smuGkFiDsfERoWXD3sA2tdJxIsMWUSGmhh7Xz79
ENLycD67GYcwUA20FZTF1sDwFooZ31ZzZa0oH40xq27TX2D3/odzse7YrcVMc/KPYteLpFfBDiQ0
B6vunV2oxiWO4NVc6C9jdy38re9gFCepP7KXEA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12576)
`protect data_block
bSKVdq4NmBSXrjR+g3lITJJvy9AGSTUFQG32F44R2jGTHWIXhz71HIUimcOQo2xL/luUW+SWFO80
tS4Si+NP2jIAuppM8v/oQQWInXdFd2uAio/2OO9NqqfNWjAT4NjmPc3Irts2QhAT0H1YUR0mAJcb
pB144ilLLGo/eKPxgu4zDVIEGM7hP9RF/HxDucWzZ6jYLOfzX96y9Wz6ht+l2w+3sAdeMZlTJKOn
mX939KCeoyOcOBm2r+6ABPUVxST4WhSJAowaNfTtKJRFNOMVDuLcGDBiX2g12Hdm97M1fAYDxgHL
hq00Q8WaiLh+wuGX4qzYeQDhBv75BFyIY5OX2tWPpuwjh8+QOG74gUhoPPfRLX+ssj6Uyo5m5jcP
ufN12Rzf0jzJYBPKXlj9PQyyY6MB6OEaNLikzMCaFkZjJZ5FpUaAEkuOFHgNX00Qnfz6QJuiGqp6
UapcP1VQ5aQD7czOLgKNPbd0nOoJ1kyMS07DQBSDY7ofEPYufu0kaU2t7/I7vJ582wcQMZZQU8dO
cfe0DrbxlNDj/jOJYDm8neqMPIUdyd15vHGYVVKX0SqBrcHHgEVKE4oblwE7KV7Bg3dSwWTLojrO
NWWA1m4JCO8WBrLICieEYDX/RUYOzE8+/sWQV2zCHarPBK1zNZfJA1psAxPLmVjhmU/6bELcVQQE
Dwodkob3EF/vL3/YTuNigCVHX/nALQev/KAfU/HoMDZpM8pUwNIOcVxFz5xwNsKh/dzsecujakxv
VYcEGlOZNUC8cQJRij6TR3ZXugTZUodA1T3ad65769cWwSPGl1vg2JErLSNq/n5lO1JFkdtqyd5b
kqA6wmYq6ew6AGH/J8EyX2sUOBkXl1SbQMc27kxcBX2zry0Eta+eFthfneCEMchU63EBNFq6UTMb
OcwoikjoXkkagU1P0qYBYdTAmgNdt7OSNpKVesVFruu8doxEYFjmSt0Fxz4aTKhDDuGS1aibQLoo
UHMdDmW9qAIPn6UeOkef/GWxPRJwGmTHDs6jKRbQIy9E92NYMwrUZdxiv8I6WGCSBRsJGD8vdAlG
utjDVtWgCz/Xw0htdz4d+tMru4rQuO0y34ohimyVU6Zhva5OB1OfN8qrhapK8ciLU/jnbetWH3nC
gQlX6P0yXsUB5WYB2MHYw6A2lFerTSjiuTHjb85/YhoOrff6LGqnrizTqxiYbddiu/MqScwGvttH
NsKXWo/CFPvIzaJ1NecoCBiVkEJa+vjRtREE4RSYRqUR7k06ZqnOSdEbRSPQKoke0YbM29x3iXj+
EPb7MvrsWu9mcm6SSxB2Tp+8unMaTvqerlQw/JQTvhQG8M5j/O8VhrI34i+JfXce4LFXrN2ybZrd
gMCWe5CbS463gJ/sT5W13a3FcdW2Qfl8Lla+xkGSr+iWXSmqDlaH2aNYbZpu4naUFX6Xr7NWwltL
hqqK0Q63uST4lWeqlrIRM5Lg0mMZwPIORKmg9AjjjVTozuCYhBrIYuLwcJebXUQNYLSnx7Rm/azH
B1WDJYtEG1VNdm2ZEZIp4tor0ivon4Y79XEEuvA/6UoLmjt9Vxm3uznPd6lbx9yswtkQN4GdevCW
weoyV0w0HH7a8E0ofYj3pDjXjTTauIxFPOk4L6+5DwKq6NMpuP2AYYJ9RYrUWPQzfAXWcg/wmNS1
iythArf4pgLovZ8yhNxbB0dzxOVdbsSSpDLdRoGTaIzdiMpkz53yc1uPgxeGx8exSAvhqhGdFHR3
2KgQiJWgSsJNXibBV03iBcU9C2SSL4F+Se6b8uaRCxZVTKUTmCUGvuTNIub+t4wiAnVnTHxpvnnd
v7ygyRIcVSFsAAfBx+UcX1S0HrvOEIrox2dfQXbZXgYiowMmtOTj9w30ypWZHlNaP9+lWyEYpBZx
LS1ODKbc02BeY8z1RDVk6/3Ck/5GTBYEPxkrBfxUMk5tOIQBhhWgDRSh8QhF92aRVLHCl3QLm97J
PU7Xxi0S/ATk4hgAmrCFrdwzBHmUrZQt94ZugiCF0JHSA/+GqFu93bvVZM2+vDYHRePH8k4nSMEZ
8cYDJbv14YftmnJaEbGIM7FojDae3msu8RcpFPZrQz+Q8/rZ9/XQiapzgxZGRtbEsSAZgS/XvEOg
iY+sp+WPMH8qgtrmOPgtN7e9Zf0tzAbYbJkkr8EqASPVCBjjhRIfDZFsMwkqwqeo1bwF8vlSVSDj
lGzQxohuDn0shngrld//V3AmPI/cX44ITNqDs3mXHDJKMLPuhmVXTxd/0J8oYAYHLHwESDJruTCy
11rb6UkmhvsyH12J6NZvamP6zKHJriVB297oJk8KPUbPGwIPClfd7uLLHT7P+Z/KM+7ciZcEHFuQ
q8ZIX/Z0jsE2dawju7y52TbnQH1MVOjt8TifUZksw3zCfU1jX3OKEBLSZdGlkXynUSbUSb3dqwze
+tVzlTXMIfeJKuxFFlpy/7A2xZmvndlJabwGYX1sRrixpjf0ws1/eLthcQykmDe7wYrjQlUuYBww
j5cbEqSRlYYLIXF4nV82VNSkKJKNQqqJKSeBFDNJUR0CvE5Y9UNHsqXSnGfN1Vrj583wRUVJjm1u
9kyGJ08judm07lzkSf9VhIQWBU2G8Ae4fQnSwjjx8n6/YOWeZe4IaCWnH3PKIhayJjph1UBFr3rB
FkyYlHLN6fkhRk6Y74OubTMRlDgF+nh6bfPP3I9WSzyfn3nCXyo+5iImzLkDBFKEyMOcJYLGS8qZ
0k3LfdZSlgZDiDYK0g9pgkZCj+4XmgFrUf3ZpzToUazCYszu4aB7G7HaIQw1sFYsAuSCDb4UlNR7
pWKBkOBjZI0THYKV5cx83vYmW+fbXoPPz6QEgzylOMVeupHUT0NadMrluHdXp1M+wzQvhEOBVNJK
hzgIhc9+6WY8IiazjmcJZyaKdMI687zXG3bbO38tEwEsYN2JiaZwaSLZj1mTcU21Gj7IQX3Do1RC
AjcZijM+Lvd0E9S7EIlHfACAcJ9zumbqMj2uexLruxSPZfOi7iGHySb3xxuIK15i3/iFKKEUwhli
XSOTJIOnllCzPAm7JkFIZbubZVIFDE5WajYI+Qo04INwB3m9JaCOVzg8jKAwsYGh2MIvmOV1lKw4
d6l+WIIA2B7lZPPyI+blORZH7f39q3css3pAMbVBKJbJny3fMYX2z4NiMcQCJLyEAqi+12LTCzCl
3iWMEjD5RikkBVbP2iXlY8J/GNUS4OzFU/4oTj8l67F+YCA/EDG56JXv7WkPNjYuuFFZvFql1O8+
ZmN+zG2n944Oa0qeOW53eiSKc+U1MWTlufsgB47VV9TslcepJ6VlxANrWrTB5WYm5LzkMNaF2uLz
Ia0i7GNsFhfoFa+Mu5lwsUD2ahKacXho1uIqouoPy7ie41pq6SvNq2sl+bx4rvlJWDsVa3fRTyJk
LB73rZ/XEqGw2U+voCPL+B2QbLbUFkFUrc2XEBRzYpOfN5JzzrMLhYA97yIG2GEcmP9KT4zOli4W
Qtpzy8WFs/ISmPNBsE8xxrV2+4WdB8b5WbStDiz+E9VKNIKiSl3pa+oV62LzbFV3uWJPTqhmKvf/
1kgdj23nW/JKg0IWpKZ/wwWZpmXGPfN2VJUxshJQMnAkkdr9IBOTRvPonogNTBinSY3GlzIpTf3q
jF/xc/byhtpxrC2GTbPlYu647B0QBZZYq8QHS/8ekXrSwvvovp0wtrezr0kFjRU9ZZ+xdl+3Jwru
u6ZNrPSwuGKscFMczpAlAdEDbNvei0wXYpV+UX9YrKfHnyTcV5TqOauuWz4v5tsqL1g+fTxUScB5
/TXD3BodVOSUHHhcy2HItfCW1vBPJ4sNFHd8pTOTM6sCIEGro9XCTSokOVg3Ynn2fxiu1p+ritD2
oqrn9SlI63qDae4/ZV+Je5zaMrgH4gPcGooqVKHX5aQYTR8whxHUcrVaRGeokXtg1v3mebbrYuAZ
/uqVDe6Ep68vv34cqnMoz9T7QfxC4um4Lg2PYa8Px1u7BLxqQrtkbyOHeeeZ5kaulUYqtu6xDKqI
VecTzGw+X6W3evHZWXFYAo6vKMJnzvSvEb287CNO4ADyMUcl4N14Pb/TXf8wAGr3n/6yYQ8E4am2
ymZfjybBnE0nUsTd2AU+B7lk5pP2tFC4T2JmM/IyPzf5ZCTrzi/cM/AxJehEJhMZE0m97APa83xK
++Hvb3R5LaakrhFJHdrNDK0srnSAaSVeR92kL4PYeVIyRz/A8IBujiCzgpA5mfmmMJ1yVFKR/ivz
n2vAAtR3X3sROlqx/Qtr5acsYkXTHy1R5vWR255KvOYt/5Z1KArkmcT9Xn5FEXg0dX5Ram3wU5c0
noWInvc0B1LbpozVbgEJc2GjdOn9o968d1qgea1oOvgHlB+J+EHPZtncLT9j38P7eZZikCGg+D9u
1WutsV9i2+dPIIeYtcU86QAlx/XT6S9P9Aljbk4teiyAOs/oE7GQwsKkUEVDVK7doJwv/TqKf378
Kiy4IjgiA31QC55wygKpmO0JMXnp0gkAEAHjzzIsh3la7AW0yLupAmPUb7PX+pF8kngKQzrYoQK0
xxYe2gykislzyjVEqR338yxsosJQDM8hWEjpkI4kRBHA4vJx1i25kTea8r8ahMM6E/Sn6My0VYas
C56xlyCWBA0Wc+7hQF9AGYexXGvA74Q2j+QPKE57dSyXn35Srst1qtvHB9a4x/W5yrWVi5wNvsFM
ovbaGLHWblYu5vSqPZ9+DFGf/n8Zg8X2nCydbm7uD+qJ5nkhRQrEwGnUn5cr5Tm1xn3oNOpPzrV5
3v4QdhCilFu6XlBAJYfdrRFG4U+NkwSBj1R89ZDWGuyqFgX32MSQeihLHcSISmR9cBOBtAfNRDtb
7iu5LJy8IreMjzf1ZdZeC62lTPArO8O0YFfduz3AmdcoH591eHlZVsgWM1HIAFg2eFC4OIknD0M9
ce3Q5V4oyWlCXexTCXS1w5r2cXVzrMWqbinAJH2o6sKNrrI0FSaYGfAvv+aDYpJgB/6ZVMAs4jQM
S41/k5bWs1yh7+nV3mg5gF6WOYy8V1rX4w/PMLl794xhvDcnBmhyCJouxZkTIO7oeVN0awc7ds0M
GpwuUr4AykmMY7Rwnjoq60ooG/zMi2ObioARUXDy/veDPpznF4F1j7i7GQUfPiHk424QLq29hdPZ
08LMpMedKfVfjaLgGWuK2c2T0cdVDsfNxODjiWS6K57duxGVd/bs1NBk4/Ap42rmxxwx7bVzYgo6
DSYx4QNBbYF0CxK38P7DdEk61hkioSjQSkGiUJ6H5azyh1omNfwPsq3qKWFZAFKR+VM3KnuYYQkJ
4tw9TGaPPJOrA7RTLw0NyrVJkHzZov5ubgKw6wM4cYeTmEvPAa7iuEAwTdSUhOFBiQpPr4q7I37c
3Myr34BlyJF1tF2TeyODSIsUpt2rmbrD+dZKnlHovO3p32djr7jjIRKs7l9PpqIunfyvFg0V+gs9
FJDfM7Zm7MtZT7E6LmkWSqe9ygIohH7KSsAO6K5RFU9RAxOlaGdyC5qfAG6jpa9peTZ6onUnTBsQ
HuWLTQGxu7K44iCQhhA/bX3o4w1IykiR5q1igBrSi+K6SzvCZ7pL+HHnila2FgkU7p2YC75I4ndl
GMoBcFuECs0JZvYWWYVQupV8DxzWaDqx1+qRo2Z0eUiyI6dkB1vxFmvaflug1e/4JGMbwjq5CAVZ
3NbmmTuGra8fPdWqHA7dxVEHB1hVXRDKj4tx1hAoWpU8rTU/d2w4x27J8AIVBkITvAyBFaWeYboK
hPdC24FlQEOhtPTIVYOwenFQ3hIWnkbor+RtMDXvtti3Ckg6KixZ5AXc5Jco4X/t4icRiv2JN9G7
AYQ8/48ixX+yt2lRQQFN/9N8GR4Mx2v+oH3nxRREAaPCUf2xLdi5myXaQgfBKIB80+X1Yz65stEq
dgc8CCUOoI0n1j2P5pvVwlVq2Ew7NY9kfF7c+0dNlOnwh8/S/VPGs84TdvJUTsQtbdUl8uXbG6Bx
XIQ3LvoLVAJy5WyI6r98JHXR4rD3VpGGJacTTGgfo7V75WP10oE5A6hwLxP0oCoSYXVhiEQBoiP7
8ZmzEd1JOIq4ZPqAoNzyxa2F/GxNUZqFrtpBaWmOXrEi16MV0eMXI5tgS01F8YCLbargjYCoL28O
dEArqF+DJAX4MJ+y1OE90BSBOr8TSdFXb+Iltc+Ppuv64NbNNg3/+CW8d5Dq1rZ4Trcu8BHJb1sW
g3dsq6kxypOawBEXNU5e1xvGUFcrg8aN4iXYJpAtYtw+h10QDgp6Zd+DYHtPYMSPkp/utMg2rVfK
qPhCAt/OhenknjdDykPvXhaFavVIOIMDOPGBU97IpHAPq8tCzTOuI1uZsL/D8tWjPJZP4awqFj9M
WOKpGLpMNQRBzra4oG/Dt9RVYeXDzEuEXyGnDhdOmvEr5Y5bLSx0wkY536/HF/2nyDBB2Wthq+vZ
cn3rBjubSiLMxKsL6oYhjsMUXfi7rGpj5w5QB5R/H6kQolj9OyeIBhHqfHa3/Fj7AI4geHnQOCmz
6AVJUEnXGfC6xsQUctQVNr8TlJQ60K6S5Wur6Z1KRsHJrqP+rL3+qTvlq96XGjuErm7XMdcNAqBC
UNzjS+gh+A3dboQDRxpjLdhVt0mvbJUlCOxR5njkXkmvN6j+pL0sx26IcPlz239vgNedNmAJutE8
IhDnczGTliQN+eV9DQHqE6XAiUJUvqUSonN05nblpJn2JOk+C30amOScO0otIQQ34ObYASsD9J2X
NgCiVpksGJ4tcrTOcpsSlrMdCjUxipZD8mok1eF6/Cr6suIHSX6juiYhqIuTQN+SHFVFZc1abhjF
LfDP6RfLeCHbjv5ZcLk39A1YW5i7Vi0mWAtQ8Q9rGpL6jE5LDR717ta7X380G6DfpaUf98lmQ1cT
ZHkIpECjKoHATlnlum9eZ6nQmhSOpyoSxEBu6VM8rHrfwFquEI0KDhCXp7tyMKihEAcVVmPGxXrH
lm/Ls0oRAQhf8Q/uqi203sNh1Ce3jzzO+78LrexnDHy4vwbvn4mGEJcow7ZOgnsx+077AqJ9oXPl
bMtl6VWSTk6aSDf8kTE8vD3bZ/rBbyv4fZCUsNNguLleRuCRUbGdO11ruYSY7mx2fUzUz8d65Ora
MghArv2GqSyAjI4jxN55gMxn7hgrp/9K0UjCS7Cg/TMJok+ZK/gnJlVUUPYFhY0tY06v03c/520A
KQJwhHkZSYRESHK33bqunkf11+2w9C7ri5+vv9qA7Uqo/BcQ2UhSQsktLb/cufkNdKYQNXnsLkiS
aB9sU86G1YkM6m4VJzkkzdtr09/NecGpQEGupNpE/d9aLOFTdpQbTm3KjZY00yMDc//THZtX5EFe
r6xXFpgml9/EXAiHPfQexoWjJB16GbAFHILooKcfG6j8bVDDfrP5Y+NMldAhODdP1/EPXoP//Mgw
tFfATfGbbUhjOoKKMh5GXm7EkhVRyPHGQRtbONbQMfVYp9sQvCv6gfKE/iAvBT2DswFtBlOo4Vuh
+Sw0gv4qUF+5fMIDeJYGqqsgXKN5/FUiOYeDqvUPnW2RGBMaMRRDrWk66DqJ+bvDtGLwPmOTHwwc
nsfjzygUEk5cicE61kQUHtrfAkSrngfRgcKKy1+mMSZfZqyXaIaPMh/WqJRxT/Q7ot6hog5Kh3lz
0vyimg0VvKNCLPc4Wx/5335LHLdNVW8rOg2s1MM68RIgp+yiO5MMhW+i/1iKBt5Vw6ndK4J85ISt
9FJwhW4nHPqPy81MbyR52QORMl1usyq1d4tKhrY/635sGvpfBqG60asZ85AEUEfz4zsOcDAaQPM3
GuFMDk8NAUez6V9V3J0U9rPPpuF88iz9MDoboetj0kkpzq13iLai85KnnCIx/LqIpPDrLZaFMjkY
GHMUeJjCJteJo/PvSLaOU+f5mgzLMjaqW3f9FImk9IfJvcbeafzn3FG+49Jsnoe0Mo2413GjcBfZ
iTH6ReAYVH6aUurk15+i87AabtYBnCgb1gsieJP5WHGZzNlQdgHQhqN3SlTiEvZU1mf69XKSatEH
ems80LwoRqvau6/3W3RRsS/G1rEMAX2E0b85raRQDG6X6bzID7mkMfFIAY7Pr6yVNFd+GS6AyXWF
PKEPNo4C3nLSFvIK0oohmdUn/LltYhHbnTnBSJZFnpdHDS5hErfqVGftQbRI1WxiWopk/jH+Kh/v
96SuVdWoqe3ZztKsiAmTl6UarFp9x0tqQbyKg+IZ8tXM312+V67gfVzWEaPqkok+/MRXiVW7Uoh0
Cav2f66UteIuM7MHSOyGtmAQwsqq/c018hUVOOccYusO6fi3SkmcPvsMUS3YUQ1XSIsKVs8fuSzb
teI1hXUWRXQ2B9W+rVS3li1T17zQb0kHC5sh4FYLMlfY3GF83OdYW797EVoVegeQElnCY8Z/UoTj
Pu53xIsfXzo653yJuqKjC5BBZ70Tq536t0rpda97acCBqosnGWsKUk/4mJY5QbHPOGnNdMx+N/Mh
tPuitNnKpUTN0q3OOvipcyZ4ek0mYmzy1cdddqW5bPSj7dpGSbvJsGXFntma0m4IKTKtDze6yZJQ
46EB7oha+1xDpff5ZjYHS71JVPSdokctBECgwEObv1m9uZGtBHC8Q3sNCjCZEtTqxy7yXWuwS8tn
WUL7pPdzEu6ObmQMkgCpIYHMVcwLG4KyYBGqJTnlGzjN5wCZr8bHzj1inumDSuYtSRSQ7yiZ7727
A0XQUVLqhusbx9zppiGUb+wXiFuKiOwS65ylzZhs2j7ShXfLc/MptrQjBgfa8ARCsuuB2MpkIcVz
gsH9H6tFJR/fnMfJcpXQdxX/PpgdW35ekz4umB3U5irpSxb7lqkYzslD8OlvFov/MzIc809//sIl
w5YjwvAnTb/TU2r/Y//O0L1P2nitfstgwRRyz6fd+OrRFQlFmni/KtDKyc/llhnAT2LMYADP+AZy
/0WZ4idfATqMA5OmMwqSw4DupUp7p+di9zE7Z95xu5aOJNbx8RJMNKTsFFJ923vfd1tZM/LDo0gV
89P5hfMRXje4++Yj8ReCiTQCiCCyywWxmnhA5MS4IOQbzVXCW0LXNXGny29WFEq6gd8LgtYuqsTp
EdRLYkidM2ZjiWpa+w3N2mTOu82Iy62xpedMyEWNklxVlD9ytmZ3cPWPjHLTL3GgArAMnqYHDxOI
v5vjtjb+BlyYEoJNaHi1gTLbif5AE2i2W5/XCSFhx6cqfOK2kRCUBPM3JlfOrlb4/eZXCsYACaS7
H9pKW/3sGTquY5DxcMKDMk+lpV8JFDas39mc4LODGRZTb7EstHuiEiJsfaF3sjE5juSUn6/koWum
WXnS+9xf7aD4OKfwlO2X775lPgZaG4eQ3n/FsyjME9boGhOZsXWVmDBSDnQ1ce4YBzLpvu4nwVkp
juqcQ5WAPq+/ND8e8zF4OyQJDrUnJFfW1sOioC0sowloEAKCR83s7MrAxmhf0HCtcBMxYTAdOTdU
RQ8kJjjolMLJsqHOxtettp7EBhi6i6YRmpqNi+Rh2pJ4Zx7Z8tr1qz5D/nYHYT7k45nlx01ur+14
RPbq3AQsjLuE4pswVLqeZKPtErQvkHmWeiHwwBQfipZ5CcQ2CMux+WYbMOmI26ICUHGTirlFm8Hy
hpp+hX2jVSCyLlHDNWfCZ0hDa04Kg84wnHP6DkfHkhYvlNtwMkTpzG5CFu4gHtn2mT+8g547k49T
SRHGcJCYDEIB37gX0zxLhbaDHOebBnODoj71g9NiEiKkBfHTahBH9HQzHAW+nqNizXhsMYQWSFN9
PEBdHwX+SrWLEcqEozv3pdzcVf+w/GJdYliqWPF0Rs4UA140gb7g1PzEILBhRxeaO9F7CK+xV/kk
FHz35ZDZbmixlAUViNs0u0rylW6/n9YdlzvMPn9oxeyOP+V8Ai+DytBnM9NRkBwIIBYI597SKB3B
6cQdibxH/+nYO9MZLmvfoexSgsjWTwrevzmzlbZrQ860fmTybXMhsWvHsYx9iuJ+aJ7360MKSBX0
qA5euNZV+iXztrRyigCSNOwo9K5ePFuJQLm86lTjOLFU+RY65nh+WGS8WSAg95oNlrlNV6AA+Ant
iLRVMzHvRO+KsYhpgvbNN5gJFPbp/NKl2OttFWj1ZLYpbJDXWWuYQu3TEHn0RVtN8S2jOxdX/UXZ
E0hfLkMBzDOfQvhiCmQ0Tsg8wDKYbHodGHk4N/8cR/8cmcQvFa85WzUUm9fuTzHymg+3mjJVW8RQ
2MvJmYXcAzy0kKQMHNL342BxqVc11jcLJURfVWTuAb1idVPyYb41ICqpRyPPk+kIA2UxXGiOFxZz
Am8CcTmvwyj+0SeruWDl0HcV4WFsiWz42JANDfLhJ+cFFTvJTDdxX9t2BE+yZgYw0oyoltisb+9Y
BtfkX+bVL3qxyJoJyinur2Zq/zdCYEGgkBzaqEycyvZYJcpuHwj6K7qh1nliBuSnfEZ7phe05Fth
ZqSP0Zo7LYlBeZEr1+GKOhhllYhBglsslb7YnvCEBfwFfReeL7/EAT6A6pul0tR1KzswhHl7eEGr
a7wFCMByXUGdvY0JXaY+jFW+nuYJpgaiee6guu3JdcHbPDBjFpKeGse64iw7kBzxl63vwfk2ug8M
BwtlL+vI8c7htQ041UXpiqu8IasJ1BCMkkKQGRk11UCU3KzGRnHUIjuMKa3UBysgX+7WNq/Rwg+t
YnFOkBOqoAYAC5ESK5dbEDlWOK+xLA2EPIgtcSOrub+S1zPdDj4ROT+mssr9bWY5Vhh9TImkPixH
JvDYDF/GSQ467rQzUUQuJp/4yZFx318UROTZEG2f4BGnNoPKlZqtccm7W6f9TStAC9HsXkGYBgVI
kPcGhFjTgweC5HzLZKT7NLcyWSip5uPRQrkZWdRltidQOPPOy25k5pGGP2Py4Hcvg1yf8VgvegO6
0vJ8d2eK7TwnYTRt3GeTGiBjQ30ZiEpwu1qgtv40yKfKaYI9KD+YmDD7qdurNuzhaiXAog8t/pfb
zXwHb1N70IxAmLDFRMCNjbTS7Kv9PdwXLU8wV94lqMDJLEoIAkI8A/u7xPq5aXAkLXfG6LONf70d
XF8EsFy5gYjCP/T6hPE7dhZ972UlfH6ufjBWlQZ31zwiayZOxBbGV98GLN1Ecs+/j9fcSTOMwIaB
lr2BuZ0jEsDrPPpQGC2sCMDeIUfumrVdYdII9id5JhhNOjdHKh4pAVdBcBfsXJUorBoVD9cb/wwG
hKAi/M+TRqO+FE/+j/AQCGdLWKW04XrEsE0lmM112xjglzIUCzL57rFlRMwy6+o1p4RAorsbjQ+1
61kfxtLBDaHfFGTyK3dpP2wJsYQuV+naCWHhda9SO9IhGcfHMkun8pHN+3vjQt9sv9OE0g4XXFfE
QRPJSFlWXrtgScMq9DMCuidnSeBElaFyHKEHNCHZhrbNoR6mhujTpK4XHl16dmlLCNoBzuyhLtTN
FU23z73EIS96XAcuOFDQXpa5IXPRnKuFVgHqMOEwiW3MLwtNxHmkALiL3Jx9ixw3QLFm3gkbOFLv
q8ED/RT3bTBbr1q2/r8ms2vgoVStei4aaz7nK6QE+w+nbxlD0toQHxH69ypKYGko6P54wm58sHP0
tQJOUkOe/nbbCyCkV9HAc8BWUXMG5r8tJQrXXc0lxOKktTrDYxXk9FFaEqqVnjEJuP7JPABDUGzU
U1EKrf2vdEEnJvE2cTwlLM/dXAXZfBe++I6XYCf65zJOtUW0vYx+SZ67au7eoz271N8VL3+WJBS2
lEdiR3CPVpIuN4WQRkYkWY2eWir7PeqPt9NWfTchlEK9XjK11KEhtLHi1bdYb7bitynYAFh8vqXl
EIsYv8+3WCDtesAAwLKAtyESipkPAIEc1qPLU7fkbrc95Ybjy7DwH1zE1I26QeE+o9TzsFrNYNWX
obdJLZZsxJ1Vmj/miOcotZoPbXD1J5g7iOp29mbS3gShg3/l63dxVqosFkXd7yGNTmr1EhDOGzrZ
nPhGxXFXvhbgM5psmobdEDMEiTlkQ9XaJ4H2h9ZUPZ8K+ryX0sX6icI197QGLkUxMhi1XSuuiUN/
aNVOOM0I5ETyGOf159HNOKjJBHb43cu+vC+FqoVTCrzmoOPXbu9TOUDMqAcXeWN00u0y2QtA8aEW
alyOqhUsb7oIvTIt3E7CZKIAff2HaU3TDHz761Y7AGyKnI+l0I80dTlZH2VMiJSq6s/Bwm2S+Iw0
2w1BnqnoG4uI0MVChyBKupxUCJbfnnifTfAT8Zyc4ztJj5NHdJs20UuI5G2eRNTCP0s3fWE41j4L
eFOKyeD8l0UmX78i1m0lctSv9AAhtYEA+Kuim0g1VkaJmwA0SDK49dDGU3ycni4BQLyBSQUE3+QN
vXg+fv+tzb8SUThJTJpeHB8Ck+rigky/vRHMzNyvQDqTUSiu9xKTdUrTeFV+yKyoXLsbfnLhN1yq
w9cxWK//LosRMIS03aYeZ0W2uJGv/qVEmgLRu4fs7Oyhu3+PXjEISzXnpfmjr2uNtM5UGxvruLum
4ZyFVOvCtk0q6rwC6VnXqbh+UHaJZfNVBzoxGC4ju/adrbEwjwqpYwm1zBb75QamW29o0H/rVF/A
T+748Y34eIetdwHqHqQnPGeeBV3uqwu0umS5Q/3ET02hBgaJN4u82iHsEnKVHc0Dd/1LhCRir//G
bgNac4gIZXJ5kH+WGXa0+LR9UtVQzq5K8emX/wmuz/QS2p7l5vCJBDiGKdFjRDGgYxEcqPpphwEp
K+iz5jseKhoGn5X/UtRe0SxDjA2oQ7ec69Yec2BgtbmrrfBIuEyfBl6PM3ZK5oaJXFVbTEnrkO2B
coea1ZyB9kCRmVblzcOuEDGm8iukem8xxsNZuUtp7sKUn4Y6e2cOzEyPYtR1sHuzY5rLrvIBtAP+
CTqlBl3v+oW5W8Tc9mQiFCqX5sdPDOIifqjSti7mZwxX84mTJgx4DlrH3k8QLjAZID8cn4+WXsMa
sSm4FcvdEjBhG/Y9b16vlmJgOdkSdCTiMe9hYgYSi33ZHj0O0Z9P3OA4cYZrBpMV56RGdxktAHgA
JDv2Odrj5y9MKEvrrqnAo1HDfI6LAIX5GYJNF7JL4i6ns0ABgvRC6zP1hwjLwT5TgwN8yCOHyPEC
PoZCMXabeuOzgvfLOKzWt8kMhrgI9nRjjR3BH44m225H8LHDHtvMYQdZU/zux1FJkqt15aMIbY4W
PsVNH7PUIIseLk22nquBlSW4gQ1hVZq/3v8YBXzfOlLEcwWoi4Py7G9Dgh3eeOEZ00ZRQMOX1E7V
00Kz4vlCAreovuKnA382CiG9C5BdEbcJl55l9CkgiNKcuL93IGZ89sCybYao0F2JJIqxUJl6g7lV
ZwCLJcC+H/yBudCKqCfJFEe7KXi+TYUlSlYiROiG2P5AOFAFsuI3ILkYBsM45lRB/XnKZ9p73uSy
XJC0G7fOXslpGPAi28PrwyOXv5zNO4Q6yFJ+Q9JBm5HSt9e3ezor7wC1KlU/d6bKz+MRpwDocWFF
PAb5pVgS22aPxZxX5d4KfshuTVqECyWmbL3dhAoQ14pwjmPDeL4h62PCl6Ny1aSYp+p09qo5uxMY
gVvt5u+AUHIVJiWGzgq43/J2asbxPC4K24ClRq+B5YVYsX7mlgAlUKxQLAlXPFwRdW7UDow40/Ex
Lc8Uw7Hes4D5YbeZZRFko5rF6J7GRt/8Y1BSFbn0jT4VH45hy/1cO45Rh+iwDFRzVaaZcm1uvDHu
u0ECWgieNKC7jjLIIaudW3SMU5KazhPR/llHLoXfVM+mz6zCD1FqKqkxor402hOgRH+mvo7xPdQT
SXlV8Q1ASN7K93or8Ruu+YoKkH5YM14sJbxSTZO+lheoKvNJLip/C4pqul4GLZ/AdRXHdb7D9HJn
oX6+OoXHbiSSsZ/2h1NltSoUd4jfe5cO9t0u9kp1FmhHiJWxExGvWKUfxAHko7VXVDqnAkFykSpT
9lmzYSdfT15ZoH/gwcUSou59V2ttGhuDDtzjN/8arrmcGcaBI+fAkwn/h7SEX9p828xk8BsNyywx
IhnRdOYJ1gom7zyj9ROYo1VAM6penwHN929kKppTBEplsK8U5twIV5ixnicHwtS0vKsHxSB6L0KY
vRvJ4PB7OSJmX1sIQnRRWIdouZB6lyuEOKuAMbCxy5051u8coIOFAA0aVdEb+OgLpprLAgLjx0xb
hRQuU4nVNeJsDWPRiFG0HWraz1faUfcJ7iGB2bFBUdE6mJySSkoUGzvGKrwLkMsnPcCym352g+R0
i1a+SAK17TSWh7Szu/XYAhOB1Sht9OEFCp5ZBWETKS3jEchU8YtcWXbPtPbn5jZCHYCPbbn4TyIc
Bb4WRHyZ/T2t4Xu5vvT3IF/3X5jpSgg9UAjLxXSDWAPX1gCdVMpkFjmnAqBI2VHiNlRNNAyoNs5T
PLCsTiynY/FozneDgWlpQ52DqHk5qrk9nYN5GtvtDcWx5SlB2F+8D58o+2CHKLhaBcZzT2D2D38N
Yqcu3sVBpQIRWqQW6IZCZtrzx5wugC/UMLPtLLZ68JCN/rNgVUJ2kNHwycFPSSwhDDxUkxrv0Wsv
Mvrlhn6UOJ6WNvYg+vk2cxbehTOdYsjxxz6Mg0d15jvQ3mveuonTqNYT4xmWDZgBfiyofPpwnnQP
EyExA86TqX0p5N/9iVphQxL9otFFPMThwuW6ft5Z0YvmpDvuu48xkgENR0EK50zTxPJEUdKYnpSy
znQD7HeoC3YJjWh1oep2O0NvUNr9G+SQckrxMYo8G1UNy+mVf+epxag78+KWp6B32CxpraDJOk9B
p7tPsrMWhGZcyKgwF6bcdG+CwdJr2w/m99Yb9szILSVTl6V1nzIb9awJcQrAu5LU2ZwMIPMV8G9h
MXIxqOgbeIttRbdC/WEIFO2xubp56mGuLgkLjtuFzsT5Yod2vgxAhKDPp+AFLmcujuI+o93AHKkJ
2/FbeprwPOIwTCXwQxF1wgkG5GpL7eTOLyTBtqKuuMMnszmsMOYToLEcliOz541zxYCr/s6E4vnQ
GAV8MTTEUbAGo0cYkWmVhaYe9mFo+l0dpsTiXAoux5FnWqObdfZvHfbOmhlboMRodkr+UwhCyhQm
QfOVWe3SpFF9LPxc9O3gGLS2UHxRwnuODVeBvtPCHEFrTxhXbew0BCigFCtU4EopuSL+cqtIclpZ
Nm/W89+BkPqX1e2T/m9il8ht7m3wzMfcW/f7UEcNLRXESZ50aYwkP+eWZ2N8Xs9O0FZ7wgH3SeM0
0cWY7TpD5w+yV1t3prvGMqGqHPrYJX03g2+M9qqNCUMSHa6qBIWmd3sY0Pc8dhrCM9PuOBcPm16K
FW0v6cQXYxC2Xgtk2H9tGDiuSq+1DaAramEFoIyjtgwj10nvfvEfSdyTAkCf7H8rRgWkWLs1SXX/
P9qPlkkCGlruXOuHlXPGV/EjjhXdTNTXSKlLmzC53X1lHSLHN7QaxYy5rA09hMzPx46cp6TSitlP
4Kh6q8sheBpNhk6jVotpeK3xqv4FFhsYhBSIF/kwmpQlgEqP6Dm5D+Av7mCIIrgknZbngH/DJku9
KnBGGJ0OiZAu2Xf9rWAt6Hgn9C2w8CrMxQNv2PsZyfQMYoHL2PP7Tu7UC2gQUPM5gmzgJRno9uUb
tFs1eAnUwrxcXf5r5pB9+GORPY5FtO+Cirmj8CC+zqm0pSgdFg5y2CEkZO83CwljFbIp6YIi8QVX
kBRgRiNPVyIwKKQK08W+VZTc+wqjwlHm0aal9Rj/TcgBNvRbcFaStN7WRcc/3n0sr7hf2hDJ2tCP
AnUPfjrmNEmghEo0EQ3mzsTYQ0EtH80yn4KNOHW37I9l+S0NdXiCN8yY/s+oPJALm+hlCCf1Qv9v
hEDfclt2pFbLS0b0nFXdtce8Eif3VD8IxFyjJnIFgLo8ZH1rP3cc7mWs1vVc/eZVSHgbvANxVyQd
ZTC0+NpmqbkGa96TDYMr/vwimYCXbnZ5+fmzY+8IVbfJJquvAxKwwrHcf5dfa7d14D24eOFezHYI
ncPmCH07Fny1+akhG68HspynIcYDaiDhsA1pCp+XZ9XRGfqyzt3eW1jk9JyTM17YlvNU+Cjpa8N8
049NeSmdFBS9bLR6gU9XbmSsh8MCa+LK8JCtfTQBn0rXwJLJFoE0Xx+ykqUvjxTNmBgFSu+Kmdq9
Eq6q0CwhMmrPumlfYQLfZYsM9lJxmwVc1WlMX0x8mzMqF+FYVza40C++h5OaJ+oM9aR8VpbcBMZg
cnONLRZZNolJrGfRtMkdhUeMPasjeWw8+bIgDBGSd5ckAfzx3ESb/mhDA711RVQx6eR5dk0GLo2C
bZzirXc0WekxYgO3Zef8PXeQkc83UNmnnhHljNwfuB9uwiYEpmO9QJTRUSx7OLfGJpHL91Xx1I2y
e/7qc4lbchuTssfDoext0VUxvlSLgqvdGZYP5wYt/hAejzo56wTQ1ryJixUKnqscBD/ZFe2XixHn
AHxqGR+ZCdKymcdZHMW5klOWpga8e9E/W0V3Riyxgm59jp7VsfBivTjohDnorTuq2AA/SV1jDPDB
frzGGn7T/3YxocxWVgWRMyjNkFfQuqausG6ANnZMa7S57hrv5hUW5Yluq6tpx/yvy70q0843rG/t
Snz81nZXknQucDk3Hy1P05pROLZNV7bAV6piLlnpScmaPy0k4PdJxZrefcLVKJpbZ9UYnYar7lL2
8RAoKRbozrMY0VHvy6T6zmif34KGWCXpdC0S1kr2xB3sewht
`protect end_protected
