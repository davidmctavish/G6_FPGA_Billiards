`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aWz3h3BVZPuBxqqTI9JSuLmwNT30skKInBNo+M2eJB5kUxYxMuRIrNKYI/m/3183iahS1zqgihwQ
4Ziuzzfvtw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dmej56WIjSlQVrfHIzLIiiAerd0dyr7L9ENmOb1Tjm64HTk+MQoP9GxNmmAAmod3YCNogKm0IQoF
mNrJCyNh4ZbDLV4qhqHjTwksxZVv4NN22eweM3flzq13DdyP5rExtAZeCaStTNrR+ncVoLMjBL+u
uLayA/U/rOuemP1Np14=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n50eMQw+zJ8/7wWxqQvDMhmm5MYLID44ULP+2Jz1csjUdkDd6k2/TfzXDaLtbXYJvTgBTtOpMjvy
ZS0k1WmTKrMh2vZgoAdRCNDQAu9kF3ArLgb8B4uBAck1hapovFx2L/O9iZs0qXJXY2mxCLrRfJrQ
LSJgUU+BdPjP2o02JVtWOnHd9FgdyaexLq518s9FEsUv/60eOGppoSqWEhP6DK5W0W/OAsF718n6
0dN5eEAgRUxFxWDt6bdDCQHW4Az004xOaxWzZVJrqJN6ZWz7fttouevuxEXBYudFHtR2Jl00e7PQ
QdiY08HF4o6ThtIYIqT4LGdBJwkdWcHkUWNoFg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ow9ZAQCcAy0m+q732k8JbmT0OdZ8X61TWc0m2KE6ehKwbOXr1eTLkmeHYsXL59rWbZ7kcAJ9wD+d
2IQpgkPIliqQ449d576zHejVgKHzPCj5hjTi0A6cQ+RdEjxmqFeErm3/oqYd8ue6SIIJAoLhLiK7
waTUV83MADTbK1jXL7s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E5jsJHS9jAm8sMgeoTC3fqq/JwFTjjl1MNhrvYOVQNUZ9jQQ3GmbceSk+9Re+CtTIGH6tnD+0FdR
gzG6CPxP8ymO2LnPlqu9Ya3SkZbiOOvy4MOnl7pqTbZQT8thE8XWk156U8avvFdKCs8falUHvlg2
7mLur8y2wqqzC3linmRMv+05RI84tdd+rTtoZM4fWS7UIN6O9Sw0fdc+h/e264k5nZJcTicAiIoV
E1pwATSgasq0PMxdRTwK1agH4SFrLAzejL5KXSV69zvviGvPNLb7Vi4fkku4VdnHH2/0euSdJaOt
OdhLSEcFcwFSzqhyfZ3c9w/4pE2KWO7UOajVAA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20944)
`protect data_block
SGRY/w6zCmcU66EFkBrMrPNbD7xVrfEHtbovGc+y7n/Wbl8z5crPgjHpqghXZQPHvgXTzMvlLX56
7GmSfEIzsjVRri9QZibGZkt33MDpxhaHeG8kA+OfN7uUnPhvcDivsiY6qhkQPm5gLIi6f4DgUUaC
h12mFeVovHGbUwriA2zMeOazcPIjTFUZS6ui/A0U2dQ5lJub0CuZz1lIzn8noZF5YGpAkOGIuHYq
Z9gWLKdBtGsitSGbALVf+9gou3ZRsWBA3ayJqUkpne7rlLWKYtoTKYpl5jevfHu2ru9d4b1SDg3H
cSN602Idwlq7GLVmbhiiSwAJ4uy/Uwc/FExIPd4r4XNsQfodTmjnGFpfPCY0lwTF6POgXEBe55iK
pam3SzF9IM1vOGfd8XA/WeCsf6ku6NkqQpVi+htBXhEFXPP5IsEonx3RqwMy69w22HYMjojtfp9W
JX+gblwslbBIv9YKNdReS5ISIx3RkxkUy8cm0ciuY681DcmA9ISV11JF9M4Yok8Y3PGNs5nZ6XAz
T89lhvDG+hVcY5N7vWEz2UIgSibmAtRoYkB6vT+GzteswyEOz3xTPxFThR/8kqA30v7iux2AB3yY
Bd7GESf6NFaziT8sokx6MOgioRDMV6TaaVsKiVb/fDLiu+JYyvCRzlt8J+tDXqmX1wqDRtZbr7Fz
ASHv+iiY6g3uYmk0W4a+c8orQ09o40ql4aFB8gJWUUApoebXSdzUVGFVfxBYvinQ8veN/pYFU7cl
UmJ2ONhol3kGwnpPgy/1OTEl9sDCTzVZBTr2OkIyggHnuP5oK8JfwzNlZ2mHx/dOxNE/AnGT6c9+
D9nyuwD1m8+eIPJ7UoXLJjw3+K03w/vOwLLXHGFSYongtT/UHio/OdCbUvT9OgUUD8m0nH2RpX+t
jcxE+tMWPRvWoGHH2EB2LvOcrW7c4WHRU0Nbcxrh4AejJBaynfDV3/xz1lSzHeCc8KlsAvy5/9j+
2dWi1ADbApQLe+MShoosyGvDfaAs3bDPgfckeQICFHaKgOC6xuELcmI+Q/c5yj43eb35m7lzL7cJ
XDeoT6aEvZoYP1rdx+2Rt+v+Ul4UMdGH7T6ae54IvPaOpgCxKHrFQibEvrdJON7ffMuHGRHn7vla
mHWz3J/m3nvYW5EpOPlu1wyGSNLDC8Z8WchOorX+EA12dmZXONO6OvMqBqXxq0cl1eCoIFGNOXo5
tfJPS6qKc4TVif8GOUNxiImaTV/5QLTocUoMqARaX8QocnC4vsr3BjDUChUC8OSuwmCb7QMBlBhv
SAhXCakwTXkT/8a85MNCj0fxYVPwmuAJOUCrOuitnMv/iozsf2yZP54qXXrHufzgR6CnyyhfXsFu
LQxTaL4z9m1KUpyyEA0LnWyyBu97qOOC7tajh3jNzy2lRuLHDsWtHJMqtw0XzkquZGE9l8xXig7j
sncLj1FD5lEiddbgytcjcu4K9KULC8W3YkDVjV3qoL8TPbUcuh7jF9bvn/+2dJyw1PLW1i+h6iGD
V77otm1Js14JX0FMuZMpc8KOBbrmyzkBek5pKyO0MbxJdLh6JRVfAEkEk5IotwxRWrpPEOQCEkRN
8pPpK13Z7sSLYUJ9459VH9caZMMJWk0Ifqk7/2dNpl4J1jqiLHaYSgkgGXS2Vw3IGMPEphpSD7oq
EOSkGrJ7oedjMxEhb7Ta7DpK364qtl6Dcb8xFRNsPHpiECerMH3XpAqslEIGtR9AMAkRTqoH0aQl
ANOHXZzzLUg7Znfl24wvNSL7nRGTYWjoS1Egb2FT/fmUS9roFmpSL6TXTQiBN9vQAEPZGFJ/0e+r
dgnlpA+TZPT3JVwnXG8XmswfkDVChD5WAS17zxMY2kcKWWESztquO77gf6Ozs865KxwgD7CN9Jpx
71BEUw5OOdBAGc2rfXIBry0l5VMoeyiME0kgQHXFb1bOCL3bueLlf/DciyA+kSzGjH13bNsO+7Ca
Ct4VI2doEVpYxVGXX7X8STSm5oY3G4ZsykBn5jpMlVhTBYKU7lb+34KI8ATfzqM2JuDtWSvdfD8B
dihPC5qh0DtfjUi1Ahqk2JTitGK1eANlFTBtDQpEBXBvf2AwZzbyTILTYV+uZZK5oRMZkUor5IVE
E28m+SY/4zwDc/lRXlJpo7jZI1N+K2cruXcr4WQz3SsbXNgXwNJ2s+q6sTzi9AACnX7dEQnE7BVf
+5DDmzrSufLT0zsmfbBaUFsnfchVUVvqa4kbIFtErbxy4f5UeqAXwrjGr1dPW+aXcZP7JeuBv1X8
c1O8s5j881JtAQFu/RMWNCHzQ2pkoCqER8LgFCE7NKuUo5hblr4Vu++LceDUnjM/olGVAJavZlzy
W11nojQqqK3HPzO6jRmQLJxh+c7lWqss8VSOJU4N90Q0s2iloanUlqAmLEv3jDFJidhRZvKIFN1z
v5VMdfFDpcQjpIFq5Nobw2meYSAh4OX1ol/qC9SNbSemikt1VbSYzkv+XCdGOgo8ojlW4t2sNE3I
QG67HujpRF6PruWImmGt4IY9WtmCH155w05bg3lggfpfpl/T4TTqTag0mk9n3LNYFJn5bhy4Uhti
jloNc6woNhsKJ/mv2ptWONeXm/kceHHv/Dtgdt/oOX3hfa5a9X9OU4OXaTlJGP5oQza3omsWpIpc
EMB+W0tyULidat/xqFc/ykb3r/fVWUOiKcC/sKjC8LIzTawlYCIHKM35G6mTD9+cZqzAdfVoSG0Q
2eS9LUww6FWlhyDWnUV8GFOKBEgaDI5uCBp4mc02O5plGb+I7CnA4IgVa/w90pACx2D3fYyfkipG
bkaCTeX/BQt6ORirHL9tfBseDqIBEdD/QL3TrcR0rZYCKQLskGksc+s4IlLj+GmWpw8lPsnr/7PN
hu0VQY64RTHwUdeLFyFIl+5pMpiY8anMJ2fwo9I20dmgKRcXvce/rWIoVg2NP5o6sPSIPiRvzXTE
wUgFoQ+7DxJJhHflIymElLSu4esaeO0PBLlGQzbZ9c1q8eDMCj9ttIWazDUtlmqecwMOGLqTrtPR
fQLKXTeRM92jRFUAPP6fnvQ2Niz9zlEmYAfP6n0IkNxxrETlNyKuzVcofHFddPFAsg66Z/6Vumy7
mf8gFUKHIsr97IdipCqbhe+xxd16FY6KYw3/WAz5hxlCUWZ0Qq1gkGlOxsX/X7+aVzeUtPLgicK1
a8+MCQBTDRoXjMwEXy9oMfLNOlvmvLQLuUVNrF6k7QTR6I96uiXakHHYpht0y4lMlGjwvg7sbGbl
6D11HJosuz87Mi+FubKQOjMFsRS4wWSoJBqf27YQIumdsu/YQSQlYugQNHyeIIYEEJ6/X1qLvQZc
l/DxQ6TGERvRuZi9ww4/ppHP+pONT7VkNMW5aF0TuSnyu/egY6pkuADA+AJfPasJICacexF2ydaU
Ove7HXuyZXqyr/x1tvnvoi6clmAsO6yJJjSa1DPO+3gixhHmWjRV9hXg/L5HRpM/qMuiIy1rk11x
Yk8mMAav0UMxLpsfH4deWzBtzctbeqL9KKwIsdI8ohObdTsqxJSPZMuJFlHj0G7stJf3kVm+rbFX
3vp/dR7tu6yK0wANhFtx/33Sb50ALr7vg48qJFRuSDd1gbDM0kkdmBnGdGMs7HTArP5tKsY/WULm
9tCD9g59Bl5k4/lx4u/1ZAChA6keWuOcRfPL4JMcGOsZ5Z6vReSnCmeXGrhs4jz6zaMAS/a/pboz
NMEmOp1GPbvuAAAQ7UYruuMISHqW3lk/Q9+f2VdDl2DNKLsfEHDZ1TRxEYc+EeKQFy+8V7Oc2Cao
vyt23vnkNZGV6XYehVx+i0A3z8CNn2fAKur7ZV+mRgvZu5YDjppumcHPS8S69F6k0oDiQGN7ncI5
TLOfSuPV2fZ6X+filYMLwN0YDrYO7xbmldNaOpPEpi+I4ny69dl2BrgoIN8etOXh9qeu41VGM3ri
5Lzia2A7xPemphD3vVQJVKrLoduhGbHweaiM4Pol8CykJ9L/bIgL81FUYtZtfXyRYdp4NYKot0mJ
rodZwaqsXWj5R4zFneeBDp25EJNXbgsWw+ImtpEyIfZs4v7a0ZvQbbGudscyNnSMDls1bp1HA4Na
RcFOCMQi8RgmegMLARZVkUM3vQKfpddUQsqI8TPar9oZZtzWuwuWkuJyEZGWTj2us/oS7Uny9XuA
RsTSsS/9x71RMS4G2CCpWx20+F5iZdy6egsSsSUKREmPQ0XGwSAm1HvkC+SX2t07P2J2FtqG2d0y
CIYKfgsSdOHWAf7UJ843qy+isZPpxhtXv8Fx0t4B6w0XYt1qL0x5aQ+qEbvnAnOWRANCn7oQzji1
wVHCZlXSri5p4+ckUssB96l74x8x+EgAMXnQtcam2atrtoDbGSrETyO0Zx3TmFPTxiMxkq9AnTxR
UV/dKSg7pBqaFk6rV4HBOyinty1mLMVnChLALsjN4KUyIjtFwf91aaXAeJfoFsM50tnIz8TbUKbP
t8ouijEaqGfnrSkrW3JZzlualLn3WQ3UVm4kVE8ANkVfPD8Fhjd+udl7IqFCPSY3ExICosHAU9f8
nQRIpdkW2T9d6DyCt6zNeVAGLXhyhk+pnMoe/rciLpRFJGabbou5QxJv5EoFxtSjSRP5aRsg4SoN
YeCfUkm7cbniK3R1L6N9gwX/tyy2G33zXajTX2LB8r6X1bWD6opeE4mmWn8JUKgMPdWmigxdzu0q
/WyOQKBEjVx7AML0Prf75n1ytMak4Fs+xrrhLJ0AoGfdLqqR9ikRToevCs5gXXhXKA4XsGjkXunp
H7ed+EIpkVO55rjYr+43ehgvpWc1spPxqD6G7HSBqPOablm5bEPu/YqEIK6ZX2VE/hMDN1DnHtyK
zx0199aSVVH6ryXbf0aqTmo0KVI9KvcMtAdEjJBpvw9/72IMb6J+4Q6EUSuzNQ6l2O5C6FVKLMLH
iwZRcCGykIsqJ3igt1YlABti8YoBLlzFWlqxFnmPHDz2EqzF4h9xZFljIBNBlG90hiMUwGM6OQkZ
EPOSxfSnT+6t6IgtRWhDj3EEvM3/+z2rbYYETkKT8z/JwRAv+uvMhyd0kp1vnT6uHqd82WvOmsBg
C5VOlor0UVpQJyVDyAXGrPGN1Wl3JOVOF8HhJ2H4h/CY/uia7FqmhifttpJz31zTWAuwqluO51Mk
eU0+modP7cOmiFkyI2vzyeC8FK+3+Ol3iVX1XbZUr19KBULjY5t4xqoPfRsTnXehBHdAi0DHUrhy
QeRxrP4FpZh0+zOf6ISRQm5RHB7SpePWHp5UZ3i7PWS90bCFbZc7lujYELZ9hAIr8ml8m4JllRuP
JNgQOlpV9pCtA/OtWhdNDwG3tUHyomLafZi9WNFjNqOvJw7c2nFt758GWG902d+QhtrgJ7UurYdS
swo1PdVrleA1YObIlyRpXzBGVHqBABVcmqMnVSe/4lsRMC/saOX7xy6HbQOs+oet2ocdqKcuCZgf
5+l1bAkJINleiONkdAhlEbVw+rvhUuDfZw/ccoEtnnocjZ5P+v7y7YMCaX2+F+K20f5e1+dQr49E
gpzVoXOJX5DWKfNoI35lWfBMleme3bE0yHm2c4M7fgxzWCl9k2fAxpv4ycXXwe6z4WyLxsPgzLln
sWT0EgxLf2DupsmaC+tyHRzzhbkA83thnsS0rVLppTdQfnBxc9wTwcdQHK/eipE+YTUhw44QEGoJ
myqJ/vWcBEqxen3hwMfTQDYQFcnaQb9LfCRuVI5DI1nzX21/q8dqvaZ0txCybLHLFXNDm4mmK6A5
JFQUKSNqI0FKOiNDHfBCSY0ZRJJahjjyASVjhR8scBlgSEYfphn4prCIVuUQkks22bqIK1dSmnhd
0amtSSZcdxlCmyjL6nqMMLbuR0tibeWJTVyP83s5Sp/QSrbFmrWvptImwryAkYIChK8imYNtRTeM
Tm8lzeN51782yVtN0DAi6NyI74Ia7nryvrfvkOqqLrfvOMXv935lz/soJyjyqzmd4pTmIpND7fgR
N65eJiGj50vSLhWTvWzQ7NXnxU7sJaWROAYaQBFYleuYAAeGV2M6HxwZ+lQvJ6z7Fi3+0AyJ99RI
c7vhHPqddPRRuk0gdZ6UXdNpfex/vQCw/Xf8U70fps4AojCB0FU8mvRTlzCrk542oDvEYeBqfbaC
MI9TgFEKd08gvej/b8SyBlUaaat3/5gKzXmNDcpRpLCaE+uU9zgH2kv65+jq+7ys7KQS36yHwl8q
7z0i6DIDLNVCopJULzT4mu5LynLR+DF3sNCi8kXdCVzBBmwc/zgGqv8DiXv7PH420tR+rhx8Egg4
t8mocU9DADElawsoiU2oh/mRfs7yC/Es/+ZFBj+ZFsYmq4NKLKcuAQ/fSfFSSFaAOlrQVtLhMr3p
eQ8Q5tx9m9tibUrbaFbWZgBOXvlVxOp3r2IGDXkSrsnYFdDaeSMF23VBADnKH2lyN2Tb2kR/ZDZ8
Q6ouH30VXg546AyJfsi054qJJ+1KXrMZYPPEwduyQ/rEMe5uhlOpntR7h2PcX+7+KxQPkqCF4gdJ
AIkfGS7ibz+y77NrvEO2BZ47qfb2rRyZenPK8i//gI3GqRuvtOxo0bK1b7ID50n1fy/nzx3M67BN
JhoF/bmyYyeacOXoeVGI8rD7aF0cpfFvA/f1T75TsCypyQRjBqsL64Fws4LFxDyBs0pj/QwpdreH
6N8GL8GvHOe2GWOp0im2igGcLcqRF4SiSAXBuVNN95Het23QSFzGFP3vmTTd5Aq3PCjU8W0gibCp
nQQXV2mhtQOI1wkrccrkHHqgjjtYkbAqZRBaA2gVCMo8g2UNO7O7JYnc41lAGc7+I44xTNIa5YwP
VZ7P4Q3hebNwSKOCUetIcqpwyoCIKBA9CLMSt1S01k0FhnxDp7awjvyueLTPXjjuXAGqbPqQofjP
lbrtR2tsIKjQ5vdPyKSufUsUJYLZ4Awcoxl7ynupsoSta9QzgOcKldJbSqDlJUFqyC+8RiKotYuT
pRCDNqCdMlsTiE/VY8461TIAW+ZIwLZlVAU/KJ/92eu1cpe2bvx9PO7FJlTynteoYtDlwADzd+nw
ht5wfJGiubzitKBpR5ZnY05xNFqMomJRCPLfVVxsorf79UJ+YRvgD/YoTwiPTXcwM8aMLKPHBoWO
nLAOLo5fdq1ee5FvGy1eugFdvsx6YjJv1//yzHE/UEJsUf4CY954G3rT3uAAg3f/Buhjaue4qw1y
fCGvaNJV7IxoXf+W9SnxQLWmRL8a6NynYcGYAhQxuQSt5mBsM5UjmcPGPi5XdAjRYuGismgiWQCC
eutWWP5TeRqodLc2BmRvjL/ftdKPcrBwuC6oSHql9b+sieNzRwhjSaXkBQO3g5DQCF7QCIBihQWe
XlXfr8wG3RGCCcp57DOgE4fpg8URqF2zyTvkceGzMmcS/DzCrb0ohCgLhxfWrKpfx+AWJO3+esNj
fR0FpqdUYL4wW6jWXQZvOhOYyphFvkk1Uau+HNMXXbreC3E1ygXDY0LVwAWsuRJ6ForGRp+QU93z
Tlk0ubk7pxH2H2DNu/zm57FhQMi2yB24SRXnlAj1rbgylka4Q1CJM6akEr00BgLh6I5ZUK22ajS3
whZWccVSPBu7RF3w9YAqW66/BmemiQIFexreIN2XIjMYVAvnwnLP738lJaDkqw7Divb5O39TXKe/
m4xI8ASgJK8h3i+G2u20o5ZW0lyJsX3rIL3wMkqLF7jOjb3m99tMyZJuJXcHnEN7Y8je1zfQc1mU
YGDDDCJd0rYGmT1OEmSQO0RqayHNUEyZ9x0jTE4HA52Mg46flXXgOSmxIspJviByImDwwfGJDFb3
4r/blaEhA3prZA8oebVOBx9IPcqY35gS2kWFeAaW+AJRXeiPxbgpNGNI3xvFaMdqqvnWGEYe3y+B
JdSYnG1AcLNCmWcf/vZV0jCJC9WMOjj8pUIMuPKJjsfd2/o3awh3dm/tgGKv1sbGTFOnBS2XEN2a
yIrSgQpr49L11LdRFk7xXLBlC6zIWRK21TN4gZgOTiZyC8GsyKcedTjigh91QbkIUfdVN7SDQ9UE
nwdT8yCH85tdjwAz9hevKgFwFILm+0+lu9DyByWesJqQgjo8f2hQvQBW0ARSxA1OHzu8vxEiParv
ZTLQSsfTp3EMj/sU28SWulfpqy4uFkOTUVqHGNbolyzNjuTrfwwYDZdxYlLxqw13RBWDCH9cxdcy
w/PcXFQ3RbkHwlq/tgdhyZGijiqv8lNhhDmQaoD2fMXUffSD/lVZoyO4JUigZx/xfpzjfHEBDmfH
haF4IHXpXZLW+mO+snxI7Rbi0j6seJH8qfSjEOwQau7Yg3ARA5IvD+7d1YDYMYhkbsX1y8c7iCHi
7Z1xOGG9ExxSXNiyJROG/IU9uczBcEgUG2NiVGp5TkRkFYy293T/LWlGugCMtXXfokynlmUZjkwD
TRWQRigeZJHzX61w69t8hz9gSetVcIa2YRZPELv4z4PI70qIIUMrwFZb6tkMhoBWoLcGEkx0lWlp
PRhMDSZCGdFyBtwHv30wbRVkkD67MfPZPYDSjzpYcruFSRUu7B7NW87qedTas3xBKVUUJTKSShdl
PjvHD9yKiSvMhzvjYynJHbCKMB2SLy0TkFq3WS1eCQRcE88reORUwxbr4BKmefvRaahB78oTquu6
1rWIes8+/FoYtTzMpn3Z25CY2IYhUYRLizly/B2dDYoDD56YZP6KACe9kzbTi8tjicWYSEPNO2mB
yxkiyiXNUhfF0sT6lFpXVzDJ3NDwc6i+X0grPWcoQ7vhVz3rcQ16+32rdmf4kK/ZiU+D1tbqcTBH
VmbRLITt/HCH+LOzK+zwyEm4n4UEQoomvZYO75ctZ4CxE0eXoSPbtZ/m35ByhcNxVy5WKUGFlOvk
jVOV+8y9cfP1xosoexjcf3T/kY/2awI56flEuUB9mmb3Wi200qJXvz4e8RPM2c/C2lbVV3OLM2KV
lkTILnAP90/xeX4qe4mkh9DTsXkPAPSFw/gWJ2ns0Ap1FeLjjox9Py6/uYe+WA+YnF9IVplqafKn
FJSZpfNxSR5zIdKCJEKj5IND0s6O/rSkGHDivBNFnVt8LffvK7oUPEfdFkr5l6v+tzReYQSIb/vw
GD+RKaJByGrqTIQTO3mKbygO/iuqP8BCsnVyF+GrsipbC6FS2oJtd43QyLqgIqWo6e7cZzqef74g
Ay5D4Km3JNXVT6LFewvcIs4IJnjYNgnSVA0heQepauAPT9ddqEKGRZzH1myrHviGkd2aTtRp7862
0f5ecaGbLh8IVtHXt0yIRx5DhQit54tv9fHOuBUvsmhHACtnTKNQoAeB5+8DqFtup+rhsV73h4Em
e1JdC/7BltxBnWqPX8XAusHbeoo0ku8XMd8BHn4K2XtlKWvNUEK1TigG6LdrWTbS/uLX1oi7TUSl
p4X3KY2q5jJgr1TDAlXJvZ1IjbB40psNWBpnopHEfm/ms9eKOIerd9AZKSX4a2jlhblGzyfH1t71
gcnNSttW/KzKV32srqRj7Ben7fC5FzCkkGqqTK2cuvn1LwDieq0XlGKYy0BFOPFwNGUhUNHuuU+S
KVcXA44KHEq/NYc6MQS5HpGD/cj9UGWCGdLkTD84Njy3Dpf+nhwTwUrMOtE0yPabg/sZ23Iq84si
UnJ5XGmxCHuD8zkET+i/dYyMZo8OY/zIJDL9Zoq1oVmlfA18OUIu9IZQj4I+LmjmzROwrTaBHjtt
2BXgtFiUevbopVxtirsaKp0/cr11UKPd6PXNGN/LenGw5nZevHgmznN6axiJYr5HvxWaBFCP+yuH
zBPK7/11N+uF3yvr2QRbQVcocKEjnG8VnoiuQOr3L+R3PPJTFHKcbDvgo/egCqeZXK2DBHWFEs/Y
e+AGc/mju352PMYVGHVnUxHH+2XYU8cg1pz/Dd8e+68XvrgcRez4XWmsHGrJDm0PbZcAJ3d8v/Fq
9M3+9BVDLF+/sJigxxQTETKzV48ZBizX15HphO+C/xudcZNZTBpIPK3WxWFqGhn+RqeMyge1qdEL
Lg280F2+EwZp4h/mywjXc4XmLMDFp8sw2FDwBI8oIYENl4qGYqowXOn5vrWjo0ki5OEbDmYX1FI5
XUUG0VaquGoZVo4fon8PCGPgieBQi0w8R4RxmYh0B/QajzpepjjvWz7RixbltsyB0KgBtpB48ICJ
yylYXzeJh9EAbGDQlPtRGk92qJ6cf+jLaBfexpgkwCZ+dYnaS+Rc5BLRP0QB53HpPb/lgvPnx4EP
fdbTtaLz+18dP2Kv8DRIv2uupYHRuctDV1MEYxxeDkqWO8mHT8qkPyh9l6XKHmKb68wtY04MzjX6
XD5E//BtIQ92nZJcgBu7068k8IJfXLy7adGp4Ebc3e//8HgJuqlMlJHg/OD005RtMWuK2XN0jDys
zz1eMYg5RSj+jyE6GDq/X9rqzEf7+VHkUnZLKoTtaPpMlHkwsKgt+Lz5MCeW0HkziYwgiypveiWT
bg6FFq50VWFdf70vly17bp8fvE5tAH55x/aYJgSckgNe9s9Q4dkGhCdu4QAXnhSGWLJh6IqltOOD
QFqjiGLS7EOHstjw8i3FPhe6ynzfgZhDjxhIkx5rQFG86iS10sIx98Fn1Nh1HYRZwrXf6hvQlZnl
gENgJ3O2Q3He6c5jA2U9CCIRr75IkelzellFbtA/NSycx+iMcylOXKRzoumz0IkYtgoxVfMM8LR0
9s3buEHlTG1QD8+J/h6LQgpl+4lH+Aav3VoitdpYyuFoCMInj0azXgfYOWCR08gN5cjD4qP7ttqO
y68eRFBnTw7syxloGibOqOGX+yzhmGLcH0kHuVp7v7ZVxg6m9aFdvGjDHKxL1gG4fX6Fmo2HowzJ
QUAuXbZ036sz6XPlwrxC94vC3KfpsJ5RJ1w45qacfnZTvT1KWo7b6ukJozecDICadI5+JZq46JWK
VMDer8RL9Zu4qlq651jBjjJDtmS5gkJ6CesJeFJeTknou4ybzNAEuH+9a6UeLyHwwH/NFci7Y8m3
UDzN3XQpUN1ynTkJitlMQJ+8qaZsWKKEnEqEbopCuNKE0SwXZBWDbCOP84Hx/Hx8S3l1Pl4z3IoO
oRCX09ZzJ2sLgT3FVxy4Mn3jOPQQ/qVTzJYLhWIB4mztENmoqC1En05Ro41IH+h/WP3vWSC4qcvE
ieh3KNMJqe9PQwJuUYY09T5Z3d0h3gCJPk/SsHACPatEnCHhwTQ66BS3HM7Cy6ZRQpAeNsvbHgnK
9gAHiPKbMNIdJrX/ofGChYW7JzxMz+xH4T0IP/dHUD7ffi8KENqoqNnk8MDF8hj04FYYTWJ49Uku
U4MStkqKnFB/rGIM/qAjDlTtvzrIHBASnZIW/yTPKuyOHrcwAw57nrTtcNi8WkfEpGAh0wrwFxZC
al6dhZ0acdRzH1evn74LKa7NKMO2oI+ikyDeGErRkAMma7/4CPBlhiW+hQBwTVD+LWhuIDY4s/jE
Pk2YkMbvqKAtO5iDeeWpNqIXUG0ZY+qt9yNuTkzaYktf+uxPl3/Xde1aMTr5FKfpwYFD8SpmSJYh
Ywdn5EvwmaTNs0YglIdZPcATk1GVdwO2KqVThRnwZmVeUgjmk4t4ZLLhpLaxgQuW4jtLPVGOBRhm
KQgmZuu6XY+7ES79SQqLJ+y+5FD+KvLAD2N17NJX/LgUlzkIyY25Q+VqfoHklR7MufBEu2qRpX3f
H8G3l2urb3fTlL7D1TQv3ass1L9GsAQcGZ+9tSPtlc6VFEORF7tmo3LEtwH58YofwG/6h27W6WsJ
yeA4sG0EN9RzTWXC0m1+EQ8RGBtiyIQAAF/Q7dk3bp3mhpks55YeYQxCKMjQWCugPoe7l/Z7Ze57
QIcGmRLSat1cGG6DCNh3L7zwfd1W0POBvTdoPioqeDOx2TjC53eLrgbThTz4Bioh0l02UfgrxA/+
3vpiit7tcQyCzJeCpkIunn8C/paILNrKPBadnHx0BkFue8NpWFEi+egmnx8Brpv5N/4QFS+dZkRh
iH3yj5vsGtuw4QJIUoM7k+e+XOkUvH2kwVv5Q5HZpjxm1R+7bN1q5jh/3kLkN2GAynMn1w57T/DJ
829PwJmtzs3DrKm+dCynxk/v0kUinC991Rbb7zo56D6AMN1WMaILdrEbKK+07R0a1xrwXkrgCh9x
N7pFOBVdAe5F0dt5K0zrPTGTe7gcKacPO/N8FXz17Qv4c/XAtjRG+0M8O3gkR2uqPCdnC/8z+eEs
qyrdxw3oNuJKcBD/1+UJEq+EoIWT9m7OMHNNyoHXAjA0Tl5Yzd5Gi1LhpW47MQJf2JPAQglIp60T
JZD77/r9/Xoc0OPVTTKfd8olN8Or1dJsTfROUERSQWcdBjRgHPHGqt23LLO3mXf29Vw0WabfE3Cx
+xAsilxTT/dCDVJbk2D3hfh2mlFH1PI9UYQXunxDSz9N/Hh1pQcHZZBBdmvg3nN2yNDNDUc6AK4O
2L0BH09xbZ4+Du6JgLKfLb7dhUSVIR88XbD54qyBYK55fvrZc1NBfnte68FM8rphb5IjCNiIFzog
y+b17CUO/kVPW9TWsk8/8914rdD3DeLIjfmvRx3R7jvqnTeDhb/tZ8nir9/mkF1y8ZXfWXiQzCOn
a+6KSTDtRYCdYwBW98I5P1mxysM+wL9wL1mrULMJwoC48VjFroH70b2LVN7F0XWtJNMSclO2RLl/
QGuCkgOgA/v9B5o3pggZNBScD8Dgw9H70aL0bPSvtX+IS/c2+OGSdtHbshHDXhQdNuLsbSEn8P6b
D2J6bbogHI5IPfeSlFTA+cH1ROmKclvsLG43NSL5QOriML7bmFspkIlE6zR6/U/eRfxT46OTmkrF
1CfwG1xmHSTBvPU9r7qlkzm0h3YwV0PfdjKhgxURndY4+Sxcd0WrmX9WVR2rRfNkY3U5BC0UaUOs
ayJTxUQkwpkvK+svekYlrJrUoeUuY+ntt4hzeqMLqhIXGiyBOYK67lXCFET5XNA7JQj6wxVfnXa1
hGnrfyFQwlGaB3QmRkdOE1nvb7+AyqJvLvoike+TLyWe+P9Ffr2E9ywQD8oNhBRvQO7iSTjWPHvJ
r5WRxHhkO00B2CFh7Gxf3GT7waq3ypaST4qtUdieZwAZMk3uQ241AeiQQHaeuXaE8KPrQ/YWVfRf
F2qSoTF3TVGJqhR5oTMTQff/WMkIsLB0KXh7rrCLwTd+tsqsd+0Fnk+mYXXs5ZRgOrJLZegT+8b5
CZlgWD2mecbqKqs/tsdepkSgGARddb0daevnBjgA4dDO6f9Z+HWKWfBbkAV4nr9FlwbcEy5O1sl0
VL31E8Md52YYwqMf4uNfknhV2ChZ7ktqt7/TLLUQbwa1NMztsGsJvVDUhH+GlVuKgV9YLVQomVHX
u8Y8IKH7l4vbA59E6zh+IWiWBxycDXjKGOngwZUrnjwQ/SuhbarVgJhzpvGHVY01jC0ltnEruzSk
Pn1qtfJMyobcUJ6JooeMIaVEzk63Tf+NpxcRevgPt5BHJxN0YtXNvmgwMtB7G6hA3kdKvdKzxf9E
LHdfu5cTTbIbV9bjQcwA3TOhon6ye+YxX9Ah43vneDab3iBlbyfWCmFjnztUomVq3vSfBC0+y3wM
+1mlOx5JsdpGfeY/jjo3ci+dNm04VcNpbdfNBOk/JJ0qSlBxUnYkPuUiin/2Nfcm7xzCRIxNyaXi
nAEpSOUY0vjUPZVbEEknMQuwy1hiftMaPxebQNC4LhReInDyfa/sPFhAAq4fowZhhNUirSaPTxlF
xtCOUzCifRaJC5hwfNcdZuwaQEkn2fwPUqTj2+Fq1Jd0Z6DuHPpFMXyAsW0hZEn6eHBEgFPxKVBC
yNrqbt+7LQkweTeJu6RSYTByCIVBSeIRqbnPTMcxPiE0alx7IWvLbojJSkCFtSUtkgY7YVupktK0
TRJ5msvRC35uMLDz4iZxCXfq91qUsKp4mIENYeAQl5xMyG6GJhs5KDEWmB3xQPha78Gp9A9RY7U/
z6u3fdb55FdW/3C3GzJVgUAqRJEtsutKU8lzDMJ7TKce+7Da5E3VhO5/xNLCJNT9sDEVqeDGCjP6
Ho9/veAhu+sOOYr0uwFvI5dmsON5se+A3G83/ikSbBK+Bz9B99WH10+un/6dlO1uMnhBqxzn+vzf
Hz1ACKUTCOLDIC9x3E2WvYhOKNK7Y1joSKqlbk9L84Sa/jojlEZreiGmuA2z2qYHhTAFuU7AxQGx
JpYc/Txup12RojWqxeaxq62iPEMWODLkUM6xR16S2PK9IfSjuunV8eSx9kypEZrpDaHJBjCzSSq9
BbQqBZg6rL5tXCW+AZjjABLembTCDASgiLGmC+6zf3thR0YwDFu1Jr2rb1Vngdl+PFO9xZMZKhU+
gj5zPxhOLY7pLdQE/SbhNQKP7V5Z5p4NHtBfDoimlB95ns4zrSC+DVLPMnDRDCwSsNIIPFI4RBLM
Hd2Oomr+befopFuYL0wQ3nZr2EKNXR5bvjuGYgyctUaCmqT2V91sHngUquPX65aihFhhC3qmwuSK
Rzx2v6t3L1zhn4MPevzCuaGXltJlK+rYnGxLMddnzuU8LGRK/CNfUaTaFaa4MMYBruozCVIZs94L
o585kO0tFZ6BQJYZ4oItjs4jx1D8xO3xU1OXPGmfg5/ubRwNRZMXqCEK77tAx5KBV29nFYzVmNii
PVc/NWsvPvFIXTn1mhfz44u+IVGkjy+yWx/2I9fuGdcqHUpNcFyY6LvkbHFBgJGU+2e0SNHrnJlY
CYRhnL2Z7neHyHzuJ2nwDp/EKJf3YlOOknDSNEKUJAMMVR41yoOlR8T/QJPjk5U/tfjh8AclSYUS
ZkKkHKlWfg78+b07H5EI88gQeDQGhc6r87PRt+n2+5x8M0R3top0/9OinS3hbPW/vi4qdBwTkRLZ
2ex/w5SW21L4EIFMN9M0mtAVvTRbsWd1bMV/6gjntL1tnE4mU/W5LJ9/a3Vk3VLsGNuog7qEHgt7
KbemlATeZByovq6ZNAlC+aJljYQZtMJixtK2AbfqMFb/l6ARP1MXyfZWm/yqGISNJWuGx0tvAAvO
a0f8E7fAVWLUG08vhTRk9as//Np3MKkR953+NAC6hnJ8//yAYjIJLqtUpTAH5C0y5kpYVjIDOkdo
KWymc9Wx6h4Fw0ipJle4RuUEQ3vXiE+0XCNVCTQQ07vsGaQ7p8XiwH2IUUSYevckmsfgo0iS3ufr
tPMFAJ9jTlQe1uIThkthQbS+h5p0vUcrjokQ+OxWRXHof2oFz8KMUvmSeQbK302phf7qH2UyCIj4
j5eSZwfyRy3QFF94FtecA9dnEYcLkB3Ml1gzmI+2Srrcavy8P4fHLmfoNAk9ZkyDYCQSqLhbBhmG
HUl/6L27Ord6UPhoXYXIr4KkcTbEOSMLeKPQYh/LhFKvktlc46N94drPmWnG2QkOGHPnOheZnZR3
aavNv5W15OcOQjHzNGwm5jxQOpeQbQuT3MLWAMjLJoL0uptnTvcov0ZDL+t8rUAK2ZBn/VuU5ft0
uUinH8H7f6YuK9ChJL8Xu16GnoEM5c4ymRCnfID0EC9w4g7tMSh0cxEy4x4+6voESbP+9lnIQlAK
SSxn2P75JwFr5XWU6PeXaQwtHW3erz4hpQ3/oT/dpuTdwfZEsy4DEtHXHROfbKZY3mWOZXgmNLaO
6Sv6UlWcJo61QA1mw6yoqsQLha4ngqm6s692BV0PaGnekrBy7CwG9lD6uzGOL4qHc8FALmR0Yrbl
hzeRrwjcCZRhvcmHEJA55QXH45N3Vc2oZW86OiGak6LtgdgIw8ZxiR1+cl/7Ba3TX+7u7TMuj8ji
evLkjgNBYaYF2MGitkKThDscA6K38DIrfdxpM0x+yRPyT/aKTX7V4LkalQWVnuh7SnoG1pxc55zk
Mrx07LoXPGycq71fDE0uX2W+TOOugH92G9CIgYCVAEi8+j0y1142bmDu/3vV70T6ff3T5pJAdlsn
QlelkYt0jddhKzJ35Nf6C2uOJAzDEH9kTpvpn413BSN+pma1VcCr3pLWJKd+g48yxWSRc+EKV1o1
56tk2vq0EUPeQlhGtQJQ30PuY/nbH82/DPKzr0YnbRjVpAMR7Z3L1NLPykvUWHiK9C+cKKsFMVaR
Hg8AS0k+6+QFJS568UPHG2KZaBCcW2SkaN7AmGfc73KU7Sj5b/1Exn0Xs3I+fTn0nqZlIVES4Jqp
thdFdw2q5iWl8l8+lIjgwZakCpwPLtLAXY9942iI4FI9BFhVA58JKSaX7IgRrsCAwbOL6p8QrSed
bO5fVmzYzCicdTQXcHLW6ZJkdDyFw+d0s2BYAg0yvarXA45gGwUxW9KpHMAI5fGIIB5jqVOCX1aa
B0AzJ71lWjQjydM2AavdBaO2RtJof6qSMX3wKGQ9pyKOaGUH93kYBcK0rlniMAhYp1xkh1h9O0m5
ckbqgUGgvMvNphwEQ7ZVkgklt/wVnTTDDM1PC5brCR36YCiLEUwm2q3IPxIORm6SUM/J6m+k8pnG
izDqa/pD4UdHylk1ipJ7KMQIvRIzTS8HyBx2AMuoUUvki4L1HPFHVVh0rjSEtYxjeFaF6/Zb3zeq
8is6De+HB1XN6+zF4sxbdDLaNmevW5uLRPCXa1w9BjmJI70qTTZv+myPs5EldraZ12eiy83oBenv
CT93A/whLUF+6RGzv0uweMFhDW+Xqt9GAkWfvFzFMw17+zRrbgmS1B5/tEpKDbeuEL53JuVUQ9Fc
d20gHRv3N4eq/3U79+VH0nAL/uSEHdTgKOGz/FBpZDk98J9m+QWHwSIDASJccyeVEY+gYox8pHkW
lQsSCDiXUmc3CZCjCFNPHl+9OFvpN/iFwqoTXz9mh7viTd09F9lwjPu6lATkF/KvjIvL+lF7bX98
2+qPprkK0n1Fwx+LuGAMH6lOQzILK5kH6i5Tp9ukCocZwNw8wiYwO7ZhEXv5u0uykLAkqri3nUay
DdTmHU9UrajS8HxSpzkcvKxGF2wu05X6tsTvgV8aD+B7MljA1sf+7PbbHVHEmYQzaPYtaZ0P5WaA
508v9ov3iVcLGsv+TQmNe1VS6eMAwY3swKJ4X7nG1uUZzuKyWWBcqtUhdK9DLVb97YJrnf+zLK+O
TTHoJ9dMq++DpLfF9V3nrgPZ9L6Wjy3dNbT+hQZh/gw65Exk9nhIgjOCA0iFMTUI0KAHxA+UZobC
tD9PxWI789TF3iTSbB56pDAQi6YSXK+pTRlAwnvtxFWjA4d/zHj/rexgjA3ysLvIL9e+7F0uBasJ
210ZZnMqa5urc9ULYIJ8KECozDxGB/KhnqT8nIwr78Q431jbdW21SYE1dAvahTlueQvBmUoK0a4s
TPjcwFfyfCs41jY82138NDoc4CW5qzyb38QRpmblHZo+wrLzJJgke4rEKgMVFPU3atah6JlN5BPd
Ztq+ti7taSF3KXk7Ip9ssQNQ4sFgY41z+c3CmP8q2Qzbw1CaSAqbQua8cbf1lOd9eCSRD62+JXjC
tN9VBVf1ipzT8VVwSHTu8PxKmeMiZceyliFrLXmMtZx4JQCPHbMGI3W4OCIV1sbjvBvbnYA0njFY
2osQlq7q7lXJsveIrZuOH2Oz1iBmG2y+lXzeGTycIv2aUJrewUAf3943Ibse1tztZAIHDskeHVBq
gNxU7Udh9dzhE6RSoAsq5Rk90k4W+20+uK+a4PGdWrNFT/qjn8OtM6xXjCvJp/oRfAobR8NVvmMW
Wtsnt7jy3DeCnzg/ujPxjCCBxDYzPvZpE7naXvo3FgvwxK7Bjm87GVXAjP8xrKPki9DmuQ0qrnBL
kpuL+/6grJAFfONy5LEuvuY06bECr/4hpafTKrkAwoL0ZPnts5AV6BWEHMLLODQiZ6Sqkk1yN3rx
oWzYCv6j2nF3nw7gP7CZ14TRN98d/LBmfnJy4m78T3ol4iZBZ66pTHdVV6ffa5RtnVFearEWfUxL
ZQOl7Fq7j5KyIPTeJZe53d1u93i41QB9A9XKFmFLv2yPaJmCdiE5dYkKwEzXnsTSZVhP2O9nNQSb
DtGZVoyEGoRyG9YcdrGaNQpL20E1mYC9MdbVqlcZIAl8vbWTQycOC4Y306N3hANStuHAwZB+QX1g
Dw3Bk3xNbsWYPKW3HNRlImYzNmJd3+YIZjk5vqp8Xf9DC4otIn0a1rlguzl7tUYP+BEytRtvkhW2
ZxMwwD6y26WEoROTrm60NHjKUaWVyt/01hKqre52t0Pv8jRbJ9cN/tlMg/TKpZHLlnFrK8QwP6Kd
sXd+JbuWzq/E9SCkKUoqlZyupe0VqDUwYVBOoOLophJCeghEpLaJVxr01Y7vS70vVx0WKDOtIIuu
690tTdB5u+k3A63fZl/eGedj8ZLIdNpGvges5Yr+mzcELb3mz4kW4qQMphx6sJiC763pSkzk6s3k
H/KW5JQISk7KY0S87YhVuiyxizDf6Q0wcjb9z7hSdiKvX4HV4Ws/z1KUqgV70dX9dGkzEXnUXYNj
1838G0SiO0KEC9pzshqVjLk/bp2w9LxV8pym9oGsHTVSjzU4XKAavx4HfY7EzXSic/wub9daoKW1
k+rqaXIoFh2HCcb6jV4ULuf9ilnWWkgYk0jqgwzLQGYmq6/DqTVCZxCbRaxvfY3GQOaNCpOqez9M
w8XKVprZsFxZFGlbmT45FMh4/dEr1A19qukpvcJndkXOp93V/T3HifkHZ3uZo+KhJv+YCo+RRR2y
2TdJEI6f5CLmLHn3JAjXmBDlDiJpv7fivQD3yLkaq4lmoICwzm3FW1NJ0miItho4y33BN7dNlN1P
CKtmFwsnwzfk4+9MHYnrGhmL1NNU6kGDlhjcAZcl7KPkr9CvUzAQDheTESitxTJtiWwXSL+8c1Za
3MHxOYJeTRNQpB+c6yZGahNSbpDLxqMBviCZnYaFlyemWS+ko172cwewwNF3LwrLTcj8P6W5jyD6
mW26z+LL2uvoe0WFdcjuKEeSp6TH6frcoTXKJf+1b6Tlit3F/R3M2zeRX+nnh274IwR9x/s/3Dkg
T6FhevtP4hJydnoOdqdMQxTCMMRqljJOj+VtNhsFFJU8eftAqEnxhw6ws4OQvq2RGl5wVX5agC0n
Ern17df7LwbhmcQeHXe5ahlI4Sa7vhhSQxUz0Z7dAvlMqq5nveWl0VSWrgFtd0Keeh0cyJC4HZzE
ZO9yMTFyZQ36K3jpA8uWzNd+GFC7gEtRwXOHTgTctctyoDI+AjQEUYWhedoq6/IQw+yvGZaEZQs9
mFdN+S69fAQ6WiPO5NUJNLSVCZWGBDA42LjzDE2IS5hlicDnqHpERmtoK+LH+babVsO4milv2rR3
fLlLDvpUCIwwEaDRSCoFqNHLIo0gYbsp0fDAIByS0jNER+biZl4mAYAuCfY/P+FtPh3+hHoM5/P+
Tf7XjDlJN4aPWktS66JGzZ2gthT0otuV7d6GlHqWBWGHGZQ/1bSDx7FRBVaVLCvB+JBl6xZ88+Au
syPjPZYefQLHyne5ESkQQ58FnE/EcTHT5IJSJ1Dgoh36FNzNk+wUBT7RzXmldE/FG0uRI0RjAxov
xv7SdnXVQ7R2nKdCRP1LPgh0WJASUo1cC80bENIpGIDwiT84c8/EqUCJiBHRtMrNu3SGvTrQx8o8
xPfQxTJoUiJhRE+1ZgYClZzuWQM1pd565r+R4VJAXyFDHGMjwis1Ue7OmHm2iEDqqc4Pq1jBvnQT
U4XsS6PwV8mbp4RDD71NJCctPDeDd5r822Sgt6J4Ac89HJ6bAV2mOf9SsuWqGhQE9LmRC/Q8LrnQ
w9lNd8CCTaOE+f7vBsrq1No8Lm3U0bG8kQZFj27yrQkRIGVBRFmjkKTiRMkBLySPvUZiYZZd34f7
hhksmQxQ6IMFSy//s2Qse2792TlTP2JYhPHwFJAVBeZyESPHbVhOChEylQo1XSddQEvIG03tt425
sHJGiN6b/p3rmxsWEIUPo1VG+AIP9kCIBI3tabMVpeM+iauX/anLdrcj1JK/bK/oqhwabMCLAeku
8G7Q2pCW190m0gEQdhv7KisQzbmN9xbhIJzbxbPHQFT5qkUpZu2PmJGuU8LUb8rq6jVy3Jx6Qkds
JwON7BvkWDeuM7gyk2+Z/7mnbI2eZQYnZDqqy+N6/hvc8O+heNPIBPVX1uDwyFYBXPWtYsgumgwO
i+K7Q15xaSnsi4mXN4f9yObJRMW2QiQ3TOigSTj9f+elGeNac+2Llt1ZeUfn6pUsNMkLYddn8pvQ
U+Eeqf2NSl/yJhQvTOF4p1d2Pd3YHlE/NVjD/+nJLMfprgSnbOc5/CPP0S98bByJGKffactY9wSS
zXWTHlXcM3IHuTTToTsDUp5/IqbLZuUjnLc3hCNO2Ca6xV6qjXLKlOB+MdifteUUFRYjJXzS+gqS
EntppbhwaEFomwMSvQO5kaT8cerYDmyi4KV0tzWuZLFHn7Mc9RHE5WcfxYY8zHi9kLpjHYT/eajY
1hDWeG42ysSPvasaj3K3lOmQ5hO85Gpj6yy+t3C/uGdI3UW8CUb2zLo7Hb1+RsgVqfJBsXoJbVQh
w3ufaeJlqlG8yNtERdMNNYBx9c5yKZZmte6VKCJkRli8DtZv7SYZew5hl7R5jdy+rhoUlBPpaflo
f1OsN+ifIhL1ZdlCrqinvzCkGr46Q4Nm+fneJyXVmlfqXs4aF/eOGXPnWpouDNnW2jZO1He7i02Q
vRBHx6F6+bIve8Bgz3BnsDfxv4nefT4xhYo2YET7RjO7E20WxejMrJz7gNvr/d9Ovmc2RvgkvUD+
salb7hIgYL7d9hF/zd9CJc467iN2FB3SBQ/7LzUU1iR17TLBXAoJ9gf6MAeQz+XLaasxIG78/K9E
OIG2nq1QV6NCNirSyK66IyGKqxI7B1/b4YvDLROzF/wL11Af0JUrqRwycrVToOnh7K6TY4/QigFL
rIMFJcmMyPqIEQvfgfKjoMcPAWeMT/pk3ncsfWj44LI/TJYdnJzFK2k5qIfMDBoFfqCUmFwplhgj
IpTCwA2FpmL7Z0TPsVY33CuGFL3OiSP5bfA7ciIzG3AQawMofEw7n113r50NMAFJUwX4wDIN4YyB
uUQr9665WTGSNI2LQfjoD626XkhTSPpj8qQ5XywWn+aggq/Uzz8xckqY1ww0ODpPdp+xXa3u73sH
8tFVhELxBPysIj2KNanFJSiL8zcHFd3bmX0yE2N4EcyAHec2tSVaQLazvyN0Ph/9bihzRJDdYeSP
QoVa3+k5dIJqZhrokBf4OhcU1S9XKYp98Xyko8Dp0DJ32lW32m02q3PLmowvR+5REoyLpqpXcSiC
InSMmguGs5fmO6p1cyiHz7/Brc927+Uw04TcZnrKYUBKqho+p+LJsto00i007w1Kw0qO2dhbXWmg
2YPlunw8A1iPyVfdSOjsLwOujiSE7JRAl8gfyMWOZImcfx+KtkghUQ8NFWgyrIbm6PLEyShh5idM
4NBbFSQa8a2iFRNu9vYxDHXG1M/hYowHaXbci50z/PJ1SkNZ9c2+ad6Rw1IzGSKh8hkbWvJTFTr5
AlwDRwXBM24SKxEUP1C4KgZ+tGEyCQBbyuE5SZ4kNNU7t+QKiBFNEX4+9DuVGzCdh8SFZOLP9NYj
sMHTnSTWsXIkh5IODlwZ6+Xmg5Cik/r+9llxbA1wEZEFhgun689YD55kal8OgL1lMxausNCo2TEY
dTrQMx0FMt8CKZR5n74ElbzpOv8TD4hY2og8x6wZL+TrsLL6ErpQb71Ru4AGNl5+IXheXme8PWc9
XwdEuRg/aPTxkCz25X6UwV10g9dV3oHKGT5yNIcm3ov7GZwekdhkGQ0yGBF90ERFcxUDQCFXRO+8
SscaRjIMaGzKIovRfEHM5vg4Bh8qz1YmDzuOBU1xtABW4tId0ZuaCpMq5L74Qn7h5SAY4XYnDtk5
Wxyw3adOaT3LTWKNcaDUacgPm0jp9Xsqhp6Ik8l1aqkq1KWhqw+aI0amfxc1kwff1cmMH1S25Mb+
AX4DarHg/bMFkH7Mm6jssd/p4oIRmi5Q7YeR7d09sNie7nbI3hK/n1ax387TtxLYai2fRKY4Pfvx
2zom+u6kP3h4iaAEBnn/kBz+r57qRG3mdnNZwoSrvDgsb8SspDJt2U5zTLT0BoUNCKRELVpcpKQR
PAd8xoQeKG3z5fF8V3io4130L98Z0Z74azPnnlmYLkkcaXlY/2X0XHkCmsf1YpK2H8g6HT6GAj/s
WRqkqB22L14WVxpsH4In5MONYNX/HilLD4n9iFS64QysQaoHgba9joUhAqCgh9SVYNd3hmyaxMok
Pf6x/gWqzlo+jaGYgJKqIxGgavtfoAnqPO/MVUBztRXp6lG8c4vHgrV02B2aamGJ1vd4dksXP20k
dY16TeQnqK7XcwuwfvAdWbFGNNnR5Vq5rtz1VRYC3THwKTM1NJKvCnHeFQPrzTv0RN4rClNAETVU
oTafSZr7mLDKxCxHxZR+g6fkRXR6AeTM571LEOB4cEnV1SrQTjKI+92D6gvW94DR8wxYgL2XGOap
sJBhHD2R+7yOXouU+i/4rPEmWfqP3fiw8lSB083PfmQ0cVChaTe+EXEPAWxnB6Ynn4T4m1ezf5UU
pjzbBmd3sqHtUIzWzSXxD8tDhcNOCgvNJAi7c5FJo6chYno0x0RX62b5w7afa81e6kAoa0kXy7/U
2h5DLAMbUN4IQ2RrwzbBL3HUV3cOr2YKEvBe4DnNywl87+sNvlRFdfer/7YjN+0kYWCdKOlapZW9
28pKZeW6P6cFMiYj29RW4ab+JEJWfgGYLgNQWqE5zOtZ/eDhY+EOKaP9zCZiooZohBUGZ4Qg44kB
uNVonqeHEpljG+sdAZhfnGPo+Ru/7V0tkWY4ghN+MTkKgLUABgDJ3hnat7CP5LeKUtoJAl2wLl+E
AODSL3gi2KPRid+X6Sbe1fRaVSzzXrXotptFfWUTa8ouLK3+lWs4D9kRrU3IE5zaMl9Hst5bOz51
BtK/o0OXI14cJ4zxxRoCVgWbjKIny+eoE7qpnB/ieGNsiRNjtnYh94jV8xtRu6SQLSthWUxBPrxG
jgv4Q8zwyzn/usM4u786zUOt9lrhiZ4VgPrCKTx1UCoQJ7aG/8GPRyUtbxKJOYAOyabJ3un/o5Hp
6yzfDhKzKYey29vb9NrPcbWOsvMcBQo+fkB8KetEaI8rOBwOldqHsSOu/whlxszHip5wujoVVSoA
fRQv+9Ep2PZI/n4qu3rw3pX6BFvLEx+uwNB8n4m3q1AcLiz+nyW1zKb59lxjCoDHnjT8s8OLeqXX
h8mamFlFF1TVy2Mbj89v/6Gu11XBM8os9WkV+ckVm367GKGzvXipafKqpHs5CvFFHPFZMHBR6PWb
97ugMciDMoeva1Ko0NrUfOylskbN4paADSjlbZkwRPa+ht1ft1p2+hCvUkBj4Mm5noEAi+M4/rnr
lOe4UctI5hCLKoU3MUUVxy3j+odNAgdWIxxQRGRoTtwheyACpuWV0osuw2sv5/eAVCVh1pP6lATP
XmLEohu1mCce08LRq17BleGIMZJFMLNc7NTmlDPhbAWH3qItB23hbdfZAqFDKecuIJ+QBRNFLcEk
u1c/+oXzatPHRK7Q4Tt2ZZJQGPgGwexA5Md+nppPxyYqG+JQttKwF2u3ZTXRR6NHJtQDWqbN11Ux
T2XeFBxF6ytU5Dw3Bi6zv82/KuHx8xcnZku+7SuGbsmW1i6hzcZ/DtgwiwxYxViQi/ykT4USGO0U
MRUb0RyP/vMhEyyL3iDV1iTVhjblUr+eTivP9+QYZslx1mFb3o8lacMhSyeFr4JkSKJtkmg6x4Ck
qspKmHJY+VltaqIwnbdyXEBPKH809YN5t8ZnOfQ11kb51RNMuscfAoih/DqruMge47Vy7N7ujRAv
Kv4jqqSA7EzBbHTluUvhJO0Hca1P7S2B5tZwGm8ySWYaIL8J9CYlWHNbntYprqblZo57rS6RdQ1+
Ykdg9XBH+rtjvZBwAvX/cjdIFjHbh8LLd58tOpI7O9jgPFojpFUkheDtlJJaqhGiZ/QlKz6+TSW1
KXcufssYUPwhVvi3xeCm4DLlljSakgTp7dPkC3hza8Pu3QWI5WqfRekHUYfxYGgdbHD9O65qPksQ
M6HqL/J2E0EmLK2ycD1ezWNP0uC2TPivlwHu24THdAzfAG5KiIfvtLuWOZP9wYGmu6dtjcOCoIqI
SQdlEiyveP1F+LvhmjdNxFrSdzFmaDSHHyFBBcJ7DrgV590/F79HwAkmmgMOxT/z/ibSn1DtzKfz
Vb4OELXHNqHn7YkrqjSpBhEIGeLUNBJolrpYZPtUwstsort6tUjuCYU8FeZHaGclyXLwZ2zVadaD
oRLqo1rCTEOYOkJ3CYub23aunSbewtfXiIYz4EJ1QpmbSbwr5f0M2XnU8S+x4RDqMNuUIAU9ZZ1R
WIyz5LHoBWMkkJDOJyUjfWPMcfSLK+5a46vV+PcNqfTBO1RDuSw9zipNETfYkcI+ptU0Bu+qUhGw
jlYUhUSWnFuI9n8dwcep+ovreQA78SsQ2808IRW43m1jAf7wFpZXK4ILXpqNwq6a2gTRQ07cn5gu
imBytYh6fRmxnPvwuL9Hp14WddAS6zYcsqW9AAqOivljBIhGyNpseXlEdLVoQDMaXZl9ZFmjQPD/
VFJMJc/AZ9862L6c8Zu7Tb5vd1hBm4CMPu5Dkp0H9rUehpV7Kn+4XF3BuQ+Xx1rlRDrW1xWPWoYZ
rqJAg4jsjjiY/uHWBB4kYXxIpzXbc31VlTjPQJauIihkCGcwS2GPDfw9ApoVWQlUkRPmE6SjV7Co
7iJ6Y1aor7OmQCT8habxvWhDtsDoNvdibMzb7r3X2n1d431mOmbD7ohHfPtLO0v43UhvnMxhxKoc
LjN/NL+7PvgwiCq7OtthH5CexICcJXjVF5pK1jKlF15ZlXhML0SA+sw3I6R1BnjOo/2wix8Fz3hL
wHuymcANW3CUcSNhFafFE8EwDT2NmnT7Zb6+AajbrBoCUUftEUHEtXu0ppVCtvYoreE0bFw6b251
tmWR/LjLNWJ8Bc3lZMZJcYMCVXfftqjy9CgLcRLFmMiV9M6ERDcgs19T1/DpWWVqbfCOWIJRouDa
xVyDh9HLbMgoRvOw/FEn2FOcY4GTiGjeqcBcqJ+mCY2F/4uEy531lj2tPn1//fkiRUsz15fAbzDr
Sz3X+0KnTWVu/nFBYvJumEdXvue5QZD87CzvI8PvqekWnJP73pnd56Lig8Rq32TjBQQGk7PgnveY
s5eBwstRVXYjrt5VlmS6oDlfXPaP2SLtumpkVZnnQG9PTNLwDbiU+aWdiCdYkfL6I5c665xREMnD
EO58e4bMQ91UgIscJu1R9Wr1jdUTuEopjbuMvcgIvj9N2DXRbFPyLBIqTtRZoYW0hGsLTjqJKTAV
jPIHBpgM+XRllsB1cErbyT2VhyAtE08HEjvL05+FpxWJI+jDNtGmFpNcC/obnsjVGTgoOX0fNKXd
la64imm013WEmKbVG3lI2a5wQfB1EVMaNQs87lAvSqo9CqTxE1PNhwWIRVLUK5oOhI/Vw3x6e34a
5mPiCpY0wCujvdHsiQX/Gy0RHpX077JjI9fBKcaASMxEY9NYXSxc8+IPup2O5MCcMbMEtFVs6RO4
ynL6Vsr1J6heju8eRHvC1sDoZj28TEs4j3+J6jbiAUWwajHjL+8kSVZn6MoVRvN08WFZ4fq0AnDX
CtRMDAJIVttFBMb3o6BBnjvcH9CZX8FbGg1kmFmWAr5R9Y8Cp3Dp1deduJ16uZHjONSR2PsVvTdF
ztJUJU7VJpm1l+jNa50tqBcXbK5tTg6txTeCtVKXQuR8ACVCv7nN0Re50adYiyplIWdC5hYfjwCH
g2aQhx+XsUd2ZgPSonfEFZZzqqjwd6nBuk2Le5nj9ZUEu4Xv8b+DQrZVbH33BbZze6kTiSJUFSAY
Bx/MvYnj4HSmLDAOCp1x0jUmJvgri1qEiwjU8p2kctTjFm3V77+1YOryy++K0MIMcT1FC8jD4KN+
D8WqNCQNL+1sQjdmUHhzNNP9n4wH52zWECMbCjfMZt3JJsEGWz8m/nLLRq+hbhCA1B/wNmjA0Bab
JZu5gBpCQcTkN9Z60sccWPu1xqZ1oc9FdezDM93DK1fZr0weprRtoZREuIPb2a7CO4pydBH2Rh3S
maMQraoy0/yUN1xl9zDNI9CvQdNyQY8vwlB0UjopddF11wZKmTJu4pB2kAYqjgnA0uC+9lBeg5Bf
KYGzT8o8wSWRiMZFepJZkXOPMa6DeSHaCnPSoJgYthayPuVAS67qpsNjIjPq76RO46WFt3V+D8Wh
broGoTyl8fm+gyb3xi1wYPN/AKRJdbX/sMHW9OJAJuC9OxXD3x/VpTEj3291tHhUj7yFfrK7d7hB
iVYldtDLm1ZTQrEGVHK47shNt8cUoVLq9jdmkyOQzEjw9XXIPjWDKQAV8jXLyB4zqtb6jCKDiVcn
sYp/sTIN/l+ydNNk2ubH1T9+eOaUEEQUpYgKJWSRRlI+R1e/2bxbnDIGxZONNqWvVHjvu5iUU4kB
CMvHKjAFVqes9K4hHTshaHvzdlhkFLCWYggyvDWK/XEgi5vWGYRHRAZ9oUCNlsWjojCHloYz4j8h
4/VWutscQhhLseIAvD21sGVBKTvUNqyJgKeKgaRXngQD3xyYbvaYZS1YVv9ejg4zgvNmpwGuUtnr
wGoJMpCFK3jWtrPh6+bQqB3BSiEQDhqIVrWvbUYEeNx08UnRAVdpd1jLuh+34uUzSnoN4DXdxqxm
uuJTd8qPRDK2Gs3LmrVXm91kbZVS+Q04rWZN3XQg06Hgkyc06qELwq2DJa5FXIl3VDg9PAw2UdgF
iOHpYDtkz/mhhPlgixmxDVmivKHf1bF+1FZlhZgq3y4RixRJUu2x0gtspjdlb2SpmZ4d4STic7j5
1ummoVTjgFx7wOIOn52/LGB4jFUAJNY2uU1HLHvqHxbagqUiEj/F1QbZuXvyNoVei+VQ60L1ZPXu
yHiOo9D9tGqmX8TiBgchKaDTVM4T9mImFlA0Au5OCJIk67li8xGRDaUoeMmjG5GEKtOGbjXbLxfB
4cXMFNgC/+h90crn/GLzn8kLQ0DGgtndVgVFCtay2DUFg73gEFsAehB8S2GRVepi5KkbzhZ09Bhk
dynP7Bx5R56Egc2ficwpD+eJ8fH24lONTcsFIxj5MiebpMjz8P8NENPetok66+lEIPjFRztUVfI7
UhzQgHZ4vTQ2qz6MeF0dCVyayOFEg2lFr15jP6xqIk51pWr4cLFgM89fJHo4MtLi+JCur+I4BMLv
e6aSPEdIslGn9y9xh24TgwNTwsh4xoCMSxQHoizvwxsOHr3zUnJrFB1NxD75WFWjKZkmETuDsenM
vLyaCrD9TZICFb5DMPXriMyLh2D1kHEiDOn9MnCUGOUWxED5iZm90BSx7Jp3cNNLlqu+ykjcALk6
EMFikO+cNuUvIJFy1IKXyDvoL6JYR3TD53WfnqfAxBMIBPZWM8dRX6c+SC8YHcqGKQOYRJs5zk5u
76WsIL6XwR3+i6yb84AcX3k/NROcakDIzX9U92c53D8kNmrCIo5tjmvy86q5gw96OW0GnhXHPB+k
8xi0O5PxxSi/epZoEgn0yElNGNMt0IJodjuQc62dR/mjArQPfaMJx5F3CivYHmnNPBZSxAs1ENes
M+BjIPO9ab2Te3sqi1k/bYU9S33HpdztZMURyXnIqeQdkeMHPxBQa6wZ3IxJqc+1mg4/fOctNeE3
Z9pWfeaNO0rpkzOPkSILNUEDrcSj/i7k61ahPskRUaBCd3CASiiIc+F9kfw7HQ72aNA/WsCvm5lS
pLVYEf/NW2Z5ddjNORtsQ7MLgsv7PqFZMDkJRDN01ihS6EY+LVImrpyMi7+VZWtxRmJn7D7Gdc3o
1NNrKIpbVuv2vzrowjz0Jy79HC5PjTHflQ==
`protect end_protected
