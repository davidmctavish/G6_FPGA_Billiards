`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k+6IMpCVIsbHCsPocQnhhF0IyL8U0R97qdHXUhgCV05bQFu3XbiMu6ABtuEDvV7BoznAvRJfhi+2
BLxeKCyDCQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
flIlMnvDeIStt6M50LIWXRQ5P45UCA9ePelHHixC+rPVFCDkVMJF1zGxRSCffHXH6Mazud8XoWzp
SMY3EmE2LfD0HdCYwIAVccd5WQSwtFG+LGe95ULY47W1/3aH0Rp8mm9mG3l9CJBzWi7HouvFiGoW
FT7TR2AKsfCQPPclFNw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kzdqmH4k5Y2x0rj5G4rZgpiHh5nTxoFetMGqdX8ksGzHVrFiWYqA+W3kau1id2Gosfp+Fij4CuXr
2+rKue6epGb5dMdjqWzbrY6oVWGWw+ouPTBsi7g0TSxYQiiJGVtsN50NRutvkthOZmmcJycbLMqO
weaY9uwrfYE0lTF1KYNLyODutPZstguswmSEVD7L8aXUaCfp41D1lz5ksQ4MfHa5oRzXUvrXV00t
O98fshGTMXcx30wAhW1tIdypv7EsW+FmzRhcKm6ZG0xPGkULZa1zpZv8yq6pPQysBPlqkg2q+Cyl
pd/1CFGIcr+gvZu/uUXADhfXVl6dNqNkU0QSWw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a4Wwj36rylSjvfx0JgLSOY2zeyblKZFZQy3Mv3iZ82f11AJKCMLlmVlm6nkqSJMpR1PCHFSFjoPd
OGToereSXqggKTFFY8RBId68LLj1Bgj8ijSb8N8GrfwtAgy0Gi+AHgoi2JHlk/1/LEidnHblK8vY
/jBOptXxkr4MMkFShH4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fzk096kLdTDp/n8af8GXEaeVYpDMcn5NSVNsMS8QV1aRODuexqZn8xGBOvNX+IFW1e+47+PRy8zm
z7/weMdiQIvbpg5HsA4f/vczEXav9yTwXuDazrElzc+o1C8zSUM5bfmJWbVOgvUoJQ7xAXmuxIe3
4hdJv54rHNzAmU36j/rtR2j9yksViur9xTdbYAQiWwxd4Ni/lShSwL8r3YFd2OKShRXSJO/23GEY
EAe8I3mHOWW38QVXZAMJrdXmpDdCvjnEui3Sxnryc6js/0bB3V2g3QfT/8bB4nmPY3CeL/TvxWjL
Jhuo6grHJlCYpVOXJzx4SimCQ/KOC1a6fSebpg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7808)
`protect data_block
wzcPydQErYGpNJrlDOJIag+amcZU0936d+8cZduVL+aQCk6QTN6drB6ag87RSUixQn0Oy4s9vZbo
Sd2iRY89HQ/eGszVcWNxQnA3h+OuzVq3oatra7h16OFCHnqq/1b2EZWf1a6qCgjgDAgiOUD+wGzh
D2MrmrBP7igshGHtntbwTzCoC41Vvq1lKYkDfDIKe9XDMAjpeKbUtDmsQezwzw1EWTTl5Ey9gDWA
t3a3pHvt9H78iIzieE0FlvEYwij5GWGy0mTJH0VL2QWQo6DF/ESBuJtoj71fZHfOnKcmaunjfoUB
DzSg9Re9zjBOOJmhplfX1Lv2s7g5eGvxcoTiGX2XnmWFa56SQJKYtBvuJ8KK2BT7JB9hKlFK0iZP
Zjb2B/W8mc8igIk/YOD7sLZ1PlX4ynvjn3Ne97ypaUiHZQwpR3onFxn8HPAojTGavMV/Couq0/dx
QdMPlUxQBitN9+WAi84o9D+JPEuiClllXPPUP6VsPidZ6WlIrV3x9Q9ZFupwest4H1lrZD2gisQt
meUkaCGAOGd68/CN0hplYj5G/xWJ7PDVQWyj4/Isk2iVazcE2MR8GB4qNsoHQg17P/Qu0opp4kkb
NkElyKHmHlmVA2Th7XmzI58miur4X9hs0MLezRqId0xKxHP6uovjgo2iNiEFP4+bVMdKT3rO+j36
0PwPZDbbU+dpeA2B8XU8qMlR1YPObsRpK0TqwNKihPX8An+nSab0B5vmC5BJTxL4QxaJjLmaTcY+
qI1V8+K1Jl/4bfXV9EpHeitBSULDU08vN5lBwFijugJF0lVhlbBaq91J+tgepmfAVAnZubRn+YJU
xvHlCbwxnjknCytfr11eJEefumpYHzkNQjMBLz6fuAlcYMD92+4ml6YnbRrzNvZ6pcUuwE0IQx6s
hXQU7sM9mMDiqvbuXcrlinuri+/q49k5AYFVBT71/LRaCgKibsy2AzjpsMbGLds1bbe+s8ck8lLG
+hiMJHWSr/LGMtKwE8yny3sNBNshSy/T9U44dTL8s4crGAR0YaJXp0nZ+BI6/CoKVQ/+yGu65bV8
otetNqnLXhmFvrf5o0IhVrgz0sud9j5PJRDRXos1zp3G91EB2EyLbFZbl8AvR558lpRhcBYQ+nvk
LiVVtUjRcE6JzDu/lupNbKFc3T5hekwfjGzd83P3ZdNWXyPQfSguVTQ8at/yS4X2gnsOIIetHbG1
DsNEKE/yL8dKmQRujUxADlVSWUlgVswFAZkbUCZLK2fR6iHypKNk3YcANppDQ6EyFau+qz5t4imZ
KEtdbSIfbIufgxvU9LO43cLgeTBLk2ne4C/AUR/uCp1SKv40ha/7JTyWFP85wI8zv3u36ZT7vupe
1jP94M9nLT5WmrHFvmBI6k+0aP5WffD0BzeSnjzC/GXfAlkrkL6cWKuP9cOWECFN8GkE2TVI5i4Y
TMPRnR1u0dIWREn9zFA57FpYABwtgVrEl/haVAgdPljEbVtV3+34eeQi9hanbaHYh7RIgGBcRdLF
bcCjDOPAWML6UhgAjQSgq9obDA8OxZlMJ/MVLkFS2r8axmI7aIQbWXL0nA1et3bo+DIC0Ag3ttgi
Ny7Ifb6BonpX1mG0g2FcM+mF8CRlYNKMRdGQTqEJX2X/+IEBPKZPaowBhEgqkGMoiNJTMntMf7ak
w73O708STYkTbNAQql9eJ0dNfH9MEFDH/GlfBTxDr2j/cnzeoWEpx2qixJF0JsghjVI3+rM/NiVB
pN8u/WzBa8/EiJUOgDoRX8IZ0ipZDUaIRbtDOp7VBwjY660tPa8ipF3Ie2I0WKK0W+/MHyoXO041
Nkisf1Ym/an0bTz3OXIudaIfXGe/Zf39A6XKPqoezb/XgZsT7XpaRb83EMJ9YhX4Mmyvh4Bm9uLe
OUn9gFugQJsTSC5wbYsOUb87+Tv9U9gNxPr5L3EhIbMbL35/jm6GU60R8oBOkTdZRdUEQW6tTZ+G
MtEG5x3j1YLIC8PJeO25RR1biaCcuedaib37i1P7oFf2yged+PrU5K4j1CXmdiVHjeN6waNB15l7
Z8FYn5XhJzrmB0vPGBdjhad3qqDFfeGqCkf4zUk8zA7gMevvXDeoclobDEaihQCJLcy3S/YBxNiL
XDh8enIS4WLnVMtdr+eNVyqUwtSR+2Wn1aOjBs0y1zUbNvxUOlQyFXnyPTQNIMoFXC4PcHrqjf3l
OGpKZwgs/SVW+quWSLQ143wgmaz1UY9YZIFEXyIb+GosflgCtiKNWF71ubQ0T2O4sLuBfQs0OGnt
iS0T9Q1+0VLeTQAAth28TMXMaaNl/6gGjFuM2eZueAdVzdFcqPX1kqTlxw0nonsxwK+9NWRR/rBd
d8peUcnUUHgek9IYYhMw69gokj+1iaRTSTnIgY2xarLytvF5g8g70jLvfR7IJ3g4v+Eg0+C2R6IZ
TigeqrMJIJCSamzoxwKP/2DTTmUo6YfVnFEjUxt5A50eMls5SH4ZmIH1t00Mx4cmOwHk0TmgtzII
wZYx1q58J3GLp8FUsHbDoS09SvXp/YhS6R15SyZmu96LoB9poxLSozGogitBgci6oZkgJkVoYA6X
gcHjvZPiooFzvG4ABvOD8tyO7SYhgCDV31Oky8C1aPbtGODvGluZLORzjxuERbB3HG0sXA+z50L5
y9JzjNp10Y9E9caPy0WVmYmO353QJXaLM8LJ/UZqxr/G7YQN4DRQYoluOR37OtwMfxdfjdPakyDq
mYigD5mwds3Jw3bpVSoCILPQufAN5h6vzq1K0Of08cwcoIrLz3LByUJGCLyq9mHuo0Ayeq2MLPqP
3IrekAa24s5VPEwNVpa36sb7h2qFjif+6PZPwyeZlzRjMFyS2x5aaHYlRb9E+jaYV2xXg9/zChBj
6nVCngZ857+vZ5f2HAi6a6C+Cg2bN/EODHSLKdPuXDne+r+bvG1+vCktN2vqVeLvxA1HfY1dTIei
bm+82HLTbv6zKvtHFnv0oCBFZZ2K3EL+jyM71ZEB0bm2bkH8jLX3hk+t/cClz7n0cTfqMiCTO7Tv
XYIo/ZyUGY1lgrekGU0uYNA1g4Aqrc7BO+4/6syfoOocVtnfRPdEY6Sz1CtttOceb69ZTpj0YGKF
90jY1/Jp7N3QziFe29SCuBHjXoPN6UftKe3rJKhlt/I1l05bUTWaalqOcLphU+fwEsdXlO2RG/Bg
j/Twk4EwvW+DjF8LaHbwnijcLCAwrHDNNvc44MUR6zvFOxcVVxK5aqpKJWPHXlCAsSbMgQ6gXi+2
MKIdFdJx1Ravewa5h8hUK2n1j0nsLmvbfyC2eD1Ob5xO/POK8GnSA25cwIg7lChCCmkjWXj92b7z
VjlNd9ww0QiGrtPI++YIzniGulzyECIJw9tVabJFTagrimEI7QcdGWc3HZYBo0rSiqIsJfca21sn
HHqW9nBysaM3BJY9BQehO+Ba1OWtd69rosFxMHjukBvRPbgtmGEq3fD5v0u/ZClx7oKqJ44XJ/lC
nIHLZvZxSW/NEkUQK1nK9QT6mc3e/vs18nELF7ZXR+j/L5NLRY7BNzJINQLLxNA8H0lpN4NQtDYJ
2N30gA8cLSSCd0v0PjjxYL1DUb6hMSzOCsg7sGDbRQ4qVCcMf4FBVIxV2d0xWsav5oKqS0forFMx
Qgd89i9n4146bwz1izoBoNZBEcl/VMdAIXehpp8/TgmzPCB08CWsi/NfEVGxEvTtFteuk7RvFFGN
qMr7ZvH3qzckw0inislp3m1NLm4bjliFxZty1tHe2lP4cdZMbfeyrejUsbAX8X3mkifKvx4FSd/1
gRDRtQ7MTO5SZwc7zZVbV5MML8iOE+pKJ/btIO7KaPr5s56uV3z9MIMYrZK+a3mtPs+DF2Xsm+Hy
nw/KZD2LIPWRt1DlCl3/ajXUcAcefiNNQWJ8L77zeqstWxiR7sxcFNSzXChGLd09S9JQ9Dd3dciG
KzvBOTjDidvBAhBg5ezoHTtc5UZejDUqOXTqIh0bZSUEevYQjxzb13uF6vHZXNNqyGSgFicbGS8L
674A7fGHfIOO/0gw/bpftldk9yZBxD8ZHiqU/2gA3YcyxIwtF1Dg1VVTpxdezKkOnfigAPzzxjBw
WB6DdETD//G9NvjwsLSohP7vAEqNVZI/b1r/Gn4RFBiuTqq5oeGVFt4T2fGWUIdJM3BtB+1+u/P+
nRT808sV+2PapwF3gpsuIATnIyX3XUPqvl7JKs1z2sY/SNu2rkMvDSdZgdWJhYa1hkeREl+dtb7E
DIBdFp5VU9SlDSKV+lsS2p4syJoOPvWWghdaN5d2NPfuxwP32EVHq6p5hHv5vOkqk3nVh8XB0F18
eO8TKeEW9mJ96/VDeQdL5oO0mrewjCDSsRdYDUpUOht+JZydSu275yVDBNGt2EAz+BUCtRvG2b0W
JYWupB/ZFEjavj6DWLg/kF/lIIYejM53c7C7DJ0lzJl68jeT/gxhyG/9fCdWnBQs8G9fGhhV0W3l
m9OFPgI0Qpu1ndFlvj/tpAiSWnkIYUe4qw50PoFKpxtKGD4x7cDIXgl7zR6yeLWvq7lMRweK/8As
RZgK+q+ONG0HlMD/TOVNvKz5yIopqUgsy/IWC3WWI4RL6n1qn2DlNP/GKL2aKxcffRXU4kI7oqp/
iaes/FS2/n7QWkJzunlSUQVyWrZwdW0OjUny9oV28tWqx0vlP75Q7CeHpCPlwxpkGgGF6i6F7VTs
mIy80YGZhx4mFVEqNEuu/b+EoXFg3fn575GcsRqOX0LLOkKtCXHxuQOb3XgDWANdM+FF0KGag838
Y83Q9CGxZ+NN/mggwbtmC+cbRsobsipK0J/MhOiD5YBeNo2ce07XFxhW7d1FK2hKW1l+5RonzYkE
ycnZeOvV3uKsLWd4nJUcGdSRPgQgVgnYd1yXYaVV2lJpsMSWY59pFTBBD4E0Wqqox/fXAlg0hU+7
ttQ2dmmBgHARW5kw+eXDPXV8+yqWJ+OmtCJ375JxaF00JDt9YIge7k1PgavcXN8nEPnsyq0a6dsZ
f9XFpYRK7/hN3NZc0m7/emHbvqxZdZIH3U7D+kXQELyKJqC8xEkcX2gj2DoW/UBH38i5aIXa6N12
C7NgnSvpTjLfGw0Oq5BO6K6mJ75YhS6eDdrVw/zLs072+H0/V4WrQbrhf0Byvk1unbmh85Y0TBnp
6NyXI3hhc7lp+RO2nLF4JC5w8ZC/6liWOwApt7eHtdh0/EM8qbRVH7sVeWnTtHFwiaDdnMdzCY4Q
F12bIhg63BTqcDsMcrbWbY8T6O8gQzJDMf64IWFxsN2Kte2C8p/IenWoJiGJbvhGP5YGaa8GBmzS
uWv6fHOU9P++9SNr/MMW3/u3H5aNE0rJi47SzLp/2sX9gZT3TYDa2/cRlkckmE5gjDplYN04whfm
89y4jlLHETsTCH9a6231QLgIAXhBCZ0jA/ibN1th6FXdQctLTjJWMqCYcyb38uTMmCbaGgbYIg1x
Z1GmCB/igg96vpD+ALxRo/X32xIyZxIxpC55Rdv2YAScfPJ9qs/6/gvxAL5SPwP6iVFJc3ilOH1d
nF964Xajtl5gWkNbM00qClFqRZwvULIAANbx0qxMHZNNPDe148CNpKO7YzaC9kA+kC0Owc/V+Wi5
XRjqsAH3rh5yCxkBTDVfp+38jYK02Bl2uzMqN7G4LPnDhRJO25TtPUpGnd3mjAfulA+oM/QilI8h
C5j6so+3H1e+C5CM0QG84o6sDLbSJtYl+cfyDRyikZyay/3I7iVCQ3LlXTC/NL5Oz20CCdIrlWIl
1qAIrhzN7u2D3aorF3fKPZa8NZlAy8cq96B+Ijn49JtYK1auKL34Ofj+ZARXadwPbP3eNgWMPhyB
UDHLGASKoKQ0JUrzH/erR14wNdubSjSdjUOFLb3XMrDnInqc/7NhXjuJ81oNdMcQcCn6/kPsMhuz
T9eATXguiOSR3wL6oPwoqi6PVg9xIKMkk2sz/vUwhgInR7z1VAATX1uI46CLLjI0H28Z5wcySqgN
VibclK8sFOG5WZ6iL4lFfGFqVGycGEhFAPugpCABBp9/Nq+dga9M/fvSmv8GiN0DBGOXIfnLdbhc
C/o+qHLrec8PvrIFA2HWHU0uvX6FqgKV4LCW1Ck0hqZg5CV1onqP17ubk45w2Nx0fnSxx/qw0E0S
bL0ugG4qLeGRcXsPv9VKLd1ws3vHo2uj27mq0Val3HQH3O+y2TWUMma03IB+NirPoaGCac5bEvyP
VAzBvQ0Dn18yvvQVGppkXWdZWxcipywwzGdlrb/Q2k+Dxe1ov9bB2vyUcaCsddyqSEBOajeO4FP7
yHXA4DAQ2gNYfhOU/HuVtwtyM70FD9L0J+OSeT8As7xPRCiti3JO1eya0v0zgVmLKMw+Ojg1QK22
3SKEmsiUKERMU6V1q+tSTTd5OCJv+38qQMh9rI1nCbRG64gSaEs6sSbSKxJatPciqNvaQwfxAia9
GQa7p0Ueq7EQq6TkIb88JvEKAUbSUj0SZhjRORQzqTT/MnJwnADv4LQOR0XF8nevphBESnhc6hzC
hILViAeuKeATaSODG8JNsgPfqur/zwljWriEN3hXaCMtOvHDWNWA0jg6m2xE4iCF5V9TOcdPvhQY
mG/uggSuP5wdxYHD5+rphUTwl8uKTZFEERprIxNOtnrsbcRzruvLk5w/iMZndz4rk7VPyT+7/DGQ
4T/M3oY9Kib1RgTjUkepZrQQtafabVmJu5HC8Ik2lkbk+uQB6VL0hYN+o7kR6ssvX5qt6PifwSMO
x+JlT5unlFMm+GLVPaV7K0F7UdcJiwjdGmhF9sXnrjnl8XjnS0D9hVTFezAN9S+gNI+cDwdvUP7M
ETa/e3HPsD3TgRPYRY0dQXrEEyTbLA21REtkeVEuRHa/glD2+73wGn1NEMxMc9w0pttVr1gvvH5F
auwU/M2L1Uki8VHOapgu99+D8s8JwgD79yzaaFF+hfaGOT6nlfepHYrsBmVyINpgU5Yyhdeu7tOm
f7VlJZnqOjhHwB4VZVO/jy4P3Pr7JBpf5vG4As6SYknpnzp/K9Jii3ZvoQ4DjRLO6/2+2kCYCaCY
vy9e9HdCGmF//aUzXcksRuQuuLMnZa2k2N6Sd5fBwrGJKlhH7HkgQVtDE9/BPOJmsK16LgCgNTJZ
uaC8bTA/o0JlbilysQv2gOyfzC3aP7XyK3CGPTISd13nqJnb6lOKb1OOYQ4bTMPcCKQJG4xlKDz7
LfHQS56txqyOeSgGk83sbQo0VSn+r/s/NpOa5Q/w7KHxx8G/DFQqZefyqir+6sXcegjJp75hiSxC
AdqY1ZgY1W4Zg+IrPscAPnT/rRevI2hz0WWERLMttNKfeWmLqouHkEk1wJvtPzfMom7EjaRQ7InG
RQr+iVWIEBD1fRWjeoekhxEC1LjrSgh+zIk9uS9nVBLnBbdCSHSszGOqSGjTs3GBug4kQBsbWapp
rHFs4k3eK3VXLO7UV+pVOW2YVveCPeAHKRvRREtuwOCySW2Nkwk8DONk82XXUiOUlqliVBHbp/AG
tqhl+BbzGawoZfdYVXo+IuD0Lng6pILIOKHY+1c2/UnymIawM6bpZW5HBBs6J5tBgcigfv+9Cr9K
ozHmwfaGMyLTVQnTCH60ec0XtMuPDSNMAA/EZ8FX+6IyIK/JQDK6yFvsZBeXyMs6S+yZXfgZZeyE
aLI3GLxU5MRg7tz6kjzTPambu7Uii86DpWOmK91F5RGeR3Gw6AZfCYnZSvOVACemn/1yXOq/LUPu
Y0abdeHy21KswN5hvDUOKnJBfzODHuw+c1QNv12sfAakckq5jEv2nnl73b3zCreVcN/0fQM7TKVS
jV5rZ7HkDvy+JYQ7JfqvjMJyW9p95gnveBczvgUAZbYFZgSJ0dF0l5PMH+B8ZeRVZoocvlgLjXHi
wv7LsBi3Wei3627Ay4/B6rWcK6C2nWCa8Q7GjHFWtZvUi7J5/IbJtjwOk0wWv14aYW2ofHXalilY
jhguX+jHxTCxyRPsZV4fQsKNJ8aEjcCdLbIPSEK508kSbMp1dgB+JCbT10ETVaECwGGnWgAdVbXS
SPO3x4gTldhw3PJnLvgChnTMaq80bc+GHbs79gMdrm7nZzCRzdhapRUhcCWqjhGMDkD3rnnhjZuE
ZLNuKGGAzQjgRCikXyqprru6K69BYIFbVD09NSiCoykOE0MX7ZbHig+91c8/ko/4fHO6u4KVH3Zp
oOaalEwxVqQ+oY14MI/SF1TBr46wwjbWxQbl3WbTV3xP+dclG9OrmwPyhhZDOGRFoC40paoa+uHe
314q9a8555l7be5tu7OooT8pupNZAI3MqNmJt8Q2q6FmQmLSb3s8D/GRSAX3O1cbRac5x4nratzT
mpOUtrRfXBcep3WROVgkZqvqE26C2T9cb6iXBkC3X6N2cV+tRwVrbUBNZl7PEB32QqLspOEzqrLk
AYl8K7k3G7Rp4U6weMdRjzx5mSv2vK4ADqmiN3DOaRoEDdpipJ1rW+gSDlRVxlQNAKoY6mLuMvF1
edasmRgt1VyrSaruii4iQ9A1Dd8DGoE5SQfPkOZIIswHggY/W9Ejyordb8xFNJDvA3znIKekQxE5
B7+A/H14rcApoLD/0717NBBr+Ic8PJGseoMdCKX+DfqiHbaYA7fDzzNRjsJD2k6ckwSORxSNZ+za
YhvEMM7TSu344+sDOBchkAogSDLXGD+58ucJnsMDRGwQQB0Uq0FzqWikKaoSgWl0G+4CbcnwX1iA
304FiTfXYF1vCHrftH4SMigv1ZWYOUcZhchVb3bkUe4F5TiRq3+IEWxiWoV5BmiNvXimbGOC/8N5
OCUOrtkfR1UWh+PYRyKstPPMUO2qPUfkv36JCxOjFDun0wjRRTZ3RgN6zfJXocQHCg3wCGmD0KFf
t3wRVYtZucTDoiAC+xT2LmaU3LSoM2s0HgL23yGhG0d9anv33DPKukd5NLWqhd/TSb0Bs9jViNQM
bMwcTjx5tG7J4a/49jMUmqTIhkoxW9EzD3EXpkq+OpbAI2yyK3uzwHWp9u60y1rIFWGMcROcZ8yC
9DAVVexoEaRaQUjJWrDdxNoEH9j60caHZDrnM5Bh+JKv1coEt+SdNPj7FGCpSrEJH5I7yQDVCbQC
4sVn9xHR5YFD0tO9hkI0HAJriEQRA1He9icf59c89dRgMXxACfBVb2hQuks9WHInFYNdiqBlKXqc
X9x2UddjM8d8TqNrSZGFrSmFeOtqbKnklvSqbk8ccRJV7NRgiEgRhDySWfc2iVwubDfhH7ZCxpj+
fqwYGemUEVOdzseMAiZ2d1K0ClEtars8HM09+DFSCbGMa9lu94mf4J5QQpydaeiVbK7rGqpcycsM
I0j6GDSUfK5azqlVwPatau+mvF90es10ULC49VlEuIs6UZxUceJx6QEKUQIpcrH24ej97ZouXMeo
v6hmWtMW/L0OvOKl+gHgYTy4MnLZhkjr/lhc2Tq7cb6tvalKI9Hh1/DllR8K3jZ/rx0pQfI5K5hr
9JL60fbjZOGV1NjYbPZWgV6q5rxcK+9/kes5Fyu/aVKwSp0kXeAGLNowZTJQho4VgRPLW0Ub1uJX
OD+s3nq7R3bj3/XEu/baRZcvFQygTKynPcfAHK4x4ItHyc2wxJKICIMfLtXOhe9tkd32s9vxzGpc
WnzBuqdRjJUpp+WiZpHp9aF5VPE2Atc9Aq/9R5fdY6ffUUxSmUDhdicmGHAP3o20rYJGNDdUfc/f
nleX1FNFf3tjcfUWhMR5saTNeZ/YI+7lyNHlk3sYqIhux4Vafug7wpVGb9yI3yYPWanwIHSjxGgP
JcDoBrvhDS8AJnAupOsrZ7XpkZbp6M6N06y2tZGbJoYju9FdXnCeAjmAh387s/JREXFcD8NeSwnC
VR923tCWbC8XiVQB+dcDrcIDkVFioFAm1OkqtwENpBzH3f8yaviztMlBFeDODWiHEIROrZ+k8LVB
6q8wX6UMYP6fCBMGUCgA5jl9d916SqSc5G0KBx0Gw2GSfy5WPM80UkZdie+pGphAEuM1LXLKfjC+
wwe1j9cTFZ+kq+BQXOQuyKlr2YUSMZdwPzhcSAae/zN88SQubQA0jYlFNiPgXuS8qhx00JSWbjZA
S2GlRNju8+SgVMdboHXmkaWsBYnck2GnFutHYcpqeoE677DK/qgg8OmRCiK/UWoYoCaIKl/JcCox
17ZH8O9zK77lP1lT5z7OCC4ieYsthy6PVurWnpPlzar4g/etVmftl0IXLVlIPhjM+339yl6KoJhP
K1dufS8OfCG5aJSJaqc8HFkE6NAXVplJQYo5xRSLsyV2dOh4o4Zk4yxz1+iv7X0uhH+qaI49JIZV
0Ord1mEb2GMmJfO/vhjNnIzk9fsPW18/sRot4h+hSbstbihhoqoqbPH5BLumeCBWjHS05ocSkwg=
`protect end_protected
