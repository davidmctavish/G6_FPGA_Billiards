`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EJqZdQq8nVnK5ypj58RK31/jiaVj44lXjMypHi70GZDkUwvdatIx32BwVlbE9cKUjJ40VFcWQyOE
NAQtkW9DHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a2BNmJ0P/KDDphubQfjJh65LQONNGS+nPDI+FEBqVqVh3llYcPm9TEnuAyovIirerrM92px3IQSh
cFSpAPp4u/cd2TJsfsLOrPD9ZnxO7qy+e2JY5FpUi/XAqggR3eAOzMXj3D5VHeXdh19yOQmdTRxs
7IQJAFlwq6g8IYGzFxI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HJfCQzlhZ8q7ejhQ5EFzp0sqg3HtFae77IOdJeWcto54U3E78SpeEDF6pEhwACgUqjZfs9yzpiY1
EUUgScwgIN7Wbwe/7apXbfFWsLRTz8x5L+Yl5SnoyXFwvLOYWAMsORan8OWr23dd+9kfG7yc62pW
BjXmSWx7Wi0O9XlFgED4nL6YYV/M8k6xPyx0GNKFeG1doQNF6Utkl/sAjy9+NglHdDzTmALPsQRU
/DJUOlU3QqBR6nCUQMBlE1kkx7TEFVvhuOJDy0wsNIcbrlyf+PZm0ruu6wGyKsynW4HQx0weUNsK
ODzfMWLQQZMUTvWbLVYZberOAXQxSc+pXIpW9Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
22ja5ZdxCeErOR7hMWKMcmpZ+VKfeNCMU6DxuiFXT/HUT+7i9bqIzlJcz/hQC0EjyB23hZXTNzfm
c92ta8uxwh6+uP8+SBSMnH8ZueZAmLNf/5UV+aaOZAkmdYvLw6D4n5sDpBVVjloTF6tV/N+f8w/S
eAJYzTeQTy5nodOpg38=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bw67Aw1Vod4+yEV0TbTFZJaFDqK8HUTiXKh6QYc64hlfM5XHhrfCdy6yOxSysow3bXzUJqJGp6aw
tAeU/hA19lI2p12pRkyc7GhOjslb1ulgnqKjCqtr9jZL69HHOpRw/lg4xsvirSgCPOrQgZ5ou1ig
NA4Hat4XuLKzqjPgqzY3V1qTaS5VxOOfbavUc9WEeh/84FKAfghw7h1KPrezdYYv7QxJHnIo3IPm
sWfq56b9MNVhEvGehHmES9J4qHGzwAtzm6NNmj9TFZrDAEPLJ3yKCvXPBT441pK5ZYogHF4H18rU
kbxd7ZO/JjAzrLks2cKgQuhcXRvNBt+Vg6W2pQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74576)
`protect data_block
BDJkwKT7+i0ggT/c5enO4549jBinzkMmeYCLn8JCaIUC+BFLiKutNf75P/gZqJHJjylbcwi29Ppf
BoRPwwR6yCFQHaK7RK/tyJSqhrHrQPI0NPsTbFt718YfWa+7TeqaOGSUpzDj8X4fUIaZ0AZ3B/IV
7/TR9OZQoniDDxlFbD6m8VatDqxjUfIWhGeXwM5tCd7dS5U0gh/3yEPB1dtwryFS1mwpql1qkH1e
9LdwcEmdvg+BmV0DlJbPCILrqad9xhwl0RHqTAjf8Qrd/aJhjcCTz5H0kqrMesUAl6OOwWlSLqjI
nhAmzslqVQvJ5AJmHWE90wM/f2d17Mj0RAq7XhphqB3qM8xczw7JWNeeKGN2rN7KU1YqsPsbZ5sl
koEwaB0LX1kBvaxzCKWALvF1GMBq/mGZhmk0fmXBSU6Y//jBVYnwjB972EVPDOF+M04ERX1DIy41
WB9te1mX3OKtL/CRKvr46PJ1Egh+OnEHfg1U5ztlfhIL72c4cLrloBo++b6tOLTQy1uDPlkRVExP
n4jcamVdET2O9E1oPB3WHwLowos81mn/faGzKwSLfM1mQ8eKeMaZHInuavtF7TXhUki9R3bdK1Je
WycfLP0oj+a5HmmTi8NL1mZxnhX/FWtNr3MJyskLhtUA3g+z+toDjuS2fLQ2oyYlwtM2h0dPdRPn
imYSmVFxuZT5ZbFl6ZNg7cBPzbm57eOO6xGLkc20xn1Bus8uRoPQAhs0ib+krovRqaFlqM1mI7Ey
ymqjBI1Cmxe8CSww5RS9Nju/j03eFrGRC3tF5FmWzzUQsUTr9L9LMXwiIvR1VE+hD9/XR7YepGtN
QisrXFrMBTR3y0xnOJBUWqGWLZNTwMRcwcdE7eUnlF9m05Ho153OPr7IqeyeRC5yic5AXLpxNABn
FyfXQl68QyviGhOL7pDocNiXZeO9tD6fabEs2NdEO8P783KXZmgnpmtq5SSn1MfQW32C9yqrru23
CnqAVuoltD3sPjZaTdJxJN/Ay4St/uU07YcxmBOL3nxmiASx0waEjt/ms8Bz5/mWfRYlW+OClrEZ
+JyMy7sec6i531n6dPa4mUd9F/4Sl8lyo+UAfyFOD1fXMuw90RH1NO790kLrDa88IQh9r6uw4hHv
s3EWdMqQUPqFyqIhsE4Iv2HfAHjrcmXDu5f0hZ+WhAmN825ah2HfswcpIFZOsv0gflehS0jh7Vp/
r6JiKY4CPlB/db6KBbOiRbZQ9pDjG7K5Uc9q2W43xA00kzQ+QGIliU6qmwpCYLpfTWHEVJtlDjXI
pP9/TqGm3aXDmjnjzCqO3rcDa+y/koppwAtDQDJLo9Nwdv4WBjmJ3C0kDbrqJUgNgmYKfKOP3PTZ
CMm3s+bxeyyum7XVw7Zw1McZ0UrzKWoJDEGIwniKrvn+P122xAsxhQ64Bpdw8DISCXm06wq53KsI
MAMScBE+LBNzOLHWXaEhcgGC9LeRnmfxEg8RMUoJ/uZIx+AOrLxe6J1WzPTOF3KaXuPCQ4brhWuQ
kXb+bZk7Sy/+05LJwgxPXJd+nAAEkZrYLUvR6TCODUitqL835EIWzC/2fed6oTe3M8yP4WSU3POr
YpZ6sAlbKBEFJEFhxCH2nm/lzQNI14pw3iwzqbtAbSRj/QsrLYFs5u1vHk7Yh1m+NlyvFz+23Vd7
84sCHgKpQ8chs7N01inDLp+0OZ7hlWclTBf6sYTcLR1j76Fi5aaCTof1NUGqYt7tT0jKbHzdlP+5
ZBteEEDMur4YcXSK3PXyJr7ljZ7iifWIRTNy0r4KSsfCkC1kOofkffLYpHiF5qJTkqECwGtRcqv/
eiWMwwIdp6FXkMPDiy5CwHEWCyjZbNmM4qh5MWnWIt4QY3uw8rJAqkPXV3JZmKSMdhpSOnbgm+Vb
RYzooF4cSoCB7TJNz0cbffBP1CycaAt/TQ7cj35zgGFPvc7cqhZ6Rc+rTJro+UI9tH4TYJp3ix+1
Iz1XF4auMIe1+vh4Poo3Iuy72S15Cc3aA2NJHgV0LybXbNAq8TqbJ7FfNCVpCdnfe8PZlFvpLrZC
2M74hFtlop82Lb+MQfeMFzO+e6rS59J5OhduNXcFH8xqY3h2qad83o93MUsn+vmj9rKxSans9nwx
R7JRuaAbxDJOQyV3C9tu86ITxnrvJhxRFntI58oF2pR55AHA5XKYOlLyHW+mPOWAzFDCJui1b2kw
xK8d305fxRm3ZQBYz8AMebSC3K/EGYo59MmxnBTCZDa/NkvPhcC/lgeYmRoRQN1ohLjGtxEdtToh
sFXi6Lc1l4QF2OEmvLa8VCHkXnl2RD3gJoFapKfWTq8jtxbGIGKkrDE2LbiF0AlZtaAyBWxiQKPt
Yk91MKZCDWn28pIjkiJImRn1iWL/p1GYRTPy7m8Y0FF9LO0yHOe8qFekPpVZvViytES+jv2jTO6h
ZO2c0lCIc1QJm9u4tyxJNGPQjwDZd6EpgnEMMc4bmjGaZKlTNSQlM7/iLpp4bURGlW4YNUsxBA6g
Ce+ddLLVcERCgKNA+L3bYY53SMvL9XZzmdMJkWfoTKeJPqjhd821G6ijhF7TKj17Ln/0z2Dge5j6
opcEUlZ3XOpYKaELVR5haYD/c+qDZTlv8KcOf7AOwMKTqjaXP2hoP+zu20MKE+zgIckhZykvtbfI
QskhD/T+SCCJA/whaEr8xsYb/09kQ9sz345lvwHyFN2r6V2JXC7NPVnX9JFY4K0/1SmGfdnzaYDI
mm5+PsVxuS+D3e/uwr5t/lalzqTlFO8/dr2bgBq/I3jKJAAc0P8TOgdUPoIzc02TUrMeqXde+4l3
9Lh8navQepOYWnNh87rJXt4hnoqDmmb9UEsAe82XnpzBvwiUIPNB2NlMqprz6P8F+zGslvtnfe/u
La8UpsYuxWXqKtmnB8wmKm3+4wS2AMzFwEs8utnfDBF9i0v8lvDB8Xj/l+v2ogAlyVxm/9yI6KCz
KS6JKk2H8WbZaU56u8et6G8rJCaNEN2CVtmVf9J5/XDF4iikT/lbEq3+36e2GNQSi4FfP44MVUeJ
XisDkiXOoiPZahsU3xS/jOf/K4kSIYKr1yJxw3Hs8GcdvnVuvyIGLLPh3eUTmDOa5qUvzeKw8gik
4e5NpaqOz0uCP+ti11WrabFInBU5HAeiSRQEVnJKBGe9BiTCZVCN7S8uBuKGBah32I4KHWvW6+vt
ZahsYtjYqlB7a8st2XZ8VNGQjdTuOB8UdU6+nG1g8+dgMHwD9SCza8L0358iOR+AJN8aLPKJX4Bz
2entAXscX9KBYP1+AwhYRAhlOiEZYZfX0RaUYvwVnEFCUYGFZUaBXmNjNAAhg/mYCZiqkYwk20ah
cxfcHw4QKNdma/naxb406ZY3s/iIu6QOR8zlDzQIZTS/Zv301165UgJwjt2h6bV0uHE1YZQJ/+9u
xxUSNOLqcBChM3X4MOagSvEtbrsx4Lqor9ivh3absBFXgZtOB6yVLHU8l+Iy+t561GVk6qUHVo2t
R6DW8atkR01kd/prQTP+64eBtxiAmaInIcxpV0I0qmG1YXVAwmjKC7jHyusjhFLwywYlvNHObziY
Fwns7rZ6F8mQylAgeqNC7xAOZaY2mDvk0c0RExOCVh7VY54DFg+agvvD7TeoHUSBylu2oqK/iLQE
ay1YaeuZ3tNlRonLkMAskml7RTPikGdWefGUztPhsI+jZ5cNklxwhMJTpxXTimnGUr1RO6QNSgol
a9LfJYDyq17MgFtopiMGGY8od78VQoM7MC7Lzg0tl4hFurWP+3Mjjoy3Gr+rXqWnb+6CJM+V5zmQ
ZzrFjuvZIBVQ7IqTbLdgk4rs0+YjR1AK1HuF4nhjc5ZBWCB2X9dWajXxUZhlB66zgwTz/uUbsPFe
FxhNJPDMNdvBkL6PhKRmxCjAuTgBqkY1ONhrmYz35nrOv1S/D4NU+AU1wmIC+NP4r87GTgvCZFp2
U471LZ7Pd3Xve83LoDDVtizPxmbS6AA0rVFwmoozDwZlg6RA717qeqco3YQ8Y2dRcP0FpIC+5Ra9
6xm0cnB8qEfQt78L6eA8bmS7afFV0JswwQLY6rdyEwzgAMuKVD9+5k96Vb3ShR6fudoZk28eMknd
mcTuWoyNvbCvuGww7EHoTXrIFa8wHuVExDlImhXAXZciv+/Ty8A0w5lwwXuiDS/rvX+6sb1HkQcr
QzxDJKBBE5WCNXrX5YUnxpiPol9Z9Xzr2lTXCBQf8yU6vcxA1PRQgG2OdnbXftAXO2OUP801x/Ir
Pp5UOuIqnu/Cdwh8i+OtYG0PFAuWvaDgOF0DX/EDTkkcifXsGPyHI4MlsOOxitkdPzzYRj80Pb0J
BiI47ZC8F33DMVbGZ81ghqq3wsvx9gtp9pcecDYFglPGTEJjV1xIaoWastSpXNMedwBrOnRxdJIi
HOrIRk/M+0bqOpfNWMlXqhRlrFfiwZFIG3vNgBaspJ0jDLLeN9alCqyPJKWhKsupXV3/OnoVFfYJ
SMDyjn864nvaGiM8HIh29P1eOlIs/01W2Gkoh1833d0j4UllwKnA0+e8WhKRGf8gwWhPju+cZ13T
H1LW/NFLl3esSBAV5nquT/G7YZnCSfsH/icUsPK3pH4rZP122iiOb7tW5NjolYMELIMMJYEJ+x5n
QHJZm/YgfJP5DuFc71Ve4EoUdssU9sYJTLYxPc7yjmJquM/DBVR/GgaMfe8OD7B+u7QGYBBXmHcL
g1UEwGx795wc3sdN/jn5C41+0bWjKxbAI2vQQDeJFFY2sWDPX2AW5TpLS1VK3zi6GkrRwujVKDMq
yKDyAEZ9SQ2KXbpqc3jmohsQ1YuEPTh5XNYhOKtGn5BVAgfnCwdLecU2M4Er3BERP2AvQzWMGkCk
xcvv1FgPHfYgZwKh9/MIwc/vgD0CLrcTr0V5bOWHl+3RFy26/gsCfcugtTOlW1cZRspbiPldDC2f
DIbhcTcYNyZa6m8WzvjBTVJV/AHSgL1ESCZJpvYbxQTP1NOWoLvu4AabHkIqcwFONA1q2i4gVs9U
/w3Oz5KlllEbKUQYNcmaln0T+JNTZRa8FK8LL5k3M1T1ngQecEiGCUghRY1iNeG+502FKYPqB/dB
/PKDeCvsbQKlO51UjZlz8cgSMhLxzv3VK1SfbzExxYcriP37SqzBIMqPdpLgkFmxFWAWQQO164XT
wzWsY4zfmqAzj4MZjTdbh64PySoIhnXwfhsoJSRLGNty+sGJ4bbJMefaNE1PC0hG3w94pfztrRXi
Y7h8EkFFqaClJ5VsLsRmPZveo/F5QJjBd78/JlxSsAOr0mKQLJgJ3Nta7tyvXdOrtYF0s1Uf5hPm
xFX7orRGht9/LzNAjiBSH0yQVSPw1Cke3iCvYi7kiDolg5ty4Y+Yj6v0PYSbdwxcCDXzk43gNOym
8mgs0UdeUFa3KDeNY+P4+8xTctD/4EQ9oXiiyaNM7Lx23bMS7ACxX+4x4PRJoQpto4T6OS0jHKDC
s4n5bFoLD79Fa3DpCFE+skLXCSwThUiwIKPAN65aJET1cl95liga8/2rdgokVtLtYiM2+n3kAfQe
g0N9E6hzTiW5zygOtbhHGcoIRn+2RMPE34v9BxdotbuXu+i+13C5FSzzXDoAp8RsWDX1OsFMLycQ
Kz00OSfH5rLY0V4IKGsjnIv2E5/vb3chew/oRdh7a2Q+dy+RpJjiOV45wKuLmjn7Tx4hvKOPzmgL
vlesYU4guafpx2dlt2Pndo9DwzMDpDRiI4qYq//hUfSGhEVP0Y2jaKWrwxz+nZL8Q5k29bqRcBp+
RHX/wHhGdkuUAen1+ZjCTqGZiFbEt2uXNcgsjZQFe5TTnN8XvU3V5OvafjG0FE3r7Xli75GusQfR
XuVkkbYxNG6ZTIxU6Ld8woKe1nshgKHZfFBduxTB1PnBRgbkbtmeZUus1sCokZgLAHgpA1AnRedg
vVYmtNliojw9//l/pXEVQ5xM/aVKlVQP0rKAVlvT85iCvXiU8qZ1MDDhJSek4b79OVN60scXubei
CvfaAUPZty750FRaooIUfXHX8/hM5Ue4FRj3cCuKqp6W0xwh2g752St1MgVgzA4ysfjrXT4UXBOt
4aoY6ZEZxA5PTCyRBocyiBd6jCzSz+NKsAXPH8iglv2BhMR0XWD0HaLUfk+fuGDgP9gNyvSPqt+n
W/cV/SfgPefm8yXGAz+TKkhX3mxb4OU4tlpqwELxIQ5wbF2CEsl31u4r9dqqNYR0HcljisaEi0ce
FWGa42D23LrofIjuYUtCSAXhI3RBdKxuUAc1aV25aknIIocqQ9t8UonJUAkzZkJP37RT1IZBdMEL
qwDFrQq84eu40YKExZz0LLSlV8ScxmAjuBfGIuNibnH1m1AnKoiEU7HfJqJaH8y8CacLQTS1Kskm
FGdgcEKHud7s0z3m/RzwALDn7XvdACTy3GLksYOEdlNi9EadtDcYitHLlFe6oDxXkXTYdKc5ibOG
WeBpnXr4VowL7L6HXIdYvHIkM1pAsEuF4MnyxS+nadUolivx19FEjI2HWS9IhiRjZBNrZ0ZrQsP/
3ZNRyPZXbNU8eB4bj1wSnWwVMDIttrPg9tVSb5CP+nt0VJtBTQ/DCxyQ0iI0OOPxTg9ZASe7zcIH
ohbLACVaEdNn0dCscDmGrBoyYRdZ/i3zW+vMJwh8AhJu5U/DxmVQu1itwqHzAjirj5nSYBmKJRVW
Xffna/vFoLm8/s0qJFRShUD7d2iKo0u2SjSRD1TpqPlI5YPvI6Jp4kaMt+URrlJR9/YH2JNsRq6x
LPMtCwMe03b8FefsgukYYamxONH9ewjJYSIk/fDOW1yjTChJBC4IMvBznHYe2borCB/YM/aBJxtA
5fOF+9HL/iAwsReAa4w3Tyu2XdXknTo6Qqzz3RsPZPXu4w4PTftx7nF/AS93rW9DSw3Un18TtDxI
8bGPL+kvQ0xw2FPWs78CxUWAeB+MpLMdIMtXKQMi+MwqKBvo1/eGbEatDnyDwiZ1lQLQgFFdRKn7
aWPeo9EasIFB3kwkHFS+YkKeRt9JeNRXlUOyFJACn+EZikzER5dVxPcipf2C+pcKKSvmK7Zg/XJ/
UbQtLHHCU2xSSfqdZ4km2ywAi51Kd8sHMpbJfSGnk2ujS3w3Tker8Lnhwh+FhOSvaqLU6X4dd0Lq
D1Vn4HCueEv1VjGm1cJ7pvVsYxbqretjbhZzlnAbXSld52GZe4caXdhrrlFTUFPkzLxB6VGv9KSr
jvh/OKSIpIx+oqoCIWfYRYtu2B9xs77FZ/S3kuGZQ8Yo/R68HOjrOqvL97dQKgKmd4Yo7FEaMeJw
dA0ErPciY8SfQIZIAGg85AAXaO1HggMa4zhHEmsqhXFULxEOnp8USHtHogBSTljUDVFJ8b6I+EiX
e8drnYXzDUGTAciNiz8Qck1T/qL+2OC77Ici6obBtWTFA7C8QYldDYoR1nx0Zpv9DCbyhlAmY15I
CAC/62zJ7nwJejWU9OF6vEteucOLGhHhmU9IJs039fXOVVyWcvagqMj0mWJd672Eh54nqTY7WuWE
MnR3L6GnCWCv5kb2kkSMW6YHEy67E0ZWKpPXeF8Vx/8X4i3oRv14nVLavLDXgiv58Tt9tVTzRmKo
CXGGppEiF6tB+YVVA+ZoRk2R2PJz0U4PeOrLFGgj3/dYLXELuBVFXgMkTKFhmC4H3fJbOo7n+vtM
9UzBkK+hzaQFRRcbiNiY76iUh8mPV2aZKDEeInn1opKfIt06klvVdnhEMOwhzALcf/sJj7jlZ5CQ
mXnypCYMQDioMtPVL1JvDWncMJ75MqyCiC9/rHTQnnxAkiYSyY5IjCH/x14wP7tK1P9eurjOK6Cb
VDNmn79QELN8bRcW4TOMUW4P2KC1UG5+NJt7pfV9f5+B0uAvlo3X9eOmnOn18k0OuJMULfJctbqj
1NGeXfF6JwRpoG/2J0khOwm8cMyxJqyJaRgGp7z8SugFK1qD3dxIFXqWvtUo+Zgp9gbcSbeXf6r5
o8fftKhddyPfv4q4hIaxfX7Yfaw8IliPgkQCe6gHxAzndNUvs/semrNUycRXRkizoblItAZwsmsm
GuTEWllndkStevGuBC6aMES8vBBMUtKgar1RY5e1izCZmJ4V7NqMx85QSnOsjXMwaFZVDZhV+LHJ
ziwtomCX6CiBOAdNmj7TMPq21OKQaOlvWT1PD7q2PfoNfIEpNUGpJz0lVhtszz3pxXonaXom9Lxs
Aooo/uay3kuYB5g8JEsDuKpvtCgg+kGass5ki8KSsq0bcadLs/xumn3F09TiY7/FwS8rUxQYUwt4
rqvBnmI34Qj5dW/YpmqxBn/tMRTsTRusN36OaWkPoE5VqTMDMbqbsTTv/qwxKsEo4RCasSKX392k
85NfrI6Jn2WaLiJpsNKxdW/C2DiXTsQyK9AwTW8B6lP4TT3FHj1SrI2OLKsq3YaGR/u4AdF7Lfbc
8a/lOzlBQ8DlaCFKQSm3kDTbk6fnwIL1ob5Y/BIhTTEfP+NYq+D13WhQ45a4HJhyiRQEFLT/tkP/
J95rhMHJBftomA/jhKAGoZRMdxekLB1kMj0xAsyF4Ip/K0qZkwoBOVYZJU46dY/XWqYQEbJV0M5T
2FQkd+55ZIQi8njAtawe+e7N3fNi6LxGl/aXvQ3WghucOScLC9YZCS0HflAlOqC+lQsNVf/udm08
yY4emEBLgP1JXIFzVj56kqbCg3MqAavAu/XR4PUWNIXBSgJtGMFFRGWQ1QVwNHV6LsESpTVxAJd/
1uqShQtOKgekP8IzaF8ugYfglzxb803odm8NWadaVZLS6hyYEIC0pa1hWB6ornKPdCHv+q5555H3
+gfyKeoVWH9U/4mGy8xB3YRceNe9nQ5Z2TvJAf57Q3drdrMo9Omv1kXAmJLfb6aiNGqkRoQPeVEv
e3dI7yVKqfFcGr30h2hkAyR3yMT4WXuLpew9y6rCro9+XV+09w0l50K3cPdnloTelI6ukmqNA8Ia
glBrsRL/SN7zwZTxMH0CkC7uQHIJ7a7m68vhBmuApziHFNQIvdnipiDgW7r9atEdgeaHykNFND0o
5D5YDc/JGWQ6fpGf7WH5LbsoAlPmEKJvDHTysivvBZhNV/oR9sPYbyYtpVdfTlFOVuDbJlBx7uz9
NnI3SqQPgsUDHaXcqqykgxNWWrnK8IV5HcFiZAmKAvvoCsHI3OzDVwvhC27vo+xphnljCPUpQYXH
rSuFaSafoaqgTMz7HJIt48+TfUQy+4W36qLOOBMq3peC8HirMBKbqj/Ifs9NhzAr0C6iDslEW9EY
0lpK2I7n6YPuNIS69vjV8mCxfyAt4ZGglNwx81AvUXSxAVZy18nDOhhPMgFCJpLE/vs07kolm31K
jX6RrN+VpKOOCFZFtcJGqGiutY5Ltm3sx7aZ2gYoDpFBlvWBGlxsOGQlZnmLy4qwuK6s5bthtjn3
1TZmv05ujxvZGkUYu0oh//WlJU990FOV2VNfdIEcjfy0TnoxJxw3vjjtMRh0ZkIL7JBkbumdjdah
PHAMsqomhe4dd0Gw8UsnJ17C0RsV3JRVsn6mPvLZQaaHgEl17sR/g1uQAMbVKzZmKeVoT+RoxFAr
DrSoUY2SoaK9k7Zi4FQyHaZwSYf3Eo8yPuaNeNe20z8sEZ3svSfVzf+qa/upTKNZUUdXG973lqqI
k7JAKE8Nm5yn8nKwWHX9zjW9OZylqsHMP8/IYtElvaZRuc9Sg6Ahmj+Tcf3p4KYclk/tMrNfj6kT
+L0sHePK0qCb5J5pVpa7J01jTCTlyHHH6meOHAw3TYnG6bWntsu4qnG1lCJQPzoySjzb4Fsc4y4g
Y2Tqj0wUx8iqYXwfvpBprITmeeRU8pq/zZACXL0Fc7ulMQ9+b2kWDYfC5HgNMyOBHgzat8rZXVDh
jJKsqOB8gq77ljAuMsjVq+yjNmciTPG13INWCx6esI6kCjM7qQaUVcpVRVlvWPky4gkkUSsGiKoc
A1PtGaapKXNtAs6IGFgVaGujcU6S2+Po8DsFotExr45SHI0Gi1k7/7X+jlcoFeXEPzIcHNoALCVB
PeOkGASEPCfHh/S6ChFvRr5Pvo6FOk4RkRNcNe/1T8x2Hs7X/oXzNOJrJx2BIONdozsRpgtHrcVL
9YDOqgNkNZLNE1C6TSoGlaYGhL/imaPVTjIK5eHuvyj9hfbUBvqumj6ALElIO3EOxiokqxCfsAhi
jbDlYyEDzLMfgbJSwDu8oJfbPvsY0YTS8DGQifECMd64QsvyBjOu1SveZFxeUdqj7vt4x396XDLh
OZK89s8095h/fc72SnlI9hQUGsE+rEPtfgktR9xdO65PeyWsWmI/V3jB6lGtGYqsaZPYmiSlBlPK
oZ8x9T9dSD5zdPYtfTZUOe5GGdgMIktMBL8RWVXcS+qFYlP7geEZcURO1xMI/8Ar+YvGIkB1TCDM
eAqAmcw+LIHVAJrm2Iy9Gi6Wu3VVFt962HQcdfZyR+YYWRD9B2w0iISQpyEOmWZvXA2HnlAk2U7s
ZdPltsg6pEbao1jYAfgG4p09bQL8/0eyWAD1oH+3U7sQYSL/U4hv0vflgdUPJClLwqVRJrrDCNRt
QJCVs3YrLKRZnHHwUhvCUSETdTNuqo3u/afur6hg8JfKZHkoJB5vRQQYtBz8OselyIoL+O+3XB33
BVJeW7+XCrdr8nPzQye+rDl/Lfsim+5ElTLf4ylPO4ZqKHQpHHgsFEiIhtYRMv6p8ewRZMPgdOXC
yuP9lEHdkS1BtcAO1HwgaOA4MHiPNdcbQEJnjeQ+dIrDHf2I3tJ94Y6CIBfcy6Vbul7Lo6zulJNp
zvK/40xEn5IsAH67a0V54iLl2sBNZ6X0r4jXagARUZlNnt9abaw/dCkOgM26NMKOvlunF+2vWxCY
9Aq6+Iu1yIbufp/RfewjOiid2iPR3vRvwr5lupo5cs1TE8nj9P1gYIFUbyAwSME2zp+aJefmVJZG
cYuL/EGMGXnf92H1kzCWSXyGQ0CCtq62lgt+yE0OYWh1kLp3/M/2y3Ht65AZPnu8m0+6rKgjmnvz
PhS4LMLI/CVccKPvKgsGpPLIu/5ncto8DEkrcRPZNOlD6mIo8h5I6ItitpkBbb5e2lkIXSig0T5h
WXCT/TjuUfPIKR3wenVXvDthYGclcqLVbYm8aQz/GnJ2UwRGrtdb52BDpnnK8/dieTQlWqddOFSX
myuA6tM1y8Zsm5DfGslm9jDc8/3sREXi+YQZNB6ghF3bR/4kdWMX3eudifhY5eC9wUwi5Tptzk0C
husdwgCVRTmI1p0jdGL96OsOKl1Hk4NhVvE82y3O9+SGAt9BQvjLwc9e5z6f2BanWWxicZw4A7Od
q4/jvNW+loHcEb0C19iqbq7pYh4KahqCiwsJVt+Vpr/ro2KkJVbt5JAkWh8g7hYg5z7MiG3AHrnr
3QDvuRWGNhV1LpnRzG5TfLcAGLb3cxXFqDtbOrbgRVMYCC/qnITaojVvpNHvj06ZU2UXS9qUnsIB
L6M/eByKuy1+Xc/+ldQAIUviimL7zS9Kwy5HEcewcqGOx6lp+cz9qmGFjbxAhRkHbZIZ1MWxB6GI
RywNArtfml14Bck7e/p11ifqcMN3kChQOSAHMpYxpLyyzD5mlqLV4ZftaoOBSIyYmkqoDIJJbEYZ
s5r2ORb6Zt89LSDR4Mao3u7UJpdGucp8fPNvm75DqHASPQph/2lVnHJO/FCTNGoAHPmYsuLURnEu
e8FeloqUuDRbO6hhCC/2r7LTmQgjVRxT29a+sCJxw4TvOtebJUOZCx0txOYZlXanURmoMkEMmWAh
0H8WC10xSnzYOAz2ZthJrnxj9l6jirVZwhev+dSiNvk5TdI25xwsJzqQB532HHOXSDYTN4FvP+nn
pIGndFckkZjvt55I5PP9kZVdRFb+qnK2HuVwxfxazF4YCSbgFccOYlPU3R4GAzbpUQi1pzBZD1t5
lq2BIMB6YhZ3ocDxtMiqfxBQLDoT56nnUvjg1VrabY0m4f0HS5Ev9fglTgEWqTbIJUbDt0bacVFj
k4yA4unaZ0UWsj2Ml5wbCwPkftNQLtmvbM/nUUwznCQBq+n7It0cPzO6wbyCDg+OT0mJNSoeXRmS
VNTFtLEeu5sNoeApi1U89WuYXpKZY4oN/7OSd7FeLdgfHSE4gJXVfMac/EoMk0Mn7tRdRKdZYYnz
TTYgbGH+p4BBAgntezC1c3PhcFGX9t/ubZLWOri52t+48IvfGkUdTxLBo/jGCLznmGgIOlPwCSCz
RBvIHQ+4G1lk/YL/z7vZeem2TSsF/dAAcA6juhEPZhh0qC095N/sFazBoWJYLDZNMaVZQ3CkVHo/
licG2M7TGWaA/v3IaoTuhDjmmLZcwS96G9endECC2Z+TJbiqy8OCi8JkyEmWzdgrKk7TLOtExNVA
m70M8nbeFBWzs0Yd+WbZrSe6gnE0zZFLTaBDQSgw1q1W3PYYsygU9bl7smGjTAV+FKrTaM6ccOrq
nmUczTlJUD8V/tZogNHFU2jgGIPzxYRC+jv0H2kItE2PHDJkHTHmyvzxxshgev9hI8X+khvQkG5G
iMBYyuCMZt5wVs4maT8o/DuXo8Gii9AVSCiCFXPNitOzebFcc29XWUknh+8Z5vfMASecwXmDpyQX
PqRyxqdeuYUGP/I+Crz4IatsrHYoaKO5wOvzCoU6p5fEjzmGr2wASworEDS0hEkogyWF3bJ1U0b9
RGz/c4kBH5PCvR34/5X/fzQZh9ku9pNBnE1siKwoIJSJyYpz9FxMBEY/t7CbWkXr/8InEyxyP9iB
pU++3Cv73ZQ3euBhZMQ0jkS22WGpKDb/kn+SXUYoDS6oeg27ZDswcSarj8zRbHIKqtW9Nn81bUL/
xihiDWyxIStrcnjbK7xT8w9ZyrKAX01WYWCzRIinuJuNm1qJJPSYW14cyZ3uGX3M34HdqGRsCB/d
+fEMHpPjF3nmA1vUJj4yirFEe4SJkQXaGadRtN9pOgtOJ40tTK4tQtEA2ManxeyfHroHSDdxD6IU
7kVJeY7hLs3Sp+RrAB7EK8IcpmTto5U2gU0F84NMWPqlhdkB51W3ysVQhMEOSX7y1VipNQSaW+Uu
1BgiM9kDpczvd5aA0AS7D3zLEQBIk6LR+7DiEKsTJpfCFb6IP0tAxNvkWZY0Nz224Gxnbvb2EmRB
OryZ89OiHyiId3r7Ks2N7lfFGHYBmxuMGjX+f0khroxQXFxW3eGAZmW71OITfso+Drt1+NsEpaIV
V259q/3496tofwFyv94VL3vgPNIzrq+AHMpzGqnwRHy6C8JEO9/iI4IOO/RElDVjwEC6l5iQ1Wud
hY/3G/T+WYE1vyvtiU8hk7jrxntWreXUSEMmL8DghIxcY23q6Jjlz2yXruwogshIFy9VOb+j7pm+
zgnq7Cucm+E4XBxgr9uebugReq5uYKKxMOpeQQqgkCXfpX7y3m2+Si7xZ2WqcPgMDhMb/05g9Pk3
S5H4FWqQRW+nyRpPnXP/oOdD8hYOeJ6bwyvx3DenqtNDFejmDnGRqpa+Z1/hdk+QTrijN2AhiHqw
VG41ZZGvSVVUN9RLcipJTg259pdxjLdmS/uwBCD5yWr/xjeFwWiyziz5y2XLV+ozkxDHpRglJQjN
jOXwkA+CoOrQZrJee4eggVNhQ15sucMJViEPTMs4MGm3EhQju74QV8NbeMpSJrm785qK7EbgKxyY
jeYw1oZxrkMxrtCODe3Q+QXiQ2SQfLm51+xIvtmiCIx/iKLEgjuFoHyBysRuK4YaaqUd3BkIV0PO
hEq6kDP03j8ZmTz92fhEMNUW0SrSXxmAPJFo5o+hh2C4fVTrqJAKqrbgvkT3AKBy6oe+fAmj0jhu
bUVBuvOMgNyssgsxqoPd90eCFgHj+VHuY8Us1SLMzqHPgycQhUj3DUCg4h7bn0Kl8vocOKeWMHIy
Nr3z9MmzJ4iywlq2Qd2cvqnxmx9Hb8iHX+EcdRZnq7hljBXfaJt9EmkGgdTDljOjFwBM5RZP2l9n
F05oJQKVj+wntG+QA1Zre0uho/IKCIAuBOilgYLqVGmD5YYhm7becmjcV/VAC8eqx+KXoDZu9Ldl
wouXplyMeaVqkE3po/G1aATieMo8Gl5LNgdk8T3GQABF0T3HbkMii/zlsnrzCvdFwCAX7BbX0Ghk
CinBhzqEBh0IwucJDDNFL+FZ1OumbzMf7f9cBCqgiZturKOHG4nncJs0MWAoO7gQIc5oAC903IEb
U8Hg+Mxgf50gWKbRnGtSKns/uCmcm5xHQNiTE3Vj9CsxKTl4/sSsIAVoVbRR2da0m8oDas8HrBe1
UpeUoF5L4ksga7FlpubiOziXkAlsg13i61bvRuK1HAWXi9qQmf9fA2vEo+3bMZo9kqoEpIGj6e0b
8DbF15T5DBJReTISOdPKnil5pGkFxECrOQWkpTOOc6v/PyvMNv0RUY+SQVmPXUwOyq7CkaWgaIOk
GQh0Q9QHziQR3vmbsI3pRRpsTXHaqD1sm4on/6sHt1ScfXILzFAjQ6uERGDD9XvzZHBzn/GnTX2e
mFtNAfvVkWZ1oRfwBK8fW7nqcCgFP7NVBLNcc2lCEuJk6+fq070jtEK9KYs9bHWG5P7zxnLUV7mg
btR5OsEqQnD6Um+GA/8ihrZ/STD+f9RthBp9VCMYFATeK9CjoR/Zy1agoN5mwF9Szq56eI8sLn18
Pp/DegyirjY9Xugnptj1Chl6aLEidBQdSqdrAy2/su8/hJ1YHTg/QUiRMLnUZN+G4PwNMq6FlHfX
95J9+j48JbxI+67i7NEPDZTrDywwIUgkC4MriektM0+l9NMDCsemdFA9wBTSiwccbpa4ptZmEn+n
aB4d2uyVjPV2ziwpZ8Foap9R6dv3nPDaplNHdrje0Hpy80/SO6fehGeoGs6buKq8ralzUUBL5TtG
3KHIZamuTsOaOA8gBSknNIlnpVi44X+Fmsj+L9ozJyDDtFpTmRWzZpK58gDpNIbND9W7XtmAUvqz
7WkClPABLD2Rn/KqrIWTvsJXYMTL+V8fVxu/ZlftNoeTekzBS85ofKGOG7bHAki7uOYT9VPIC6KY
UnVNCS+VgL1nB5NsQVpBu9iDTK1+/L9P7pWahkY55CfdB1k2kdHW6ijeOb0fMfXI6jrihBnKafZr
/Oyk0wEmBUwCTzgQ6KIr1hXPOLD9uRxblrB4W4/nhsu7I5vBtjmkCM4xKWYM39a6bbF8nizAHtqF
1CmGZKsKYdUxbzOq5qGx+cVmYWC0f50IITM8718hCPyDuNjn2n6wCw6VdzZKy3R3sZnukyNGjnzD
8XPMirEafDLdR2HKAIbDEVlfX4uXyLjHYnjAkHZtZDwOZk/xQDZqevdtk1PF3YnT17QqSvvoD/83
v6Q3BCjhqXB57UFsE/Ewf9RKhbbbbJSdM2nmEL/5N8Kb9mUWmI2GUbd0n+lpB5dItdo93+eMa1us
2/2YvKBZmQgBWZyASrEKEqwCTQ2HhVqR+cNstucxrvRQmwAJMuou+dRFClIVpL7iGbpZio4BhXFL
yu0+YqD8un5+Zu2mlDIlTPPrGXlxFtpYQQeeBakDe3ojlSjvU2vQ7ZQfSiK5l3pMFdgm/oPK+6AZ
842BzO3wZ9UMoOeNKPeXZ6AnXJ9EEoEjpjsDzIvFNMaz9J8qMji2aMPzzLDUrYOlbj/GfnRb5sON
UjTUMYd2fy8mxnK1Mn02JTxNivCtVNGBa6/lJcC7QX9DoD6BJvRKRCuHyFVKsHD//0ghOOiCU2NA
9dq+w10WVMIBFCjy4SjGe7dTDnrZrsARYX2gGzu61nQcmqDb++sYc211n6QM0POeOwow95aA2dWQ
A/k8BbuSGRRQcVZInSCbS49sXslr1/APRmDRHZYnwyQXJMSV1uh0rHEhldejPw+IMNxCgFrWqIzQ
fT8RPINuPfwIw8RLFpRlpUov6m/u/o5uJdoZgZLNEx+bQXTtMaZPRemUeDv1N6t/LqeAFuq93peD
2Iv7Ng1dCrMmajF+43j6seXcR1NFRHmXFABSKx6G9xz/nQqSbAjgmN5dRwBM81q2YIeSE3953qQm
YLpA+eCRdhYaZTNDZlsLpNmLbx+c5kiHRd76Q5taVycBbIthPkS2wlz7+un67dFIU8VJNH897Fl0
hWayOaCnV14f4AEaHs2YN4jgMmWj52hG6W9p9gHHR6HWF8Hh2Jowu21+VbtWIGkQv87Kbzzb187f
/ns7C/04KNGghe8HFO/7ly7NYPzZI5CFfxIonBqh1xf8NpkSX7zG4+ocA52/F9eT18vGwQTU1YHI
7RwQLWgLtyjK+UUuPvZRcEutwwL3fzbxSibSYtrzyYfrr5xxRaSJSg0PywEbgvQ16N7NK1utmXE4
WdJqPBNMf3TCa73axp2vg1KLyqhHJ1JSRKRp3qG25pkIPP7bDvqqqztdAQKCq2YPjiqLt0SePcdf
1shZiHwkusnVhiiWDQA+hKfx+3BS8LI+4dXYxeQWkaEQ04MfaklsFczDJXJjacuhzBXKDpeDMcXG
276h9mXnWH6XW6Ql5+JMUPaEkCjC7Q3fszlqxR7Uhm6ach120geqz0LZ10EZcTzKAyBUV0CH/wsj
LPtLmTF/J53GPVYkCT9L6+zCm+nw2Uy/Gwl05wU8bGD7F2IM86Ad/sIqsCj+IbConWnz10NqjSHg
DiUOKAOqOKMji7Gz1q+g791hIdsddk/2cM9RchTWR1DfkH+B7FRA44BvIhktWuCPZkvTmpvpbzO2
P5TzpSHOx2XxSqHpW2bwQ7BfY1naRFnZOcqlJr0+yYLmvZps/o368poV1pjZZ6fRjp+0/wuYptFy
Cph+rYdc3IY/BFpXB/i6iu4BviPNhU8PRs90RwXX+nBaDHXY+oRy672bdWay4/vtZOZ76gFtbNU+
/uPHDudbtlWpN9ynlB4SqwKlQxnf3v4K//ttlWaalOaZp8OSvTNw5vJ8/CZ2OaPo0e0ZGWSDw3Md
Sj7a4SmdfthYqINqN1CYGZk2pQDHhO6g0tcWPCw7ERPjB7nDHN3lbHENOndqWLSTea9hH3Fyql1k
TvvliJaiQCTSaqtyPqC9xarNnfYk0uXngPZ8yNZcCadrGlfWt8C0x8ZLBuWcrq2i42cFJLNonu7M
8/UhBgizhz9y5lZqduUQHejGZ3EuHWPEMssiKDUqxoKaEQmJJtYX9Y41h0i15k+TSnv/PnvlVVFs
kePihP360X7S4lR9OCi+4dsVp466ARLfhYQzLyjDm7Ma0CUOlCPPjHog/UqBqML5T4V5Q2UYvDyS
QF9N0FpciJhFSSN7H/vUJP+3XtMRQPAUEu0jVvUmpAixmVz64ppmP0dyPDR2abMGxjgDwuejHvQX
Bw36YXuu4+jLfbpOJpn9ZdsmPXKRDS6f9Dat2jvQ7+DGLvt2kvNYeGieqetDPLniwesTHdkTPEpq
z4a9PZQg2b4xRNeviysB+cdWuGaKNify1rqjoGDGbcoIiExgF7ZayMvZydM5hbF+wEs5fQRHBO7Y
5NhilM17YQFEJp/5du8QydPDwRzqzW3Pt86cXB0yU5+3tsaAgNGFtBpX71zwXVRzXtf1PWIyb0Td
WO56LIx0+XT1mVu2zWHytlybciLOdooq/pD8xUxdhIikOkeLVA9mVc1F/zAihD2AnPEEiyqLYmww
OCov6g+ojPVZheB1STypemgMQIWY612iW7Yw6x5lJ9jFx+oyZwG1EEadIsqj9JCyMr+dyFGQNlou
oSL7q3ukZu5LAYxeTAQHNl1jPv2WKeFqQ8LiONLlUEB4cBiSAmVqbqeJHS3DoxNQ+DaMab17YOBn
5libykss/Gld4Ozb596zaM01UwEc490C5bTJbpzlpknkIC7oGf1fui8Oe56Q3fSufxTrRtzsHv4p
QqYNBRF5g9tx12YCBU/gR0SoDGb8EhC6ix18zBeXo/F3YgisYPLs5v+Qk27icvSArJ9j4ZSt9v37
24eMy9JYjUwiJI8vdGUoa8ryAzzaCPSfQD5utaEXg9R94LaND/ZT6Rnp2OV/+Tx/p6dtsqPIV8wq
F3qxVVc7fnsljDgKAdlDj8ACwZrce6NkW/m1roWILb3XKTozyWo7yvjD1LYLv/xCVp9LwvTXc8nx
PfQJQGr8hCJ+KuTsVOzT7B9Jd8q78OQHVadjUtppmceKQdCV6I4Kovs9KAM8Pq3ZXWV8l+0Q3uO7
HLzQhlL40HP3SFt0EJWkKQVOCREWcIhcDJZ+h+LmDxI4VYXTRGkk5TlWCedtz1jY6ehVG9rdaraP
Gj7N9JzJw1azTivfiq9kgeKs30d6ks0DpSg92XG/Fx5sMlyvu0N/HZFkw6t870+eM2mTNKKJsJp7
ypXpEY42X2HHzbqBRkpah/BQ1QTq1lOYZdBIlv7uyR63fishVRfY4BWTynSL3OMh3+5tCdaduane
5sRWhoM4MOB/l6ztHupi5Sfkf6gl455ggAjkc749vtJN24GSsbOtm32XTECXBRyI82AphEplZeMi
TlE2ZV892fgD96le/tLD3CTexC6PQbo9LL8wqeOHo17gAbh14XvFWRINywuU8EeCFsYGcD1sDkLu
U/JQjI7xLdorv/fAZ0y/kSlJHA5GWh/wY3oKfv0aIA2jNfXwb4iTsaEtybZhFueJcT1CsviOc6pF
BA+Rehn48w1ipN3UqKiaZzaOUhwkfJpu6QfqjXKMB07Gt30YpbGSpgmNaP/VCNuImA5epvsjKM7Z
z74Te6uFHugJ0sHDQKpxL+hGQYscIscW2Qd0YSEQKzcHtPMuEPP2l0A5mhrtmbTKCgVhpGDKtG5X
7inL0eiHHlFYXZmhpHuNkiGaBo/cban9HP9cBn2PWTiA41H7TM4a4atG0ssV7uMaNCv0mtKs/qBB
ZSoqlR+kq2U6SEWxronA1GFeuf1c7Vje874aU80B7g2hJ2k0zyrf1gHUIyaNH7SmZr/wanttFr8E
gRnKQTP7oYAJPPfjEp0p75wZSIGy5SBqmv5wIe2Okr0T6hnR/EtVCWgve2/YPlZVg34OZEGt8nrj
6ptPbegAvWcFh4uHEbgmkfkdkCkY/fdBgkyjl1q9izP2O/GNApKIU+jzSNyxHQt2uC4g80LmOQ06
tc3G8K9Rqk1+2nyvC1xM10a+vX6ZU/LzrG8OPCSRc/yuxUKTgPn8q1EKmdsrq/ZdKCZ1jRNEg9uL
e2NzlQDW7+rKcF5K11QxfkKdKEfRUsH+SS0MHpzdpxhLHk/X/Jo6ANzbTKNK5cb1ZmyQJApKaIjg
6ikzjSTCqPYq1Y52DbCjCAu8+q37pUaGgXb5HIazBirTd2J5bhKrVV/d+s5uAHUXJeK95R3/DeqA
OjIUFvelfrLdJsL9lWlgSZjPKuuFocDhbGrcDs5xmQfbMFCVx1+kvp2ed4ouzwyoHEHsaF7gPxvy
Bs5PHGNktdzz93C4057oGb2qWi4rGRszkJSeACJdyfRFgepGYRYfP7zrmI/MtQqrMzoajkmDzRuP
6UShINcAmLqdPS/HV2jwQIkqOa63ktbKxT4wp+uNTSvpBsTDqVZmgU1bw85gROfe6XkwaSWxFeRY
6MkmZSz7kOpq4r0NrboZSuHypBKPpCrUvnZTNFunPPNzR8ip93/MAsy60X/daJHvWnB2qAUj9sMF
v3jm3Hry1S/ot2vqVYNWoRXlPaJB5cqMasYJMy9nnf6ULs37rJKsC3AwK757uQ4qHX+GhAYJ+6FJ
vgv7qWRpoHqBWy2PSafuSbpCbakhYLxaZNnH+170HL6OEw17hlM9oVSSPVP/EIvQcLgv/PVV1EGJ
9emgfShRoc0OVvcoasuHWq4o1gSQGHzCoskpkF/cJDg+5tP3BO02PS9uuXJa9rJPvoEYxjEZxxg1
qHhM+lsgjsm1I8EAVDzNNp3RNKmaN0iE7htUQJMudr+sC400hc6x6JSU4y6vrrDRc4NNNaB4T8TH
yT3mjZw01sFF+M5fipoOSbN6UMWyJRrYzHJObEdMUuqN9qqx1/UPSR+WJlHhDnfsxVV5Ufmn766l
GxtO2r+VBDTw/N4CoPUncmZg4X7oHlScR8lpvNlzSp5lnYFHGg9/qMLNyOWFoH2S/R4Qga1ODY3C
LKkhorinlgqAhyqu5KS1I4xxiGprQ0oLalYB+dngYqsNafix+qiUsbOELdx4kJvjflvN63A2Y2qe
bckT728OetwgtF0l0L8L/9qhZHIop0QDV6LW+698eZETImGNsWO5H+eywFveiKb/Yt2v2eTz17Tx
C6Ek5ZAxp/YJMKsp1CDL4YAZPQR0DfkckX3KKKy+05vTFTHrQU8+kYGBfQux6XTKEl5Wl0U8YWZo
y0lMMMCKsjyTNcJPiPcNwVbSk0OolTKvSxJ5Uq+/s2DIqJBIVL9Uyc/NIuOPBfYQpxEqONCmJ269
4vkxq5J1lRvHILpKS6g9nUGFrHnCBse3GeDbWlXEapIcizZksN6RKxY1BG2yi995GxCTNDSHVpO0
uat2RRgIp+SSIlHTTPFnj7LSQ98qkCjkxuGnEAUsaGdoVObLm4rXDH7hAv5ZQYHtAD0nhppIzFEv
d/uF2yphdil/A7MlAiFUwET6ZiTyUmMoLr2NwpMLFPQTXg7kap5etN+C0GyClRInERrXltP24vvD
xS8DGrSatMRCon0ySF7OtDj8w625pb/dIN4aqr38r1TKM3mKBNMKPRHm8kintTjct9LKLkt53B7A
BoBkBcQlYeJJxSFvzxSAfsFkMpuJKOOVfnirqitrH/VN2LvkHOWgeKUE8/drXHPUs5/CpHgyg3yr
+yOUfDly4bPVLf7FG7tMb+EwgFSl/CLpQYF8johczZpDJZOjBuIVzJifHKOULdorMTQUs2Xak8Hg
Nuhh3N/2LXm1sXtU/I7nTpBbgcwAHdjBX5oMc6sVMrOVwEplGbtDR7LzO3WIlB59NsVty0o9hROy
YKtmv1aPSs65itUeyCsM682TBRMK0XyreA4A/bFx5LOiQVKTeevCwyvQL/BSbsMHP/mGnIbdN5ID
Jdi1Sah6mI/NZcCrNEyGyJjOI4yH1EvPshxtHLeytgIu3A8G6OXwz5FHY+zNE3vQv8LEzdnnnHix
d23MkX//g0hG37UxSiOchQbXBg2MUyN2xwJigRr9nDyNDhud54Jr8s9ewjy3ifR0X7o1tw0/g6N9
QSNIoOwAwtXITp3/6mNF+jCP4ezhqgxMCXOnM3yLvg/HrpNaAvzxn/hJUwv4P5UamDW2VvftsgFC
vZ929NuGXWdOO+Ogix5JTbBlZtF4lSTEs8T20B/7ztv0nmVh4LBkHUI5Iwhbt+Jnb/UMC8Nff9F8
A/4DuORgma9FqsPzyPTX+3h4n1u5Dc0a066nauafcbTF4iNwFvFkP8xLTHZvCjp2veDY3kimN4iv
7njYBQzCqRuIuigqG44XKFg2EsTYJMYkvLVdLjVrbUigu/EUNI7V9eH35EFNZWaBYy0P6MwOKOLt
1RSklkhciTICYOb4HjWyUL7mrWCXY48BchoKlNNjI+q/0Rspn2BlV1iddg7Hxc+7PrnZumg2ugas
ZKVIVqcvDdaJ3e1F+HWmi688+UHNFBCNdI2wLJUmE/QLOA8UhdyFHGHwGTuWXjUOQ2i+YOsq2yis
NRsAbTVa8MPCeTY0T1njPDLOIB4cgA9yQ3yhaoM//a97bb4u9PZaz6YdwpdvWKUG9Wc0quLPjvnW
L+qkD4lmhrGPbcjrt2mPIK3jY3PTLg2C8zkMFatGeTnWUzNLZ2TAP1vPlsgef0OLblTaEVxu7U0G
cgdtgevwoYfgaSfJDqdI45bef2C/JgrRJquR2osTkfQde4/SxUaxDH+3b6UpXteQMCjgoEV8wpju
+ZpmlKAZklMzYMqkg7xdyiJRoByiSUWLtI58E6zbEhx5v6kOUzcue+UEz2Yd46DPS0B0chVZuKpT
nUEwRdyK8NxJcOXE+yJEG2QrXLYXGDYoddR89HRJYzMM4fmSTVUJffd6ntP8DVfNmvkrOvKiGuYc
E+OlmtCQbum8g7W3s6kGOWGw3WH6Xeu7w2pOhPwNnazZhqZSMAAfuq/J1hvChgix6Ov5+dB7EdV0
kAm4YGLCpM66HEzWAheRkYO7aPqq3gxAkZh29FFRiatggY5j0enCquoVeYZl8MK5uWB0fUvSVFqL
DCCV9D9uxeeDt94r7hYf/7dLXyqrsqRz7Z5BcIIDcdQxveqbuPdO4+JfVrc6zRAgQ8yXyntBebBF
NA6rY0p1ZSKJRbuK0oq/hWdW3tzXheZ682Dh2L7GbwChASXsYKumA/GOWzDttLQsbR0nIbUWddbz
iz5iafuzBfogbhbCqDEFuU4X7E1f6BPGeU7RQfX9o039Czq0th/36G8GU+rEtkwp3sWDQ4VaJTK+
qjAfMl9AoXGbPVaRBEltrXMwY/quBUD8mcgohy4YNy7FEZxdqBlk8dfm17FCzYUxwJMnhQUZeDWG
G6oPoKNBzK1NcQFyIZo1wit0GZE01a7wp2Sy4IROcnRwiRwyO7TduO5mgMzvbaDZICpeBn5cxzqR
OKAd5RxTp/FrJ1Rn8rNlDJ8SvKqL819TWN0Hl15c0yVuWMiO/CmZSgHmVw55YGyffJx0oBcn4p/2
iH976kvXui4/HyKl1CC9OgkbWxAwwXA6CX4h5BP3FT3sn34buB0CNgRtnfKeyLrkTHKOk5kMEpUQ
uPcDlRf+yH2QZBPS17SdhxedJvcZFJD2NLQdXDkL7sENdL6a/55dbmmOm2nfzumM3Xud+mZaEGsJ
rVS77AHJSG3HLF6mP17CWjhdeQBJdtGEOrK5ZCCAoCAHOsaGsd7NmdXgAuoE/WorLJy3yBrTB2iI
+cEfdKPhoYxaj7XFvYfQ+0xGGlucS3S8420Y9nSJnwfYP2CTrluyyGThWDe/RMJxUHF3MPFjDcvj
Qr4rP/TVndVGBkzaU7EZZryXjUT06z6bsqzZaiAr3KW1A0MtVQZKFHwx0qK39reMvqGw/grEZgaX
8zXWyNq4kRb8QZz44hfJZ2R1ArWY4/roK8TkF/NynOpWWBIWeqyz+Uk1vl97+303qdhJ374OAMOx
3xIQW6RHlp72ATOb1za4ozf6mznqh4zA31NIa+aRzyaPT8fZpz/0+oACCJIsoOSaWZ0ZkZNMWqkT
/U/81tTwI0a5g44jbk6/ZiQ7Mpiw0W5o8wLrOscu9hNGjsKZZBj43D8yrMY0manbwyz0e2GMKOoI
vQjovnyWwsezAFbfHOXlew9Gg9aj5AIafjL1VXM2M/gCpbw2LLEeyH4ulV7slgtnRIJgsK0Bq82r
PWaOEROdJvq6nQMZZl56D1en/A2myKD1v+dmfHYrE240JWTQMG1lTo7V1YM+3NPAYxg3xMkri7PK
KVyfG43Zu/KvhaJc/T5DdZINjTeULo4O3VKFq1JKDiAGb0fDTm2Fi4UC+UlpUEJpCXxrud8z1Z/7
U6o6z6u/D8RhgE8ow9LuQ6HpuIyQ4ZLUZAegNoKIF5HilMdbje9gkHwsbDKkblLKFCtPnRNbJX19
9wphpTYq7wl67Nr6t+ZZQAYaH68paNwDVu8GhGfETyiI0kSpemh7xMjaQsJsc9mBVwgF8QXxPp3a
aPzgUS0queFtuJaBUUaFSEY2YHfq9W98wI6qmqrjIH1ybHEr7AEOMAQf6bWQdXf9jdXEr9iXvOuw
A1lZKYpqnbXtc3Yj6b5P/vJCtF1VehU5HyZvSY7ADPtirMhdgHz//JspyrIWB32WnXEUST/O82WP
/FWpqtWjFvqrrmALrvrpS5wfeMSGVfupKglUYimJ0pl5pxmzGyjRbZ7daBGWKuJ8r9C+i6dtlHjZ
rmg0y0JrpiuzCsijYNMnHS3zfhMje8cDoVgrANN3tSGrDiAfths5afAqKTeR8kO5X3pYT1ucUcva
iEkb17UAH7E8Tle0rRSL6jN2D+/TvVdZT14ok066PzzcUKVF53bX59XZO6IWja1JEJOZtRMrgjgq
D1zoBd6qyHYkYD0HuKghUa76/fCw/jXBjY8nGn93pgTKkMm7ZzLTfr5qi+BZ9Cb26yCzDfBf+9a0
Wt1GX2pMGmxph9wImJU4mIe2mnFHR93FngZ4mr7j5i2e/fUAyzPbT/JNzai77Kt+NhcT9TUQW/FV
zi9eb9RqFFRz51/HTOLpBehL8Q1jLgjV9LlYQtO9diad0sqELTnsQS2ViNdLN5rjdhYdbyWKFuqX
Anj2oiongjJF6R8NBcZ9+UvVTNBjUXoSgSWbNc6rjISK+4TfMOgSWIWl2/UQEbQ7/cOTniKsU2wM
JniszONiOMT/6Qj2I+q1hNUgZBJKx16rsnl4KCtnwr/IgvPkGIRFbHmY2YiZRC1VPNf5A8Ys/OUx
6PBAnNt3KybMy39lpus15K6HDP5DF4k5q88nSQR/0DQKUi/4lFLw6q8R+ypwawU6Ui0PmbE7qDm4
oPP6JkeJEjjeRl9yZpRkTMhDcXBQuVbfl1TiKNHPbc328ZWDS7TyqIPEQb6mzC2109tbPoSgUQp9
ZuDTAQUlnlzLWWiWIPr5rl6Ijl43hc4W7CJ1AFFHMPW5RYfYTHg/lG7YTkVDUScyWSxA9xpT9r8m
VCNOaxhPumA/hyrSZlcV83/Wg1GqqJQa2czWgTxJ8zYgiEaZAPbA4RD3X4dGAUmWwtdvo85GYbl1
0w0Ah/l9t2N6IvvSvTPBZ2j1oJwAz8/r0j+vo1b4u+SEV4OtebhLCvAmhgTvTdZMrNv93foTyZm3
DwWE++L9PTkY/5Zaxsvg7G7OU2/1vwIrAPyKWmLHfObV+zAWlJJ6wdvHEAIvwagXxN+d0RVmbPXG
NN3/GiJjX0pRvA6HGGZaLf3FjqrjdQo1mS3SnK772hf1dnbef5mCqVDdQPt5DAj5k+hiYJLnLnbW
uJhWBlndR/xaqFnxuvOK9/fPn8VAJSSUE00dEvwwn7003NC0owSlbiQyEuYgbn5MMaewRSXPqwcA
T2f4CI/G5AUPaFBDq7zEVqrP3rgwl/mRvlyK1AO7h9vvEjG5iU7FXC7/7/9u41I82VyEMjZKYF0u
8CISKZWNS2Jhc76pp1/wW4JVV6vUT/8WH7tWtjcEa1LBLhTtrnFFGibrTmqIA3z7YY+S1vvG0Nnv
6Yak39jtDcszKcPedJZDW/C7SUNNhABqtvdCYZ49px8wxOi2s5LBnObM/nmXI9tBfC8Q2R4ZDJom
AKiCa1GThjk7w7V/0wvkJ6VufKYNFKB5shTpSPs5tCn/VMCQJoswI2+BH1PlDVSpqog6eQhRE+u8
NunGntd2ArnCR2Y1ZbJUk+9It/zmG4VJGDnGQWz02jGfuSKxjAMHLNqvdADrM5wrl3uEhx048d49
njP3hldrrrtqzDb2zh84n7BsmLP+atCplIO5pLnUrB4eZboTkgq4GCfCHmKrbtBbIOf7kJBnFt3F
pTG+pAxTUIOm7INPR94Pf/XpsK36eeYyD7NXChO+WeD+0BTuLvZzxeXW5bY2TUECyJoqOQ3b0zKU
BRVG8Ts0gonfnCOURoCv93HUtQEYz01fM35FnV4AbnPIFIaaI0IEeyko6PQO995zwkS0hSQu/oOl
isXRDVcTeCcR3fupo2Z0u56HpmfGE6lRtg+m8VZF9weIWsg2WipP3cz0INQpFLLg1z8AC3FnCiJ7
zrT43cQZef7g4aqJvC2ahSh07VLCIQ3DsUOA87yXrvgUL7BVB5CJ6bA/TaKS1X9BoRx4LfjUs/ka
+crgB1Jd8UzafXJlaVU+j8TrlS98P0nv5Jm1Umpy601Qzu/fI5VhtBAlwXNXRWEf7aStPjztGg18
pTkVNjcd4XjEGBBn8W3vy+EsixFnFgE1t8uQfK3o4JuUG3Z+lnpj3b9xbbRLZcGC+yYU9EkZI4Mv
NNPpGspQtZKnQoVGT0SrMM/7K/34/IBBJmCFUqbgBduy4kQ8tQodM5hd9VzoqlGvdIcPo88OWR/U
N4f2biLbMhL0V1M0lzhOCxmK9ejl+kWQUYabiktnLC5UPGg169y5J79qOgGvu55WQSLS06M7ySxP
7/WogJ0mKBoB3oeBbfmoM9RUl8h2JOrSpRsUVTNGc++mv8Ify3QEqAoWOhxHyLumR0AXHcwNTjqp
H/S7cABmn0yZ8boMiRuiJ/9Vz2LrN+VAe7aBAKHyrqOHTDlfaJq7a2vUMxsQl+DsC7w9w3OuyUT+
VQfwxXdiQBUWJsjJtHz/ZXexsguKtOjTXe8tjxn4rK7RwWShjE4nQ3Y50yG32TeV5Yj1mIZxLrCw
fFCu49wDebVfMbP5h3rGN350Jp0ctLRC/NdWGuQWJazs5NPQHR8TOo/aMncxHxNfu1KUrtGTZvaw
egcWrCO0/JpJGllcR/5Sph/421JI5lRaBC9dLMJtQQTPsVRpuJv/p08IkW7mkjabUO9UlAChOd4r
2HS6FMkdDKcVJVwI2FlFXToSk4egWRJZ55KWoV3WsFS3+VkGnQKl7uuG6c3Z17g0I/YbM2GuCh+E
m5EjOocZYlL0HkLZf9fx/zd+x2giAVSnSKnuzEm+xd+JYUaclNkgmUif6Ac3+fM0BA9J6GzXgXvM
+EqwWLE8GNDcAuzFgGZ67oM/YKMHgNx9KKltT1DMb4XMv+EYYB81hEvfL9ejyJ20XXwFdXu/FFZ/
I7WCbm0cc6tDQ6YSKvHCFqPFtaRKduT741JgRoD16Cx6J5CZzobQ2zQptsc2MfUElzPupOBFgyZS
py0OIDo3r3Qwx+Y9tyRXnyqUgTkNNOSIUIXHrLVKj/t3kuHa5NS4XTWiYTS6hOskbKu2FJjb+RUT
49lUnmvIGAqX1BBKYPduum2pYd2JMAgVviWbGzsT9XEW2v/jCygIJ2elaBt+Nw87184r3e1fsV5P
l4NPeZAKPmvjQ+iPpCdhZTuW9PiTgEUT1SyO8XGzUcdiiUPNfONgT9Ud0AA8mkmU2gbO8eT+Az5U
esEQpACbk+50bo/HfcJ+bIin323tszbBWd1deqz3QaOhvrkSZ0D/1Lr3B9eawLcXGAfeb+Kf5s6I
8bMiu4l7FCNnuCoCpzCvppSNAP0eDbJ3Gxm+R7YvZ9sMU4sHs+B7/fFnSzRsY/SeV8WluzQNPODd
Y14dGsMjRcn7g2afgv7NIY0zxajElssrtfkFeXgXr+cn5zIwljZr5SJRn+rRgKnXdfxvLHYMFMTG
/UnbH0YtH3PfnTJhCATjOzT5KEj5RhCeRg7+lJ5+gS0nlpDtwa7O+v0+G71b5KwmYYntTYxztId7
pc0zDyr/kDHIaGwa4Cm2GFL9XmT2Ep5y+XFAIkoRcOh2T9HR62cZukloJQ6FLk6aNJ+lyyCBuCx/
NksA+gJUNSuxfd6yWxqsRA4wwCkGOZT1H/tSlGRcZjrtUK64V4jHwOcca/e/a+90Vqr/9E/9ygRc
tsTMbTWz0ATtzDMLdhJBV29GqT+ytFhINeQAGScz0j4zA/CW0rhbDqKzflI3cd015G6V+WekekPV
fAh7cwmrscOhFO5c7zZBQlCKUG6Fs1Czi7sXzntDsWIrwitEbM+f/RhD5tBryu9/jmOY8n6cuD9N
6UkDLi9KmaJfbYFdFg8AbJivLZppc+Wu0Tv0fhRJ0gqHv96t1DufLnCRFt4lKUypVVSe7gW+uBLm
MICDb63kGew5gsKFnGNoyxx1G1J7iycccA3JzMN4FK2ZJ9iyh1HgLSD/PFoqyTGzHKGg5/z6HGTS
w+kMcB0HMNVcccTDiGkd0/IM3Da4WweTGrhcGFQ2D6HhEG5onzG8OpIQVtkSNPpppYJ5oMHGxNjt
JxvAYIbVbmtFgqsDnEo+ws7O5XrccFQUDMztTkqUjolI2Xnj9GO5i//RPXoLt4eN/C6GqFb8gZlK
27Ch1IJTi9SVU85GTZJBkILJ5RhwH7Fz3B1Szqj07zxeXENgogOpr1aDyeSIymnCitGxbNLdgV+1
p+uD3pjc3KyLi5D4r2fH2rSn9sosS0O+88UqiG5rroOhzaC3lC2w6ha6F1IDAN5ao2DRDZz1Fpil
8pTgA6GbBjsDPLEWZPqvqS/XtYwnNGZ2N8A8MV9/EZ6Es+B/rD9JNyfRs/FOI0lVc+3ka1hg91M3
0I0WADIAtMVaEEzG/PYOrIW5kHRQDpcFRBE2rSqWiWYrdovMzvCtW2A5A5iKo86xCFhNTr7WN9EO
vqw9Utb+EKXOpUzEICrlTLRmSQzNEB/wK92kDW5gyypb6yj+RibeAH64o6ibc56+fiXFxJ6CA4bb
xyQFt0fg8WhNiT4s1wPLVtKKcn1WlMaUhnyhQD/klCXoj+3AryZiOYQMhapFqWmyf01O809amOPL
NbnnS+Nlm+fOT/jBd8Nr7pnwfxwc+jhr/ZZoztKsMd9eYThH1n4Br9wG+0fOMdB9DtISBlXaHn7K
yu9FMIdTU1d765ootFo8pDF0/R/a1dLoNMcJRzx2SMIQ6WNFxWxro9gD8tdFVTnsmsWahC/taKsb
ElXlNsXPNAX0KjtP9EEr44dUVEYIOCJvMUD4r87X5BZ8wjmKBuh++pnYwjTfK3+Xz/Bf+fk/v5t2
brLt6mWI2p90MHK4d6cIHrxr6Jp0NL0BeYOXSb+aJhjs1f2Ut9i6bsdlVJYgj7R8fe8r391LPX/X
qQogHq9OD337nCJxC7YXwnb6WOD8V4tzY3Q4c3KCiiDm0H64fw+nAqpzzVDTX/V1dfp/r66gk9qf
RJpIfUveaw4z7lzF640+ZL+MGNAKr7fZs/QlpsdXo2CxnO/t4i/XdMs4PpA1BAMwgSFHmonhfIuC
I1EwRd7oQdrUiNuW5lwVlPblb+jKeH40W5l5myC3mcHWGNYGOy28/D6Ya+08HWySS6cBOcXxYEGb
LagqmEuilo4Os9bFWEQumcWAgi+RNep8wehyadZjYyU4ZfFLuIz5yg37puyMgKEZyczwkmUu50kO
NcKkQmwsJLgDLskrocYpaHAAGy63a8/EDou3OLMTQxcv/z+rbxC9egg6/s6tGYJkO5AcLgCO9kuB
+SLIl7wa6qnySReGnOUL9JD6c65UupPLPm5OgYPyqy9YnS0Paz/WWYjFJ2I9/Nu6D4C6bq1J5GJW
ag1l77c00wk5Fgy7m9EyDe7lXBT1mn04DEktB7vj+qxTOYHiKAZSLeB8PbTY16U9YgGkDNjG3pVX
2oDAJZRtsSXnPniByAm2i1VT1JYdiSmmmkfq3VtEQyuOyQ0jQobE2aYYaJDluXl0niao+g2wAems
qBdq2RXkCzfQrZpAgnqWh/9ee7MFVbWdkIZHcZDMxC1g7nO0e444rv/7kFE/3qjmiF1HdTEWjLPa
i+26eExq34T2/Py1qKN9n1dRVv1rO2EzVCWa5M17dr9BBLQCuqIvfjDjFO5tSzv9GazFTXSznEXg
iQt0mSHug9+prM8SVmg7MBzcoPAcgZgRfCKeBcp7VZYHMjN79Xi+4QTTGKWJEDXwAo8Mawda4gOi
nMJAVO5sY56VkTO1F/48pExzKqVBHsM0dk/II6CRwlZsIl7XWUwnC8wDtkoHZzoRjSpMx3z6qS+7
cWotrwl8epCcoi6+0KbkyNs/QDcqBgCZIUe9Qsw31O4XIoa5+Cao0zvt4AeV4qgIGQ4rX1aK/g6d
v27ZDU1obUM1WR3g4XIcgs9BNoA3QzkL2Mda6wX6jyEhfLiX5M58A1DERey3lQZowBBSePdtwztZ
/UYvZSZpZ2kmtLa+ZVpqRWrnDzxxLaftVH/O59bbsPS0VI+xdNYZY/XafhNXTfbY0Y/y6GxukdEB
PGxLYNn+cnfyKLmBAHOcvU0EbEN4rxrRScvYJow8CFKwNAV6Rtyg+XI8itgwrA/Od0JxbUKYI0MU
biehd7rYAMHmjLjjcHAitLqbOrOKk5vD0IQDFXPRItk1pJeylFTfuTwfMvW7jOnCuQEhMImIdWAp
VMFaj+bAfm3O5KndLEpCTws4bkB15vCrf63nny8k5pS9NeLUdMKQT7I/2/iadWcEy1S8GjUzcPFE
MpkFIk5C9YO9dXxRlc+RKXKmOpoUOYZH17S56W6KithjGKeJxiUqzNmCGj5lfZ3iLSTsRL2B8E2h
rbGuRWf/gY4f8F9QH++6o85di2hbsLdQ+gscz8BETWeSHYrjWosDCUFqvFZtKmFVa+QdNPfq9w5b
45ZlPPbP6HBBvaUQ4jQP8pxoIh6NpPUrqTiZQm6KaScU/WYCht2rhRbWup+B9B77MYoDQS/O2ST8
jlYN/v/zMwPjyevO2rIj3ZzSvl+vioF/J0X8WgAZKhCAG/ZjamEr9TrieZORd4G7NrU/rxDYOs3o
U2/cvHIZ+fhGZGmkFwm6YAmyDA5dujXVhsPyO6OITZ8TDQAFyXbaB3S3qVVgpRlzZPasgRsVPszW
o+q2lN83A4VBGJqU1U4PYsjvgewLPbZL0NZsUe1fhM2DOijiJQRWevreXn1xoS4cncAGbG+vk5eM
8gP2TxnsJ1GXiUENacr7wE7YSW4ttpp3KyLo24vWmxGeNCysPZgTrZrYVFXAwyIDfJIUS2+ooZgB
XGFSKwDhSwkxL2LTzN53AkLoEnY2mA2hMA7uO+Svv7RcJATK0unER6lEWXVHDW9aZ9bgI/qPtq7m
R8CVNpC1bdCvfrgaOhXxPHo2XGVNsYV5S6oMJCILnxZNmJI1ri5WF8vD/TZYKUtN1npdVCnuuwDa
ng4ZPvHVWX/vA+dH9xtdlDdBHCvqT+awgK+ybggpUwnJzojG5qY5Vo33TR8dftMdFaSC9pFmmLYw
HFa80MhaL7tnXMCl92OzoW9RXiZO9OXbjFyn+RsSrz2Vz4zTkM0NJwVXViK40Qrj38H9KRwLDR7E
TNCEB1Ek/bzGgeIgklng48G3YEaZqotJP/Hbc04A/OpVMnbvu1I0xErQbBCR/Tnsqoo0ANznj8E/
iDfVDRplYGv1leY4t+6pqIIhVMdD2gQvefHdjd2vqutZv7QxyES5TjIblscpp1Yw5SZSF+n5ZDZK
Se+m/KrqDUZqcd6KvoE37fa11rP0mP3/OWZsrTESo0pjxRcB7+41su6zwa/KBCrW4gxhehHukajA
7//5g2wJw5B9zOk2AEFPwNvuOdc/2Uzf6VkE70Ajaw+QK5M5KaKgnfk5aoN7ZYIWwPQaqmeYTecY
YSxcR8Jb25vlVPu86BU0PlwnMiP1DI9XJj3PVumV+jPgVx94W56XFHLE6KoVMo7Wfk0ecWaQO0Zx
hdO6Refuyf/DqJmQerbCvbZbnohRw95J0iwchf/iuZEIGYSlnsTdOmx2uJvCH0pvWKgr0krwXWMK
rEh5gCcpw0u/F/M3DElH2DXcQ+Lcihj65XVPD7FrnG57w5FiGuCaMbGyX2Xim0pbgagE9McDYSp9
bYsGed8P4/Uqv204v4kttjg8im9pPK1BTObjMulbFiYm1CCVv/v2eYEM5SdYczGb1dZQ9slx1G0S
y+ZmWFobZ0ON5KkWsd4wfPqtodMkJ8e73tiP3Be3NpG/hsol2OxnUNar4c0d3K6P6ZH1RR5OdX+e
z5X864lPAX7vyzh+xfEeuOTLsM4pErxiLGo+9Z6UhQPfAYr750zMpR/kqyltX8ShL5blK/uaGkfl
tPlswIyeQCDgZo8uLk+smyLQaRewjv0MqYb4RAkIP1aPSj0aLbTDIacgYDmldhi9BMJyV6cHXNJv
E5RT7aU6/auyDPzqkU/ElVN0s22WHV5px5f9WWwbSYuZsmevF5Tja2IVk/y2D+iupcD+0AmuJAXH
LgngZzeOq789P6aeF1ykz4EajY9xhB+8aghHoqvySYB+SDYLG9HofOJnVNRbYzfgwJvH4BO+GbCi
Puu14J2HiGhgx2X1ur48bQ+Ftl+YDRMBS64Dm1a3tAl4wUrmRcyg+7OfNwSwYuWgvOw4qbNuwO6i
dBZ355jQJfOwzlPRKImvaqIrazLuHmfPtY0ayuESjpxi/erK/yieXHs7jr351+UhwbqF6XidcQ3X
aUzd3XnkX9Ev0lKnMoJ6iZdJMjvxM3Ry3BcNN9q2FPSCXp/1yR3JwhlvPNkdX90VpsRjI+MaX62+
/rBEZuKvItkw9R/7eDviWE7ziY/NMb7QF8A1OqR5M4qut/42l2wvpOvU1GjncX/zgJ1Hn3ZsM1Us
UstZgKDqBh70CNhvrHtCKVa9pRIqhgi87Vkiq54TYHjRccXMU6bZK/wAAImIV+mGbm3nJBf7Fxy9
ngrZjkxVeo5eUsnOYbKC6UAOEkqJdJbOKCKNICRriYr2w9UFAGyeUXP31hBNpmydY9x8vH6cUQXD
guNG0MqLKjn71N58puYstecNgp6HbdPrFx/Ubr5nDTrq9xFnIBIjX3IQPkQUN23lUQ1pNoEPbd50
hPpjorLU3qwP6u43A2uZHOzkB07tEKinH9mtRISIYNSxD+d3DGTx69pd9NsMUUisGW1BLnfTZHx5
WHSn5e+UTna0p4OV1G816XHj17M2goOQlIvfklPPTL0OZu0afdlZQRhLHH3VPxS+Ss00Jl2JuJQq
XsIrsDIuIb+3rnYbfGfWk9UHxcdKFvqT7LS2eMvr3iYZJ6u1ccrYzngRA8TOLpMGpUm64GP15kKB
JS7zWck7XyJ0cO2Qh3AET+Q8vCPb226yDiVZ/IjTjrwitrMEhgXetxxDoRZ0TbjvoMvrDYU/D4xB
KjK79hV9TAdxYYQ6w35d2RTRhn3F46LCZTUDFDIng9mnQV/eeLDD3Qtj3+8UmyywNZYVjFyf1OGG
Us1Xfui8dxjD3/uB+QCYDZo48uZ5+2hQ+IDwsVt09zXxBrqIaLLQ97VSxGM4QZgsAdrC760elirG
cQ+PSq9quKH2AP3kFqi4am2zV6cd1xaD5SUswHKB7rqfJsKaXh+F9aNYECq8T4l5mS1RbqNXAvIN
XF1TpsI1Zy+4OYoH7F5KzJ+gQBez2Gt3loDVDj/PGyO8y9hevSYlsbuM0H282qw2v83Cj+G7lZjd
Njpf/anglCUv9zLlKRRyJDd4eiJeSYdJbKjUCxfLuqvoCwiHLleOEPMxAtagnMPlxP1GJetSTol7
Z2jjkmDh0/qFHBNkuZY6vNjBRbguPx9p6LnRsxD5/VI47WakNDIekuz+dxg9IOr4z3I6hNbriFOm
MlKbZQ2q0Q62unerTZD+Ly5hAIT+5en7+gvv23aUbGSX2mQrecI57JRvkVVlTT1PZN49NglEb/hS
6BroFhvu0QlptGlI2tTucXyWwVOQaAwV15J7lCZniTLgCbIK2E76gr/DvkaqS/tJqF4iqc1mMoQt
der3aotSAiCsDxZxR6v9dOsF2mbiS0sCFt2egMyvEJ8SY7h6nozub3Yfkr7sGZ0Hkco4BIjJ+0XV
NRXmgmx8BCVluaTCO5H0dir8i7/gfm1NolniRii8B2FE9DU+cy5aFjb+DRtopwHDdLsZ4tW66LQA
fGurvzlDSKrr3v00+FbZLcqZVtl9yM/blUfWv8AGgN7PrsPJo8sbp5Sxamnmnl+DrvFE4VOQ1dE6
Gy0dcpVFFIuOLv/MEV74kb7dfHHTJ8U9GaIhIsKMn4SCNvh/EA7MBTljDCPn3K6rPOhKHpS5LTff
8a7LvTNVB595tHOAVP8HOgKerwSgpOougne10chgdELGCuC1SuSMvpNYjhHYaqe/df1m2cPh4x1a
EfTv/5mRYmsjqQn9ZQ44F/IDrr5ddviAhR2Qu802/a+59U7Fp9yuXCJWmhl+ggPV8tEdhCZqrcFV
UUd80D9y9vYR/N/4TrDRR1jmGnPjSie7z4pkXltriyZZZwq+JjHRpMc5gJBOvNFqRxEH1UsbGJrj
/gad3AYZMpvQiOJAnBayOP0MYrVSTi7IrW1QmgoqDnQNI5+iKxwjTvht+bwb40z5yMqOCB838S1Y
cHLnfPX2svyDDDF/q/bjiUlf3Son+ExX+9VI+UrWvm0J/5UW/LBG0QFQnGgPvlmx/nATy/tAb3CF
n1Q1facY1LKKuiacngcs7U8j4M6AdLqORMZri3BCBcoT5AJtRZEndr9O0eFLXJrfAooSgwuID3Mm
UJRP6KeSuIySYS0W7YBWC15lbVmI9XpgHDJdpybPPdF49lf6V1BRTP5tRU7xgEiOynWRaMgZLJQb
H+Cfri1W9XtKRlIGg4oyFz2oW5O2l1UyiCIZrSp9NELKVnbg4wVLkT2P2o5yFTiaU/19bd+jRTVa
JIqSYaeT0Hd5w1gtUrezJTqrfNQJ5wuXAthXkYO/y9+K9AvGikZbqk/OmGn6iVPJ/1L+JYIkMdfL
ll1abRVBwcKXBvUKVg3tTjW0Eo+/tzGsX9cMfH7er7r4ay20l18PXAq3+/GWwBnALkkt3D1PfM2j
EiBmnzpuNRU0O19r4nsIAI4Z/eHtryEYHj7h/IFtgFAiwvCQ4I4L41sB8ny/CcrimggCtHrzq9Wk
V3RKgPhOmszsbWDmt9RcEgy58FhHQyyMWUZGinKABmEfOA2iA7RdALz3xfGWuZhAVngq/OCfdf5g
8JDhboFhr8MggRwBFGNSiwuS0Y+x49Hx9DfU7r/rStA+JZi+fYfH3O56qIr6vHQJ+00CtIXX/mEw
a2bw9v6QRFB5ssjsOZFq46MVNwQz7iD8QrxblBNirCN8iQI9ida2z6KEPiiLyMlCtzs85iZIUght
T1Rx9tGDE6x2z3uSTMg1LDgjICWt4EQfOYIf/F3SihiWy2GLHeAxuIHh26me6Oz8MGnpz1FSuRA5
41H/B8BcfOahn9KKq5ufQb1iwPYCE3FDu2GsOPmvvkPQWNy8Kafk45gJYrCY4LmtE7FOIUBBrnPM
MF9qLW5YOmXWEr5V6oHSUhNieyhXzMF8UXBCdTwu+JpINU5vXcBW+dUiCHFYsLM/JMNhQA1vyhAj
ZLFXw9AYm1Ra5cTeZi4Az6tAkD3dML8NsrLarDhi0elccM39Sp9qWrEORNNQKtSyme8y6Nh0/YP3
fBbTzDnUXsuEIDRmoj6uDyY90izLjVC/e+gY0XBOUpJDh3+k9J1gXSu8NcvdbGLHjAAd9qrx1JB1
b0MvpBHs+Zz4lCJYGniSk/qTp3YZM70wFuSHIF0Eiyx4nwzWsauLTJzkZX8Vd/eeuA3QABk2GPtU
RUuGvp8Vhe180fpfKEu3lTpIc9u1QrWfrpq0C5qXqPLpBs/C2odGhRToqp9ba4SorWGwnpWaVZl+
Zs05POe5hKX/taQzSTZFXHg9nf08GQhtURR/d9yLKYYKxA52TqCliUyepBQ+AmykwAh+U1hS6Tbp
f1XeSQkfc/kjtKOEkzombE0gfV5Z+dNki791X8f4wk7a/JOCp7qL7n9BuhtBywWHytMnkGOpo2/8
B8M2HrHcmu48NbeC6yrtUGAMtc1/jaNrIXDwBOL1kZIYaa3ZXb00rd/n5xdmAsXwtkZ70OpiOWIt
YTz0zyzNiE7wBYfY3ZsrytO11mPl6C+kwdkbRdnckm0tk08eRCpPF/B46yxQ6OOrm3nmbF2pGBbv
ceyS1FF7kDDnP1vCO1jvGYTjvhbDugzhfN1GTRaiVHgsTh/PbXPT6zSxaTNuNMezCty52pqrnfAe
irFRDdTMOJ00sSQTizN6IaJHIIPuos5ym56mT9OMKrhmdXqEcGKwY4aicY7pBVpTluqSJnkpzAI4
LVxQPVVpmhOcnf1SKqq1WMHkWQ4dIww/yayQO6W/WfeCwb6lKA0X4wCZNMcWZIvK1ywficzMpLLh
yQ8qfhyrpSI3rnN0IPhDItvDujDbmrw63L3QkY7NhZ/3rbB1UUj5ohqs8buiUB3CeyMog7lXs7YB
3L3w2QWy2Jor8rDQNORHaf885ZqCuB7KxsgE5WBhOflRZXuRwJ9koG20nH10ObJvJX5il+PgTZ5M
P1vXwNyNQOuy9Hmr4kZ63U2euiIprk8I75N7Gs3WmVk8CbE03jVwSbxWzJ/QNaEjGHoJzfxTjNPG
NU0Bu6JAPu6tF9mEoxaCooXEaYbkxA46sVInOWi9gbG83kbTkyt8gq2jIfQpEInh45hP1PjGkZHY
/OzMpbUv35YHW8YnF3/uMzC8qn9seqUAnWxjd9UQP3vLnFK+3WAXJELqCwk3FX6/Zr4qnHXD36ao
U1N1mfuB75Lw4YjZR0P9uQ4UCJtKR0+ZXASI7kkhlDHpWVj6QXnzEIcNKPuY3JkcsJYhiQlHwUoO
jwEaxuzv9+xkrLw5zXKcp/Oie4b5dxAiY6V6jNUk8eC2ZxJcpUO4PBwAQ7J1IpcWjLIlOuZ0IscP
P5BsD08geKTAeXRnrRJ+lXnmDEbQ7xi6rWYkRKrm/nydemJVwaTyBtNZJNLjGOf49IPhE+jDYbfv
HjukiPZhiHWE76da+w0UdK8sJGPDPKYZB/miaQ6jI4Co4ga8pBsy9HFP6PaTvzWKf2nK3tPdg5zL
svF574IXGQ2zZBOSsyxKOc/+uEZYyDyGWwqdwE3oZXpkQFIIkcA6GQhvmSK3iq+VPGyJRyKJFLlC
/pG5b6OoLVS35ux9nKf3djePTDr1VmsnWWe3lgVbVmInjieXK1YtPD6a7YesRXGCcCV3QHiTAXkQ
1kY2U/+A4qJGw6X2bHmslIrN58eu3FH5yEh6dN4uVCOO35Xi1rN7KVgnmdI3LAYjuPEmKeSBizfJ
ow1R0xASxc0U0HuM58yZ/OpQKRGKtYPYGjXZLGkbtiEmSJ8KrezPAIZvABWrPLPtAzJh5pg/3yqs
LwSj0zKW8aXKs+C8RKCGx3BEPIOV9hioPxnNLfP7O1Ud/8FuetrGjupe3tf6c1Mlq/Y/+S4CyW33
SMc1pkThzK6xIZe+U4sFl0L2ChsQOr29y3DbAW6pdpuVLt+nkzd64SOeVrgA50sg+3lh/CtpdDVd
M7jz979e2m4Mepbspw2zm3vrPjT0tvL2ZjxY0z4yqSgSc8HRF8kKHetmP9LUD/FWpoP6Gmzu+KFI
v30jC/JvevnFSWRuvZYo1Ef1ixhI5WcitLoUHnNLnk+vrZu08fuCAS3jWtlxe36G6IB6iWKZu2VM
lcup4FwToZo9beT7hJp2XzXsvyAbGJ6tnGWJ+AcIW/DhJs8JXTwNXUiCybb4JNz1esm0Qj791tQF
XpjUFPLWalCj1QS4fsoFJItpJLN3IWU1Zxok9OrnwyXNnkmC8u3y+kTotm4i99CRpj9WGOJ4WNb0
wx0kSvDWyq/jNXsBffnmPB7Gq6ZNs64Ob2fJtJu1eTzdv/BS96OLdOLc+GDg2jPoUZkbRVJS7SZf
cfs/o0YoM2EQrRfCBMPSrxFWEWEJmkNlcaXXK3x3MqpGCXlnLg+uEG5o06Lhb/m4qksgrSzLvcMc
YJOmgBILMGr6wmfCFAbImKEXaUQIslGoWlrSPsnPxAUdvMR520GoBQvJmwYQZw9jX14XP12+Y0x2
3cHvGGPeEQAls5ntDaFJ5v4VQoO6vLfng+DkeiXaQwm/HBxf94ANPqJ2cuEZOLzduC74NiBGjEZE
XtegkCJ3Z+zwej71SA/orYcTclf5EOg15sShmPBa13BQvW66hmj2dEbEOSeFPj9BK6T8TWpRRoUf
2o3BgWeO6gPy5r3JjhSU6CyLc9J078orwV+o9soh1T5+7v9qasMg08bzMSX6hbGsjgPfgBIxXQht
Xk+C+dBI+bkoe19zKRbtjpMZl5lhsDmwtz0MNM7Z/cgeW4UYlA9VwmKs8oAz2kCiyl7h41Mnhnnf
xEixgUU0GVreF9Sd0d7M6CLq7biZ3tSQroDM32w0v+aRRXIwIQG8Ld/yv+2OyTQVl2A2OwPMrOJy
H6g2fjLkNPk+SE0Xa4QEpo67qZtQqO1cODfdbYHFdGz3PBL/OCDS7fznKJ/XrtfRY7Zww0EWpfEv
QCLdY90/B9xUSzvZuOsLjXdY/f1gGAufEWkxCD4Bsj1r+ro+Fr172NrL7SUhf8qSugNfWIi/AFw/
fVlAlmE+2/m0FsM2lHsMX8kQNBfBiOVr1uKLMJrWRQZLdCtdYfhV1sQzi6rblFVFNgWDPs51UpBm
SsauH9yWmcwd+aayPHHZy1PMo+CvXrv1HD6C6dV7dB8r67pdZ+madV7AHdFBa5qT026ImO1gw5u7
tKKKaxcbPn9dlufilX10W7LS5Iam5ldnD+4gSkt9ptQsRINgTXaA12zt1gDbndnM+qHEK1Rhv4Rt
8RaOcpglfBeb+vsTSQamEy2m0YYgwqfhO+fmGxPx+NJ8OeOmiR8/8mKtffQFDqqevdtQbcqh/e6F
ekWrzujKKyihnfiOZEdLTWVAAnKCzDa8TSREOulE4HVh7BQhN+ZWu3cmhtLt8M3/gkzw/VWq6nMQ
odq9BBdwT84AmN5j2XnshfCMLqQqcQ5xs3u58oZI9sQyYVGXca10EKPnysKUMoZZIH0WoSLIKz2z
W325e9Mb3h0JAuE7ejc4jJzzkQOIeDLmFrZw8wGA5ISpfxvBb/ZRDot7iDztyX+za3Ie1GRyn4EY
2Axa2xPZbvtkPrJzmia6qLYZcCMRrCYGFHPf7iNZXu1A7sf10h4H9mLPrzicyN2Dyzwth5ExDyiO
Io04R0Khc3Y3E3IKKERT0WG364Em1dZolYRJSFr++mselrPcNW1uYdjruYcmEyHB+rH2iEYp+ppo
XoF5KT9r9I3AoeqkuNBnoqorNaid898LCpXq7bwLFf2i9mzkveJYuXN4TN3AlxRNu+c+Q1DGfXYD
EsGtjz4OnlXlg0goVpS2Hu0tSS44pNBzWHmhJIfJkGwaaXG2IDvWot4K2RtnBaIHkCZuFbXWbaP0
P7nXKVPfcvMqb2JUxz/fcNYxw6GMC0Wx/aRq0VdwWY90m+t7qZOXCMASB0V3sUHKLPFJfWLoQ8+9
8IiKz71gCwkGATz5n5mvTsLO3Z6xUH+/X02NjKZd1gSHrsWC1l4og+Yc15Djk42rqanhRYks6YwX
ck9VEKxv+pq17KIcm/iX3vqtwjQnYwU3iOGIRSNo/hJ6Vc/B7fVjvAskO0OWUoogOxhYtl5U6wu8
ami7ukubPWijKtoQZX+r/488WKUWBuTevyLsvjaHeqFq2oszeaoWBSaJMYYAPjc+4ICSIHcZGlmR
Z794Z/r1sXlNdKItLza7gs3CM7BEBcQwF45+KU8ZlqUAO253UsMZ6VMv2vrTIikFbXZjhvbjy5Xy
5iBCrbdNEX8Ib7ZFzRtt0vimXu9ZqTnow5fDAaj1hk0Jj+NsvgqaOO/r+zR8HVxwhiQIqczuKoS1
RajzU8jocqTGExqL2cuw29FgMWENvJei4jyeAIPOZ/M831MD8dmOKqTsUfLgafSgCWJFmSgH38E9
gS2HVOomxFs50+Bn0nnT6eUdVjkk8uvT/5YgjA0Y8Vu050OXy5p1P380DxK7nuBcRH7u6+Rd7jgU
kFPuK+f5JwUiXl5MK5t4eYQh2Fr69vXf74UzYWkxdWoynoZMkNFT+uXgKM2NKjNuoZPRtN1vwlDn
sZThAt8QRmC02lphNJeCihN900jswwmrOKIja6FB9kpmRnjhjvmQtWeOQySc7qaa1BqQgIE/213I
x8J8nFi+enyNMiHa8Ijlb8SWtLFxEFrEx18KrX38v4OjvdxW69ShN4C/0y6EUNmFBUD+aNMSWgyH
ASoAYBQY5dbnO5jQF0aDQI4iVxNHEXKTHKOfbXAvBKYg8l4dMWQpDZ7fDjjGLr1hRzKU9FboOG5q
uds2cpL+f3ghWwEro1jHtPJM5dkltxHgO1kRvCl9U972GnAOcaGY65S4SOKnMyy8Oq1sCO13girB
QwMo3KE40uoZpRFYk2kx1pbX2raHVdRIqp0uhD/S4aDlq2T+oAa1NC2z941gyO4+wHn4+XyURnIa
Q0g337YvcPNEMZXY4DD1v7MiUyDsYyMNr1ziLKcIH5oiU7I/R4gIE6Hfqsz2xSRmxYqvxoiZ3c6G
z7Lie/KWYcb4I6HCgovADkzuCzGHT7HTHFdyMEZW5C7v38ET3WI7nEDyLWf0b4tfat+tUHQ9XNp8
WeTrhZBJRUXg4/BEa+4st3F41O0Yj5Gmjp2J/GZXTYaKi9zGrAzGQMj/hnXPbcFEAq9LoQEDl+u6
BV1BP8Y2smn0fUMXF4QkaCLqR7edm4NAm2d8DWnvASSnLrA3RUgoZSczDot6QZ3pvuo2jbDc9FdA
h2XrR7EBkWMjjMaOw/PVSoOz4Gl7LGRritLkyvbmgC+WrF0rO8kISsSAsPKY4SRzYE2y5DTkh9/V
R+lGbpCc5RQDegQFpj59NmmZsCfJSfa3ORKiKAwq+YvdpvzhW4FR/6YKYDM6I+1LT6+1fLvav3Vw
1ZKUpnIb6CNDzapUMzw6BuPJcrQkTJsnC+1Qql5WVmfe6cY7ScgfsVM12fm0Ay8Hq5FzbmlX37UF
EYOyT9r9HibjBhTFLRXJxDv7JmIqLcBdzGGaxXlTohaM8XH+Z9/6alGlJb6dj64Z1IXaQr1WfENz
cYICZX5vg+vr3YX3CMCx8OFGsOtJIfnnboX59PMjjO4gTDcV3ukJNc6IZMhiC7lsPAXgVoQOAHpq
ckaFz42CZ9VQI3VSxFOqmgfxFn9cr122h6PmLKQcu9LkiFDGS/MbeuQA2vejt1OtIOUEa2yDP3y0
jVqJk1MDg92ej8Ea1kWeHOBDYZcrEC/1KIQwNzED3nL9CxednddMdXmJNjzdXrC7bMQPSkYfavS6
qoLke6kCpPXSXVb2CRwNGRnyjedNJynESy0yHZnc2cGWjKDWj4dQN2y8lizbpAMwJvlK6hd+Yrr1
1+E2en0k216+3reX9NvwZ3NJYzZ5LDMyFVhLDqTqvZUEeZ7xsCb3R2nUCTAdEVL8k0o9mmj5QVVz
UnXoG6ZhSlJvglGxBGX2MIQSkSF5DC3Qcz8L4irECX0rs4OLzVPHYh42XqU/olRU7S5AyU78FuC7
ntRReZ1QtLPNXTEWwlvcRuUeulZ9xFznagKKhQi0QKHuhHfyownLVXvU3I4B3PGeWTQ+bEKP41j9
4G1p2gN/lvccOSF5hVBGlTxa9yFoHktb6BUccLMgRoxvoJT6eODtqiK+kJYW+H6D+t79cZ3HqdtC
WZndHbcMu3fUL7eSt5EOMTE719BlB8W+XgCogV+sXNgvVgJA3QJkExY776H2Fkt0b/HBAlUodCod
xk7sp+ldDTAR9Lx2KB/TgXIFoS3WiuDVArE1yNQ9nleDu4ShzQowavyPYTdo/yaOrk5g2+LSHOly
50ulxJ/8YRRfaCd1NbT+C6CK4KpVEKMGr4ogbwIM6uHxh4S1ldUAhHHp2UfX5HIgkP7Zzcf/ZaBX
ZrmLhIlaE62J84vp4l4bPiTLiuceEedJimmJv8RvDw2wop4PQ8y7KzSaf0qrkoTYHTwAWgMGG+R7
WXTrh96Rr5CwwPeonxLfDHSw9EaB4FBy3/GRPNQabc+ErqZnlI0J9nbJuVXy7zEnYgfQ7B57Ns32
BUT1lp27nw0FBgbAUuiaT7ooAJ1FQAzcNpzFUl2udwMyaKd61ZngUXxp8oL6pv3U1nAvopr+WeEf
7QLYaMIibmco7GA4uuv9Ztfb+xVwm8llcGZPcnJ6vdLcmju8G6IbACZTMcMTmZ3cVW4sTz+BrwkS
mNzn5+DrUyy2c1l4tbQDrqdxg7F76ePumpmVIPp/2mXwZDCvAWwqSoFfBF84adpaiQmghVOyqLZM
rADx1RGB2V5+jmHFO+rxEQm2KpyrNIiN+VTy8dNUwbBt4ZV2p7Y9zbep9vmGD+lRHuWXJucSiSEY
Mgqf39UqXegYVUdmefWOozG7gt4mR8ZtdCcpQLt5U3YXtnfxvsJPKgdP7KcIEC22NiOADGS+ax+3
QwS4WHHL2UF8D7TRMHDmKvmam+grtoMJllFQDY5f2IUa96krNroaPJLpKxGaJ9n6vTmEXSsA30F0
Ue5MTnewLq4grdzL0UU2tXGCA65nuSeqGpX9mPLabDVaM0Z2FY1qf/Z6huB2/eSUtdsv3kQLWMTE
4b7YyxMo6ZVb6Tyfa83e5RX1B/0mfyilAuZdb7IMtonr3hx7k5xrxbK04MAMQHQkT/+80z6ey8x0
YC+JkP8tb1dWQZ+CN9DK2jZHByy8jbAjIqmr71N53TV2OUhTcKUVXxrpl26/vRK27FsGeOk5WypT
yvLj5wKTvdjAogpgZMSAdmheiraDrtLnrh/FO8FT5RMt0F187v4q0Um45oWYIKAjbKLH6E93+DCg
FTPNxFRYfUJqNP2Rs4io8HXQGwh0StpKBMixifKUFmcUPb1JnQ9e6tNZRUACP9uDtQyOdFfft5Ys
rQsWIdPOSf724ugA4iXqjOpjF5JBGRioM7km0f+T6qHXe10542yUgCCdhxJ4vY1dLAWE67K8SoVG
Q7xUi5uXjli7r8hc24BeGJSniYTIfZiPvLe9CG0HlXPTEtUhXMZzPxV2mewkZyfC8IBtTCf3qYQm
+dfYG0i/D2FFrTWsJz4Z+E85JDLPRtzE2oMGs7SR6sfN3r0pV5OgAzATUbQBMXRhuHxkGzuRX6q4
nWMu47iRUY3hJtYkCWdGsdBVSbN5ZZqlYV1C3Htir3nb8SXvBcWUWOG93lEsWH1taCp8lO1AZg6j
X1edG5FxEgz4j3rh6E8xdpRmeiNaJZXj9SV2yIYuBzQcw/4QwiibkcDh9EEbR2W8r8qGCzXiEz6W
Im8v4MlQRNkFm60KBb/9fEzpx8rbLQirwFwQDdkAXJT0cIsZMevnGSKUIaC009YE+3eX1eyjV9EL
4uraY9ktWbpBGhIKyua3U9bB62BgRDBPUSyGyvygCef3JsoHhg8M/PBpJ7COJgoiP1bc2igA//9u
tSprJe1l6biKPiOFiD4l4drAbJ5d5KTgeELdDawa3IKCs98Z8BlU74HHN0Vjcc5Bl87wfZPCjDuJ
/8zAGqB6kk5gCzHz5xM91YSFktQVmg2SKIHHu5Cux+HK1pLRrTfREpWDFMPwnhO0QP+LaMsfxF1/
n9Mk3LXIF4YoJI/prvXu9Bh+YTcaW7bpXDbYRFD/09Hca8MKCQF9z+KTKRBG571YB9Fmw95Adxb5
blfU7MJqt5SjnCDcTik78pZ8fMQXWUwjFwrCyhRdk7C75jS6p0Jn9xwm+8psQJFPerHeJgsKvczR
zsu+PYSPsvJydMGq24irDU/gtveGsGOmnPSWsSpeUuHOL4n374nw51w0f3qR3bPA0FINUwybCs7i
fXgeE1+zlADPc9kkvp2CGirluNQ/MQxYcm3rUnYxTfpLv8jGqzsVvzRXiJaHgtFXzh2evzeHoHzm
WyBvv5s2iVvkwmbpAnbNqm8N0L5dFDEuRI4iL+RKl5BcHKTJFEOC45MFgp43v1A3suQG98zvycNZ
mLcPRHu/mVSDq4/B2Jkzk+xHZdPxzcVF45dh9f+Pdey4T5l7KxmDz6Ak7dCoRli6Oyhs3IaAtkJA
A3+jvoMz1x3cLvRRECrgiFENxupytvaiNXWeyRqqlmj7zdMfYo8Lrlp/Sqy+IZXDZTMCWw0daSSH
AEz+1sKt5d7nrg7QrvySLxuYCyPXWH9zIifkTBqxJh8pUaZ0LWiCu7Vx/FpwOqVH2vXUF7G5qGDl
/4fNBzRFf7f/bMa0eO58pNbvA/LPme2eHW7GuLHMT7fC72AMf44yu71fKztdvAcnOeY5+qqfTqs8
vetY4HW0vMdKuw+4339J97slrMVv6YlkTnI11G6eEAGGj4SWYjqo303OT1FlNK2is/cS6yKeQADb
rtrGeBn0qZV6qiKOYMCgpASrkacWi3btZa1dG0dtvzwEuUH5Oc9ueyG/ajSCrbrnpZ7dJJQJp0Kg
SYx6MCm582wwclQwnlI8Cl+mq2NPyPXiE4a3E2EDx8PA9z5TJUDA2FIwsvKUcrTrPvzmgHBSNdtb
WCC38ieVyegNHvs7hlAGfWfg5jB/lIR6AosKUNFnOHObyJX8CEukYr3N5wj0pZpLfNoKuV1La0xb
on+Oc6XrF5zlMIVb6ZqfUhBFXIoWufQVUx21n+IGl5fLZ46yo9cgS8cJ43vI61290N5qXNMUgi+R
cdDR9xRzxO1r2HZuS5FJhAX5xjHft4N92u+AU1LgG4XsUeyLuThPStZYiDcXoR6faLgHezRcmEs7
nt90J22putepN7WxPfZ0d02WkiCMuaC/YmyoVilTI/xNqhwDkoc/0610fp9fDLixIQ6Gwp2Q2wbO
+4BL1HS+MUKSQRspqHSYhUdlSO3NzM1PqH9EoFVvsdxBdyALt5O+mhy/TX5WziEemyyXOmI81sPA
srdpOhYeK4B5HMOGDoTBjwQZFffM/9JB4PLV+6G/hRcpXcXSu7iUJtmzbNiTcq7Z/V0Oah4cXyna
6Fc6pZ3q7zQx1n+hGVv4ZN+E4egishxBqRvu3w2L7a8aDH0dnAdpbi63GO3O4xMW4M8j9rkUyC+o
pGp0gxrxG64oBKxeMcHy57/qg2kgauN2W1YiTiBbqGzQ+afFR7Yb1VfJryJoHIdIjgxQ1YyUQ6ss
+rCKnTbLa7HIKWjuoqrnM5BbrgZjXlLnOZt8dGz01nTHK4Knv7e6SAtKlIwZjJFzI0UdcwRTybud
ECx13ORDJzr2+SZt4dUPSVSpeUUBcT5lZHQKhOCZX8Pr9p6Yi4CnBF3x1DCx8veyGTzYpFqGTB2T
AzJw8pa6AopKobNuFwGmJV1lojPq6xq5FD7tPykiMpoT6qAo5te7hAlmb2/FH+63YfL5Xmz5swaU
oV3yaU8pdzwmb7BuDNhV8FuZeHoKvoCPEaed3/VHNyhQVoTOS8NowHe/7m/CskXQ0SJytSxRYXWs
SZmKaG6/mGI7kMbIKY+rTUDRMPywxMWBJRt0ichLCgNcluHwXJDGKZH40v6Q9MWKyxXMwYUBJPrw
FwHBbQUTAZ6KcMLyqr64EPTDXfDa9I6J8gwhojgYph/gOtRut6yDZd+scO/wY1w6PjJrfmWcZPds
CWkC3+MIpUsiXnzZBKOPumshpm4o8aQtZ09G+8fs3RGPqf/GgZOXMpkCLuTyzP0Ix0Q+0nEdBhWj
dYx5VMbZ/hrxspZqyoznoTRPY3GZo7iOW4zugUkBbuOXDOH8cWXbtx+Vt14TxAMkJfysS8P8byw8
enAJb4++Vjsb1EFpRN8Bu/OU1NFWCRsX2hnebKQJd0B3isE2E/IxzZtdD/9ZVjLUBNz1DXY9Pn12
Fz5n0Yf2vHtnCmaiEoF31Uz5A225G7fHP6BvARsabAbjyGd2Qulpvk60/fTw99+IY6+Y8D2UZJXX
D0LMcl9AXhOxY+VjCgeNc48Ab9AEjqh6E3kPeLqZp+NP1CypX1hf3XQNej9UfFa/4lQWcaBZA6eK
MdUdsZ26VKGefHT7mEoPgECXQUHHZMxV9+eFJn4MSSx3aFevY97FIDeTeuWT0/Du/+cL0Fwt3ioo
qajuV2EheMQJafro7KjqDJmwdi4RimLQxrOJbm/LOGaAe0TkePewbioC6q0H6lfpyzP05TjfKuqE
AKkXLW1rCkx2bPK50T8e76Pldj167pA/hHEmE/obfM+YVUNfK7YQsmeNy3OyQi9PiaD2mvhkA1Qk
rVhXAUyzDtyT4r3U9JfBHrnM5BBO1tVhIlxf4eTDWZs6SA4/mDZfArTKou6SZKQlOSnWFprd+Lkm
nY2B74MNaMkusclebwBfB9ywErQn9mU7Rxp7F/I7amlZ+3SgQLoFWILmQaNgw060aQWGjpcMc9RY
nsYmPFOSjZMY376CbhpugpsadRiOGS7i8gJrcwCkSwUIjoxdOaMlmZkAtXhxw3iZ2Bp84lfHVpdN
JmdULpHoKLbj6M4/RNfvxEGC8dTZhdUN2IUuc2W8r0irjnz99Rg0ibAKs4BgKShDVo2VYXhHnT2E
IDrhwQ/8WeOokslfQEvvhYcPpYhKDxoNC36xcQCo0GSETShq4+D3txJ1NRe2wR7k9kdAXQfmNCyr
m0fOQ9U51OnfG4TSRnULcPKhM+VMuQydQVk6rfborMHgUyB/oUGACSqLYm2jNX5wPPuzFw93U3Fs
gWlNtgG0dZZj46ELbb9at9wroPGrxUWBiG1Xy7hH0wXIpYIKmi8x9FRVtoAiIHf5HQwo+zR+JhwA
TRrDviKdjyusMolrm1kkLBPc2q37baapVBXoLIbslUHnpp8Kch68fHUBwUSLguPzHN9NHmZqqPJo
jVYeuX/XXahh51qHjra8/wX61wHRsJM4ir0Y266U0fm7fNnj5c0hm7a6U2FDsjjsP3mwxhj4g8wm
OTp0PJvoPvdwi1leVVJUPY2pxXTjMRKMWFFE6poA1t0pqRP7EKED4urNYJpMXLiY4OZItUV3mtIX
kgS34emZuA0zCN53yhRJ0xEsZ19H8R90T/YkK1mnwsftQQddbOyZn1KeLcGfvqhHeSufc7UTrsnM
kIDafSlDPsJMF+e4OGAkNk5YJhchCsHXYxdnEtB2NJnAkJogWjek6lnJYeduZEYiyATDxWQ7UEh2
85RpPWhWRN+UORfDXsjbGuwqxL9FaBugbOpaCNH7jfRU/CKGakW8giHCGHKLRhG+Avm9GekSgN9m
6RQwNW6f7kuDlyrlE67fXPPujz2BRQ0W57Tck1hX1fUksSGQwyBNHAPfSsPGF7LcJyr62Jrcobth
WJNwaqg4b2qgEnsHxHgMhLYYwrJJFU373XB+NBZMSzWG6IcTBuQPBuHzYNbUz7tqQmK+3Yf0AL6p
A05h3ViKQRq7FaZGn2xVmSxJex/AkM42a4OJ/ohm63E9eiTDcBBMcrncdJI/rsqL8P9IjrTnwJpF
lYIp8CkzRqxV4AVFlYS9GaTzfrptJPT4LMnqJqxeNLQmCLM8cC9Oi+r4zmaClWYixZkBNzsqKgOC
k8CtKZTMlc7JUPgecncz3Fw5En2LwH15rPTVjsF8900HjeYcJenIIKzrKl9hr9GBQ2cgcOWBrSfj
NIXydf0RoC/TjmH+xR4DjVjrUbD8S9oiC7+7B3BbXYZOaFSoKJdpqm+dDTwIo7RS2uz/AA150u6c
Mb/zdP9LbBNJRDqrq/zj2fvNZyFUyoK6XHb3arBkVUjaPVZwOpP3eYx3tgzLKKlKzB98FNdmfSnW
ITQI3dhmcPisCBbR9leFoYU7Y67n58brlPdN/cZlzKfOTv3Is6EQ5CI3yVpJgagKxPmD1oKL2aXP
agI6Bgnf8RiVDun/tchxb2ZAUaFhPKRdu93tpKeDiDrSNS7ayPQ0s/ug3HQQylR9yg0FoD3EOAEI
qrVpFizBj8EQ8FMAn8ANTs5dUKAcLUiOS3GNLU/cuTrSwcsTbHGfoeEmvyHQnnDiPDAJeO5mGcQE
D4yISSc9woYwWNv0aHZydbgJ9pSOLEN65kJpeA7NATU53EY37S/5ODr6EEVExkmRL5s0AvxoI8K+
EA9Cu6vCudBx3Wcc0/eIcd8wdExd/xGwmgt4NtyqyiRubrjcGjwvTFQElEBk9YOTfgtTPjWtwtpH
kjJEwJJkt+8HWiNmsu8Owy8+Cj0brlqrkf3DpNjvoHrk6yoBJJTnNbLR1htNFLtYzCdZSPHAEQHB
WqDBl5dM7aLwCn8pw2VMdZUNrIp/PMMbgkefvC2GkRNbuvTS7Txycb9zJ4NlSyT81maGVrMz0T33
k9EkLbg5i5rHbL0Hts8l6Rd2pAre9K9vOJvUEwObqVn6tnuy749K4V2JkBB94Ad0no59K3/UyexY
nzEVVgfwO5V8eXdSB6mXQ/rbTHl9UJeab0gvmH/gKxOtg/KqPNp46cpcpYmlw6eAHc3EG93ioSi7
A+IPd7nrlv7o76YMrN0+m1TACVMNSvXsphbDVEK1HF79dB8LWxyIet4hsL3Wzi4im4nUDF2fzl8T
8g2HvmyIEE6tTC95uaCM+4gHCjz1S5TBtWF5NQkDc21U4J3/RO+1eF/wXkC0cz369g5BYApdwW/o
DUOugQnp/7Yw8UeOk6KGxCSa61pcR2SNjQFbbOFrxh9jqiRXEfV6VM+IuTRfMhpu7wQV4Y69V+p6
vNYFy5uI2QHOkT57BtS5kqNrQvh5KOeSnnC4eUt/DgLAAZALhFxGlY1i5XlimExu4BKnkhZxksGO
3+jNgEnY8TEvkhCtRXQcHypMyT2b2svCF2UIX5GOpaKSIyByv/virFe/0SldYF+7hY/GaliE92R9
LrWsYKBOerGUPjLMEDt3cpeXJREExmXSC+PkOYW3c2XR+/pOQMRp+vhM8WoTSatCUguu4hOK7fHs
/RwHaRaXVJPeCuTfl/6QEl8xEInqtb3MtLX33UcsPkNVHZTkLSFl2aCG+mbVbTnqSL8p8EOtazRp
5cRq1FpRWoBdBxXE7DRokVgnm6gfaMiiKwV6NTB7BRlULCxOnMSN8h+dCRoZb4lMGJxKf5CaQf2C
BUEoveNnllPEu1sAkdRXPWIXtMy980fDvi/qA3gqzg57+kUUropaRKvFCKCmKP011AIkfhcHQNBB
ZvhWmwI1N4U/tOCcoKmAvrSW0JUg1c53lMJzkfiOMz0CBwLjsxahRoLKaGBvi+56DMXY0NuxSapu
E8m8+myAWdp2Rj12j+piYib0jQzKF0MV8fEgtwBjwHtIz8mJ/2NZX4fTexoVaKljEVpqUnzMbvvA
ThV9xi2cEpFJ2OGcpJMGSL6WJBYBlCGxN3dPOpGEirW/sjgq/2oVcIaW6HhSjsMdAnQygc1yL1We
FuPQsy+3TKAsIjnn1TsZOFuhqH1KXmnBSSRs45VxMVpNO2ftLA226EA7PfACAp3i6G7mfw8kkdO/
/IOYtLuONxchI9/qAHrI0IBwLc/TjmHbJ/p3zeTSBGVbeRyKD8g6n5FgaKPKTM17/AnXB4o9VGHN
dfRKifD029GT5qBXW5umQ222huJawT4ivMdEnHFitOkwghC2YyYN+TTVR2FP0YFlHRbHfk50/E0D
1rnahowjmJ48DzOuq4dbWXXwJtFON2GZQwGkPm1tGHWivzyH4ItJ+eOOP6CU3/ZftrlMiIOnDEBE
PxxOnt03tZMDq59bTIFe3cEZvpLo3KDc52+LBrea5vQGdmjf6qzlrRgZml/YNt0ktvA1XRumtAlM
ioQiIy0J58o1MKvlhdctTtSzM9GIdd8qaiIJ/gaTDfNnB44g9Ig09AifvJWolSeQmZdLAiXTM6xs
Kyasr7UzZonP4lhEgNYNrkhWZmorfoOoo2SID1yjI/Q24WJMn3A8SLpKclAUD/Xmw5/bfOqEe/ux
ar7WX5GOpcvaLbjM3RYMrotytLdTP/pr+f29RiIANopXMqqD59yd6QY28A4Nt7uf+MNqY15g75RP
9pZhfQn8FOgzOCtFV7vgCc1sIHN+kuKlRp5GfRViN0wkzamaq3SKVDAQtT0hLIA/3zgqQ9sZtfhD
SuULWm607rp2ZFtV33xkBcLsEwnoDZELYmQ6B/qVzwAzKlc5W9lbI4E8YCGCfJitP5lfJ8UVi4CU
X7/buIywF9w8sS1Z3Xb9HJcj0UgewodxfgzNu+bFpyWdX0hmD7lGXfOwbxZ6nN0FR7i86NpLiIH7
0IO6hCSExiKZEO054GrT/XReIshfWnkV9J8Hli4spK27lt/nDjj2dCy7YgjYGw540IA5wJpDXeLw
ISZ5YEV4NEDCND4Qqc4gZ587EYjpoJsEREqwuTMEGXrzAv08hYKEOL9yokmXCWtOjhrp1O7i1MA+
U/IxhPMFTk3Kmg91wugA9INcKHjBRUUhzkE5gps4wEM1R5PuWLS8PISRHN/xnZm07cK6y3KkcL2O
/HJVIhdwkQ/KLGJCOmTpxQIo8h31EXYj89BYzXtkNpr/updosojPQpByyj41P1rbt8LpGRDRm0QD
VhniSz3bt50K1sC2aUVePBKGpae5P1cxE1TqUZZRwIkMJKoTO6JTkfnsaS0gsnJ2T4sVrpKjSEl/
bOC4aKSeIQmivTeWvWoomi+piNzaG6WPdd0q5aa9Wnv91inDz+cWvbbzygusgbLGo86X/VWdqUeY
lWov/+HU4zWT7duPknVFNfIe4HH4PQ/yEQ5N+eaJ3xJXlQ9hIYkaCms+ps8m+KEHDpcjuJy4BbKS
vH+FgCTjrBR/TVBvXjq0pJvSc6xddB2sYYvNTeb8r1L/AR2vxBar3WxE0EyuXTQLXpEIC569iiKL
XBriffU1b9hBk7qjvjvheZHJTW1sB1NatMw8HH06LMMiHJ7z20zvor6/KAaZZ0ttsIft8Rp+Hk8z
9lVxumVdvg3NR5kLQQLC8RvU2mCWkPPgdK9JREDq41V7kBQIspR+xESRN1Osqzud16TlRxlLRbx8
APmvF7v7J/yd9nxlRgjUtsQ1KjW3jaXrhrLLzg4lu8RSi5iXSmbRFkYrPvlCIQnQJYU/evhLIftU
Q8DTQpL4JYo6qYBXBpcGRtY6WoAYVOWoT7HQ0x43ZWV2G5u368mKWHXdyP0ljIg9uL3bqbE/3l+8
Gdl0CQoBYrRL2AHOPsonYn27gq/mKUJsaHuAc+xXHV+j/6PhWHlG6rR1sPrVmrE/TRjZqeQtRdQX
gf3jXi9U50TjQTK/uyqvaNHoTcyiWI6UK3rYDi4WQMvdxQnAvHAYZ3bJYQA4fDjrA7c79bEX9LQz
TtrY0HI4di2FCIZrH7k/juq7LHxVYyEJblIsp0jrp+ykpC4jrIOrPQGHtmpBJZ28MLpNeVxv8MDJ
cVGSV6IlGqvhJizBBWXt7M1guEPpiqFltXvZtEYcJrsTWftY5j+GkpT5bz3katIiLhsFi/N9vZMv
tlu3D08km8IXYJOMS/L2dB2uabv9oqklOQyRbrjU3LhhEEAaCRnktRdL8os3pAzoyyfLuKXsy/RX
NiuZWlXV6AhSOZfuqGzkSK1jvKMLdDv0ru+A6zq6zFBRMbvZ3dS2ZKhPrA9s+WoZmHXEt5eNtXtn
zrupg9qmljxBtjV8mfd4C7842eIjFwmQXIe/RVABwP01CDiRYNnYtojFfHeTcGEGY3EcUumgIDN0
7QvRAvWI83dHpcoO0RE0ki+TpCNMNVsZ9lOq3NLDmiYNQMYICxZPuX0EQxmN93wl8dCFoGEak46S
qQp8wzhfpmnv21/5R4wlqLd/AqN+oHky6cH4zt3VSYFetXZfrWUD3YWB3WWdEk47Y1/eHFB+Zw8E
DCqpsfxzXibFn/OdXzWfVAD96LsW+6EGYPVtYS/HFc8ljtvWGmd1nBZktK5OjVyXD+Scs02CKRal
baH0xDTTr9nHz+Tk4LPhOiiOIiIutHThG5nm7k0HaWvdbvjD1li6H6X0TQmOsi8mnu5vfYlIF/6Y
hJGDdofu49WN9NhQ7jJ8N7K9WiHxz8lQTYaS9n9k4nFRlSHB9e/u74ZxdF1brIX8wE4iQSjRE196
7/N3LviAN6MUynAL/xPDabO0RPQWs9M2L/etIsut7n3mu+Amu6WPvOmKz96Ek6FlDWyaluJJAXko
C9JQpTmIXwGcdh1TMg2exlL0yQf2mKmcbSBOPKF7uujr6UlRJ1ySgKSzWj8abNqLZsVvI/xNsOdo
c3Yclp/BtylcKkORlqaXGDdO83VfisrB7/0QyjWjD4Zb7TuEL58tjrzSQSUdTUQWEq9LYfGwYs9m
41yC3a+T+qUlg7p8CWSpqKLwZA+QUVlvvb24/mSMnH+1q0xaFylGylMb2KC726lN2IfgIWPgbaPO
hip8i268o6Jne8N/46RaLHm0EypwZzROhVySBBcNmZAVhmyeH4K1jSpSvhxdifgsWVvbX3zTSo/J
k1rXKF4hkqCombmsBvnRyNuB4baD5zUo9XeTn+U9kLiiLb8qo35MXnru/QK1Cyk3G/dcwOuNUl2B
CZVabV5KLax6C3JL0cHmY4bGkQuI2r7y2EtLorj5yFzKYy1tBgggSuAnuAQYeMLDGowM3K8HqCwu
UMxGMHoZnE/CDXb0oyFLCXk4STEbsCzTYREjffwjfFICJiIjbI2njiXsmGQX4Kxlgl2rjqE9Mmid
KiefKUeThpDx8qCibh0+CHQT+qNYe8O3QkA1dHav9sOICRW9XCcHuC3VdjGM6oXQXIVq+q2M7gfg
tE4Sz3QYsAUhIpH21NIZB2N3mYbElmyV4AVI1BJG2ze9s189aquw3J8LfIoqHTipL1yEeJAigAUy
wVw8aOlBPxcwEOMJEQnxZEN4DYPZaEQe1s/kNfuN7XmrzLz9/N6NcWSw0BRuqWMYEqIygZC4y3G6
hAowAqs0EGoIPUnJbBp0+o2qElDLb0V7cyaHljEiR1QI/UrkAGeyjMgjUArcPF6yLveUzjO3T4Qv
XIiE0jSt+Hqyp39bo/ySi4sMHDHU/64p2XQW9yQ/YrWQaL+sq0nGrIWGlczEnDvRLAMCLS3ikzCX
oislXashkI9/S0RM1NA/35eChCn8LocyL+X3gZ1ezOmGnzefiJ8m5CwP9Vj/6QkaD2ix077WdQ7C
mGUmL2mapH2XkJtlTfoRxZZyLFhOa4qwa/hkqmzTke1Iw9fujAfZJ+IYTWJUnbIBDn68/5wMmNLC
CTBmzCGMtpE9k1gVBBMj/sdMOT1ZluckL8av3Jf16qXCN3PxhM4MZPkMKRQ0lERjjKAhRuHEVrJC
gS2FWxF/aeIxk+UOyJQ4uspdki06oVbAd8STeFwVetWKXBMJ52/rZ4FwFrL7cn8CXjobw1qJnTO5
e3t8mSGM6MHU5+ay6cBptXdihHVjCT2j3eJUr7Aq7sm/Ebl3tsfGPR0CErqHbM1LzjWkUXKNd4bH
FpgjIuRhX9DKyaqQ43MJjpYL2W5r2nrgovghx5gifBlgkHkkaGjhc0jUikyFBlPmTDMAfI+66Coe
njtlgSBPL9kvGseBvCiYsUfYIM43aJRYy5lawY1nKmH9EZSRmpnV2XJLyDsgcJRdscaBds08F+pi
F/As+Qnn6dbk+bWNXKQKg7itIY/msP7TaL+kN1HsJGoaXYPLHDzvEFRCQWWaxFGqdsgWdMTYtfEE
GJXm0pCRaGVyQ4wni/XtkPK81zSmLKUY/+dMPmGfl2JY0/3OJaOzq42BNHDqZaVfGtKP6F99GNi8
pvb9eeX3HZcgIgyxxR/BOdyabs9J2vUbGjR0qUCEzFO76ksKPJrCwiRALcYbnfDO9OrqDlnHFV2y
rxjI0j5DAgx+ONAmPdJ2ftCDEhb1gmsYWLcySdGbFuDXiIj0zd+9tnm/WFnV5YygR6gEF9xsAMoz
3IXMlQPTE84t3V9UKZO+VjOyGSsa5F1zPdSpTO3xRWH3MtZPCppX6RHRpL9KZyknYUgGb4VBauqx
0vzn/iqnyt37oARLsMSJNyLgCOL0BfmbJeRX0qfjsaJj87O0RGQ9O2ta0WgrowJzgrj6isRFjZzb
DOBT3fhevKW2koJOWVXKufGakGZnV5UYK9Zm9H/ibDeSf+K+7583/bkKHZIQPUd8ExS5o0mXUOeA
+D5nqsotku20GO+RLs3NBOGqXUF/74qbKBwv79N5u9yiU5bEIDCWbU5rpsJAzoFd4IkACl4dYcx+
9non4sAwWF6np00M0gjOzB07hwnVDhimUmt5ND4NfoJCEK928PFFzR8ZA+QVcyS9Ku1XyfVIjDOz
WfjJkqpCaX5MquLX3x0Pa0MmcJy3TYGSBIeXcs1X6Ml7AUWto44S/o+2eKYknzwWD5SaJnC8Q8Ew
9wSiSlzR711vtdYmyppr6jTkPYmLbqxUxkeIwKmPyxVqrnw2gNUa7Dbe6K+0OqCfIV6bnt+Aj8Yp
ecJKpGBMWq6bP5u6aZODgrHuQJRx7HpsqinHbYQ3LJiGrBPknI+q0aMMRjgD6e5JQYD8IZDanhTp
bOGAHr1ubcTSUkJzsZqHQEMnI4LpDGff96le/Zkp4ySjAEp42wNcteHqkDKWrjzrtw2Oq6cHqezM
efkISE5fUJXWwphX5jPehyU3C/hWErcBA/9sMraX+eGcMz5y4F87+L/SKNzHDygOg8qC1WkHRxoz
z3eN1hoY+7NYp3OxA3bLCQBxkjm91NZ+34Yie7GlECnOvkwJzLEsmQI2dpX+uHF1s9tJ80hWdNmc
LtGpHUiG4wvMz9cYyAOb+RVFfodGdqBKx4Lgnf1phxAr6Ba88Y1OIeBH/PQFqDVABBOPVmaaSSK0
xSziDrkar0JQlxXXeWfmomlhQ7Xhwpi64gHulCwieFbtirHG5ycL4sqQVvsTvYnziKIsRJS+5ewY
v7Wru2jsdfiyUgGJBfiV4XSBLhtpOqOrJomAFGXmuXxhFn0n0hsBL/yU4clOmSZiEFzQiWaa72bD
PSV0T2pxXSHtQ4TqvQceI8FBLxQtXM24ew0Ecqns+eM0w1uJElh8BqLQ05rG2CMHKpuX6XaFtDxk
Pn4umJluRFVMKT3ejRsvVmCd09z25mRNIoHzesPwMvvIzgvfi6dxja971UBQwGiWSNvWAlioAjKA
+K9fiSx/bLUOOR1Q+RGTjXNz45QD6Tl7Y9BnHhNzrXN1bWkfnGJy4X8i2dY1Mmj7j9+Nz+aSvblB
RkNwqe30j2nGlLNoP2sEwi1xrmApa6WIZlSOQXiKYvoBA2G+rID99KTS4pFkqjao+g4fUUSfcoX2
MotZa9UXrTHtL0sNxXl7YN6C+Gg3zSEeCRkb5h5+vk+WZSUpeyRZ36sN07rDVI2iQTIm67x123Nk
rVuSHLRwSi3ot6ZCOJK/HgaGH/2DUTnrxHctUmnp4CzAx4JuawBwbH1lBYLZ/BPXIGMw4YPnJ4FJ
vr6hVhnQ8G5jkSL3F0jUGt+ZvUSWUFqG/Rn/qshwkTCtG/5SMNjTyNNBuu0Y95v1G81MJ89csmY6
ix9VlsqPVZzQe6Hp+hBETVyXxUBJltfepz6LghFfDfeaBNJ9kTgtUZ+ovOWWbVOL176vCG98mVdG
fst9dUH32WTmWAvAsOL6U5HchAS5Qzc18cMsbjv8hd/8HiaL+QxG9TWsiKmw2esthSZDYMpUWiy9
lDcQGrxQKlUvLY2w+XUTybRJ2DyuQB4PX7CsFbnobcq7//8rx/L+yKHLvBYDtl65IjLnL2aYrovI
A98wd6Y3yZva7ORs93XL4LgxE7helWOZLaF5kLpb0dnSxL4l56JAj9p+YvdPi/c4420ZIy3VNEWv
a9qX1QfSk4PBVdZnkD19tLQwvZ9airaoe8rXps8MSFE+2Ssd+efwfG84UMD+1Zc4/qIT2ceyXbRT
H7ij0xCHwmHYO7POvGli67Pda51WSQ2GYEtIlyj9/il4JbwMw8YvmkOkxh7ai9VRMjC5I8hoZpab
ZvgvFDDuu1hEiQ0MSlZ7wAV9Msvkvptc6yZBJQkKQEna7hwtljxgBZbjZfNWnov1Q2m3+gl53WrE
11Lr1wNXY6YeYt4QPXcFDleU7CBgCh+9dMAqhboXBzvMDRY77i3OpopreLlwIqRCoftSfjPUeCiO
KGpfDPfEa2WYtG2dk0fbStBFACtF6R/hiR98/ejrXE2lp3xyUeQpZoThdCbpxkjFJ7EiV28HlwFc
lCWCisRYdD0QjX1ih6m7fnxF2isrBU9JlT1/xd5xHb7L456buxWmzSupx3ttUWjpx0TXLSlvLe4t
kTVYKtinX+A0vBiBqg5YVmXkM5pC1juzUia6CVaX22L7bfe+KQFtm35De0wU4L24j6UbbUuMPbzX
f3R36a+yn96v/QrsSBxApy8YsVjtUnHfwxrrK7Ob02VEJchoWAEMi3QTo85e+P9NeYfeiQg3HEar
719OrnyYkT+rdhwHS+DVVoFNK/ZgcbjMCvdkBJNuaH3gHyVxF+eSURsQovI2Zt7TmEwicGkLETk0
d+OytkdUEt7oyG1wd5xP24mm/S/97u5JQN3msYaJLccdK4M+O1YIo0gLpk04K0kZtbb2DBfsUnoq
mFPQ+XRRSwBh5mJU+YtD7/Ve/XxuIGaQgNe6sQTPCZBb7Goz9Rvj5RtPrRG2osoYbIHAXVjwgfkn
PgmJFb1e6tOH1/ZUataPXoL8IrqUWZCv02sy4tYYxw64nIrQU+I7DYbE2O7FTVyoFXgnBD9oj2J+
bZss4mqMel/1//rGX7zacVIo9p9JaNK0cQ2sh6pItoR73ssqEayI6L3Q3XfZjwMxfuBQ6vhbUmbm
KGxNLXizwPMTV60Wk63kbud+6uMO1hxw6wnR2y0xUDxBNYwTnIUpZJcIqcf8NJBM7C8uJU7uPDEv
W28ieBqRVtnN/7ozqJ7RjzhIwhhZTMknDqgK0oCnz1h5Zr1bLUmD7zxR7wxBYYnF2LOAqm3XXifi
oEz/se6ry2q1FZ5gsYsFhpc8mc3n9DFkCpto3K9jHcU+fezybV061GPpoBVpD+DJaGCZXmA5HmbO
ZWN8D3UETtogQk0FUy3+Ltrn4bkLaSLmxPllGaQlSaaK0C+4FrIU2sM9Sta7N3s5+SMPEBxoS+rc
Bdh3w/vSYx+Vr2MM2QgUCrKvkjx8cUifXfcepmsK3bB/O7MwRmvvHvyZWV2Km4aWbKBwCZq+xPnc
hH9TMNP3HBq8GyhAbBJO1Zw3vIxxZmOAZZZ787E1TOqwJbBkEa4uJid/+jzCMRTJUuEtRZ58fSU9
1bBbjZd7w8bgaPQ9sflHLGFhLA9HuiQDYB5OY6zm0KIQoNn3uG2YHd9iRYgUdfT+sgYcp1j73boO
2boO23t0y0hoxM3SFeMpcq5dQYyJZRXdgv9CY6J7X6QzzLBhPtYZ+mAMb+6jKD+rmaa43L+O1ae1
H1J3nh3C8dJaEadkpgVHfydNYEJmwLLEzERXJrLy6V7vzngiObBjC60wqZqo5IJG4b9DLn4jflHB
bL19OtL4pWG8ZytuehxfAYFUg/QhnWgO8pMQkQkmysOLm1lKd69fTEKx+yOzPQ3EgxgUFazG9Xj3
Ezgf/qs2zoJVfECqw+Vy0xv/0KrNYBxCcn6InfxkFj1iooHEkB7Pfe7vd6+97Pm8eVWvtvCoAzcV
qVEA6/u8t5LgkWiFgXaxOswDLs4fmHd7wQ5Mmc1/XRDNVjFZs62/Ll3cjTcu3iTcGQywZgpRgT1P
2vMAFPm2rGLet7aaognw2IT2s20YZG40vxsy6aZhC0IchegAZZ0bF0n9t+H83+N5+0fQSrMXBeKB
lQWvSvXlUXBua1a7FW3ti0o+C3y2qptyO1F/W2wOKETFujaeb8FqrRa204/LpiYHs5ybu3qEzqPC
8QNFCMHHuzCnnnFhcfhWHcfcjjtzp4sz42oygIlGoe3KjCzGgwXBqTMbB8TLMpUhiwfp25JqIk8a
k7T2d5+acaDvN7P3nDLVXfeaycuvWKUGDja03G74Dbf/xXOfkIrADDNUf/14CCZ+jEmAT0HN4au6
nHt/YsWPjIYkkgY26VJpkdIPvy2i60F/e8kpzouvXhZbe9xezn5hiX9Tnej0NfjYUldHKwVQNc2Z
J2pzaxEIZsBqe05idbT8EIV/qE2aQwWLRYCoLSCqpE2bP55L+Frun42bdpCrFipNy8fYJxHOePxO
V5L3NVDkjEj0plr4mQGvQL2t9qvws8pyNlJ1Hzctz23u0OF6PJQH0Sr8nLJ+rJzbHcZkqhXVyYQF
HVWzyuJNw/HO0tEkpSM2e4GCEE5ZVLUvb324StuQSA1WEF6/AfVoouQ1NonZbQIoeeDo6kMl7k7V
UhgrOM66ZGdcIJPeOaADccrjC41s14y8AYIbk9KUm7FhRyIWXjLAqY40xND8DMi5H41bGJN6S9+8
l4fK97UcK3nOsb3scrxIif6XRPg2OPWGcCAxyI4NIuVmXD0T+4wQNxRo80u9gLCEwNk2w6wrInNt
wMnK6denIYxh9YTsaICG6hDnt6LO0xrTpzJeYtfehw7qQcQGaphccfSSal1wVoqvCYLp2NgpaAn/
M62vjvtoV5F1uYxDPLcpxX/d6CRBL8pIEWViyPSrXdWfT+tj7pCzk7eic/U0NnsYTH0e3e0UjpoN
3YQdfELrRWcLQlMFvQVC4qZRsx7JNbvNylp40LDcLylJ4IJ931O0dYTUhmHwItl4gHX+Chm160TQ
M/KhW3FGay4zKVC9Tgk0ItbrdfNQppS0mLC2PG5pDZRmhpX77V0iXHBuEZA6KE8xhpBAXnuGm36o
bgpqlkydwihUpxvIzA6GrfgyNyiBsX2vJR6w62T4GLP8bsVGy/1z/qsPhZONFq/SUZy5PdJdLIAG
kYdgzfE5o6nYVRfSKFJ9fWePyuVYkkboVMTc/3uFyhhd3+9ZYLUoUtZt/PZ5t5HI9n84GW7vnp79
JTQXegq9q4WDWXIMf9lEQxQZ5SRuUXlJiw2/7eLpkm3uN4rrhja2mF36IWT2fRKv3LxiBpaVRVp9
4XyjuJdbeAix3ZnN5gaPhFxOqlrAn/5VTBADk1jixdJqjDP31X8RVOzr3NsOT2B6/RcecdZGv+Rf
kcJpa/I7AmnLGueHzqQ9XbDCItFLTuf2cUevWnHGWvCZz5YmSnrsecc1EUj3MKDhpFOvuGhoNNar
JZimuKkurzQykl6FoDcub939GkQ0amOv7WxF2WuypRXpV+nGsrdGv9jNvY9uqoLsRQSkqZtYMpUM
IjrkpDr4V+pbT1ARqUnZ3rCZPiP4kMq5G/r4WVs5fGN6BBkf8bVo8mDwSnq6OVFujTe+u/KmYtXW
6Z/ml9y5Wpg1H0pAWZ1p3UojkDaSnJ1prZY9kwW9Qv9nvbf3lEHsTlQ86I9i47D2RDv3m4n4u+Fv
Oz0vSExZd7x/mj1/lrJOoDiXsDnHheFA9Y2vmsuZzsgnxgSlocRQhCpsLXb+sYqNAcaAHq6tjd7I
rtVidxPxkQFD06Yx3DHpQLgA0bQT2C6+Z9478pyKEMKYfP4hpp7G55pIHPnfZA23wmkCvjS3LixS
D7KuuqKWDW+8+NlJPrU8UzvxDgkNQX+M3y1bAxSTbj/0Ch0HqS1dvaZL/YvGg5MTypT275Ptnyaq
pFSHlZGmKwWhf/DT04egQPwDx3Pi+dYbtTi+5TEFWWKUc75FJYdQyewVyd21XnXvX8nk9EjU9a7r
xcahZJXDx87vVJ1re0V57O7cEz9JidXPr5picZvY6gOPh7wf8JSHtBBKSEfpMFgBpMuqHuv0gnDp
WIlfATILvjjwyihZnnLUceOt9FLr2DeF5Q7TyPbeYLTJatC/34ebA5iUdZLs6gPUbdks5NOoR/5W
oncYuPq92Y2Xk+OEda4iqKMu14UEEgXyaczviU89Qia199S54AxCieEskzVmstBocsZ4e7elAoCT
lCUFHr76dieSww6nS1+EmIsgeMjFEqxm88Wiafpb1x3c7R8KytUxeVdHg7W7n5Oj0LsDFNxeVGOl
PbmjgfOAi0LASl7IzpsG5Bb7pm2NgQWVrkzYcCyDlQ2wkBiljNSGtlDImNr3S1pjDPvuk1KAz0GH
W6BnoY3ww7QDyZIHPxmLqgzJFrDxDi/tGEpyJFcjnw/r9G5YE/D4RHMg9X3aZG+V4sWqvpkuRUDe
J9DONKT1A58mTG3Acgut85cPdRa1+bdczHwyI7raHAsGlzuJ7gHqcxdpFESPYP8xPpP/SO87cyiN
xXmTAzQOq0XA3eKMKEd1O7ZoB4tHSwbCBpN/dHDioe0pv5B1GWCtGBKgUvncTojFDQMJDCm4WLb0
05pbDxVW0Z3nvVjq1QxBLxNfibxD4YlOi/xGTzzbAlbRBRud+zcXtyjyGq8kCsYZJuCr0KLX8jFc
EQ8nndWv0BuaYnN+t1vYpV8+783wMXZGovHIaEMc81Au6AwY98xQ6UToLMCL1/Bw2bbySxy3BKPx
pO4IGs2NVGRsa8+X6w7E0LHWMfd5+JqQDNBlpYydYhuq0oTKi1wh8B04W6S+y3Fc6el+G+yRPy6I
lrpwlFO3lQCYJ44v1h02mCBcgUUI9hmqmN8YMpfdDKq7En3jRXQxCOiUWHzoREaFkA+5XGXnRMnY
IsDSsMKDP9JLflBl2IDL25OjfnhZWgoBvt5mXMCmS7gUBgaeeoQcLPs7uuh6NH+S7POW3TJVuF19
pZCqP/uiyVEfGPgwYFSLrpZlovlGmhnq+Xb9e8VSONpm8gdMIz9sC/OZ2mcWJz765tC6CaDStWXP
Ax0Vizk9EZUVC0HnfFGDmKVmdCVfzFz0pR624vXMf194O5kh7tpdPhOZXR7QVAPTGq+JeL6Vqdiw
3X8YoSxStKa91TAOdUXiDmjxj/i6FewlS3KeNCQc3ZNGMELBc2b42K5nnB19/u5bSmp5KLpL46yw
r6Ksb4FflTMPV3/WjLaikjA/q2ZBk3aX8HaZXi4RICeytiBCoGKNnOqoFSq9re0zMqRQGxI5uitf
+V1+d9R6klBwuU8m9WGa2aH76ffZSNPzUxwnwcj2WUkE4Vi4VAgD2zlIp4Rb+eE0KKIq0OU75bk0
iFFLeWn9HfP4oGpK0fqQhhck6NZA2GU/ilXm15OVzHA6Th6gULdkanIquBMF7fK1qd5QtQ3J3pj8
35DnSMv5971xqYQfTcy+QLZb7D8e9xgR5NM4vmylR8tXteGhTR6C4Qs1UcEq2688/kK4ZJ2VeA/R
uKFLVniZKKtd+rz4GbwozBLsRDuQSCZiY4cGfP7N2Fym6fWugK2An2AeU8wJw3zz6d99iennc35h
Q9sAuPKy7AIz8GHhDhWdy8grV2EUxUVT5pY/OBndsRAnD0I73ZjSImqi+WIlQ4uC+aYSXbSvoIXk
1Zn+1eI6kdMOXf3Mn7n0OMKB059HU6fuEv6sVVp8dwbOyKVRCFYHnhlb+xHeajvPpciIGzdtGk0U
TCKtzrFWkVkG3+U1XJpkN5dSJbE3qyyiUqfw+KbgSbe913dJOHB5pUNo/H1sLm+XBetaUy2Gm2+l
X9d7Fo4rNycKAJqysBfamGRGLnozqh7SAD6fGRZw3ZyDsabExs87oXuC8tk6ZW5DHuu+m5tug5qn
9JApOMQWMSpkK1xMHx7w6NzwVQwtpD4yqIf+vDUTRptLopGVJY9eUXlS69VcegI76PAZYnYP2DZf
Wk+2eliSjAy4BJA/GwB4kz0J+fEdcD6FdwOydhlFUQJFD63BJVUrbdV3SylqigEqqMFuunRRt2mb
s0ETIIxF3OaLspHJTI7vuQcHNsVpCRCb5Dlx7FLkIGmLrMGegoYNuwZ8FF3wUkNJ3Erht8IqTvXd
kyT7AC1N4ueVf6vEFMQppx6J1/uKm9kc6YsFC9wAaUdXsd8ZFmDlVXNPJLM2iuwL/pnzl8S5B2f8
wjVwFkYYrywrn2JktLfjSs5cARKRLDN1vddiIwi4TyDRTWTv9HgCqubN10dApHNJoPZVzG9IcWSN
8Ov1acPRxtfoEG0vQ9IpzfEGPXOXQ051UwLo7C1p/Il7lcdOPqZghc7e1vbm0/oHR3zMVoAGVlNg
HkYp7Dl11AajwFU3JJMDAQCfzfgsaPyg5/EEs2lk1L4z8l6SQ2b4breEb35/nGN6Dt4VoyKTitq7
RX9kd8Kcn4Rfw/Igiz1jbLpveAXFMkyEHExnzcaCqwNvVoazse5gfGzJg168gaUqJr9/odHUZSUJ
7ql37YeUbcdJOUQaj3rCTGm6NzilqL2bBY2a/6V/Z6ViI7YvyWbJjzk0JUtUuHjvdurQybJHI+jn
zT7oCyNkDJB5/RyGO6MVbZcNI4ia+vY1wd4+AVOnKeL5rSNoOIpMcNb4NXmQ0y6LFzkR3EzGGD81
y5+HFWfS4GNQUoTXchGqVPNw2AeaS0qjdX5wE8LeuA8Btaot2OnCHrO7fd2EMAloPIe3rrcYDXOg
EiwbFrCXHcLjL4v6cD1ON88GbX28pyV3LqKSDqK8zckEDbOnDIc78gwg2rLoeAke4P7SP7ajijiA
YIsw6TJNdR564uXq/oo8KTD0KhIvna5OjJ0utWle/o5tm5dpv4sf9AdMGoqwiW4agpAH3C/FPgF8
XOC8/egKfc6BGeyoNKOZv/QHGVsXswEl4sZP7xgM4cvTFRNTB4mUGUt70QDaA1ddoH3DqRoDE4Hw
wtgSGh2i2bcMllYSg6SWzMXYSfSVxFw4yThynfFDZsx5l/ee2fMDGaoc4NlwTMQEEDcitCtKSW6k
voQFkLoOkP/kIMFYNZQlmPkgOCf2+QvMDpDD0tlQdfMQ8L4KLMQ7TbY5Elzvc1W8kuWogzRZeCv6
B+U3Ul4BNtBC0nx1EshBihzzo/+Qnr616zyOnB7FzJO8E6rK3O9lPynePb5TaW7VU+9W7OQ5q7/X
mwSCSieBR7De+kARsXh+yHCL8i/BK86rEyBxtJ9+j2kz78clIIdDrthnK86AgdQMfOM754IHqQ4k
QPPvEEQvjrLwp+1YSPVpnCbI9xzVKz++EL0O/IsQN2dLdz1A0OsS7ButImfnNrkYUnkzJtSeF5sP
ZIwvPh/HxuMsV+alV3I8WjomGRS19gHkpAlcQl1kU803Mpe3uqNyVhcjYHewkZ81+HlOSok9zOyc
DPQznpogEsbjBK68paSBIES6UBo+sJ9qllvw1TELofn72BpyRtLhRoPSZtdG1k5bj1+FKmnaDHCX
SDE46JddYzDupPvSQD7Ks+yhzh2x1FncfGbr8PJcdZ68xBPM5Vo7Iu/cb4OdWBR1LEz0mB3urMmZ
qoG//slCOdjnmZPCecjoE31vcOd5I43uQkkI4oJMn5ePObhbjUCYYbsikoHawZ2XZRBj5l3IcBjJ
U8BKLVtp8t3i9KY/SHIs7IkqQ2A1zWNYuTg52sRrUV+T6Te7B/QA+CRh3nAC6NU2ImbqXJlB1B6d
AyCSfk2uoeXNBtVLqNNvu8I4E/+fd13Azg7vA8slGVpRjqblRyVzfaCZnaqJg+XH13113lDcFq/W
uuBraTV3BqLUH5EW5bM6qDyEojqNMwGo8/yeXFW97DAhIJWU1MQeEB3n1yyPLBANnzCgo6WFz2Qc
WXhwjtRhZyKgvRbRLziDHtZvSoV6iZzRl07hoTW1jiNTxl7tUxU4/j/5GOVCTLIG59AH1ESAvxVj
nlXlwc3P28hN9yyQxIb+G9GcgnUnQ78ACSvIRswVjGEMnTDW41eAXwqAqW/dHYcYG4EpoXivbU2j
SBy67o1FgdFpVK6PURsckKHGzPnXni9Fvb2I2CTutW0U44/PVFauo97Nv+XeaIGa/HiT3hbja0Wd
iMvdDJWLON4X4ugUk4+VtBfHpvLgq4pRQ+Np2Zzk2VbjqKYshN7e69mF+OJ7Nx7WsXCGoBjf3fw+
1CsnSK/BSiGqXU/zlj6fSXc5R485sRgLWncswBr57l41grFlQwEL6n+pUIrxtKPzSags7ZRoy8eD
PkhZbrhaga8MBrXUguYqK0HgVow6VYDD8gYM1TalXKN5wKXMUtUBex4XZN4SAef9KyJ+EbuEMVZH
D3adz8ieiQ3WnaDrqTksG/yBubyStUeM1X9e+ye8gbZiwD/eS2BES2US8rKIUnOep0eNb+He6iCM
7SHOOW+1cu9QI8lTMO3hkYE5UJ2w0UCRyIyiCDU5nNZGH286i7dgm1gT+DZ3OoE/qF41HOlxowIZ
U7Xxk6YotBaoPO9asQhHyzi85yIJP9Xmf605s0agmqR405xIZ0vc3Q5DFt/0BfC4/uDnFfAKWvKn
MkiifP9mwy/GUbk3Z72XJsJM7YCbE5lpbtNQzZFwbjXK4CnR9dNYSj2RLfqr2FO9B8hLhJcLZhZa
XusfEahAh8tnD53KnM2xJ4ExkDt2z9hoObdVvhodKvoxIxCkaHsrPJpkZtSMCF21QXo5GDsi5LU7
IdNXcNdK7g4sLM9mOmLCSt5NVMtYFJtM0Gy5xRqSIvFxEnrzm6B3YOjeKujBzr7nmgaLAXozKUFJ
y8kyyEJBkcNdLkaG0xukL6Hi0oN+jjcj4fajwD5KAs7DIF2lP7t0ve8Zf3jp1x9BXtQwjyCJJ2nl
gHUYGCsoK5J7hYyuSsTlq7Env6udJa+oOYvaAnhZ33ZI93DHZ7T/vc4RCP9vMcLtvR6BV79gwq9B
RmJQmSg+YSgLurku3en8oXBFpoi34CpmczxylGAqEvKCSoY5ZaO+lH2sXgphy1R3QC7iqWKcFTi2
0RiIdbArVKRztBguS4s3gdzWq8f8dQL4XKnukh8V9jcOAtRT7HkQAMf/oBS26sX6oCFsHvz4K4q+
08zBUE0i5jVZS50rt3N73JSWNRzQHfPHykFOrQuRERWogXnvz3WTvJ6haeTdMV1VBICcxSXUcPUu
dAmKf0m7fgCNnbG+dZl/Jp9+cOo8Eh9Ts3fOwnPRCVza57srrlkBtwKR0VJTO2k5N4JJkEnGoQnv
ub5jxFHqAGkmTj5eu2FeXGvbP2h1tHdyBEC+0bXx/fM/XWEYve+iUtWKpstHmCjrzw1Xus8bx7zd
6a5IWz4I93JZtdGWh3LkXP8j3hDiyDIcyrRyERuJq5TokkgNTjZxgQXPlaTI/qFSBrqJ79HaH2sc
wqnd9cvncWXVZaNJ6Lo4+z2nplz4gjHcgWS7hmSYC47a6OgTPYYAVc0Bcn+YKT/KWGPKC8lTm8A2
1Mj8iGQrUvnhCGOftsmR4Y3lgq/Z8kIkF/aiJ5dP37lhts739o301jNs99V5WxkuyCH8FxjFnevk
ZhACYC1yD0FdLRuw2WLCQ1OlIW8XxukcGjyfr8Jrej4Zm+NjPC7LQC2WLlj+Nk0D2qezfKjvOEAI
boWCJsf8r9rY2x9rb2HXx2RwmofYC0xzQkeB91fDn3p/AU47EDANKWsVDxiuKueM9p61kQr+4CTT
gKEV4Ib5Bwdb++LhVyd77W/j+3Gs3yL7o5QrsUtlKszEK+KKumWLyHBm62WJq8CDiULrj0DxQL0b
L5RPeT3gO9xDBCWiw+4bCgBcIGrHQKt2ZTDZEEhGyDrV4Bj9Npp/WFrjuhPJ4q48rN5DlsnK3eD5
dxALGcqnLypY8ODvPjD+Vm6cak8mMoMq/VaJC7gp8BZdWsOim98uCdnCPg0a4NcEHpDpTUG9Hxbf
eWIGeSQs/aALQNFxmdykHbOdT5naKG8eBJqEQk7U1Xiego74tOWS5xo9fbtJ8SPPcG4Yz5SxPryo
Szf8Ss7JDp56aTqhVr57DPvUPgl580eZUKnY3iggTlIyzPh0SlCfCUOFQ8SfVIkYhQRmWsYbUl2w
Ali3eTh7e359eiLB/xuprjvd5ObYxamZjyLx32Q+nzrm/mlBAtvAnU3B7Gnr5Euy9oPpQhAkDK/3
dG5phO+BFD3qa4Mkf49d6/ipkaxiUH/7viCNOcADiAdkDyJIVTslRDfIHQU4ZkIWm4NWaY6gktAP
JI8Q5UksqYEhs3VVl0VBZrROjfIva32bHX8s0bmZOkS3LfCn1LqtGWEHVPbDtE7Qfd7E4AR3Z9VX
o1WRREIea+P51lUSfsEK++40RXfHZ025yfYa4YauFp6H9/IvY7lMOkKa7e47JPUXmtIdL/3m5zPg
l5i9Vq83CKbig9nT+ozM+5lYc473c0r14O5wPtkLHHIOdBzzkD+g337gu5o8kEodN7woFGxfq3v7
Em5aocX84z0eXdLZBxuv/okL+1C50OzMDLnXm+R0ym//ILgdFCNgGuFWmAvgvMyZvLQxGXFVaRU4
Zh2TmONFsqzWIV+YsAhYLubR/VQM8oqO6W7iOCKGev4BJtfPKSR23ITZj9l1E8lTAHiTh8XiDM+0
zczr57pn09KKiFe/lWEewCL3XWwYHmE6dm0Baosp9dY3mVMXo4GZZxnHa2x3gFIsnEQqLrPSIosX
nJmsZXon1douSGf05j5AT9ZPPXmXejN/ev2eg4FB2mK4UQY43vJiiIAwLNcSIf8WDKtRyjT8FwkV
qTLXy/Qsw0/DQR3A71SEzDasBdyo7+BHdA20lYqncskaGeSKpfJgPyDZyUBNXJ57YS21+Vqli55k
lgDbLO2nFaCzupqkfEE4DM+86N7fsI3le8yxUowuBoWp9867e4eMeprmZvcY42CXB3tQqbfkA9ok
B+d98jGX042YWAcYiaTaT2eiZYnje/VbXmiwABKTElahh31fqW2dcQ9JE28k561t2jetmMNbdobf
VBmfNhnyUaStE6OCQBW1wJYQHtlSm8KPgZvZi0muuzSIi324oZ4p02+KDwJmO4BEpqGgWKijMFt5
l8SdK+b7+jud49VTQoz36QjMjrV4NyiEtMiouHiZQjdHU2Bhak1vUETRB5ERNhWJnRXcJy89lwOc
AihdCdAer/CrkAfWgPnDf8KKhd5MqTM3rFDgrS98euJBAgN14lTaCEw1oKkq+JoiECRW5sVQkjQC
kAQHuqEuSzovhuioG+d000ZuOwIP6rM2EUGpEXv/MTJQM7HK7yuT3GWg/SZZmq8qwt2K7VrhzXPq
dElNCN8yrWNy04xRgpM3pCOBMRBdf0+dnlEMEDIjpYdnF+tLgiEZ8RNRrVwFCuS9YxFbd71fIkg4
6OR5C9f1jXzkNZicRCF/p6NUd0e0oLQbEZzSUKAP7yAJKQNsYhsJuCiwyWWXsRrHchIik/8hioGl
4zysvvoE3jng9iwe3zlMNQc8VT3JkKw8l2D2lTwnOjO3CKHKr0tthEMb5FgKoQnfCEdt+dFTOdIY
dcyyWFzTxGjL3zNtvArWSmUCUB49seVmNwU68ygR2XwiVNKBJyl2EViP40je+OwA8PZ+Ux1/gm32
sl9wiEODJxuj+8PuvPRM3mC0DTJKYu4/7dtsCYtGQO4pYjbl2pb2I2WPSpeYKhrAFVWoSUqlsbWN
Xa8iSlF/l1+P2rU6NorIKpyc2s9F6j/TjThP8O0OjG2jo7OlYmgFv3O2S0KIMRDVm+m8UMNA9OO+
XG65l8c0SYRpECR02Xlh0PDkzjexLoYC9RI9SQ0HN0qYhIt3r2rF/TSwXzLGL4bAsj11CdsM7RWI
Oo+1Q6WoiPusA/otrD9FjLomg98hJ4CpelWbtWUl+finHvMSpUntB6UvLC/fJokfbOQshVV5Pepy
LFDdh46xI89ssSeGzQhC8MLnpR01JPltIqTqcyzXllXgRafOOVo+WLJz677jFpDgxJKtjdO7VWhX
lYaloVUsqwDW13JFpX3bEfexQZW6AbrA9lIjpmRU+vl+9IeVvjioWmjSEkYJbRR/KYOprEFmeZDd
j+uVTpdkFD6Fv8Y9T2elLtTt3A7IX52yxpuUkeeT/FGL8l0DTqMpZn3lhKu38U8JloyDs3DMi6nb
5NaDNZNd8JiUbFkc+QAW3Cv7zkgEBOLQME7dGnzrVVhidvUVwH+i8p/5EjbMPt2v0TMF3F1z7Ahx
adByAcHFmMh6MdolFgJEX4dfx7yhar4Ge6Vh+t0MgzM7Z6IG4bJrmSTgRrnmsLy3n0ZtVaPO2C5G
Ff7P9GPZQpeP9u+cPAXWAzJAzqGb6dK5hreqncStgx/gSUL+/ygxquVTp9AkkuPssWuc5T01nSil
6yn89PFjd2NUgmfJjTTjislpA2zR5WzG3c06dZ0GbPGHc6YPUMHc/Opy8UJqXufH6PZ9dHxggLkT
OulDhElM+BLd+AP/t8d+56vNZTd+v6EBovp1nvu7dNsk4gd8DFHZhFSHa5o9yAdCTUP20Gsg1jR4
Bi+3m/krV9EOWK5/6KB9pxyM81A4va57mSLHxHe4XiF8wXuIXTmMT6YTHqtP4hmnMXS6C7mgy30P
u8wNglJZh/8CQkzqmY/hOilyWDZsN7PhAYdto/G0Jo2SoNLhA5q35k9WSVZRpyphsfpOzTRm1s5I
rh3yGRTAIgSOffIgzTFkZl+8MsG23cKKjj9s08DWL3T8uDNvQhZuv8VA0HtmYD66dVYOkMEzW8JC
qHKG4IyzsHkz2KT58lSKAxm/7Uhb+ZCfggaxh+DjeFlPs1RX2puLN3t4eoGXuu9t96m6pynnPuRt
ZtgS5e2OSW3Agh40DOtigvts9q0dp3G7e6GSNyPZ3gxsPQlep1CpRKtu9UWVPiRJDNSh5s6zAAc2
qihs5sk7xpNFvw4vHufVi/xQ1eSlxUMiB+Rpc+b2xv2zSa2h0Gsx14tFNFIbxpHIqDbl+SrP9UEd
hxQ8MW/wMCyGeRP74Y+3LcpFqDiNdVjf9JqhLuWe5iSwTuKaeQQ3oJBnijLPkwXJLrMyYT9EOxTP
PuHD1U++oa8spniEHuXqarFWWAnfqbCc569KzhJQROk9AEsssS6bqgdo5Jqp2XP/JBn22LX7QR2G
WBXUDvYODjSS9mOQ6k/ERVcw+E4MOKpYfcIwHhtHJNmtCArZlLK84BlqREaDRdN+0NEANoVN/en/
JDYfPQ17knoUbMVeHwGEj8EZ/6QxvL0/pNVjNR6lvlR5/Tz6bonxlWEXBsQtSt5c2pRRqPprr+gC
3MSigftNHyS9F6wfNb2wVyleLH9vSEIje25/uNO0/F7QYAGqjkPgZ9/+QSz0aYBsYc945TQqGpIc
4+VdW/JXrcJbKB6mklxZcdithsqPHDwIXnu1UItCOyeifmQeRyUNu0dXD55NBEwOsIRFpOmRwP9S
lbBmr+CcHdzYJ7UvNxJNcQ1g4WproeJu2KVJw0wsGaHLKCKqlVpyLCkIgXodQkHaQHBKaWJ2npbN
c+gZ73TKFT0PfhWsFqwixqnMdNNpH8oC7m6qjNi3zlIlAEdfolQrUJPF55LjuD7Ln1/lLfVd4H75
+sD3ASYpkUXxfvBlCZeBGLbWPh/Cupo0qmLKctZ1j8BocrsfBsL5GeEdmb3cy3bNhqx/J0/Xqi9z
oL35NoQsJ+s4gVkvg6b04XSCQ1T6aV0IcHO+9or1c1kCnnxqZFW3MavHW4D5EXuGNCesqLY4PQqI
CAxX221wzHB4Tmqr/LQNTQOSryCUCMvlkXwqzzb8A7qGVp+Jl3vCRAUl8mil1THJN17GtCd2Z/52
krAFTyI+f7B7Nnyd7ooLwpwcozVkHZ9/AJBG2iHX5VoQ1xWDomcWC+71alUZjHk3TAiEfEPgCBOW
09XjpECd0VTicHAu45H/8qrIQmDDEek5KdWoyuXwVCy2VPmRJyJ/XDdguTQK/UPjet/1WgrOn+Gw
KiYjQBwRqLRzyrxirLIRWa4Kf6uyrCB2LQy+br70uowgChQbzFL5pGOgV1zJk9uWrXD09Dki1KAx
kApEvvmqdn5p6NUc5sWeyNpU7hemcgmdfcxokZP06FYSph/kR+gSWSAW3eNl4dvgj2QbVIMSGlig
zxTgkSV1cxfEMvqhWPK7RRy7xctArUUaSJfy5Vo1dLJ6oCEe8Au7FYAT9Xbo0JFy9iYHdbOIElb0
PDKDJaC6p4x5kMqyTPMk5ltVNEekhmX3Cx2F2oK4JcFI5YFtpd34GCnKoWZR4buzjnRgbug0K3b1
VmLTCHraUhwtS+/M8z0gMaugok5gh5EVmYVjQjURyA8r4XDELDM7IMBe+5lvs06vNnqgy0vRK9hp
WNPJv+C2ULNJXFFFh3UfKmWfxu3qtHKPglrs+JuSZulx5drPFzVaoaqRrsz4QMGjv3vyOqLzHxWJ
YkNlVZv7L+34RVk7WytqBBZRWtzMEco8LVKU1w3S3BiojChZdZZS+Oupn58V/BEVHXda34B2L3J8
muhLyK6m+KoAftQshJP95XoXTnBvD2k+e3ob0WbGV7vpHLX6/pjKPDoLz3oCVwIkG4neJlVtHJxl
ViWPnbN3MH7qDW8WnlVISea5mLYHv23K2mlZZcUq/FNNSmy03U87G+9neWgmPhO01Di4zIlqjNSE
45yRByowWWezQCpL126XhVdaue0DLgl5UhvjLsShqbvb9RxMrY0RrW5+Bv+IWU2As4UhNi5MQVrX
IjR9CPZ04j8xB64lKiiwgkEwRQzzjT5QqKXKchur2bMa+WQClUkPkQqCXF5LTS2m5v5CqPw2EHpZ
TMpH855k4/veC86xvi9Fl+LCx0LZmqQKFUoBggzE4lll5Wkx8lqZrlEiNbkUFSbdb9j4j0tNRdlV
ty4iuawMt/lvEUCn7oyvkJMvV749SE0zkr5mGA+ArDQp4EDtCKcAwkWF4F/1x87c8cCrNI3MViYl
G0gPaQQQkJsOx7npLrJhLs5P41EMJb/84rvTye1pi+gGud8+3/Eiv2BMYTAdeF3ASudQCc5jztV/
4AjEzitzzI5ggutrrar3FeHgTpJyNczG73ZqJcHZHLa0goCpKzaFQ7WzKLgYa5a7RPrgKe4yZS33
uawEOo4zK4gqJaJfxb3CuEmx/eIbdd3onJJXyuwIx5PJeNx5ftVEt5Bf2SqNCae1VkO/JmyX7svZ
PzfXpVmqEtipAJk9GQRHgEDCNNy50NLdSRXUujZDaTvO4gnGPtoWR41YnzEx9ERrG4E5jtauEPSZ
IESihgDZI3+qK3Fqe9StO0YG6J+3HkVUotVn2+CSA1GzJTmDBFAsyewSVEde1fKc9dhhGUrVEqul
Qq16LrfnyGklS5zE5AtRYq49qZzH9evh4P9TEYjPlSuk73ezYkZb8PQx/mZbDANYsVHKeaXz+aYn
7NaWD6gTM5lcksDebIeLtmYPfchiYqYcMr6n6e7icCikRtXY7BxO/WKyzdo89+W0BcoDZ0JnogmN
sRpJ3raC/HchpiT+/tyxmm6MDuTljki0vqQrfta/OsW72FhBsQvaZFdlFzB03RX8od1N5k5wnMUq
2aEE27UXLIKtRodQ6a6sjUN9UY2lUyAJtp0PBEc7k0arYok6F2pcZClmoH7OzU+UmJ9OeMf6j6aV
42vHZn3BLsdSSWNzYQgWY9rf6I4o3BOFEW6ZQdZjCe0XJ+BXLO4Uxp3+FFqMgFrOA2DX0jNhFgEC
FhxeIy+cGS0x9wIOATinI//TbJ2R6eNHCKDa+I5nTycN4pFRMZHaJxmlkU8ePYq53Y2R2+wcpeHT
Lc0AB1WAMmCXPu/Ep4hinsT6ABxcrKb0eUQQ3vncMX2tpv0jGzrDCsJWwBWWTptTA6WxT9CAxoTj
EB/PmJG9qc4UppsOEvuZGbqUKarHfjtiqV6Bd0KTyXJ1GrX0em5VdZKRTGPQoC89JisuE4q4//xr
Gdl9nBEUjlwjHFRQtfyDXZXZ5tkCPoN94dZ5Ghi7royNPga7FAEMJVGUcEZuVbnqa9xlS7AYn8/v
rr5wK4h68reUf0dFjJzkYSrw0v7o+NKXhjl4onHzFo4t71hxa0wWmPOhU00jssOFR5s95aO+NOQU
zEYiqPmBcS+FcmZutyeBkZGm86XqzwaalpO0oLn7rf0LH8/E3wJZIa9f3aLRJ4Yvk2V2xSwnaX/H
3Adf9z8WArVAnVNdaNcmv21jvtXjLEcEhOb42BnXI1DyZeLfbRpw0UVV2zZoE9kf1t+6t/rAGnv2
wevdLQOcNKnrT/lhQdUr5bg0j6DnUsFlHst7aMnEjDdKzKvOo/pt+FPcs6sEJQZ5lGS4Qgbz4B8I
abbjDFD1w/5mCf3K9mFsQeGKh3Edo6DUl2UQrF3FRQNi4F6xNfkFSRez3xvX2d8c65t3JL+uq14p
LNR4/SF8INkCvSU1ZwXJeFfjZY50V68CO9Ks6h3I81yX5nlGFPt+tqCZxp+oFcg46w7p+CkL71u2
ldxl040hAOiXWuopGFZJ8RpFfSMxiWTNOi6k+dlpgOUebmcaB5ng5ksPbtmB4ibCJXjOLuwisHCl
LvERyVHeTAs5G5dqPmoa1dKTSVJsOtVmX2Hl6aubLenhCbTI7zQ0dhKkrIRlmFPmGMJ5EZ9lJCx/
CqWUiVMwx/fSgzyzxAyB4LGrA0PpZVhjPjpTuHMvWQt5VUvZSiiYryQs/cs5OicQ3QWvCQtm2cXd
o7d/rGHh8+zpH5gFjnqeftvDXD7zVoPLJxEuop3Jhjz7Z0HfqGhmAyHcjViWpOzoihc2KCT3WgQE
MNSUbWqd/1YXGz2QhRlsQqRAoqeR25Yu5VVf61o8UlLnpDEJpnKRzQHOPmatDWkc9lIpS4I3KJCq
sgaSgoAWvOeHdR025BWj9Hs7n7qDhqiivaiObZSiCYaCWVWx9QNd6YBnNctxsPTceBOdDUkevuPc
fDNRLPMUk+JI06nB3WTdMnzfajhYcAygVBruK32qCJSj194R/XaxJ6FMQeKs7ZJdJxvuaFbHhzI6
XMhBVm07nQ6v8/2IhPMNUOnS7BLSrgfJDcvref1vpNh8Km1d3z47Ic9pFnhidfCl3D4qIbEq/JjS
w52MdbWTQn7zOwCMxpZyQ74V06h5BVi7g5p9UWl5m2l7RoMGfqjznRGst2l9psp86ldbl+pQlKFZ
5i4ZG4/Yee5Skxmm7GZx5XsMpio5hGLE48e/5htTskHviLZe6kaWOHISOET/nYFFozLT/Cyl8RU4
gaVnn8s8hynRJcAMcEkfoJu1daoFMzR49K1LyTDH2nK1VkAhmeQR35odq9ngS8a5zdf7RNBSs2jj
AIvHItpWV1FSQbrUuyv0yLqZnybsVN3BkQc5BkbVZuN7/LbyKQudE5W8bXsOHow7EeS/dElPA9Si
wFfA19hNzl5fkeKo5emPqKjzCOA4oz4NqbNjp1682XYrJZ8WogfqSbjk5CdDbwGBpF5b+iBr62EC
Os5EVieQkRUlQQPnP703yEwSdYziNX7MBjEboatF2tnI0Mca9ygxxxd4k59fPtzmDxnE3sHs6H+Z
1TnvRa+SmTQVe70WJG7PMLNidsR8VWR9CfYl1OC/I2aj25hm+awW3Qki95R90iCKZHJXD95JEP0t
s6enuYItQUCMFI+z66kGSvcx9BD1BR9fO4tBtYDudyYhMqHbxvNtBPip++WEglwiw0RMdbig8frG
0WciTi5u+n6LEN919bGDLTBOUDil8jEiJ3zuO0yT5QHyjcaZRCKut6DOg0idcvBy5XMfbIhNIaq/
B77HCvxV99bqIwS6oxv7f6UAk4AZWP+ijIL3qkEdLTz5FYPCC2joGG0djqkjjjORXDdZvkV62YAF
5TQwM3GoIMs/bK3G9zlGa4jO3AGslozJJsYknngtDIiKDMnSoQz8xbZsC63CErvVf+SuFE/uKPL9
p9dhtRemK2H+Pt1ZxbEoGoUvJW91MINCFWDqemE/vNb1eyFZaGl8H27XrbQ+bK6JFat2iVxxFQ4V
OCkMezOx/1FQtQeOPWzivIO2qi/LKGVrmdDeGbjN9Ww1kmMzi/cMOUWSxGTk1ZgziLi8Idmano0F
D9V6S31G4oZVfbFtfeQUaNn1aKhODm8m9c5/sBPzssSTreMJqTXvqC3E/jXaHljLRfrwhtMti/kN
KxLbCndZX6ss8eMw+a/uHY9xzAhikhUQ+0gkOYZWzsARHbZsci11j5EA0+QscB+Gu+pjCO1VG4ds
chLIR9rII4/tX6pMXkbRtM+Ii5tJnMSLCZmA8EhbtHzeHZRl776i/x1bvQ991ezDeeqqVqtQPTT9
TgyS3nWcOl9fOUItNf9uftAZ2djCLqprDv1hadSJWq+Evy+ScRrs9yGrHOPld7BWaleq88EjchrQ
s0KwO7ZOfBzLfd/Q+Vf65a97+nK/xZDqtRuhg8/3pFPEycxIOCpmBlAFjFi80oUGuwh7kbgESaA1
EX+8rujWM3PniSv9540e8xftKC8ze6XIFbxYFDgWuxDVrvJQrCWr1xT+B37/P4MQcSIBA58aeVDt
Gkfcb/JxTFW3hA7tNWtgfggN0j2Jw0f+hndpwq+ZSczowrYgFbQ/NaHTcxW3eY6mUgljy9HXbfxQ
DwqEHtRYfGnCnjDFoFpvX7BOirnu0NdpyNNhKK1mzVi+/t7zWCwMd1NTA8WJgIJzXJcjSe/b3bP2
GIvD6iYAwTgac8vSLP86uOUk+cdzju6cQiBK3N1c9T+uXhifYo+hGaAkyT2CzyN7bUmUIa0qU872
0DVRnqgmpVo+BF6lb7LWWNmFOV5sVqRHbb/zgDXliocWNThnW86Q0u6VBh3o2tTGkbgy+peZoSDA
QsS91p9nac0QBiyd62VPJ7e8IUA1fUllpIE8TvHr/NaWRTGWnk048neAppQ/rJWflcdgVA8KVg0A
tMIN3cv/GKP5yh50jikUfM8EJRttGezP3P51wnSxXnZHkb5D1NTtQQYJyjAZRFPc9b6zCdT/vSCN
VrIf1t8/LSGRGoVGcYAgpBEzgezWwXpMr/jQvoP5EqlXQl7jlSpIOac3HG9kyitv0Vbp9QyaaE7l
BG1SLowGaq8QzUveYeMmvnnYQRtNLPBH9bUFm5VGdye8I85cJN52FL61m34mCuEToSRjUapN6BTJ
fZ5Cim4WSEA2kSMXk8tpE3xHbvCf1HcK711h4itAEUwJ42z2YCA5DcVs+MOC3agbC5PRISnbL+k9
9+kAVC0RYaBaBqs0ZSKE1CJ8dyaFGnPEcbATktGqU/PlXTFj2oaZQrXC/1XFP77vc/V9I2kpSZbH
BUaFFroOTRxXGeHB6kYipMZpvTjlVJQsHU3iHsjn9y0mCtjmUpyxamkz/8eDDEmDFq0Cd0y3vaa+
O93EXx7aFML346uoOP6PT6n3QXk713oPQgkY3uu3NU7Pa72ncPCSGD13UTevbDB4XvwjVHt9UAyI
xgGB3M3NzkE2WGTFghQW9431tYjcZELAybqmA5277SjmsqKVt6++kt9n5uzbXmgS+ps1668CDFmG
GXdaWFnW30j2pjJjkFrhbPi71xe/+kSrVXFpe+xEALFWvyRBUnEMIklTXN9IqQ7KzjbRHMTnZH9m
M/Ove0L1kizwRibcum+xtbRbGYHlJetCGriL1GIDqCr/XU6GGpRlzZALpqdzISkj95eQM2Ct0ljA
FBgXt8BqSBUf6QDCQwpM/FR8tZ4/GwWCQ8LXPDuiKGi+durUqRp/7DeM4F9D4QMS9GoimRj6SM9A
jQ7laUtiS/b8HNn/0F02MX2ib8sYLftxOzVpmlv9/BKRuxdyYKPnvNu/x1c6wC+zUJmRcq/kxi2e
PW/oE5vXrJX0BmcjBtnkGobSLQ9DN7ioU2HNaj4Cb2Qk0/PIdZo++skROEjojmL1Awzb9WxSH9BR
bBmsHNQh+YiryFtbanBhn9r0Fq9JfDbsD+mYfZb008VrnnpdoiG/ITpfDe2lD1Z7JK/WV3ahwD3y
hh93ZH2vqRJKnXM/ZZEN/BqJjRfO/ppenpyeMml9Z3MXETW689FAYGO5BwH4GAljjF0G62TM5fC0
253ItHNxvzGoj31F7ix71pcGrFHvmPvaPhZzAV6rktrd17ZgWMS357p3nU6wtYlAj7wb3h8xufDV
JktqiUWM8bsv5wciYh3RZjqXBgfWyWQfbwkCg5+RTMBs95EOTvCMVGyHiTh4QhM8JD7U2TRTcFqB
NZN+M+ekk6CuCPoWzwyCunv8BeXpW9cdUkWvJ6srG8Qgiw9fRV7m712H4uAy8owz9+LhJ5Kz5TCs
5+xm7X0byXx5r6W09mqhnHyRNMEDuzY52nBXga77oRy1XUAALYt+5GZR25A7YHhXtqrWu+Uvddva
PKwcekTuAfqK4fVatXEQrjTD3NVimK4lu/TsW+QhDIzYYmLY3e+TSbsTtjujAq+BNoizv+Uc5JdT
aIAGv0XQ1oqjPzALEtskIVlD4gmi2LiEfbAZ26wRx6oDj76z0wzGnDXFj8kWjgaS8bbFcCwbd4RB
7C2jCFBW8am1CIzj/yeJFa51HxUD/3HSLmEissLtVwpssETKLxKCPl1OOaGGWqN5If5Gq+A1LikY
zkezrWPfTugfwQfEhF79JSSefoL3N0dx7rZYuzDhjHYoEUaHMEkSYYNqpBH+DSlkSDunr7v+YefH
UBGoGe0ocMv/UzUu70QvSe3V01kMSFwfEBf48fjq9dqI1rFo8O2tt9f1WRrf0uu2lvEv2imOlbHp
ujHQ1U6wTeSFQcWrojgRKgoURS/mPnDBoDXxamoFZRtfiDZ28p1WGDTIkgNydLJVk9T1fwbCtwL+
u26RdBnzy3QwgEYiDRx2hnf5YG+kRIeVcpbH2GI0fy4FzPLlQBTuN4vIs7xecnlwhkpHCAhZOyfx
TTGnpXCscs+n9dpwWT0Xu8O27Q9OFEmjQWXJmPZa2mwYNfAtuorT043spMrJjUqoFJTO/ARyFcCj
eqgq8tG2k7BdL/tH2MzT2bYVnIie+EIZwbs9K6eAFXYlLlpyIKRfBu/X4DLlolKaB/jnkQmWoV5A
XxbyYKI40yQhKtbwvT3W7bvKlzAAFZH6BgAHpdL3xtmkibi6Owv/k/b3gVVUubNldIJu+fTJ9mXC
JeYky/H2vom14JSG+eiMwbk5oMXU4ZnIjRV6Ws799X7W6oWz0HcmdsvrUZrW6D/RmDHb6npgfET4
tE4UsNvYCZSEGkVhQ5xDw2WsOFqpmElbGxMddRYR/orE1JHZv6JvBvS09Yy3t88aFxIL16zHMIOh
oKua7KnFJy35j88xDmhY1cwq9n/Bt9tQMkYcf3dH/25viKZnD59k860X77UQxX53UET/q8ZFVUCE
yrpW2bwLvlsNax7WxVO7HjEzj4lTATy0Vrdczx7FFLdq+1mPeGk83tphSSljFBMrYVOQy7KIYtjz
N+zsSfFXqrx7qeCYDeruLtGJCj7IinP6Ns9DMYNyDAJyF1ADb0xlXTSRis58i6ZzK7uzBobNFuau
xkx4/LRwsX6qVHKKmiElTQfvK1Z7fKQXqU5G31z0sZMivq1HlZP2SON4CN93nBP7VoiVAL7WhP2q
fD4ZpYQOGGu1IWCBgmocQDmSM4vnVWJ4qo6FyzLDOIFmje5wylJxdV5CkMpbbBfIDYWjCfeWCnMG
4PJy9R1mHaTdAkLXzMw6VehpF52mBXtwb/YoBBIz09TerYg2ebUZ8tVN8Bpjhg30Bbp+JPgYzOGt
mF4vb0oMclJKWPCvNOGpFRGHmCIubyN3v5aDwoo8q4+PtspQmpx+OEIuOhFWqkp8VZNPJ2N96CZd
gBDy42dF9QAz5DUmr+9VLiI26E4vPCRUViAMpeWq0lM4LmuSFNf6GuL+ZJG9G7W2KAOSe7h12y2J
0nXeo7X0yrWb0agGGvbrOteE0r9p5zlmyW5uyWoY1+qGvtynOTOmxfZPLMSl7peJWhUQ45yGIWB+
gWpaVB8sym08BOl4Oq3LjKKAawLMrsjr38O+0661k744uHiYX/pqMWhUtpsQwyjYqPKJOfO36wbp
llqmvre2QIKvxQEuMswTev4oGdg2GvEgI+atSRBXdeGzBnOP27HiwyvX43+lQKnyMrqZECq21Sdt
nI20VdRIeJOIwe4xtvQPZE9rwQFG2FqTMxcL+e5fhg3c+w7NdQHyFfUdb7yPSeagn9UwthHhQBsC
XwsEwmHr8gqrbE1MhwFoeDuRl5ACmK0tjMFAm2ZfKqbt0O4k5EkzXVraSBkLq4L4wi8xmC++LTKO
0be1UMu06+7Nt5iAZMTo1JiLRwLnovvQ6rm3x4FE07UvcaunTnfSDCp1Ue7MlqZ1E037RVUyry8i
Nb8FZt+LVXhTIPhg94eRYXl204IyCHk8aXcMPIZi30Auj2gh6kccPSfm/tdp7JBqnmeqIAxm2pys
9ZFRc3Z2UiGiAAnMDmv+CY2qPeawywjiIvSUHKrv4Kc8aeS59h3EHrGsa4WyCNZThLSU6+gBmalU
TvEoq/CAy/vk4vHlmUd//HjMwOghEniT1uA3OWTZS+WX+o6nVJ5opzlACdX/eDJcEQDpL5PAteLn
cYGEMVMbkpc8ycxEuU1//8ZUh4aLm8ZnM9x008AaPL7pHP13PL1em4OwIGJa21jO6ju8cI6L/7mB
ctmyDfFCl8ggcgZ7bqG34+oF8C5DOfhwVZvkOagkL7SVyDxz7+buLrsTCgtnjxaeu6V+3u/UlLPP
pG9VrcNOyvFSSNOJZMHrtVNtpu3p0Pm07k9gqalI0hdkAYdLvX9rquh17Eck1ria3IyyPMjiZjrQ
bjpTT44MMUbEAJiRoMRh0VObVJt4o9Ej9OtABVfY74uFmL8mCd5Joe+0k3mo/lRzMb3JpckKB1ha
hl+SrP4x61yLc9wk9Oc96PTuk0ZgmYljdi+aYIpY6BFuTJYS1FtbuI6tzW18XG6VdRh34+1PwlTN
qVmRdUfbmv2ClU4MH2sq0P5nvwb0bnCG5BHk3yFPVZUHdnhbjyr2DmqDZuV6qd2V64qd0nzvVYZi
zYseTQLxz0Kn/7rK+FfI4aoDyXrr6MWnBsULcaEKkitXPDkVQa6NgYtKt9n4k1ikWGwoqkeqdKtE
MSEdSOVlgekx0X7globIdhlIBj4uvxL8sbVtGpgRsakjI/TOal2t5IoLJ5wNb4Q1zOHbS8oynQom
zC2gMwwAXrH+gCwroa+5QcaMSdA0aCtxGDmA9boeGcUmnctKyKn4lk5kYxGZCA5jp3K8mj8oKtc6
37B0Y1+B1knbBzwkfkZd78nMXZj5frSWg206lBg9mEPuMTVybhL1NFDrF+sPOCjQHi0oXbKJYee4
IQSVau22ampPYxlWe4mxJoHGRrCsDEviAfVHhdxXdzyGvwfINxTGFiiNlsKVVJg77tqFSLSfJNEO
FMQyjWuxLLk0QfyqzI9fRqt+HWaVNIAwZthF49Y4zrVW7qldkKAb020HCfR4WSbu5IUaZhJ9N5PV
+ZXDtxknjLJcGFxk+bCr3n2hGdKCfqIl2Voquz4ijCMYIdGDTYKAYxa3W6vChtPJ1yixozIfcEzL
8XHwvkw43+7NLTGjVQoeyTUoFHsQwh1in5MkNmOqLCCtrz9qEhn4zhKkY+FHuByaitV54lWWGZJm
0QXzp420bNrOMRkrGpqjGNfGC3NgwLL8ZwSekm9QLvuBfAm9GTnh0wlvv3sTu9bLe6tSpnvmwred
VD7qtCrcmg04hfQjDWEbKrCr/0w//QThrp7/4o1qgmxeh5H250j4VHkYUaPVgFlZqkbWWsjbvlD1
eC/oHnGGhDB4ramVy1QEYlz3NB1KGtkMWX/mcrtfZbppC+9nwEQzScSLieTgaYRAQ2nZrtOFt46Q
9pOOwnA/Bs3ONOFUrAlKtql6vNtDmwXWah5diaknU3hZNly1HkGpVdI/NbiA4CxhTMs0PngrzKpW
ZKfZlEnR+d4x4hbz4lA990nzOSN97TOsYFTDGIJKWTU87un8VQEuTpOO9xkOJGNs15ZCnc0aFUc8
ZWY6mPgs4XP+kT3oqPvORjjjvyhbxR3FGpy85CrW06eYDywLbJhOW1NDVxRIYtrYJRENReBxpSp1
HiAOt9lAEKBffnM6ew8iQtpwksjDRXAs+pgtIsXyJugzntpgxUo4xXNixScwiwWPIjhdlsZXpUse
eRpRiUy9Zy3oGT8lSaImcMXhW0epd6mYnLlLJiPaxMKeCg2mxxSe+ErEEJbyn/ySQ3dortWJOzWd
xW4a2xX/AA4K1ecNkZVVdKThYEB8wTGxiX1bzghsvND+Oat5SewLJ6heFouq9MRm86iCTUDUHcwt
mmS0p3tq4m94JmdxG2P2fxmJ42WTHlcLGd8So49ePYpqfP+lpB1+A2Wg/1junW+VZr+knrBfkxxq
U9NNSdE0puaXws9mC4K0RjR+YniEIjyLO5V2SVst7zHtwjBfmbwK8DUJe16ywxYMqQH+npklIfuJ
oykxvFMYTFtuvSRt2jV/akoeOlw+i5U0qytmdI/M8r5ED6V/TYLmb67tbPrMGzx2yLbzLo0bmnMB
VJVs/XvGWzMt+wHoi/3SoKFz50/+Nt/ISYMAR9R7qAotzPzBFgKcGmn3rhKyxGVhwZeY9AWMuhSw
yF23UDC8MU1CfqiPkF1eMjl6sCzXHU2vkH2ZC4iEPY4LoLgG5IDfQz63bLrJY+/stdcsItMk2f6Q
1jEJJ1vDCOGc7U2CWCnuylcwGu4JKg1676/30iXPvPC30CR70irXGvLsZek48SbeBO3TdKqOXB7O
KTiM2sM6SlKA9Y5iM/NcWGhkHPUCLhxPe+er1lW3GXQe8MakV0X5TYvijaSja6mTaOLpVw+mgyS5
fn59xlFm88Sb0QSAiqb8++xnCRWwlwBPAba7tALDrptTs8S4hyX00FwuiBvSD7NaLMuWL7ZvD8t3
JUrEUloMXSc0HJNrCBT4KbJ58ci0FbEcr/1LjM43WbPaHNKV6JAnR5RS5lbYjnOzdV66fUbQ37V8
IWV5T6wcWDTU2oP8LcaKLXw3i9JzFB1e4Phsq19xby5zy20PHW5x3c2jyV+35vys27qCzmKwsWA4
1JiO+6U8IGEQIXv8j+uO3MB8xe5JF+W81sCdcSEJigqhK/h6sJGy+NZ4jv+3IWmdkuZbUQtd0pLM
8EywZCWkQXDCBwToRXNP6kmF2fB9SVGRduBmfV6PQE0hjAoDqOKXa+5/mB0HQuRysult3pkqQ77x
T27h0s1d9cM1ssqLLDYK7tg3XM107d4KQOWsJN2P5rfSe88UdMHeZByw/aT++BQC7s0EUjdfu8MR
Ww6KAYKGlW6dI/szzLjbrEt6pCHjBmtiSt8nkIrFDTGAriDCGvPIAhzeBKJZwrPzmJ6vi6i925/Z
MZ7TBfAfgpk/CDj3Q3xr4ZAvOf2wHbwYz13pRYH/M28NDxQGoYMHJQerX6icZ5etbxEKMN3hKPGc
5FdOJlhVsFJ8YIlblKSZwTWiH/T5sU8nzN8uZcGEw+KEiHb1Gv7CdUw2Gi/Ly4C8ny3PtGGpQqDk
bvrVYAg6w7fgmj7XmSriQbipC77cSJJXo5b/TaNE6OymkppRqbc0JCJ33WwlRm8qqWwoz4dm+Hwk
r0AmQn443JINIYcnDpZSXpug2M6f0N2jB8GbtUQjNgOWAXtEjhwJyPrE3DraT6wY0IF53wTezUgA
nxSRsn5gUaYKYyVVi5SM2U/cUv237382QvUVA+RQPe1Uy32FHcNa0F6najpHon6UOaWr18JLWlF0
UplGylPNGAdrMOgeG/hKdGQDyGU2GM6J6rnBcgfze7eo68tUdmkaYQxERBZ3f51qS4IPF0l48Gig
v+1hbZgiLxr0LII7yzfYDSZ6M9UvhuFI0PsZLU2buEz58P5fz0pRQOl62rRIxFYTY+4nccB1tqte
/txrQL6UY9lOxkB5En+LgKc+9eENMgwy4kmSI7bSc2RrE8FfWYyE8UdU/XhNvI5S8leWGSaqSdCO
g9uIYuwUFWyKL9wizebZFKmlXoqsqumdOska564k3ia+NGQyYps8TE4okPpQreGpe6F6OTxM+FYj
Ka25szg2hJd+TxLVSMaNmw2x/e7z0sw7FAWhHlT0w5QxjMfM8jCdwNUR3XRNQ/fU8k8V+Gp43Oom
pqECR7kvVVK4eTUXhNtedxLL3QJNufohmqdsM+pdIUOju6lpNzDc6Kc/xn52HTjijN2C8t4cEvop
xhTfCfntii+/Ld8NsAiZrOHv3LzK9JiFW0za4+2SD9FL+9+Dea//0LW8F4Nnmc4YwPJcghqed47H
XqiK+ayTEyxihYZpHWnUwXSUbeK+vT61nrhVKAhm/5vJxC9Sg7TuDqpph9bFFSaHG9EgNaw1G8pi
C4YYfgVCIWgNwvoxmwakdN4n7NiCQ3vdfVw70fWX33yMONFwLzPUdHiUPeEAA+qPTooNEVKa76vS
jC2qd03bcUNixX8ADUfyVNf1E8FaEZhz6rpBCGhayVCiDCireTIPPOKCrKt8EODMEHE96OmroIbI
CmxV0J5u2ySiA6efed3K7wb7uJCgewqx7ZdlXfNHg51hg3jzxFTQeeUw5AWo88ccVtvovzn8Cjpb
8FAWDFYprEcAhxa3jrn8kyoqv9lShuEXMVhH1o5T2HHkbHOoaVgGXSHK4vrGLWP6WIz0pGGPfAof
eQuJ0q1dvMU1sQrlA3po3NTGO0cAnRTeEmu6iGS2yfZRLLZ3VXqMNrjJa6vA9la8N3Jw9S/pUBrt
OoID1p7WF1FMdphjHxq9c6C0XO+rDZ8cVRiihFnBhi4viFGqpwV4qDomh2qiI9LNIJ0bfszYvDHf
//PiEZuEeRigNcz54K9oOvizKBe3WJqiwGLYzkOElU3A7pyvO4PKnZzyiYs1D8I6fo7wnyls+yLi
MZ3i71L7yTXXH2W2tvEKq7MHyxPHSoakraVVX7nBRLENjXIDuk9fNu1uoNEGMlNlW1doHqX+m8Qa
KOuvyU5qvpXhie9aitCC/zuD6FW30jP8lajE61fWehKrndBdKuKTeaYGDQCtWSzPcyRCbHHTZxS1
7FmQRxVvOzFTRPlrtamzvsZEHHZB5frtBwcf8AezkMfUNesINaun7JYg9Z683R+FATpVELJmSu9s
ICjVAhitXYwiyQ92zOhvY+TBLJS9oBfTtzmY+Nu1pn+O5DCLL/hQDwHaUft1DAsgRd8UwG5N8yxl
NWak4B0hBZ4djg58hJqxIwNRkub2IMfzBx/nJMpo4qoZd3+WQueRry+gUYglv016OAX4aQzI2dqZ
Am30j6dvF6QJznMXlHrKTj+bG3QEb/k0Mdwdue7IavaUmkYU5ttp8MXWqLYmO2KZQTEX0eUPW0cA
frzpZg2yPOBFhTOWXGHusgkwG+iXn643ylJ0K+ioiUExhukxrNaxyH5qs2cJgO7V7b5u6ITy3CII
ExK8eecJC6d8/L7UEBPrFggLPEBw2DchZB0/BB2DscSfhLJ/H9q0w6T8vRMXldK1g+JEC6M1RPaj
kkxeNbU5+XPDsbx2Y3+yhzkB9Ye54pqshRXTNeZBFDzhJq6lMLG1tI2hLX1dVpRNfznPCevyr5fE
8MD0jleQUcPO+YasqcZOaT5zZzk5ZimrNtyxFhbwmX256zXowa3/mlhlyLHGB9QvoPlKHhWTM9Bj
APJvc0ncE3ck1QBHF98xfvVyJNFRNVowCT8NiMvCOfjOHWaHaL2B+sRTduWwOKts23Ggvibbx8oP
2AzGiIX7pGl+8ERopOO+q3xY8xaKTX3OAU8Zu2ASESvv1CQPvE0DMABfr1nstgshrXlBUOGHjzxf
CnhLy59WR8Pvu2leHBLLYGCONRE/zuLHyKkLKHGBk1wPKMIF5TwYaLwK1pTgjc+pNLysHAnRt3x1
ZqgifvmKTUOh4XciqApdW4VLXHKI3zE5ct5LJKixldntm5v8ozeO8Sp6euiASA1GqSAO1kGhD7BR
tNApNgqkE3duFwB5rCflLzWAC1QbYnRuUHSkwxj5+DA8IikE+vh8z+VzSQBl7rYKH/TgCfIUpUW1
ZqdkVIv8HDY6F9piNpE4SqWPh81Z/RyYqtN/qy9TQMfNyRQvsthhvWpRm+aOQu2HAZ24wFtY/6Yh
Qw5zlASjkN035RHxHFpxP0200w/GOHpIFRRAIIMBQUje0vk8RwwvDOHTU9TgU9PDf2HxUbHCHsgy
3la8PnLANNq4bMujodde48LMSBNdmyF/+U9TqaXayVd3uakREil93RDH3OoNxa5WNsF6muhz/oDq
OJeQaqoM9aEE+Cv2/kNlj7HLEO0vUhgMLrf9GAJecwTT09yC6r4nMlkFWI0FgKewCV26P9ytvn3G
/37OTJot4orqT+3Y8RCyv0g1kMs3Jhisf9YoDXaSqEq4+GNPRBWWU2YW3c9vdK2lVYQWiPm5twsq
O/dhdBnm5UhkGRHS2ie7Z3D2WCi/b2aZ6oA106wlVLg44Psb/dfuy8HMA+it3eD/Xmyr6RpLkAb9
D0/vpiUnn4DY+jD5TDHfYzzFCRJxCIRlsEZBNFLv32tSKgdIfJ9QNSXXRrOh7/pdZzOAS4fxy/xA
ioOYBIoXJYnS/ygvRIdEJ74f3O705u93jNENzJq7dvJfzu93pQgbFvAksxAanuo/bEoPP5MI2Cmy
txkWK2MnY6zsTg1jARROSrVgCM9oES1zJ7F6FKZGIJ/o08IFe9z4aDmcYSxjAeeh4vAlAz6YTWdW
WTWh+K/kC0XkcfgfLBjXNWqTwbQiggvjGgGY61pHHDa1+PlucM+K9hR1mHlfzSXgqJ70hqpQKmjX
xz194YoNRE+Zso9FN0jDDHxQpfGkvcitpX0WLEOqaTPpoMrcShF8OCrMN71sqk6raOC3ipHvThsR
r8SXsdagfcr0OkNhWHk1eoNXJ2LNQtpSlITCtYwxwCUJmzm5OtQUnT+1g1QSEaJyYT5TAEA24JC8
16sfqAaEGR0xBOul7p9eAMUJUh23ClTb4ulXR9oCYg7pwelLcmMnac+/9iXmsuHdZOp1OkI3k1BG
ZqhhbEnlOnZYKyZBPw2R2m7yr3oALWniD+NxKfT3vMzcQ8ffb+XRLBwuzSUuBSwyD2uMXugRs2QF
Au3Qs50BoULJfXeOWGCmiGo2KoJVwLDvJ423YSr7sYHkTVa6RTWZDfIU4sdcT0xnbfVmQJk+oZ/w
Ai+JoZiVsLnujgbZ5fs+nra7/zOxy1lpZL2FL18NERvVSy0qV3IS/c6TUMwnwoO3kOUPCzx0qSjH
kd4/21uUEtkH0Kc6PsY2EGqiq2iHT4LjriGuW1Bwlqs4Nh9l/3ejPaWN3ox2J6UvgjB5JHf44ddQ
JR7jHDeYGLYonRc3GtHoTas0nrGrM2PfPkwjr+f9lWuvowFEg0+ZSA4dy9IpoaNrS+zWJ8vYuCQY
5lW7UHeOxxnlMoZVUher1EP5PB810KL7xfBsHJy8oDjD1Ooo3mFam9VXCsZT48uwXC/aKLZYVkWz
eKNXdRddDbMAjOcw7z7yWpXzV9F0RL6+WSJMzXnusDIDvyrs1/Sv+lrCPR7Ax0ibtMj590DWkP3C
ou3I3bXCQ1Z58WQP9I1n8ds/+fqWTkzyedCJUMxcc5TSZm5cGgoGlxYPEtFgAO2UY90zR6Xh3MLx
COZ+BkwJDLRC3zxjjsHZg4P/mnN/V4SGsWpGIhd7N0vV4qighlh9nd/lg2OJ+RSjK/ASGvReFg+Z
6Ti8XTZf/LX0od3SV0y9rgnff4mu/4kJIypYQEk9QH7h740dKLQI987l+Yp2Pk5+JzF6IhueGoh4
HCYJoBdyd4P+xxN/saz+smL0rSR2jL1/HWmvudC/fc8gTiIOIDUIzSYoD4paQjICy33BD/tZC2l3
BJhX4z12oFw5Am7YNirA05fywDqBD5iwr/LYoEOIcYwDxGrTysVLHAEX4BcHh9VxkYqFLSh7Ofln
++5edoi8ln/W6hXoSvTE5BLaN8kLvpvgaS0iSoMPSLLeTG9v9PLWJSyqsqgVUy3R1WZpyiErzjTp
avUMNH4GerKZ7GQBB2QvNgQpQWIuSRBzUUIgzolR6LfEgyF29bNlyMZs/UspGzVVKF9W/hfXkH2U
npo5neZzNnf31icab8BWcuvYo+8i9QTPi5SioUAXRun82OR6ZLJ4GuDtF6uP/tCjsBRK4eCQMmPP
eEzzILttdLGucc2NlajrjlpL3KwGdA/UCsJyZZMF6Xvr7vDWJLARL/ke2l1L4pgCAA6QpxEHinO7
poAnsntJttn7w+20G641TrF+D2q8dhOM8XDGEjGNv1BTPTjk9D3yex0gHEOy7IN9J4HCwT9CZFEE
mn/aVaKclAsug4WE89YBIxUdsJICvjantA9iOtvGuLSDtCsYqA3SfGWAAuTyL8ZyJKchHQFcmszc
G55Vb01Gzmd6imZ835zUXohgUYa4iDB8b3L87s5rbvEcn3k7x6mXxcPyW/g19afxAukSBnWrL+Ay
KKVOisvgt7ewcravWfjsBRIahqYn9wCcHB69vGO1y1lpyPNM3G+pWit+jj1Te6JZ7Es47YUzLNhn
Y90jaEG0ewNRA3WI6yVXzPJljjEkc/kOrMZYa/b1xkzRIrY5jPw2hhg0eiN5lAZYW4TilX5jNGNJ
XilLP00M2zMT+eqe37kgZV5ckCEwQFbSkRVd4XThh+wd37J2hR8BDrxALMnx0h0DIZ1XLQuEjY3n
l6dRb4Mud8Bt1Y5ogGepYaPPn6/Jn2EMv2rJ/UUoLgBL2O4elAh4G0tVG1SXvs1bmhhE/xJE5JAf
x9CFLqTXzLkQ0JIrwRYO024zPXvta5T2ZJvW0bto7Qroslh3TMC8m0OrpfiwSjFQXUx6q4NSK/Gd
AkpnYoQvQpNo4MHG+OC6iFY7ysME/eyYjDEOUSTdiVXCTbqBz7gnw7eT1sQs3VFs0REPkT/OeZyj
SFOuo298pYXmPBru8WMidcSUGK1kg7+tI03vN5p1WuH4nC8UceiCW+KS5tjAEop+Ayueil/XOp18
Z2E0rgoWtD+9H3Olqpr1ih3YulenFiHHuLeVqQlF1bf9NxQs/7oNNVNdRa/veovcPVZvNZj2XENO
zcZ2tb/oj6dfFdwF/3Kt3btRVMg9BJm4zSqbfYkWoDr8XP7J3dycK37UgvKL16a5G7H0fiiVrT8U
gy2gIdiOAezDNEZPu2J1b6KayoM9G1e/huahIP5VFKBFX9o99nq+9OguHi+IBt8CQ9ilz7N7yDcf
OySyqpqdEllCOqNLrcVPdr0V5jja2itdsvF9i7kRSHb6Rue1QrQhiUSs5JkBYEmxEDY8x28wnh3x
BXZTAurcKR3GPaJ7o86CgdXtCevYGF4sgkrNITmulLwz1YPmOsEgwn2vZdp8/e+nb57vQuosVMlg
mrik28o+drn6LgOEjCBjC/fEFFJUOAi+oMsCEjDUL7C8MAkT6yE4LTti8T16QsKzrX1SqiEuH+ud
HOJGa4IokzZ05cJzR6BfwJ4TIZpKR9R9hDiN08AEe1euCn1dz4sRSKqLGhXZm4dxpVK0ROzNm2a0
k1epCbAjEjxhcF065/eFbhIwryBkjXOYyyzJDI7N5oL/YVzXjYLLZSl5u3N2pBbJ4x3HhkrJAEtn
ltytSJ0HkWSEMXesHic2UYKt4p6Ee7eHOVb3cyVCWddWlW/H85F9Sc0uxiUsxVaZt1uKCirBbIH+
/v6AtGqlWdhNPvEsHwVhqelkn3k8NEQEYs/Yb0t2Qlgd+a/hhOHUV4HtdRFUbB1P7XsYDTOZ4tui
NORbERskw+FNyG0UEuwELL6s79qdfh1cy06BJyM5U3UOwHSnjXE+LnzF9CO8UpOaW8z2nikWtNPL
razMZCaw1Eq8umdjWd3UVm78nj91i454xYdlQ9e4ysGSjQr+viv5loxnTN/0T1C81rFVNXrOgUEM
1aNbsgZ4pVrDNh5EZlweZ9pQC18KMeXBTo0aS/P7OUtjC4lQ3x3eLij0YfGvuGzvcX1jwEE2pJTk
1INF2KR04KShuW9X9NiVBflzxlAZSbxQE65T2g0OM+yFRixVs6naF/s5lW60IY+gj90sNN17bQQM
87cX1ULfsZXUsm3g2yDK7QgXatHhpmBJ4VAVq6BWsiXxabIzlCA6M2CZktm+1JcscvGrsNMy8Usw
6jupPaOIHkHAdpK6vYWiYhBm6BQhqNVa5JxuULNiN6ekzeL2TC6rycmAPhU1b2InbMgQvW48jW19
ZST4mUxEKtfNyf1N+jdVmI3LL79gVivLNKs5JLQcSSAp+G9v6kxyiFCISu7E4ezqBsWxH+6INoF1
CbOuUiwi+Vt8c3eBR3o+eaMR+e/yohMF9UizZjNk8L5LQeyUeQJx6HWDoI1goC2eAxgLzURKZ72i
686pBNTxKIcNRhBsqPyCVGPRYG60bPjg3fm3K54+a2wrOxDgnxPuGy1dsvs9u1mchsbgz+kfH3zC
kSpKlsLoBtRmAbgivDCstDM0wecxPfXhHME53mUsVwZSnHOqrcOsCpQc+Pl1v10qxryCgozEpC9k
HXFn/WYWB64Z5HFd/t2nPKLPHpTOGNDxIE4Nanj6nThvcjiF/ZxsOx4QAXWopr2KSSLyPd5OegDL
8ZZDNle1WLx54uTK2tZ+p0niRTrDrgGMR0sOtYLCX2oAoTkR2y3wgNQIHluoteLzaNz1voMX9xwS
Oimfm1wSw5i4VarUn8xF1G+cmlo14EdXVW+r2DkOnFelA9j/dv9Fmffj526d9HDMZDWAJqdU45qn
t/mgnwhrZoYFsdKqByhtZY+9A4B4FHWcG8x6mRpW9Ao3Leoix6mNmJ9g1YvqYL2Fd7Pzzay02XKQ
YQ0hZOKdpoLmVF9Mkd72InVFyYv56s1vide71sFECTshBen3f2Lc+m4DwNqPfv87d+/No63W0xRF
vKIz2YAEB5ru8zzeKn9ooovfh0nP3Kl/OP6E61pgLQNd84zAN8Xvcv2Nd+wvKV3Yk1yFjgMulim0
MGi36zx6emDz0pPtheurZghJgbVKM5JFrwSsfT8uHn2eNYJAOdft55XWu+dkIxKtGP02U622ZQos
F+8mG6amKPXW+OByiUVVjh/iDm+5w3QP4tj9mnU1sVt+/kl3rXT/PTy1N8pJyP8m2tkqKJyYjGr4
SKur7XNZDwLLF6Shq9DuGjGakKrRAxxKKIYLpPFpiWuChWVZhcqYjN8jaRuHi9updR+OJfoMva76
WMW+XKplTVh1/+uF91glbUc5hazuqvsRRAwJGSqVKzsCYB1FNkHfA50ri8v+5Dak6ikZdgrlEW44
Mpg12tE91vj6BizsYzDu7lAH2LKNnNLOEhyh5sWJeKxxamSRr8T1JFT8BID+6dz/KYskNYIbugvb
btRtAjSioWzKjYIdqfqkyWuqa578LIImMg9V+vK6g+k+/uHAoZqrNDucdJCZPI91rgLrt2r/dTvf
jjr+sQn0L9s8dPwgR4tYvLn1Ywxzqog7M/hQ+8GSjqiwp4PbNwbpEVpEjPlvLP8HnhCPM5+QHYlC
L2T9zgce2bHlr2mEirgs2nK8Jl0Sndn7Z7bsJjgpSfmT2Vy5tq8NUPAroq03YzpmxXaM3KN/L+z8
7zcPMNn6pFqgyobpF1e1RaXgNoKHwWUNfqJ/sRipVljvLN+gZkIQuEHBticZi8VVjn4WSwGG9Zo9
0N2eFoRfGV78xdYxJU8ugxffBwwJwS4qhsk3m+ZYWPQ4FiAZ1uxB5MmEY6C8NHp4z8int9lpqkBF
ckz3zU+ItKvew3ECXT60yVZ6DYx9RiPnmK4c3Jm1APpv8GJyJ+5DZvKt/dHLz/gxnIfejV8kZ69U
3oPdoKCaaNy6DKF9kjxCLHttwTFMIsBNvgrAuH82Rorm1cdINo5XeSRIZtan2TTm/Stp5Yf4r6gB
KWbYOhGPfT456OyTBwrTvI9ddtwAb2PYEIBnvAdLJL5gKWo5iJEsmv/MlOLvwA1LWzKZPB7vH1aE
C50LhIzHfXOybAMPFYLU7r0H5LI3BWAHAqsFSY3ikV0JMKckTLEuvpnM91Csbbz+le7mpPlqlsAs
HN1fAuLEPaw000Dwxf44uH7GXaTbIr2b5w1zQFbagfaw1rMbbrHfQ8tXNbj69gEJGLdwIxGf/vEK
ijbCb07jqgmgX29nxffBNz1wPy7Hnv11PU+csLV71GggKcZiybRhAM4MN6r0oBkG/IShcXxzwLB2
9TSXtQqWqCKXpZOl2VyfWn7gmevdHaXPAwvhFR2lzxquoC7T9uDtFQVfWL8ihloDSHffhEP+0JMw
N1gZaLyifCia+nxFkyaum5q+RWMu02ie9m85+roiL6zenUx/Zm+rZmRik9xZyy1HCrquOKk7HsiM
W8p6fJKYbifFnXgeAJumfvl2wZP8peUajTua9di2GV0F7avEwS/BS/WwrgijYv4Y55Y6jia9Qk+V
u1GUfxirdm8M+OpKxbSi+5piNtGRD1iLMWgZil4suHNPBy4IEm7u6JAOy0qN4i0llRCI/G2a9GJq
wL9iWDni15782vovW1fUBNftEsuFMFaiiryzNlwdH2NiLmxcv1bNX+3axrrFIl+Xsic2cUCRFLWe
Qlk4ZQpsc6sQS6O2JvVoKUZL2mTwGpvTlbaA/7hUrvkO8LN9L317CYqJpFBnrcHoOtnVphLzoJg4
lXqFojUzFrUk2uU8GcwWoN+5/B+G3niTc5+cnPKWXYOdg5c571MTJAXlz9lGKoZK1/UBVdyBeVY/
3DSeIuIpnZQXSJXIhGdGjhVvcu8bbW0epn5VQFYnUnLC+qWWqw9IzCYYcRL+80q9M4npEIiJlbLa
1jL9uKdKbaFItTs7BM+anrdrNx5T8vf1+CEQnbUd71sH5npxzSVSnqythlUYHx1OfGo2182xrBPM
v2Ok78XquyYhk5alHnjQoFv54rkSgxL+ynpS/G+2NlE0Sb9nkjMI5LkWo5PE9R/KvWqQPX45IZPn
CxRBcduMCbwBsBsS4y7/KsxArcYjf7WP/X5KTwQYWOKWJbivmn8agvKBeQQOBe8+d5JPqhbEb+R3
s82cerHqu3wjlWikMiNnXraj6B3cEvlWmvsF6fBa+dojKRVIkHGd8o9auIMaqyH5Rua3sx3IrAsX
D6eCFM5ifznCjGK4erHeD/N5SqMFcoTZTMKVrvuvA42+txe0vwSimN0omTGvZwdmqkGSEehEoytG
MAqqrm5Rfovh4rHw+1jYRwObPIp5XOuzCVjK8r0XBa1f/nofVgoFOPdUE/0/vYe396U4ky35Wy59
n1/DNkPz57GqLm9hF0q1RByxIrL6Cb204AWOSxIk5XLX98i1Uv0Mlg8BjgRMnpSvMNR4sgVg5wIi
UddWzPMvPgbglSw1lpAARzWMsPwj7VIVospXXavUfYDFx6gS0DqDLA+vjB/kHwZlKR/7Qsbo6/jC
MLh3pgVELPLSy49XB9rI7hAU0ExDGv4VoAWSncX/IBfK2/9LvbSN0XwSj8XyGPdNkqkSXF47ZzSx
9cmlQ1pSgMhoxnvnuxtfqOi1KQ1yk479yDVGlmC40/kMdrYPL9CKfk3tHIJNKEt/fInPVEEeOHIf
yZ7J4sGEHvQhyY0PAD5opEer1BTN6JgIkETP2NxDr0michgqV5aiy2EG+sY6iHs169QRmyY+QsEJ
o4WoCyN5EMvSYi39isAx5+TiWNb1pR5RqcglSg8NYtVcVfkBrqpCfCCjGwWcomqXkecvLP0xPVMe
CqyIRHihb5lyu2270ziVL9tSs3A756P1rvjWM/uoxbVu0RW1+agBE+Ezhl8I72+7Ni+C5cjo1SWz
yIkJ4xrrb24gC7Ff9+DYenS+jVsr6vQn4fPVs1bwtnMH1+GRwg2Z9gBQleTU7nHD13ZAnMlWRdl+
6QKItJXdL4gp5wOF1nk5tyJAO28IlAnI9kx5PzlX5W+zecrxDhN1ILI6c9zpFhIKTY82jrEPVEW3
mmHJsMcyh9kkMdpqP81fBIf6FrLAIvTvjS453HMIGBz0hmR5MA6/0RMWPmS94ouNUIxJvwKj44f2
kzWsaM5TtfHK6FF2CfBbvKmZyBmiAMKB/iL5kW23NDGLUA70mwWiQNMSGxkCWp11h7CkQPz4WnWs
X45FJPZLErIcHMyuByXvAninMDWhDCZoTjc/ppD6kEOPsu3scWOLlhqESLpoRzU7ZTRC520sY+ja
nvzEUcoKEKYc5Ml6GArhjUYGKV+Q7PWqaJdQIrJEaI5WXu7tw901DcKm/HG3bZpWLIMVWukPKCQ0
nmFCbf0MOdMqx0xnRu5nxpkQOqQ8/9RPvCVr+3t5ysbUXlv2kgKtslACJbg5z/yonbDTVHbc1gDW
YvxK3UmbzAtGP1+YFqitSqMlAqooYiC09FoZmHWcnbF5EWCL5c4MLStF/ZigyPXY2YUIrkzmuDq0
9SX90IRc0U9LI4YmcsWZh6pOWV0KDKMvWwn0lMacRh5PdWOdSQQeMXE7OiPbl7689gqpr02/0SSR
xDfRBm8URigHrSgH6Xmc/vBzXc8cvS5LZoO5nv6uf7uBf+WBnTI8H+hKjHCbgc5zDv06q04Du2KN
kVtmLnK/qXRZmQuxedMcLh87/9g2QMQOo0cWoMyGH3+xYKj7C6SUNnv5Wid49q7O3ixgGdWRqUeh
5i/mKMtNIierj5CiQd4rh+2kfyzElCyQ/fYhdzZg1iLG1WFeGi3TUxeweGsu0NWGetV/5X1zEg34
PA7jtqJvkjWl20qfgVsbOckHFHMpcJrCi0Hs3aOHDI/p5oQ0gAJBgZSDEVPEaG/x3w+isXygMi3L
4OOhnQe46ksDnnEtNwVVFCk2MyXUVCRsdz7b1tU7EbBgpftZ3n/p0DeXeyovS8RJ+rrfaYAtd1GC
Fqh2+Hp6YRHZV4/80WQgHFkyDcj9aVkxYecJ4g6iSIoK1QOoJgT0QOpcnMf60wbNgippFyodliMT
QH2X5g3exs3uR0k2udEtPXUj1cfyVmzoJVVjIhHrGSFne5ce76JuXQVkdfnWub9l04UIMcd1TVg3
8tyPzCbmpfMdjMXhlNF0lb3QlgdOBwLiWPU4hl0/JZWZPqaj9VtsHWJdwncBXeZrQxy7myH/FLic
uVF/E/e2N71lue7rWE7WEjgF5ib1A6buoR9he38u1P68H445vZAkeGDxgevn5tKbsnmYgbdfZr/w
Ci2iLARWxcQBnAZfRg3ESMifsPe24HkWuvrd/85a3wfpWld3Voc7CYxrOmheRhUWBl4+W+uyIDTo
I6XaqGmHLAgfmWafsKduzIseIrWQ4CQJQHMcpMc/TFCnrhOJNsaMFEwMZPfM1RefJqtqSftNxzBl
0C8YJCLtcZeANdwey5K0ls7cBIiGMT2tpGVctAvdqjgvncr3bg8REqlu6+yHXsFryQ6LMxA9u6Qv
eDkTAc69EeSVxyjW55XMAKsfdez+sDnnmNAWzkZ6RGjG7e7ACJvGfslkNwkvTm5djcyemYN/oAKD
FHnJ4uukKMueC/KrZOqcIOd4scAbD3uLW+A80niiY4VtoU4k7x4+PjaVUCnt4CEq/U+p8lehTt4l
nCrQP5J4poEP3ChNeJ+azOCx6erEqESfVgSKSpGtLfpUwrmWpU2x5si2MQz1o/Hc4ipc9AxvLFyo
pZWcseNEOvw6OS6sg3nlzgXJKgtXRPuggYBgel6nFRTOmXsywD/gVs8S8FdTtELimxkjpmJEltLj
0R5r1kfKypYX5srcV7yFWFh2xLhvFOouePD5Th7b3WPOrkhH3M2oSKstq7f6BwpykWlgMhrKPdM6
Zdh/TqxuUGqrXgy3P0ay+br92B7MX5WQRJzGCjSuR05fiOXXji26nuz0/+tzZci0DsTgItgjX9By
F6nUnNB450OHgsyNx0g3CqNmy4hLROoSDFbEVRClQJdtlz2uSZIxQBsp7UgxUz27x74WFweSiNaF
PNsChQyUaaolX3MHXxNbfeq1uID4nEGKHG+6abY5VyPVSq9Ykf4FngigyLcfZy0XHuv9CXdT/zNo
GadIIUcOqku2NFSMjhQrM2QhiFPLxESnlcuM2kMbB1NVHYajainzi9ugMzo7YIXmayciH+Pvp7qr
YVye7wI0eWr9iUB+WABxY4Ka80cBP9VID/YHsbr+a5CYW7jDYpp8yXRwflVN1BvOgLwweR+GBHCR
Jzn0ItvgXl2DJEpcR5Mpj5waWDQqUTIadVbEFXLcZg91tvupjvs3Dpt7YUkf4yVpveyEUNQWYv5E
/BwHipuyYibWP+N7HMhVUYtbdu3U14x1eNancUXwgFoCY4aKNPEejBBXNEmG26VT06u0I7x6uf7s
M7NSsEub8mktEa83wQJxQyIE2O/69MDm995fqT+1o4kohGPp9lGII9BzypuHN4QcjX8ErSHTbJJR
dm7SvTU702waHVBTj7f6OWjLlhNalwCKPXrC1a6FxeXy/q0U+lRFOxHGDIHg/dHRfuZz5oMB6G/X
nKkoljFqE1ahHZ4xBnXbf9Ue5sviPxvgRtPUQlVWvldcFGqRgPTi1RBpohZ6UU/HjIpQOmo9gjwW
9Ft1MOM+DaXfImT0zys/TU7c5yPL1odi4wdoZJF0LCAPJiVPg2kayRKLfxJ/g5oQICUCoE11TjKi
udfXONvWMEm7z4t+wmQqX+HPopMgXn8ZaJtqf0E4Cz3Mjf89f3+UF4yncK61ET/5D1Lsm1n4j9yC
wqw8C9wjeOWWX/hPuiOhzTT0ZwuvivCOIHotTpdGg72ybLIyKG725EaZeLXnoZGRxQS82qyO9HP+
H053dxSVoaZn1Lg2xNZY8krDsxNvfid3f3NL0J7nRGXRwXbR8/J2SNYvFRc6TpB+gXF1UlI+Pe1n
aSv+H6Bg0HdRRhVCZC/Iwz0mg6l9y1lBh3GvH+KANV83OmmJJemA3BBLohUG1pTlHqZZ0iVudgxk
KsvP1QxnggP9E/fjxGphVU5KnrqoOrtNTLkJL07YRQ7HkhP7pG7wXL3hlm8EacLr4d6Qo3L0YNxl
D+04HPE+IgemEsJwaRmBFCT+00XX9H7QBG4IPNAVX6vAf+GOhvqMLd7x+bCg0OPzOK9a/wUixRB1
gZKjJEl/IN9Wh/OgrmWgFyDKNWnLXh1iwGa8fppMnHW3TQs/CkIgjgOQSINm/ZgTDnp21E60wADV
N+bTX9mAHrYAzi/ZO8QXHbhIFwjADKB8sS5Wg9AtP+TZDLPob8QmiD1WGKyuTaxKg92L0eTGKG0d
ajXRUW+ZGsLF0QnxAgM3cUPwXy+Q9Ne8LzxLyc7aWG45xlGC3Li+bhVRtq1q6Lji4/StAjPmQKlc
Scii8++Vf0l9R8hQZZrPv9mSsLHjyrwZv9gkT3Tg+rMoaDultqU1OclrTIwr4b21yeZpDZa9MUGR
iRf9PFqcUqxPZuCuTIn10NaXbxcn+mKjg9VkQ2LCYP5ZALeY6eosLEaSOAGXE0dx8OS9fhoBeXPq
FjNfE+/558DBi7Hj2FjIo2duKcAHrpFFktezcv2pn9eQKdzP4DB2E6ggtkgJGDaaw2j7cNRZePGh
J9im8TazgNOz9KzcNVENFrqdi8f/awLZNIMk/Q4xQngLE75qbwwy0AJaW7tX6VIQyQ1Ow5+g51DB
jY7ytXwwHH5SjwMCwDUp1pyhDD1xod8loz3QtnCBwwUM5xfm/t6wlN5476q/g61HnBjuKeyJsslN
U1n3eVkIzpyi7uJRPbNlEgVUk8vqGwuY2OTy0YKFQ9VdCCqPtwFgktbfu962dK+J2CBqzK6vAJBZ
IyHDZVhBlNbhgrG0fESdVOrA7F1Djn5bTkym1tvOBpWLmLPHAJ2ztFhz3p5Ch0KvG4+GxL8KtzIY
KEnwFbhPTlZuSk8/ofnbPIEbXkptUIzvDB4zjaysuwiYCmIQ3FOsigWNQxHybthobAJQKUG/XByf
fkqM6H9pq9gYc8ry+2WkmHp01fLKJEJsYoIBZjMMutURPoPD9+H+WL9wtJmNdp4FHP/LlkWJF+m/
N+Yu7fYO966OH73r7uYO1+u10R6rvEqqLA9A5qS0y/vkEoChXFmC2HhAtQmnBIYRfhMgXQwQyX6f
UvnXwzMGZKyInOjOzyyWqDPBcFMtVx+kKKFc7qfM2cEwcaCs/VsuTLYNgdlBeC9cxlvXjo+mb6aA
zePgi62H2t/4+i6uXTFAGo1m4voKtna9WntQ6sBXA0IbJbbQykrWPt3RQLCsnizh56mEGODxBwIH
QO8rUqf+rBGRdrHUOIvhYumjJt4RTIGpgPr6kAXf04gyRz5J1UGQovJXbdMNW2UiEidA6nU8ZLYF
VXjkxpCJQk8ORGfExHP/v0LAOgLBouYZx7avimtSPHz5dCm+BaV7b4QoDYdSKuORS33HFIm12Q+A
jtgP76Fv0uN1YEHdsRBjZNPAfDdGNaS3vFVy0qSmFX+i/DAW6bSxgpWKRJX9MhYWAcF1LmRGIcAG
zd0ThUDtaBTXwzNTk2qlE4Gpch7/8r94ph7lQVVsmneaUtybyzra9OXSURpccriY8FicVL4GaEW/
uUnYaW5ABEeXzQGNgwbTwtmycL6TkxOcGDyUDMLzMHj2Ahb7HYGPuW31StlRQb+htxTN0o1iVSuy
TdGo1tuKRfO10RWwlv/jE5jY34nwXcnis+88UqLTLnV8b13t1zd+cWKzyBvgfbc5yog0XXpGAr9W
bCDeOo+SDebfhvLFb/10Fg0/rcfr7/hEcowzS0a63gi5RrHEmk7+k9Q2zamnpVpfZ/0Qyusk/IR+
XGjNGcOLTvkmFFlHaNDYFstF01UMYhCd3UC8eEnDsuFz1LIr8su2QCYo/Nhjwrlk5wy1LgM4m8KF
oJrdJ7PMT1guyIHJDSHsg9sO4PhXa9l+l1+lXHsXBSBxSvhBurzWSyXQuv4JoIhwmlwBCFZaUnPr
T2OAWwAd0TulZDnqd2zoSzcvL+zcdIt8fJfyRhMdGbbmEGplIkOgt1WQXjRHQanPgp6PLQSZN8OF
2xYn2biEOtCEydwz5NZZPMC3PCs2ie7i20mg6wPl2rCJuh/f1y4SUHs/BfTw4wjUnUA2qBTvoj2S
6oXMsBD/OK4Eh1gWZBElhFo1IQz169vRAROopergmJ4LkBllShDVBf1NSSfQQhaaIE+FoiPXwoJF
TP8bK18OiZwYFdTx1XlMKoSeolXYGqehcTIcY2rLeEqY2EllN8pfUZQCLQncTKhkqEE/cPSes+l5
5sSGiZxwHO5rfxQmwFD8pcHoCLD7kHB8/fY5FywGBI/DhN+GpzLJX3fZFHV1K4SYjXYwhAusXepO
3JYhgdVN8BLxsRmAf+kt4TQx1BCn2mVJ3CEvK6oKkJb7aSt5bXCH2FKPy3EXDNI9bOSECSSIdhl9
8UloODnQp8TvQFf+SpXaCP9ZVHS1Hpc9LnowaLzPhjEkkyQUk2NSBPjeNmRgnMz12/ES2d9VrN0u
ElxIOtNVjFaZusrogpP4J64eTOwbDCmf+nLie2Z3WtN/0pRwStcc7+7Jv0M9gMtbtIX6VDjEu/RV
uzLXmSBh+hx7hV+fNzkJpD3/vhN3WvI/qsL8HxwA0Uix54ujqOVm5t76DWenBFt0LZVWIB2k2EZh
exhTP+S+Jr2erVnxBp6ribKuF5QUFK1uIE6Z3HE8ceWavLwHCiFrgdOLv14Ucy8XbJqJ0/sdt4XG
ANC5pi+AwuKbex1WYeuR6qrlp/9SKjbqrzDgdW3JvSuS6gAy/s9AUxuSR8p4k/S5Cvmbk9t0N2UN
DusqNdLtQn8nLoMbGrfsqz0y3Eqx5xTyFErunddbKfJheeXouI4JMeaZTDvcxsaqoelYmxtrTP9b
3apIBlG5q8JsJIbM7QVPgui74BADBbT8UFpGY87djNgNCI65OLNbPZo/WQgRKBl4ehFjLRLfDcBD
XGs3MfV569mraU5eFQFx4j5nTXCLLGnpz3An4L5du07soJnJwoZqw4fjA/KRuXPkv9v0Xn9sfXDr
evW1NIbj1NgHYv2kceaEHDKMwTIp0q2TQVw9ULsWLVO6JPld6x9DiAzBiv0J0uYhIuYdewAjRLCk
wNyO7ifhG+Q/P1Xnf564LPM0GiCyC7tFYjyuTTeqhLQ6zKbYYYyj2aWsb4sHqhENSMUX+JV5Xkqt
tzUOuVb9+M4+U52a1LavSg8Leu3vzj6F+hU6E8lOdmLHLnld3efLn3uV5+SErXBsO1Fa8cNAUkY8
K38EAGLXFwjvRjWJD9dgVFoHsdxMfUamginZ2lhYMnp5JlcPaiQi9tNYM0HlcZjw260QXm+iMVDB
iEHfbGpyPsIkx+vdbMYW5QgTzIfr7ExMT3m+msX3XN+8ZI8Dj+KuwGBhUX5a8gTMzW3t+TD3FcWU
A1LBoTHDPvOhUHkTKhyVjtrIs8iGSoO7AZvKgBpc6CHuddL9hyyt7rCr5pTAn+u83+x4D+SPkKcw
3VyQUtMRTlzympC+MZTO7YFAWyxmDu8AZFneQa3nwgSP5jnwC8sjJyuIEdGMQwmto/GvhU+Ib7gI
ohyGPoGudBn/DesZkIGV/GUgWPxpz+xqAFDMvGM3Rj/ZNsBBb66ZK4fEESkV97bLqgE1PHN8998o
7HSRigyCQ03il4oWyd6ufkWvCxJL/5N9nl+dTloAQOJTPBLTs+VvYB+nPV3Q6op80m8PKrzHHDQc
BM+RWurk4f7O45C0E2awmUluLt1LxS3jMwdIoLlWGf12EDh9np42MMHi500sppBbxmy4d2/3Zbxa
vi0VZ5mPjf376PP1AduhYSe8z4BzFHaFQkBgq10QkQOdNuv/mb7ttVerGIwlW3bwfqZMySdG9qPj
ICjtI6yPtBnZCwUv986+dbEY/gcI+gpRoV5BQR77q8mJ6Y+UdRg9cK7AJ38HsrkDFqr2kPGcIbtm
KXVf27Hlpa+hBpiw7jXffP3qI+QLXU1iDHbp0yeoTLQd11iH240XZN4gf9OT2DXSYaCiiQFhDDQq
H4jqD3TeDAo1U0h22LiH6pviRoGjjvcGxaGeZbLiipIJPC4JUQX7Ib0OQre5x4HdvklEazYeIY3v
g2W8fn7j3Pu9FMQwgbIs58D7vZVKJ2XtGISITxltXRSHJgvNKQ3pAeUNnGp8Q8G/yFPqIT1wG4Kh
O5rXllYqhDlYDoqIpCIw9V4xL/v2U1GsWOaQkrPo8QCWJMdhUwGbTmUtcJ5cXiGYFTcFNCGJd/sv
WZ59vfsfzMnDYGyei3sRwUDcfmAXMkPQK23BKOSu6kee7Nm+vSPPiVbrRXSQNnOhdB0CqqQOVTFr
uhbEu4lbNlByOIUNiZphwuMBBMUTxvvsPaNNkhV/x9QxGI4r0/QgoPMCh/nSleYJYTWatJuHppbd
ZLzt3hffx9iQxgInqLTVfQ1g5MZ5VNgvD3wAcp9IIMMHOoYt5njrqBhJt1X6DsDO5qmu6ucPPvmD
Bn+PyQIi7lZJXeykRj/OTATFGdmYmmdtju10cd8bartPLiThYdPCj0QIqlQ+EGkKA4yJ3ZFZqudn
G0hbrwIncmDft/SBefQzPW6y9Ls+A9D+O5QUM54MV2ST5dJPa8VbBlm3B5EWo3GLyiWnub6oRDlt
UmMDmX4KhuFpB93p2ue1LpwGB3xigesycfyK9oGVWkPyhiR+6b3ZEua3qg/RxRODqUcoo53hh6CB
XgXNr78l+XF++uRoyfE1VveiRb1kZVmBd6R4IhYEldXSH30V58yM0BS0aaa0NxNC+YiSbEX/50+1
RsypA3EFM2/a251nCO0BxnproVP6KnBGRSpQaJJBzfo3DbBjvRV+vdIV9eRm0iFcu9p0+hynOqej
u7lsFolblpF1xEkrzslc80QN/Rt2qh1GfnvQZ9v7nWjgOlR3W/lXXIcPf/r6nBrT9dGFe1b8hE6K
dy3JCSbaKVAL3ulX2qxS2EIAq+8fLoD5HHEs4RuOCnE5PGcfQEsMpH/KojeWUqT1t1QUeD5CRZy+
N0DeYLuZEo+LLgGfnrADVvuUdHadqesW5IWR8pAb+3Z8a9puzrGaLlkDDFSq9gKKJvJ5NfX5dWkn
CumMScnfuwz5R4VNAwuWS11FsZsMCip66d6bwU4b4xhCjKN0KI2kFhYEcb2kQ1T9Gt72ImgeWtnF
jp7R2rQQz7SyAPBCq2oDgUOebsOgdG8bnOm+6QvFlSw5u0PpCFbQ08eleNwakzUriDrMEA+vev5b
AV16HAUS0Mtg2oXPVJcCeelHXYSqBCPSRnj0llirjRpkyeVo+ntHtitabcWbWG2wKCFGzzbHG4ec
h7pf2eL5BAClLc6t7vkwWVjxBD+okHHq/nF3E1nVYgaRLPMN2d9BV1QpkVIFI9ZQSSh48duyV3Z/
8/GmEOygl8Q21UaHyo2Byd4RkDH2Enpjxkfh//6C+/3SEtANNEJtQbBIZvrRm4J0ZnM1Ez6iWoyz
pRPMXwMLdpz5MKbUdR9si4PST09iZpi15VCGL6kejTuCmeEMqYjGk92ve31aLubZnDOdEwtakliB
Oe0Jz0J/sDWRoGwL3lq9gOKU1sD4n1X/zgiFlAoGPnUH3xqojQeaATGkbsweP0exB9wGhu5l0CtU
phq98KqNCO2oUdCfnd9eUsrcmLjUxJA7SwTjBupLywX9md0sBqS3Dgg0Wk+W9QqugRn6KNOS32nU
dgo0XPBZeY+SRgqJK01oDv1o8Rg=
`protect end_protected
