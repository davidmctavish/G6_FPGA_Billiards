`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RpZLwlI25/2k909uynqlHNk/cxrLEpTqTGAJZoEBoAdr1zk9rDp5whAu1Tsbp69lE4QFx0p5iNzZ
xcHsB8nAxg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mfhbb9YWd7GmVEV7LZxUjUcjyF4cw0kTh5I/odisjDxzz3sJuaxtjvwetCzuyniVi5qCFu8+tLrV
fboK7DKXGOhtNnzmBQe1291iJ+nPJDGvcpjKzF9u6vDUOLfE4IqIZIF4LlsXQi4daQhB698InoLy
btV2OVwIot8NjMcTVMc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RGCZ2gKG+bwnpfRGUkAjESOhKuK7T8xFPvdZjrAKNPad0Rr4qwz/N3dv8QSFUlCSHn1GIZADJ0UZ
KipaeTaFxEzYNN0YGyls0NB57NCE2e9KuqtyxJpQ345AlspvtnGaFjPw/FwqDzCR0ZsrO3oOp6qE
tC9jrbpKVwhxfK7dXVriDKke/u1zjvNSsOsEZQDHGHFraYu8akm2qy6WoiXezKiRfcVUz4NFVhJR
nsq3e7GH1gIn8ce6DwfC8rMi92YiJz82xM8ctB2Bcm0uyy2ucGSIoD6/DnkZKV0RMy3S+ujVGNM9
aCj6dr+3jdhJ3I86T3uBOgBUtsH32irfoKzjaw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yLWCxDZ3Sr2Tl8/8Sz/sgvzyf1XhWBNCWNR9/qbZmtpgeJUylJZbg5mjwkF04djaaSBqWUSjtDjj
+q48mKmCZhK8qWgeCeTF4YW16P3QGlHxD1qzbZ3EYlcbdbvLOhvipyLwvHsYXgtU/smFUHZghwYX
uuziC2SW7WhSzFxbGBQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VsPi2E1pm2E5F3iqNYf6pEKTeu90TwB40oLPuodyBcdevvo9usgELYXiZ1jpQZrc6PpQi/TSeLAO
N/hntrguQrq3l/1f9+MrqAFfrS21Xt2eODL3jT/WmBuxkcu4QIvJ7MAmJYp0sY8nrYnlvOY0PcgO
PTf1O355+NudRdvZl2p473GTEl/EpU9p2n02sBsGtSXPCc6fhDRjHA5l7IpZbbHlPDistGGpstCs
Qy3NchCKFOYacPUsdMEmUeJAE5gp0GhAZiipUG/PepEfOoQq6f5EPpY0sawuqI774KQ9U0ZTyz6k
nCFBw2szMG5hPfxQM84dw8ZPG0Re5bimvQsIjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8352)
`protect data_block
lSGVRvLpG/ZWEVpwSQ5sjo4UHiDZ8b18T56OUh5dyB1OX0JebDN8WCUJ7JM4dfaN0mLw9BSWd+L5
FLGOb29CqFlRyYtEqsPZ0it81G7NEd7NtBir2r9NjhygbICUbspu7d7NAAenOaozoA2w1FPOs5Tq
M10spFpKHmsoXKNlOMCplxKCA0SFHT/P8PQpQt50qGFDsxF8hPAa4ll4XS+HSyUfujzq9dxQzlgs
Ye2IadFYgITiIVJi4k2EA315ZqnDEIVlLTU2YFZgHhWC0k4v3xjV4225BAq6FmPblBDXVl3rfRVR
FaWo2fT1xk0bQSu/IwaINfnS7NMLMFDCyQ5xW1aloM6do1jxHXxyXkD9+z1Jn+VPSNrlb9bRe0il
oZOa/HnLazGHHTbi9INc9d9AUCdf8tMT4kmj6fB6IImWjv3OFuN6j7w9VqQL4P8IRbvxcKV3+jeU
RA8dFrkzEw2gq0dBWnUgtmQM8Xdefs1btTIcdg+e1LC0jL2Q8jDNpnRkP5MC9YSXxZUCf+ofjCAg
UE1VC0w7d6EOtYKVHSHkXTKYJs59BCydNXNxDw0Hm/0Xg9svlCF4UvLvp3jLCZfwS8d+9RMdZifW
I04htxhZ8hkjifgiMy7lvAXfmKJ5rGHTBO1oydLM/1ed+h5WJNw6CicndBkK9TUEW57Jpl0iq/n/
5CmDhT8KOw7L8HJTD1ZNLIjSSwEEA/CKR/0xKPavzBsOAlYvO1ksO/B/Y50TtL3TUHWcdQiFhosk
IdJ+IEqOtXzKBp5qIl3Yx+zdwTgDmieU8JYRToxV0opMFEcVuFBmEj1E/FyFJabgMl1cs7LG9zRq
uTMcbsLEexT1EMalosPIbCp8utwSjyW35sppJsMg0JIpo4cLXo9ZeNpnfTxNWpY+I/vdD852J0rV
o7C8pJGRnPCTpK6/qAAqQiRAo8O8Iy8ujT8xXmxzrzR99QTu0ir4cZwcFK5rh9TVkRgKQoKEjRws
yjPIWIdlO8yv8IIryNtXNEt3cRHkCYvJtfIZ+obaVIhZKDuWOcDWJG8cPKFFruN9k+fGbWLrOBT5
73cNN2fpxvwVxgBHmgDMWQ/sMyhxOtCmmXe7ceiXrc7uiso/vlyh/aCL+kh4m6EiHyYnXF8v3rSx
ZiFouPJR3BjS8N8QvjmKh4tbWDDfxm2U0Z110JVGOtmvQXDpA8puytakFMg9uKTod/aoDiHmQSZd
EpwTtB+OcRkq0fi8L7hVlATwhG2ziyX0hZ+J0NnIrV6e5vnmNRZ2Qij5C8qvEzvaLh/o+Vg5nO3W
t2r5xyP6RJ6xyxvKDn9cx0Ge5mx6ikf7QVjVj4hD9EIfCIuHhDmzB7gT5TFzMpcaag6u1a6EbTzZ
Xf6Gp9Gd+DZYwUMpt27L/ZztWub+tdkHfclMxBOOc03I/S2ctpyPld+a7hHW+yZM5eZGcrWmMBo+
7q99MZdL/dPqftHztTzCjfMqdhecPa4at5TKGxH03U2L291rH6znL0hkUy0ZLLWw468L43P3Cae7
swNgkikm04BUO7sP5Ow2NJCTBW7EPOr/NWyRDRRUWxaY7oZxuK67jdZR43fQ8IcIwJ4JgyvqL6qL
4Yxe0PQWS2RWBS0Q+eDFS5fbxkKk9fUD54a0aPcy2BFgLtEmzvMXrMKI4S4EexmXJGtoTqRNtzuK
DDTzqUya6wkMHeu4LKqmDx0DndqBhJnU3akLD1Hp4zpPhCk+NHc1BHMy5Udg+mkC5/XPpjIMGoj4
soQ74T9VLrZaQjSZbfcobXFBvnPOrtKvpE7zONK4BTndHLxbfh0VI2sh5LS2bgqg1UGBchM13NQY
puEg7ujM9oPvIzU2Syt1jZI8QByew2WL9Yk59opo0KUhLA5CfYtYkOrDJsPHY0vPOsmf2evsXdZk
9QThr37ttwcdTubmFHyQTqM112WHsHr/HS1fAV2hBEQKdVAYstafJsAHXv1AnaM+ANOpw9q3GASE
VfM/GgwIACukFvzTr3WWYRvASesP8hj5emX6DMpyBgmsvf3gWkNseeZDaLaeDF4FjmPpnjGmAnMf
I2dxAduWAT03soQYuo8qu6SNvV4kdI0Sb5V7CFi8EcFE/TkVTWSmILWwhiBqg9Mhb6vmqeA+4Rqk
0rlW6kFcGXniDk5YNq5tit5G9fC90Rv7ZzQjBnneoq0TAgLuQ1bE6GkNN5gmU1XyOGKCY2ct+sKh
ebS2vc3SI60NG6dAPiY3BafZLS3/OYwjWFwnb8KGhNG9SUNOTwu1L4Wih3HNzaP1zQKYNrD0rSDt
DMzr8jxN/Yej7GU9ktIiopJiWNXvgqRY2+NPpRJ8piuFzGq1FLVuQSynRRe89BoaOv7SYHrm3870
qu7D07P8xkT1EZzMf4XRsUnmCzBzdiXSElpQL3lc7lpE7ZMuSvLqECmpo1rAOhqm5fNrZQ9vlCPT
JrFmR0usXCWS895Py0Y84MOxl9CUHRhBWr5kIIApusyGPYk8Gtpr1ZgSGcVhPIBQj589HEpQLg+t
Wc4DU8/gwLiAL+aRHtuk8TlWpt+b8UTDF42O7AplAmPxmvX8yGQSvRdGtZYepaTdzhDT6Fwu3Yfl
v5iaZGv8ELovgR/A2oVUGnhI7eDt7lfbAK7HWgDk7tVibptxSqSe7hBcY7J7Fcm0JgHKsPxHCAiv
iYVLXPEgDYKXbefD8wsaVKg1YhhqRGEhmBVE0MMOxunoG9jCoqPS3k9gL3ETWs1kxiv3rtPIrNSZ
ygkSeziW8EyfV9UyXD5d3wSCe6P9PJ8Mlk+ERb8xZzw/4hVuFtKHKaiP+bFrI+jT1WKEaTC5kDGO
86gwD+SHqwaYyKtApemCJfngr6SQckTB8GVMoThQyRrmGr/weH2tfE7mR7f9CfD4uCwzywH7Y5n9
fctxzzHz4QBYwe934+vkNaIDLUdltXI+VKa1iTYlWi28KswOp9G3ZQ8tEXCSpgotxAXsA9fBcDwG
9ijuObrQ3KoieDcVLeQWmOcEuSa55vshudE/1C8WCVvwy+0dRdP9tzK3NpryVSf7OWRQ0VZG+/JB
6vXt17D/HSJeFYciaAgPdG+DqsF372g5c0/t9LqzFbLMR7CdvjYud5dGYCxXKWtC9G+V4kwp+BIQ
rPkHP99u558tmSrJfW6sBDdO4HCOtsQmr51+1RPLw46O6tHBxq0PK+zOuwalNgNByh0qrDoafXQk
V3k5ryYzd63IEKE7KjJyyAQf9XUcYl+dRCRGxI4THowQb8mb77/0JP6c0fCwmOm7t2DK3eGbUdH2
LZekbFW6OUWJ7/R3NApBvVxRl9wLZCakkk00kpCZohCw2U94NddeBbasxZrNS++y91fgiy9xVIb4
0V/gfDxJd0IIptrQABTSyj8KqQZr38poDQyopkr+I7RldLTk5iLOvVWmETbzu9Nn17rXkXtk9AfU
c3iXNDmI+Q6Thf6zDoDpfei3ji14ATq0RhdRgv/ra6musVuV9vkvXv3DvvdWnXPoD3g7w4yaIXBk
1p609NPch/6Q45wIgXBeFilrNgNGxADq4MZmcMMRqBsiIHhfXVYoYFywRlzYYUdbIbKINK7elK0Z
r6mxC0LKuAj7L70f8ktcJD86DBSa7GsUcD2cFBW7rZwmVXEenC+6wtaBdYzRBkFB3/PmRBZZvmag
z60mddscLo/fpS5Lbkgz+BjSH7elDeGYIj9ljw7mcJ2rHZyEMjIVQU+EQz5rPTbQHGplia9t0nTp
bAntSbhnSQKLOBaRtp1PW1uKA0J6IIMGkB0wmiT/pCzOeXiFtnSw+LyXzadBNX7cjiXiTdAeDy9p
5xjDsKe/rpDmZ7h1TkEh75KFqq7+BHFcn1tbAW+ZNiakl8xZlJ5EhqRlZYpGuXpt67xz3oQFkdPd
q7/VBwMVO+LkOqp/pcPz1UzaN7pdZ7RpL7s+p+Gm+d6D02Jcf0zAcp7C4BT7X74BBp1q7D1Q+82p
NklLwii5ya+k5hrbjuUKl9Vf8NeGkiDyNO6jXvp4vlR+ryT2VSEeR/49fGWn8XDrAfY675O+FzDA
cOzTz35+3pDu0dJBB9S0MqUwxKGdooIiZIDbN8PU9RTKPenGyAxcBi/ydpTbtjoXpuMT9yHpGgGY
o7pPPVtBZ517fRALRXV7huZeNeq62wGx9ahV6ygU30XeZ378wxx1LU91gpkCri8+yd8/Kp5gQTxy
5PYJ1wERq5S/Ee9wn5MXptOX1fQi+B/Fc/9S/D9QaVXwfv+kb7pMg2qZMaLy8gCsUf6IIVSFs5DW
OcAnormfkwEEtl2burV37R1jXHK4bvUHD2ulMtssJnnKEWhx8N6Keqee+HRvpYszhQAwW8jueRqF
S3Iwd6duCpxCnm5Dt2NdFSKSenAYPViic/J4FaaSNEyIxWAusphxEBXP197NI1iEnDvvYlaqUcFb
L3DrXEeT1AfqDGaqcqjpWzXs3q5R/RIar0D04rOCaNBJw2EiFLMF61xqALoQhjqA2DHWVC+awyQ1
PqmH2G2fYYzd7Jee/v5Bm9vcghAxj+w2Mwxq1zlkBDzWq/ELpyvHFzzxd3YeBvMcUaFoxMbu7S/I
BN6u4agdne+GqxMlL+AOAL87FWJfkugTXYwiu/QHH9bXmnjK3OxEMX2/9A8cIaZ+Amsb/TndsL4D
66/CVUp2i/fjVsjgNXOjPUk0EqBuVvPvN/XUWn9PbXNC3Yv7bKKwLyl258txqwLWkTUj6DWRsxXF
pn/h2D9QIZn0YiahGRjHIYkUVc9hpWfCJX6L5e2XyoZsb4PlY628uU/059piHVEi13siTYoT9Cff
mMh6CnFJpNZgw0TQPXUd2BFoZ6+qftj/PKKJ77AFe+YVzSDr0wyqmMU/X0ulys54baBZXIi2oBJe
0nDoDQuOnxQxi5Yei4iH+4zIDtZ8IOmTPQCg4LogOlZa37a6IKItJFYxy+S4JLA2BHbMKfXt009E
CIdGqmuSavh5dXnbQxZkVfM59v0JXwANrfSP8/LXMYSnaoQ33H95du9L+oUWV2JctjgF985VhgxK
vqvKXnc0ANTIqiPFoGoxDYuXuQCyhTJIO4E8LBBFuxJdNSemypi97AxJGNFyvP5vDtaGI1TLWpJV
LmILDlt5DZ/gClFSUHBMle2jU4Tw1A4CrucAgYMOyBgmohc7VrVRA7ddoegYb9d/0E9rS5hcuDDu
1SspIBZqbZfMiBfbAywpKTL9anvfyxscqxEkyi7Kk3fxpdCGaYMvBAs3BPDQy5vTE97vSiPk7hkC
c5aYxGDBWeg7LuimIkm2M93VN5uhYA3wLY1Hveoqwbxp4xdh/7Zq+qHHImfe0ZgAfzyk8pprdrzu
Zgvr0xsSAVl0h97VN8295QGGPnoUnHvoMNfz5yHUMrUJEqORf0Cdk1S/LcRBapmHG4MBuiM42Rw6
pepJpEdBrZYWqJPibTf1tM4dsJyzwz0+b9g3UWJbD4EdyT/KxuWHMnEbExRTOspb11FnHMgs0cBT
7/HKBwhQlpHsMHKQs68VGezikma7IpXJxu7FPKqP6hQcsKO3o+QbuuLzzF/QlIAATr402+JaOeoD
yrp3BMjyKDxWEOGKRnwCJRQF1IS7SQgNxf6Wg6en4OeuRkSzd1U2MvSDcs8QXFA59eGC25oeV2eT
I/kB2KGxdmyGtxdKDDgoSfJTsuQ4m6p6UJLrOHJppJCuT2Av5Twq2J1PgmuTpJPH8EAWixwG16KD
0yZzFGe5mZGY3eWJGE0jCDlqczPQTIq0aG2Z6SOsMjY59nD0jHNpODo84eN74JX9wp3+t/w4/b8V
RM73xydBbGl4+aKyMeFhvbK3mCy/IozgyhSGmd5zghEqJCKiz7wqhiOltZmEyuIH7In9Z02065yV
eefzDYB89MQi0Ia4wmJeBXcsDRtmsBOGChHbO03Z2wH+Oq0+wm8TaqlcKwWXmmZ+pyZk/x6jGUH+
54Ckp8RXJd2w6bROHzBHoQxrQvF8fCAHf7Foz53dRoZnkkNT9cT3x6oNNruK2Kw6XU8lGFYkEgfg
cTDTRK8qUBRyQviyRVU+DYCcyjXshwsxayB4TNEhMa24Eci6BlKC6UwbKjxlGeWZuXHQJU4ZBn6e
0/Irh7cTgnRcNZv76+rvYUkaITlOEVqKfgICxzYZZ+EhHTHRUy9u3qDwvUfcgPvRvnaTrtG5QKtJ
agNToaWk8mQQkCdmFzzHNqVlFdq0xb+ZPvCsJEOt2P90H+9NwaQ4tiv0bc8+H+Uj/XVg4o39Rvaj
Rjd78WeUSW2GJpUjVc4KtDBnmQREgNN7qR5gKzf2eO0rlSm26jeli4CobDkfqt0bNQYHbcyELGve
XtbIasmVRQvF2YBsqXLBkS+dVl0OL/FOo9syvfV2Pz0iDMuXodLHZU+tbR9bE2Hk6GXIUQjN4QRg
ua2wIDgzW/S24/AB1jGglsqnDMYaPCPrmRxKuwoJQd6PRTzCa5e93HI3ktjbCGO7qcv/PsF8X0KN
f3h0100skzFI17T9LvTAruUeEssqdJVn5CzY3PRdGuA03xe+MLwJErOAcibQzwMs4387/Dm1id50
j2LzlAP6HkJeUfOhtCCo3EWmxK/rLtGq8RVxPhUrVIDKKwUBUauF+0sE6J2LK9SJv+MyR8Eg74DS
98w1gRvlIWklEej0W26OBvXcul+WIMWNNFqz2PDj8VG6snI32r4M58ofWE+0reBgoA/2wDz7ZIsX
uroQj1IWKbtEYx91GPqrE7oJEeCJuFDD/yULuvi8Jmh15mvVbdfUSKC3uNsXvxSGP9XUjgHzyVU+
6PScafmL5IQRrmK8a1goM0jcMkp+BmbXlXl+8UZTIg6E/pBRA6lHrJ7sU7lgoIPoeAqpEy/zCEPy
Ay4wE3PcIGiIrlqM8Mgr/6/IpCgEDspDNBsx5tflJgRnsPMwvqfAzrR/U6IQjz8GspilSmWtZGIH
zYNhzwrZCNBRNeRRWxi4jeMgpp7pewn2PWMdf9tcfGTSbDwtw+gCUkqsCb++qtyB1fTK4FoxrHyA
SsV1CPuMwIUoAXa3jHg+6x+UYX9SmQO64v6auU1FdazybSpMYaqhZuckGC2yaIL0maKqJQgT/Ih3
Lq0G1JwSRgVr9YoGSjoPeMYR5MjXRLp+dRe6J4A9Xayls7nRDkepAVXb3UwC+HopeppMLJdtijfw
WKJ3aE7nu3jrjF49IxUmP9Yze5EnSe03r/K/GMU4yKjnA6XlYn1+ItH1/dkb12F1WFxmrUG2tjK9
SYaW5JiXm5DPgzaBT+zrU9X1BNTdSkP0SK2Z9uhWj3+hf2Tj+Tqrh4dCRoq/fAdwWubiv/UKXpqj
l2UPjjw8fPbDcESbFVj8HcHj8cOHYk9J6a40639SM7MCx/QPIw6FGTVhKpkJmhozv8EKFz1KJ6WU
f+Up3mdR5PTGtDiAO5kGSoF7IPa8WmPxtBI0eubeqUduQuaZ6L1PzNDiAditP5iumLAWRMOkUvxd
EabjvZ9hB9odRZVl1ZTY55bkTGsBVcPS0lURYNL3HprOx1IDWZv8WLwpM+x9xggCFhM+WRPR+XvG
x/jdgKnDX3yEO2LbCZ43jAJZkc5i6uF+zZqucHAqN4f1kHC9Lc4Hs0I9Zw5SqLh7l9lmptjMoHpT
SnRoBqHv2TJdG/qHNZvKrXAbMkKgyj9Mg2+N6OJCCgSzv7bgr6EoSFRklU05Uu71yVSjfxp5eNRK
RZTht+Z6g8dfoBOkGSCylseBZNxNaooXJlPRy8UeJXd5aM3uil0UEhQRBPCASSl4PMgnLcL4SLMW
n3mxtNrY5uY2F41evehn0xTM7Gp+Oxo0r5AjIDJhlx/aX2SzVmiY4regqZw7k+OcdvyF8jOUt5pv
WgRopIcBeJb7FUydlHI+/RlYmTkpNuZVlw9G1DCfXrpgUf2WLjC1ENPx4pi+D37a+cE/q5DgXs2A
x3akr38vk9acO6tz7mrvdI8DqLX6/m3CwpyyMacVIosGDMO3dko3bU+oAd6A9X3dI1lriFg7RMqG
Wag0NI2mUGnebL5BDD215O0cXwX2SsmW05ZN+P3xwoQAgtyYbrVjynbQAUVpnSbcnJurvdP3JGy6
yLJdYRe+LNWNm3//oem/fJtYaHTF9CNHNR5nX4RbPTJeNWiXGPAJDqYwxq/3rSBrg4smSJNyPBEP
my3VfC3PswnfoJgEILQywuUIsanx2sAwCRdvhM+ZrszYtA9xh/eZWZLk3U9hHIjXHW+jMGiwLZdZ
t7LES+/EwvmVl2NKK6UzN+HrJsAqcmVifskClvzTMG5dEwl4w287lpPGQ8r9+Rc5TVAEu+UC6j7Y
+hPThBcuyiSihZvGdj78/IEJ5hIR3qmJHb3pnGK5sDio4oGt7lMkbNWch/XabSLFwugnd42gXguB
csCWN9tgQ6Mkm40so7sNHHWg7VlDZHl1Rmr5P17Qdbxf5CvtPM3djHE08HKvB+FfUVNzISUuo1VZ
Ybb5bYDAvyz6xN8/7vOHrJhUS0HrfS7T5aiPzIlgYi2ecB3SE4Nky2wkLdaHuSttcVov6C6RX1RX
qquY9rcAN7IJOXi4ke2RQeLUOWgs8jg+MpdkfDSKCtxXY2cWMXWZlmFrxD7MMu6Fu/TBtrTziPO5
JI3V6NZQ8fKcTtanXVNalDG/R10SSV03caL5wrMmYQgZYS7q43Rxqb5SolspypnWOyMjl9JSr0zv
iY8SLOyMegT7NKv9vhBLZ2F+Ln45ErTwKUQhgmfJVoGMgjiD963mIWJILjj7mFZGHQ8h7q7hCe0P
C/bsrGKufyoQd8Qt0IqcWcalIXhbByTCdfbHJ2DhHBYjfCuAUvZWOkyQ6XZ0RHufJ6YrUb2AvYxb
yY8crPRTiye+BkGZ8lyw1DFT8M+3fy4bCFDmsnYGRwJIKUtVcoUKpG5S7lYAkNbeb9Mvja7JMQ8r
mcNtMXEg8XB6Q+n59oOJsJYZMzCStsXQKAHd+VFw1mIDDzqJxsZWea7LhLRUsrGtSIgh6gfK1D91
MJ6PUU2XuSevaUrgxmDLifHiwYE8RC3/xIdLrTm2/PhjTgcT+BYxZ+AbnlljCC/q1m3IjSXy96A6
FgxxjmDjvClRbil2pFL+zorivftnCJYWJAnu0VAZVWexB/P7MdkQqddFOP5nU4JXaghQ7aeTMyVh
gww9iqYOaCo9PpXcxlkWyc6QGDdb8SO3no8S4CxYYozHvgqNMIr4zsyby0ghYEZymZB21s0HXL6m
K35Qs7paiHHdsiUFyat9dZsMbbMize3ak1pYq7rF6bT19nhGcZepZu9qTc7MvBaKDvsUZ7z/MWOi
vJs9K5q3F/vJMGxUQiy8GLCdkSB0P31nG/Z1ldYN3pAchauSBjPPpCdvcbzybceO0VIleRJOhojS
Q0HunFfwl2cJVLDoQzYPZCGjslXsZqK880jpAVmmub5CufdhfLve3FmdQwPZLIZJOndOVuX2Yc19
tt+PMPrP5PPEEiLXEFIpsWZWsx++ipAUZm7XM+nleKbOSVk/Yh+p1Ci+TX4/HeIj0vTCASlnfdBw
r0iqrVdW4tByfdzUUK7bXRI7h9vp87BsPCaoJZTtfrp00gHL+YdTNO/6lPU+DaOfGiaIr3D0MGMB
zGCTPNO9eub66W/Ahol6VcnvtlcFqmghgeJUJckH+SqfXe0qtLfFW3NL7fV7Uc8BcbElojtdKKBH
RKDzW5NkLuw7hA8qFfQRCxmGDx/4mHhJpRVTsuVXpzU0FWurVlxUFyQ+nexc32L0hlJsTTqcaSK9
Dulx32AkWDzfb9m0WC62NrxMCczpz7+NnNK8l1B57PUKAn7QI0ly60pHo6B9UW+85d5LyphrOWeu
BgkMFl5TCwCTqhCRbk+9Kg5m7UUn8mCXh5w0rHFx2PObAwhLy3Ey0DlBWw2syTj6F7Duyg3j7ga8
7McXgVP3HBjPSh4oZOzdGe2y4uDKnP1vLu5kH5VaN5k7p0Kd3doLJzLAmGvykPh3nxi6qaUK+iHD
Re3DQHakOAQCdc7Nf+cZ4/4Pb7oDQRj3omrqfE2/XO9z5D+zHrqsUn3shDuhduXe8R+gewuqvKdJ
dIS1+9TkamVAF+efbwz7H/Ntms+cgBDO+EjBWJ7tBn1hmaf5ad9TuMzk3xER0TnXmUsitqOZx9yU
7+NiiEf6zC+QbPGJgPKiUER/L3winzpfbegegwkI7fHlz0njM78zfUUHFYBGF1sdITnOoy2fFTDW
yMr+MKCh0cBZY8JiLGBWm5FnMVXLcxK3bTvooULQCnycC6+3SkZgOnT70JB34PkCleXhtUpEp8ty
rBZGG7qa1MKgwwVwJPvfevlifTtuzd55P1kqi/m7JUVHeSSncqxJL4Nwsq+pfLEJj6BE1y7/6vtf
djiuhELTzqh6mYf20GBXFXBC0nN6M1xAC0JQXhPmZ13oh9PQkM6lu6BUJUCTfZQ2rPWHlM3xSgXI
a/fvQq2aFEPnnlQ1CCYwV26Sk5/8r1bXpd3rq+ZBwsA8iLNvHYxMKhJEEwGVlp72icLyttRGZ3fh
RlXbx5AB58lpPIQeO4Zo3IxjgG8CDAvuo/6rYPmmZlyfVeZs51PML4Ia8pJso4x/2WkrrR9lEhxB
q7DPiAmlYkeNCiq1W1vwnvXYelDzXlSsTtt4FY7w4oOzzxmUUjdcGQMx53dQu9CzNA1+HRZ+O+wB
MW/FSstr7KuWnD12IsapHJInUlPAk6n0nZU3HViPoDttHtGOJ4YKWpyXMbsM5UX9GyQuVkqPueoT
yOBggmq1v3FvDQU5V38fv2EWTCNARSqV45D5qS92JPLly4tecPMUl2FYmX0kQSTaCN7YexRkpGHi
18j3ir7XKOAmvd3Cm/9VCo/L1dxAoLEmA57qKFBwlmWMQCMAiYx863Hg2sqpH8+3KjEx1Dv0rnil
q/IX9RgyXELuzjCAmsrRiPPlKMe3BjihASfPVx13/QekyIwiAfvbuoG5b17fv67e2K0fRY2CKsuu
IXYQQsBsOmulTXI429T3d6oWjBs+TdSFO5Fn5D50+ORCysRK2Ce0jwwPghWF9SmDL8ZnFGUmIJ4D
JydHfa7qKoX9rKTco66i+vece9TUhwPb0mOraN4sLxnasobzYQcrOK6E4PjTzhnvRXRDNNyea/3f
KaM1Ya8DnqwvC5Olih0OY4jcB/kOJ0EV2jAepK+p
`protect end_protected
