`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NFdTejwDVm49L8EGflSeb7XcHI2XkRoEEd32aVmkoceBbRvVvwreGBunFIb4DZwkSDmXt1PHYAVc
zKD9afBYjA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FaFSREoc55iiEyiMvcmk1NJWu/bLAmVq0TxEMJlh54PRwPHvX4zQGgRzjzbjCiVjHsy7cwgk1KBi
iORR+13ZdDdg3XKc80OmKEZgXtjEUYhGQEvY774ZWSJHzpu/NbUGsvadq/pz0fTedbvpT2tHsQ94
YFM9yn97zYx4Vt4MQNY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OsOaE8n3U5hWu/vKuACZXx7sY+XepaGG5kL0KCdYk1yPhqWe6PgrFEXohPmimrTXmLbLSpo6HQpi
GQn5r/Nn8lIHvrFO/JAf6xawCPM/djc9fCKjbDfGdA9vISFs36mLiWBzvheYsZ1DErQaiuQJztEz
Dm7/C6GTivt6k371TBj+KsTUt0svqvlBwPaCNE/sre2Zl7AXns39ubV0PeVb6G6BbvWrKb4X5g4o
5sFHg3sD6Ztxd82MJscAy+8TFS2So4pUph6253zMDEY5fcuBRGupjX5oKppfuhhkWi1yNcWUX71J
rx9H1fXW9Fc06G4FEnHWBJYSBnB/qW94dz0CKA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
09MfAZkDeKzhs6lrm51ICk1D2w0hyZ32gp3fYfj07JmZoKRUW7Vc5j8dF5YTAVGf3MQGKvU0YOba
Wurg4L4EYAOoGejThIScude92VeIVWLCB5s0OiSh8h4nzjcKy0ASSzlvPF+HC/8TltQ0odXgdKd/
c+114bX1HNR/zEp94Fg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZsyB/LQoOe5hU/jgz1FbOfv8pehAozorYmeds0WxVJoPmhhKjRJ9rn3cpDwqLylBxMqUzqWLUY2h
UQtRO1zZbnOjnBHiNx8AyiJjiHL5yufmOL9IqrNrS8q2TkuxAg3aJ5YguUspeyUcRaDhrA+QxygU
v0Xb5y4KWz351xJH8ssQ1vJb/a4wGJo+XQadUVipfW+jRJ7I7vnJs8c/gVKj9gEbDMIiD9KG5ss9
RbAuFcgxcUCXg9k+RDebUAc/kr8XRoCHG2XqUJSFxJNpTxFBwwZOjSb4tB4d37UDjxEsw3cEQgLD
gela+Sw7JBwvE4jH79NRIpzlLZ9AtVElQ8rz5w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15232)
`protect data_block
mh6DzwMpDTZ468WxeaxdVbgYGrVHw9OXHkX+U6wgjI36PvJaYKZk9DfNq6cqsnMUnO7d7VUbC2R5
nTPY8LKThXSXjC/dZ8M9sTDvWzk9UH2vYkRpWsJk+ZjJVFYpm+zRYlvRvAkrUvqlhIK5oNzMSxJP
r5z1Fo4KGLRw9NDhvc1sa+YTTTWfPBHOHEkMwFNNBXZ/K+i3Gx5bpuFq2G75mBdHlnL8IHjssn4C
TamDnat1yO3fRQMmZia+A66bbNjvgC/uOk0qvKqHW/FmrGokVM23/276Obv1tnepAHGUOk1tjVbQ
QT8v3y3Ah0QxZScoQ8e34DCuqaH1b+mOTxgI0tyOtFLkUN0NDIgI3tnQOwXml1v1oLl3/nf6Jt6v
fiujfxN0kNX2CkBg4AEqveXetmzQ/Puotw37R0AqfdH1dtJ/g0alOhXKyA8RSYddMRXOHMro9vHR
D23zRVdgrdBCNrEjetwjRywb7mhDWSz2ahrVLNGvBzGCTmMfNxUgfjGdk0rt5uXZCJDG676V7eWf
EdPqo45+fpbBwBerHN2PNafAaaNtx6dzKVjCkHYeQu3wDzu8XtjYC+cICEMicUB+GGaf27268pXX
GuBqZE/aX06OKF3nrQwHodi3kQpQYwa37EDEF2R4WvOTWBeAvXt8QB8GRkGUZvKHRjkbH+uyT95Q
cxcvCp0RZ6CtCqhruQhv0UxXgjXhxlqTXoZzkrU6Syruh7RKGuPDwuBNJTCab1FrGxAXEtqB/4TP
bO+5APYYdRTLSJd/RYNZOhU4zcEubuMc8t/gyuc91g8LxridFQqMF5d8O4H78yCMyNc833dTydPX
2QCYuNiuvVQ3Zen/8UcVewd2Z7ST9kdfhYvyZjOGNs/nLxL1ezhZEXxEcOnL2Bg13U3iHgLjMveP
pS1wnXIQRu0i5SMZC3j/pYCqE8x+wjf7C40XVjb+lu/9/3IJFfUEgqpk2Ka0n8pI5mN5COqvqfFC
b6yaJQP+MeZlBteAepkb8azwt3V7AdDTVoGsk2jl3s5eZ/hIETFNgp4PCQIzOSj8OaGlLQYYe0Yg
TdR5dFe9VK01Zn9wiHP3t0IIL4X3ht4VaMEML82XJwrG5smrxBTiZqQtWuS6O3f4x3zPFoDmSCyz
ip1Z5vn+SJ4rS+08+Po74XyIgq6liG6vKERxMdYCGVTGeIhtu8hI6YgsO75s60OIiXTV2Qw8MxBK
XIvSZ4pxPxGPmZ9LqHlv7BxQVSI0QqJZGXZylxdmtdCuv/x0TCnS9p05MJGWCD/YPCUQWiAIBmVS
UVQblWJ+W/7WG/svDaVdkWEaPOuMtvzvmJLHet1tGrLef39uhv9+INpVMmWCAWJcYLk0HJjuywbe
Yvb6vqsRzRoiWtlRpBeUGz7iV1Ufvi/N/l658qJvUkTXARx7SaLkvLPgVMh4R4ipF/P2fWZtu7hb
JmlmisDY1wTZLB6JgfKPNOiXzQydzbOvn2YluQtMra1+eFM29C9hJLfaFWq5jj/Vz3M9DtwdZgFD
obX5VUy1Aq1oPmIK3HIdsXSnyk+k8cbFAKfzlqprZCgbdlZQLqepklnwDfsW+UwiWoO7FVLGUkFB
S3wyEMM/9TlYIIiuld443N6RIP/x0D3uBL/iEW95Y9Yks7aji+U0L0ZYxgO1j3FlpEJ8q9Ey/mF/
4qPYfwPk4aTQZbTduAKPeTbIaTrJinzfiOuFiznCNQTFp2rFjzheuIXs25Nzj8IhpnWtpP7vIy19
FNWowFzdAG4yR6xw0HZP+1nv0MsiU4nhKFRwf+H3ijy5AH2CfiJZGhzybkGyldOza2FTJg6hdojy
jeBO20RVImNwFefIpvnAjpKBePic20OHQlzdDH407ZELS7CQhhN0ErlH4OlCsfav2Q3yCbqwLF8j
ogOdFW8O7NMxtG+gBXO6JQ7lanKeokLAREhNUW+lkHq1QtmrUmYBp788C3k/op8f5xPztMXGsjjE
nEvwgh6Ztlrd1rmOLp5Y72MaeE/nqCOkdAB69J/QOirNB2OsMQLgdAu3vOuko9VIhpYxAdYF5kvb
zeZxT3nnxbDFc15T+VyOTunXWyU1egVgAN4E5JOxf77bSdUCKcWXfScGnKjSpzqo7iACnOrOryvT
qIJi/BqdWFuwzrQnZdMsJ+wgcO1euJilONXXr7BVB7j7m9gFSWdaE1UjBN4MQmDjXlNZSRLp4sk8
luUh3dC8A7ow1frPto9d6EPHdogDOJ1wZYwB8ns5frekjoMi9qf1g0T1xc7Zx7kcOCzGkwd5b/FK
nkMzLZcKk8jb0i4E0BAMJD/u/Q3XQMkIWn7hNnRAh87xKQpaCpHiB8S5VG97TKxA6uiOJV/2KtCY
rMMLs7uy3jm04d5sBUO4FQKa8TuwDG98KoAXgO5QI/rwMTaX4Y3NV68hdSMeKp410I02QMzxwCex
JfTH9k+O2diDbN3QlcS07J7bH2tiv6NX7MAvXmS3os2VSRisA9xXfnCE4l3YXOxLwWn+0xt46Jxa
NRZYkRTWFJ9WCdIkJKIR6/i2bngaKqDjDnyuCFkhoBrydxAmS6aeKXD4kqW8B1j6AneFPfAzNtOu
yl7Z6zo/u6hj3o/m5oGFek9COw1gs8zWNg9vmmxc2z7BE2wGxOJfdH3V4FMMrDvu/T4kk2Cm4PG4
s2pS+IXppTfNJglP+9NO0hXtfdy8VFEwZM+UFoC8bNo68U/FOQsmtHCJYGlf3JTx0x+LugLy9Ams
f6MG5RU8y23pKyWBoUrTPTk5eRnije/kLrIu13RsWwck+tE1w/zYOm8ztpSjKRtViNG8kHLU/tVE
Nr6tCsSUgJyS5bLXWAhL7NmY3fCkAzE7Y6a9JtTh/6Ew+ngYevXTxFgguqMYVRzc4hiHDxQG6Zw5
Eau2zyd4BVZCt0AoYythxV2hF/n6vZpeigtiA2TBDAq7D//htMD6lmgd1w3T16M0VYYTA2b68X1N
XBY5THmC0it6dmuLoLS8RoisEcXiyR4ZWBBirg0/LDt4nv6Qn8Nzjd/QtrSZ9Y8uXLpMncJk2Hua
cADke4iDz5Y/xKOPeeRprLXXYZDbz7Iit4P2ZjQbwwr1ARckL/zup3K7Op64YWnaPOSm/JiNOML3
RWtZKm8jSYyjZv6kBNvwMzpFS7h0gzFxiMptcbEbJdW6EtlZSHzpKkBmGlh48E+qogpTUxmCx9eu
lgyjQ0c504IpMtqAOBcYkK/7sZ0ERuxk6cTbM8JrQFMaMLrfXWH5m8B8sxkDLsSeDCx/uMWaNO03
xQBsSuWfqz+KIKdzReIYQb6svpJu8x6PhErPceVOen34vzLV95aROxQk+Q2XeWsnuTowRZkEboCO
cqbS1+/GeAcUIIUe1760paQhH7JYB5970nlIw1Z20t7gQzb1fAVJyHb+AE1IwyHqojn0mSbF4zcc
z3heZvGLI7gNM2LPaRWRPKLypTqBKuHW2l4EH2aCIHs0LKtZJLiG8NoVtnZDGrlQgonYO+mumrdd
7fWdmidUcXHLcIcY1U/lI7m8dPhwMFSy42M7zizqeD7lxaThsdiajgQBZBq0XoUeDLeQoGmYygCy
eCcpOgj54L5HGqmiBzkW0CDnGiuCqr4iRD/m5t5O+BFFxYd2Rt4lJ0R/m3hUv1LWa61kfkwR6SJ9
vPSxZ6EoMLhunq8cBCfpUWCc/CYOB7/B274uEEw1kiVe6Iov9RhS2Hk/5SC7MeiFtF0ea9CKDG9E
QxnHxWMmcx9qJ4Rt2TMrIFPr82bsfADmzs8+fnBAxpQHQMag5CcF5IYKkgFkeG8h9kSciIPg45KG
byCpLC4FnNcarJj2/wh9eSS8XZC23zIOmek1j5+wKET0VCj+gBOHFh5p9n5Q0b3cELS98e98hdFO
tHqIimJIK1lrXFZEs0kd2oSNd0G3uAD5w4dVyRGNZkOo9addNgehtnPjFnHtyiILZK9YYtam5cM6
9fQBC9WEcufCAkerZZ7ewNWpOHLgdPHVjW1EWBMU3LK1LA6xDEJgp/JsC/+NyTRv63j/l5tVg6tl
UcdvifaFNL7Ov38sEeA3rNjDE2knpjs/SzZE/4GTxaUv4CceZvrAuBkugGz0i4mZxj+8et6UyIfE
gyqrI6nKl4cUR44c8UrVkQcT4HmeRfD9KeGWeQ9ESaXEherxkpqqUG2JDHTWLvYeHm/TZFOKIXaj
4uA0TMnXKqxuKR0BGAuv7VmxJR4XgXawMBPi0361YSqzgapki0Ye3mxUCb2BTESxbMrE3DAYTNcB
jVdWa3DvsRwA/dZ+X3NJrnJ2l1vZhlEVHQD1UvL46A0xH4YCZvJNGWC3RRkVXFKR9QLLswybp8tU
LB4Dzfr+2s7SfuorH2h/IMY1bHZUGitsyRc+g3TLkSYjTXz6kIJpSbXQrS1+ZupiEEL2lfwMlBPR
KJLFc5NZU+oLv2emUt/7orutstm0tQqRNZiCDoQQLDlVjwoYPHydw/tXuUNTVoFzRu5SFNFErPKq
8cGFwEBhvTW6x1bTcv58UHMlHyg35s3+QhlN0tyToESp+4wzhZ+qPXuiOID8nm2zxIw/50sYyhLi
TYPCft99NsVUoHCcJI1Gsf/I1ilAppAxc4HO2sCJ2Rrpr4cZHs8mIkqiPz4ciY5jdND0SakR5NK/
lrNlDeZbU1s8TdreJySH1eBiNw+BIGlKNCVl8Fat/Q6LXdCnn9Ua3WvaH9wKaLesa7QoUNf7/Tzr
DFpIQVokQ3wVdUHcHF+JINK3rQgYzo2GyTJqdjNujCEefyU/CTI1ra/tDiTVWRNgU1c5srkww0SX
ojJLn7lMjDYZ+G8CoLyVuV9Of07YdZBdg2+6iSmuWN+Q90HSDBXdTSBUcJCSI0/6FefpDGEbG6ZQ
kEFUpG5RITFz8aCU0WwCFGLysAnGjFaNCPcX4kDstcsbT0R9x+ViwvICgS92LUn9MeBL0LFFGRJv
sOV8oukZ6VmLztRnbUAmaBy5gXUF04OaJzW7uIvyQAGTNcoHG5ASN/fB2wL4Z3G5Ssy5kVuXX/mT
ZZ3GzfQS5ZIbFvqkhJTUhR353C/1WlKwRIUrWVMYeThN9x8s1TJcYb5FETbnw+j2BAslQXJezuQo
fKFIgeYKcYVZ2Tji6A74mOSHh90l5CXBSuTtDFdB0fgvsR4uIkF5QO1miyZx3W8XkhhmAj9/UXJZ
vEanoAybH+vUU8dyfi3+P6R827fnkrTbSOcjA1Q1af5uFHTGfyxJaR1qMMwuBX/xcrjS8HJG0yIo
NQHFUfuN7BoKREdnaBTjGzFO7j9WgyIRO7psMlJq7hOqQwESHZL9fEVIowf9ufcm3ddY0QhtDw/k
tDGfFgWOhafWypFfz8KQ5fq5z2iR6vtPt6lcVRmtGkv9NR90dKBxxc55WKuxGRFxhArLOMbaNOcX
6uYcv89kXurROdUY2wat25dwcNgXIaPggw9gGgPgVqG8NVPq2f2UuRX1Z2bf8xhSd/M72EzyzsE2
R0+3ER9fG/0L9jHTMcJDs9sSzJA4LbRow+GK2D0r81mnlvBMWNMM2vnDfQdlbKwutVTs4PWm8ddA
7utqjsacWFVrDo7n0raB6TRNWbUXaIpEXmDY6u4pcbY43fLqBkFbDAA9f2rvekVwGTHzGTQwIaRg
t/VnUtdPaVphidBAfFmPIIfshKDbKymJrZywycoVVARtKHe95uJx70gGDXJaDdLfnUPegX0w7gBi
BL1PAiS9QQnJnVIEma964PoEBn3CPvEc6h88zWyifOSBW7zwt63lbAaXdjHsKd7jJAgCO/YiZ9J0
gMyoNsTtxRrV2Pn00DY8OEQYdWXTx4C2JYYzudSm2AUssYC3E+jg6mmq+ZP/5atzoXpIcK3ttpj2
S8F5n3xcxZvdsqsFDHU0GWKFPvRKFATDbziuUIeGXhEwwM2oZx4dtgm3IR/Gzbvivu07lr/tXPps
1DpakImNg/vNBFll3WG2yWomb11x8h3v5uiFLika/L8F1KrObv1dDHJas6pKqmtH9lN+8/VvA9gq
HV+zjhWuWW0n9GgxZIeHlhNEjsIf1MMUEo/K6AkgsIjHsiBu5flajcNwXcC9pbSB65i1Sd7JfH4z
aUopzNZQePA+ItiFYqPIAVI1k90Hk+LFtIPSkZu35P1Z+SiHHPhb8bmpbWK/VDrq2QuFoNY1bEjJ
JD5vmhWtDjNMzfjNVoxtzRM6seeUxbNHKxGHF2shCib95TtrTp0R+Ux1EhmGAfrHa3riiuz+M7cr
NprxujdkryGUXK140Tr8Rzjd/FG0lygBbkyYNQ1n/MObgE0jYrO1VPmfM2iDA9le2ejFQYQWlFVS
JSq5kBYYFrGzIKop9hXRuGdNiclacc9NIOAWaS1ThAolUfUOpt3nLVZrx7TSm2akfYIVl01MZp27
5xbKwDSOCb1NHYEtSBSyyNkeO3spJvw4bQP4vGirvwa+KR+9ntTL5fUApcznJQpTD1w3OIxG3JXj
VLTZYb0hB//dI0HxeAqjKJA5XXJ4Lt5CNfn5CZESpptCOeusrhlMwbplEvjgYKiF8X7oY6V7YUfa
dCrI3dtpDwXYw5PpRHWZJvD6xDUvJAC4s+X2agTn/R/wuZXNEu0g3wQQg0+1QJWMJN1W4ccyER/s
/yoDudxPUMva6zj/QwwPX80CziDgY63w9ogWiLeADlZUALEkTbY2PrCwWS+djYdo96nzF3i/84X5
yOCt2RKI22EiSzAS8mdEUoeVmXlb16ihN/ptSfwbfVb0SNah9yYXEUa8b9X2fHsCSSMtZx/V8JZQ
SuiYWGPkSTxUqgnx2U9HjuAhuqqja07v1O3kCO3wgfPNcf5A1Yxy+4kmz/aRWJtGeBfPWQSjJ8Df
GiQjkeUTe9MMe8rInrfctaEIRN0OmA4J02omeonGprsosBnlXkQ7tKQ9/oIF11/pkPu89FxdatBk
8o44eJtiQLm3sTaZ0/GnbhCvvkdYB1TBGimnOtQKqMijpJuw520sbWd/h4KRCLOiLBWj/+nja/mA
ofsH2Z1PTL/2CqDyTfcMkeEOJes4gX/2xD6Y52RMcVPVkF8YTTjkcCcsQpJKtW+R5UnIKZN1pZoy
zQNyDSmI0QN7pAwRx4Y05VYP1+LiHUt4np2KKrWq9p0xAEemtTv4MNBXtqKPbf5AaZuX+GzcdMA7
+bjY7PLQci8k036dlrIFcETy5GTZ4i9z7e0iaEzioOe0AlrANPygHQe6utD9ezJJSktUA90xCtD8
ly96cBkjmwo+9+a83qFM+xhGXlSEFroR7m8kY1seTj+OuaU5CuKu0Ud95rgZDDuAif3U+kjzVRXp
XO9ODtGDzNnRun6mGsd2lfFVXhtVZuWp0kt0T6FJtfjY+JD9F+acc+dYad3mri8NpaG56ctaMOGY
wGd6l05jJyIDv7v1YnbNDrwbUPGfSRymcNfrhqJb8vLxcAgY2N2/QdInru9BZKlJzIqayeg5S20g
CGQI2bd8TfifK/ww92hgTDZlxFHPYPdI/bsGotNBzUeTXhr35MnoPJDT0NbylBmK4Z1pUAq5LQ6r
4shNe34/F9IDFLAwsZGaoRYo2/MUWs6eEObLVw8CW882nRCOQRlXcivCisRV+bYPklwzwsPgDKnk
5epAmpsy9UdnvMM24nN9tkvgBRdScvO6VXdC0dobP5rKyW4emocFme0BBDdppOKlPs5k+jfnJ0HG
C/XZVBYKkHUzDwXXgQvUfQ7cCUyH/e6ql2B4WA5RN+g3gQDvIjO2vmy7UgWVpWU8xglZVrTuHD25
9THCc/GMhje1h+qJJ6y4O0JyylCS2F40Mrnp6j9nADMQoIKMKrDo1I+KHlwE+1nGgt7AZ15NUWK/
ie/QiJP4vgNSSNrOuYOjOYnZvvv80BqAdKselHcngSaC5U6Oeb3FaALh9r+NVNstZvH+ljU4DM1q
xI6jyUKxs3lC2oXxwVShUjyy8nk5gfoe3st+u/ZJ9mzgBsJoGlMxXpShcQ/TtRXvHHxNggS5s6AN
fZQKVTrtR84kKKMceOCUHOR/9QZCGZdoEhCuZ0Mk93vyRshXc1o5sWsoYxFzGfH6ICukqD/vCof1
qn8Gxp/kdn5kxd0K2pCDAwG9N+STgJrTBPgfIYRMzPgfTGaHTddibXtp8cB9/eitiyrkdw8daJob
78HM6f28D5OanlyUgFaxMLqy9YnKiXmMIWORtHmqef1HkTZRC4ssLeo2bX+Y5UAY8X7sUOxfk23T
2lVUh36iD4+XFjYouAxZfD8+jABNleGJQZCwCTMZIpS1zIA+cZzbYYXCurmBIvfb58T3mMQlvM9N
RRK7z1egLzT0k//nJ8jWydg9TpRmtm5+s1U3crsQSkbp6JPW8K/l/IbyvfCbtggQ4ABJ1psmoLct
uX/DFnTBE7Uea8f58vTGK010tgrSH3pRCA6nH++mpaUH/BUwWefjDev8nNANFDOwhAI9XstzdFIp
skT0S0qmYHawK2bVwytwnlKMEY+/Bwb1+j0sPxzK2g2ckRAfFi+NHGPpYvC2vcYseVwLutmRvwXj
RO7N16z7glJrWbNBDtu4pFxbhGa7UTsJwfS0yq3PQ49QjrgrgRuxBz2xN4TWFc+AskuUmlwNVOMJ
+jEdH6Z2JEKjhz0Cy7Q38w11IWKY1LI3O3msV//llEgksgYRSlUaE3AXdlDugFi8RF3PrP3LGRWX
ZcxQn34b8X5bMYbpOCJqjzRi0EB6SR9hp+2GrffgKR4+QLJw7Ag6pZ/83qHE7U+T/BNC/jz6OmPX
KvS9/+E+WXZoq8C4EemWzQmfb8Q/ryhvcFDNSBFEMyL1hsD6vKBsOpFqSHHVUqUH/ODbuirnunYm
GjAP0u/WAGxzELHC+eUtRAzQaNr+9gG++W0nfDZQwBSL2BWR1NVPAEObklQUyc2CdHIkcykHJz/C
b3cg8CwKVY1YblZYGtIa3yu3ynfx8UjR4oUgwe7IOZZ39yK8DtArl5Ek+WxYGXduOVvwIYfIkhmJ
nvCgm54G+A/S62sJya1ZzXvCYPT6gKbSgYSfbn0k9f08vNGIlBy1+Zannh6Y6xv7C9J1LsO70asc
7lNieDzdhfFzsSrVKVQDQDSQido+s60ajZcD03PLkIOs9UMHA1kLTJyKyyM1udfUu7L6Dy8tej/0
rbZuRROHrCq3E80NIihLIiS5ZMWh13zJqyQeYhGwssDB6GqDud/R2Al5/odmKzZpQ9hrm5euD5rn
1d+uCo79UpxUSsWC8PndGzbDv+h8mfGVYysRTZB03q1/to4pL/qYFERMJySozw5/UGnUmE6jxmTO
gwdj+d/HDZ7BhiIOHWch4z+2u4P7MNQsXHS8M8Nh9HY56EMCTunqInv2KUm+ORYVJer9oINV4OYY
smXn4RSuDHMrqbO84g3b1H1cn/JiZPyOKH5nme6xzyrATFlM5GZ5W5RUXhWsHhvbNsm+a+DwM0zY
gNRp+EGnQZUBuKEx9b4N4KxfN5p8+6VotCaB4nLIotTpY3QO+UwJqklTKT2XGgmpPdtcdYhbabwd
X+I3N/6Nu3JvzaiIR0OAKzEH6lhTLbf+CJWfbgwI/stJfh9YXCn91dOBqJLrHkTuO0A0rwYJrAIs
RW33BdP+Uq/LigMQitocf/UdQtMdlOprzMamCyYn/BvGP4j4h7n2X8KJUFtrN2+pOlM8KvdDbwLt
PV0EO6pFMHouTYRQjmop1ol71wTdYygyCV4fDzgubxZ8Yu5x4lDtKTgaDKUI+FGU5atiJbGCJP6X
cSpw2uCXnVaXpNbi+3cM0OiXbtuy3Jfs5p1JfMw2EzqwYhbQb9IeGuD8I6njP71pxhH5WWHdMK0e
Pvr9N8u4gXMI6LLivaI2iesIUC4755aGEVG+4z2JcRdaKRYT8/Zr7uwrOt2HzbkjNlstiMKnCNxk
/is8kYXMxEbm4qdm3+SCpUKRPWISnaSP/pQbCzZOF9SQHLcVLk2KELFnZQLpkmDD5ivVuIaR7iDE
S8SDxDIqnuGrx8iP3BrL8MHoE/9WB/ZcIJpM9Jf0OosV50xOvctqN94P98YYW8WG0OUYPksTSa/D
ZMw2EJDgs2gL60IJhEteSVrvIm835ufZoonBU7OIZcTH1i7GTASjilKflDZWKlg4H7nPsNjpJoBS
mfBi1fbLa64jWfKzziOMJHl4arMJA4cyTHN5Wga3dZbTb15P9p9v7bd9+h4pIRdnsMKnu0lGMjgR
xLIgt818vdcdBNirx0FOTsoo+fROxI0S6YlLlKZp5ll4aTI/zkzB0VqWsSW5InPVeRT46QlTw0Fi
h90KL4x4Kh0/gLm/wk2brz6wZ15uEq51/ygTSxRHI00LU3UYwvo3oBAnfiPJvc6s48868gyAuXnz
RuDoRzQYTxq5r2jSYneAxocBQPeP3DHACtZymlMIYyAEDgbBdXwpuDhTiSm+n/qqJL7VLX7k0tUp
kUI8Cc5EPndGtWdS9YpTD+NwDIdGY3Rgdgg5v3MjkRMSwh2pitDVbBQ0/mSfCZ5rUZRZ5bYGJrie
PjmMTW8osdNZcBogqHqLmzY9t9rpn9RAR+ao9vrNmbm3g5+9AJZTOaCG3pRJYOQvjBY8KV9DU2SA
MGmW6qN0Q/hnhFvfeOjs99FMnfzmN6GUwt9Qy4oPjy5PsyeX6pAy5shBCPmRgAzgKdn4hDI0KZLv
gGBGdiEvuoNIkGOsgDk5iIMbtdTCXwd/Pi7oUwhrSsqOoZao+eZPEKJKZAKwjRMoYTeYZmRwop2K
hZvjiGsUsER+YrRxQlswFiUKBrHi5LjO+MwlKdJtSvFkZEhM/upSy4NaLeYAwO8bjbz6Vx279MEw
D2CH3RXgD9wG4mCRa6SlbUgTOW8BYIod1Nk9L40laZl3B2G1fVv3Tj4WNUtSi6Ak4Q6IVsidj5Pu
SFRlqtklyLi5hD2n606SlM7OdAd1UgCQ+SpKSR6Q1yTBv9X+FI44qZYef99HZheBZA8hrcOJq8xd
GniBo9iYNv20C2JJmIUWC9M6IWOGx1BNF5fiyBJmVqrYrfsnhNCP6tMGojQ+Nvg4Niq+Vi1KwHhJ
WxBb8Ewplhv4+EW4H4NTVGOBjt1tNnmHMaUuTPy59zMO75hBGcaL8m5tgZo4dI/9T0SLMfRtOJdk
zeq2hcbjWZiZdrXQamdbAxQMJlDVndOS+90b06TAiQ/TFTJgW/7upFhAJ1gP1Mjz3kiIp4jHkd1N
ZR8rLY5xONxcj+Ej7ARVnsppJRXf6mJY02mU01CbAwaDKaHwcU+nlWHXzYrweGZDSN4YTKyxmDU2
XBysraJ9mpXL2MctWq42Rrd242DIjpvdNIf3CFVdRnSuusw1t7A8OO2gllXEwgWxDIFyJP7WDJyn
6qDlrCNJIa80rtZQ3FwAKiJYFSQp2HjwaMqz9V3iaK2y8qSK9UtXuTz0kUILemSIKstI610ranTL
WDu+oU6For7Khvrb7OGNINbZQ5MkOgtiAtmMD/b54P+7aPftFia4v/KMmb2HRwWBMB3OI2GxvUcv
AjQFaROKbFfmoT0X4d9yuxRZShVWQjmfCHU4TgI5xRPo8cMvBx5pree41JR8bTzamvJ6kW2GDQ/e
JSyySTXJTNWZsZkUEbL75PTTWQKNjl7lnKjwb/fDFMGbeI7X1hgehf6U68C5znEoMgp8+gX1E578
IJYu2MzcN9fZrh1IbuN1AEDZcILVForyJBtGyD9D/IsQMzWJygJYVZmW5eBEDWprTV6pbrk1Hy+B
HENNH3mF9cCFe249j512zCxF8jJheziydw/xKleoGORJV0X+FCd+1VYXXP1iwkprwP+EsbilWLJ3
EkPEmUAgKkm9a0NvGy4wYCWv2Lru9Rj8lV2pploP59ZhhSm4K82oL9d2fsdoqhiFlPGe6G4mewPH
SGwzkyZXqZ9xhIz+RXqVDQhHNW0DFnvTqBB4j35M7kSMTgfN3/jHpqZzGQDFAgyFPxCw2dt6AE7I
EGvJzLmMo+y4htUGh89oTnu8BdbFE+CG+nj+Rivra7tVzvRaqYfGrAhmCJij7BAG47vdrvJmfi7S
T/AVDoBJJ847E+1Y3pnG+AMZPfccq8Sq/9wd+E1BMrSEF7s40/VMiohbBZseQlBYjr5PGy+8nBym
JmD+D56uCqDTsiO+UGRE8vsGPVtfAJvaGse0e8wNGoK1IY6Ojb0StY5++kpommG3HPYO7lU4uL2V
IoGdZUemiS8OKMjhlMtjerxLKNaYotpDL0ZFXpJVnRaEa8tyqKuuh7gCJkoKx6f5ywgK+t+dIqOo
Hh54/bNEh10zlrzBZnl/shlsixEQlfh/eZVLciM5GCYfBjYGldNc7FRPiQBlck0EiA3UxZFlIgbo
6jjpQGXC6ur6SbwMNBmQ/JrOiRypwAbdiVTcr51j3QEJNeadNoVt0f37HmiaiLUe8ycPzoCjMcq0
E+mNmnC/AkE0QRc4d5epOlTLEmcEhtZVFUz3uPDmccFIEpMmW5q4mifl0rMEzzpvhFyQI7QWX1Zr
tmC3M3102orUBVBbtCB99NLIlLL9xMwFta9Tbt9K76UQ9DeGp/6MhN7hxAj9wdyEH/I7/bJu5Xvc
DEFVPakzzxI0DfTUH8h+LZr9LiQHWz6nAd8akgzhnnD4UoiDaeoUGdD/OIYLa5KMaf0QKtTjg+Zn
6FZQPhaXST/7gD7hJ01kSCY5DVlMOr5U6SxS2X1TvDgOSBMwVsATwcx2445f4BUeicg9R1pKW3+4
NflcznvZxYGeCFTNGtyscOPjjYU3rxznBqJ1D4ZN+DlWftvMhjFp68dzlHtBhbuhUEDbhN9PrGpJ
PwlcnRSFPEhzTapWsTq42XYhdfQdgHdEGGC/PRgDOzdcK4Zwtz4wFlkU94gsQ6PSEEne+6oh5h6X
o/bUjbrt1jfvjxJCmxQI0qVN+9cXwEwEVRiV0cIWCHpXmMELQvPw52IQj7MqD0VG64u9Z3zRgASi
ta0yCqnJPa6A5bnxkSP2TFjoOKJDdXNwqgW/pKEm7yY6xenYsws1Oqm9Qoqur4DB89yTE6tVqhev
0YkXxvYD066YhAGRbbN7kTsvkrpoJFNdRUq9fHOnTYu7RdF1xVbMWyo1O/DnrroGyOQ4g8smo5MQ
djP5QrThPTGIfNCFxqIQLZmBwByhkyh/efaSaEHU9Ql857c5E47GbOwIrC5Fggj3hDFFtT3vH/sK
GaSifTGS78nund+PMsuXlAd1+XrrgXVtlsEoYUGPcWHiFVLMnimR7GwC10x1muH7vHDtwXIQAUCo
DKukl2/URP8sOXyp1eZ8s/T8dPpEcvTT6QpIFZ7l2EgevhLB4+9tr2swqFS+vyJZmaRwQf7rVsw8
jOTxNDEbVfgpzM1nPf8sOp6+XWZ4WE7OPaUBjHhzHhkt1SwTCEf5oUr/2zkSSL7kGqKpMUkayspr
eJYaCC/UzF9koUfxw650s2EYBwLodmjMjGpHOiDyZ+8b5xGqcdd8Pzd/gz9kmlPXeS2QQVxuTJs0
v2Gr6nMyqKSJy6Esw8PV4SK6UvMsxY/I3ijgZFNgcmrFcgA1lkaN7OfZ15ReBoEZiZsRtv/3g0YT
LoqdivikFWkDXCQUDey1baOcHgT5X2eWA/ijVdKvuI+XXV9S7IqyOMOksyX7HagWiGpoRiuNqy4v
Pc5fnz0yGO9+17A00TeMeV3Si/XjBWh4Rlu/0bZ87Nv8bGDaTi30uB4SkgnOWroEO5Q6XH1xYMHU
Ifehp+Eq/dtA/OpaIo0PhHjiqZHGVb7txRaC0i6pHfefyRTAiaFMefXED8UycYkL4Gmpq10oBwPt
T4Nc3y87X7Ei19zh5U3J9ANjWDeBtvWD/tOG8akQQTZ7Y4UnhwefNQlXcKm4ql66nXdqxl43ce1n
49W3N27hCtMM2IU6bSVwLtpHas81+hoXM+czx58aKlSmtfKvrbQenfAK8afP/+HPaTQGQAO6yYSv
vfvl3I2EJdqZMD4fCY3Ns8fMcKvqQ98m9H/P9kR4YlOFSYyKUCEb5pyKh0T368adETTFpRRTGgll
V4CC05tVnAuAL1zke1YmXRhemTFCcyiAvNaXZ6QERc0mAkS4vD1J+bS7aq3yFjj3jBAain8SrLT+
ug6WlkkKk+myNQc+z8UhAfqPpFfvCK0D0ALThaAVpXHK5+HTlTwjbF/mUC1Othv1Pg8ZTgI3bqvh
ifX/lyP8bhvYUI+pmRs1GPdgWt8IKfZoSDzqrKeHx8Nmfoax8SsmswH8oTeL01tvpL9f1eLC44/5
XGqDEGV6o2fC6vy0yqUpSu4nO1KM+6BON0fezrwFpo0E3hH/UWPTvmuvTIJswunWd8mGWyYe0PuU
213Nx4Vzh5QH1UF045OtdAAWS45BQg/G4tX0m+ZKAF98eNs6ehEU8F4KO+wOFDRgrgfD7bDsdGOw
Im7N272s1kLE6RhjdVWloS1MeTQarnXifFe2Wz4sUijJYmRcp6j43dxOuu3yXw3yRjYKXXm+APHL
iFBTV6Hf7K2m3l8zYWQSezQjDeqyPmnuubGlAznoLNYUiMV3cY0UUw5WmmBF241F6CnBBEyleoQw
zNcWvV1sp/1y7wjioKfmy2LJ4txOasdEsr8f7IFHAXxR1Z+8sVvNzXdeUSizYGXUyLGZAkoAxQLZ
yR8Krz1pj0TL8BA4AWW39zIOgaRNxkfdNXOGX67m/Uwzv+tdIyHwN5xDKHsfdGVPIFa5BzVJgD7o
4rfuCNaO4Yx2/bsOVB3t2JqoTVb5qxdQHlRSiq0zAC67/dZtNYRaoT2sIOCsD1DNP2u83SBbj/vA
++1ibLe0X0nR+bh2ZkpYOIFul7FaidnxKImGoVIrW89Gv2o537ySoKAQWWPX5HGHMU3mdksZwaCs
mIzMuxqnSIwnMp8R+P1VcHkrWmC6UX/B20OzGO3xILBQaK8PkoDJFdsxO7HZ8VuAAV87ilHnuf9l
1lQxcqVw3JOdmBunrJr05IBdxTYAoIA+Orf650u+1GtPS2OErUe/f0+TXh2apkMFDRIJdr2QZ4uA
/0F0ozH2IfQRMh9fPfEM0OBy9pcoLUscvRF8IyhKHPHm2n6fEAgZnuovz+msDoUYdHzxRoWgxZWL
PtKtyTVB8nyPsRiSw7fH3q0kxZ6rtO5B4PVYmlP0iJ2PFbKrdFYFED/lJPtSaVa/sfLJ2q0E97O3
h/wCBxbalXZrzUhmjyguGLS5Gf9GLJQzeW6g9gqvZEgluKXmI8oLPVCTk465/doFwZoHEH8qdLt2
wsvBe208G4cgIzqFh8xELg6klz56IcHEF7YfExdc8vEiLGvAKHnpjc5y7Ywk3PcBiF2vKpNRMzxW
RvhzClTsGQLvUY6OaG6x9fxWxVYMOTYKfTGivR9GTSenqsnTf2NzKyb8oFw4xVcvQOaQufQZPTQk
H9dzx1lYUaoNFrSJpXGJcQ0bfInyezHdzlMnk1EOFcP8p/y1zt+xYhTFNKdkySAFdxh7aP/xcf5q
QyYWTigUf/1e2DlRkrH6tZSfN4kp0i+25IPk+MCE2TKUpN1DawxtBN+hQMXbElt1wOHTXzc0q6qb
KufRZoGA8P+Wfmi+/IPQvraNZEcxzFSU+Qlh3ErWx0yYAMhslUqQIS6BbJySs4SbXIi8AOpFVGgz
BaVhfXLzOgxzJzMvWv605OecmFNGcHRuhyQCSVfVm21IrD2Eeye89Jy5k/mLE3MwFOJANy/ynuS7
a8nt9KVbR2z6cZSKyEJa36yNCvzr59/uX6ZlSHYiZHj9dtP0khfXkNpdjhQTih4vzZa1FdYkHlPH
U9L/xWrRAFz6ghjy4Oao2nIw75zfPHNh/+YVHTHgX/j5xbQukcUrpecECnKcZLKlqrDE5OI9nBs+
oRVYjOnRg9nRkH5+6lIyYApX0Efle7XrqTxKV4iMwdYFbYOaHaaF1DYmtYyvrMrCBPT83e5yJG5b
EM/S+l90P4ZqhdIbbJ4TbqMCQ1Z5qe4OohvFn1toSxzxDTISHNGihH7QX/LDIfa3lQjvyZaZOuZk
1oA2egNpEoW1hQkaBTGkWMS2aRtPgLSK0iy4iRDQX9WNruulgUyORKJMUlxkWFffmFsujSOCNHma
ZBadHxTt9/IehOYrs/MiqVGFBwiLGbwBkdGV12PxggBV6t6qW2MkMNsVoruYIxubmxD1cnUAPh8w
VSgUyw+PA6B3eWcp6rQLgXR0lShnE41MRAJIZvvUXRTDAQBHu56xkkd2jvblQ2Nc0WqkHYLyUX5w
0eZuD8OIn5MQweM+vZBjRKtFW3ylP1ZvqQn4vPgq5AFqW1spnATxyIMv04mb7dzCOzzFV1W7KIch
IUWabaPOl1yUxLWRCgMqil1yN9dq5K16BHUYOP72scAhEF/UO3ccy+d+9bg+XYDXLgQC+iVljSkT
iuF5uEK8uzVIUWsQvGkRT/dpg5xyf6H9JF/braxEMsvsW9HB6Df9OZ0eRNLAFxPOIzp0WUUJdDzX
yICdtsu8vqK17PB8kyU7NL1NV/ssulVGhoqg3xpOnvDsB/Yrr+XgoauQmssyt7lvrTQvWuihDq+l
507XXUi0XRx/MSMtiiTx8ugbh6x+qCmaRM5+DK6uiseJiRvpcktaEzOHqh2UZrRvVDwiCHCC0BWO
fnYoRaaer8wuGJyfQaME7Iy3gbGzqfmVlnDIBsDoPQveUVUKrLirqJZ3RW+bgCURx6Z/InKM+0Y0
ZKrQzy2m0h/cQmSdvIqNcrULz3CeFWXV5Ir4OzQElDTy5Xe8DRs7BXRynHRBybgQmAg2Fqxo7rrO
Ph4BjvYZAkTh0GCphGrk5ZRWQS3iKNl1Svtt4LG6GgpSzhjYvLAs/IEE/0pzdA/obPGVn6Fy+9aJ
bwsVKlmD+LeMazctS7rV0xSv4OM8Gpl5KvYbHzURFt+I9DGoqposGJmo4C/tsvEhdt4svO+FoenF
8OQB1gdYYjvKiflSVUyM32SWHofTD+3if1HtTVvj3aOA8TMRaSvq7cjiTlHTBsDRIEuD0z7SeUyb
5+F1SxraJsFluQn4/dBVPy0QmYmHTbhQeyAAzxD/ab2EbKazp2aQ4a4ht/Z1Kub1dYI1CEaNltnW
h807rA6h3Xgg/pM2Kw5Amr5iStLioAdRoIXlTsHIkSxmCUExjPE1VpAl0B8Fw+0tyvpCG/55Ic5G
Gpi6+JJxclZaaxXKzhYXI0q/g/mOXbZ/2loF5OIieeJwtlARCWN+O267ME/i3mfxHPt/R6SYSmmG
AztkDEnwPgqoOW6Po2LMiBhZxmyOtZgwxBkdvxBGJtYypMyIlEP6gTHh34rxo9CvEliRxH9bcXAf
4/FULTIrI9fMKg+ZILzdqHrcLF1llgqdxewHcbCzepjSFXEW1a7PriJAScRt03gNlBU4VBKRAqtg
E1jmPqiq0MeTk5ezva0bgLxHoUkWvmZfTUbJVSEMN6ycVQyMZ/p5BjQ26iCZ4Av05Rkbozq6GW2z
6c5ysZ74bC61d3Ed3xnjbMEQCAvvlfBJ/v2MDNIqKkxc4AN9f+OMyUeOy/WUJ/4Dh0UbtZAo+/QO
1lei+F2jHQNUpPwq4EPEEa8lyn9a5UMB/EL0TunOloQm+IPrywKT+b7naXjr4xQk88iSKvZtxU8v
1BddYF9yTIw/Gf5Jq9jUV2DkWniVUZjTkqBIQrg0Y30l4Yxu1iT/shIaw0tK6NSZBHICjk2+4ai6
dmK0huHP6txoN/F5XjlLsVbcvI/l8j9qXGN7ulaa0JcgCHN8zx8bY1JEPOQaQKLvgv2k2eyeFycX
U9vT6m3ROvMXWz1czBiM+3qeCPKPt13ZM3DrzRycbP/nmxd9eTIxoAxZBdAbrkNC8eWdvcy9W2RR
I2Gb9xKrWnHu6EPzSkw0YbhDcYaIKLYLd53wmt6EzzwNsjcgFBPI2d0akB7ekbjfNoKQRc8NattC
4To1tHXQMnFcfGoCvpsMb+jts2qL7MK3G2SyGI4ZOiBkl8n67aHtQUFw0t2c5GcJuVGuvgd8XcWg
4LXxdPPKi9asn3vOt4mHpUg7pci1e5QLrMIMQZnj3tTBb6lQjRb0upf+PuTqgbHm+gG7DiFKOTCw
1biYatYd9bS+p5PWnDjy1YJryuQmarAqzWxacLUKCB4FZRYy2UzWHKGQ0e6PoScDgEpogM9W3g5F
d2pTtAcfA+Ch96niHGwUr772605u2HcrUOjp+YXo24fGOqa0MYRFiJyVkF4gPc/diQV1DmF7Zz0H
bBH3o64XJbrfZObAMv5yJfAcZLPK0EJ2rVMZMLAC/SqD8L2DQ9kKCu8QZ+W7B+Z6uXik0/GLltVB
4gCS3NSvE/YrWRhl8RKdOJeDjX9wofJh/cCU1uJZv2lFtxMPUrhIVrz7hvIznGZQvthuXmtg6iO7
wfzq0D9oP6FCMMpp9sXkEEUDY0Kuy3EMQ8MxMUre3HwZQ2OzrpxdPtGk3oTnagu6qb7wJJRkZYsN
XUWyMMsbJ7CJ5LIEBW2uyHlPdz2HwFCpn6tLEpoBWScHwfaCDCyUmsTNvmZbRW12XsuqiuYYAAjf
/TzirZsmmJXCp/mtO9H8iEEKSm8hVlJPvNWom1KKgexnOFsikdqRgmMILyzMfSw93ulihjj1Upjm
EiW6XfC6LQZznbu/0xYDZntpVM8JS3uKSo/weiN3JNZV5bRk7BCYHKccQ+0C/O+GYNgk/gQw16I/
+kXlpKoqoW+4kU4EdYH3uvQXA2N/ikvu3pSQwh272BEZkzWCD/4TWg/kPknA28GOT/Xq+dvqOCze
CfG0Ksce1/Ua5zeZK7b0fwPcWp5/dyXOFmeKxzgPZbC760Y/dU8tKoboqy8Qx6uK8bt8YQ+WRHEP
b+YJI/F4VCrnZWWpkDtcvB8EuK6yAYqBFQNSu9LJCRVk7edTdOHRzHNL4QRmLyJXjMRnSUG3Cudp
JCP7r68/yDu9Jafr+wi/prXT83gVFVwlla56vMSKzkrVaXe9YhSyL/9IKkEkI6uYxpQJ+BZlr2DB
K2szOkm7yCb47Azj8Ds42KuIznpn+rs336/fkH0Vgyzzf6drbhRU3DohnV8eO7BjMYyu80VMMcZt
SOQkUCPDNGfGqFAFBy2lQx5qsFk4i9L1In5tmxV7pHXkzcz5Y26RJH8YktIyE68W2ykDjM/kx1KJ
37+A6jt8xEMU2JkH6k+MEXEQC4CgoG0Ookc5T9VTLeXYbpozKURCCi15sMBH6X4WN8FmH/fkHBMy
HJc7RuaUGAa/cfqLXRylog6tXZ1wUmF0uaQTsoZCqNjhhZFtosqCu2utHTFdkFZuswUhDko/Dyxf
rn1O5YzaDG8q43adf/M1SUPPWzaKJNBmP67ESG4soomLZefYXSHk/PP8aG0Ri2LRmCYWNz8qoVXx
2nizhrWgAP/ZzjpHW3SFYuz8vNyYXuIFzkgSlil552emaqlOXPOYD2vUiNWhggrInbkdk6L7Fia/
eixnd9zQhciY83PkuhN9C6mEoWbFtIeJw8Hg2GC1S5G9NtgIZIrrp1nDwo5ZYhoWrxjmpK/IiytK
UXpenEpdW/zD8JqkdsDY6YiIw2Mv3VA6mk2ycIZ3Z+wYHeRh1kKSXfQEAFhqokuxd0cKq5vk/hyT
+isGwaTH0xDNVblcctkOrnMVgJrjKvjSja3809amPnnNRra25a1IqQYVojoO0UA0iF0gAFqHdi+Q
hSJjEQd3/ISP5BThLeYLM43GHV+NWwiOBQkltGdT0J1e7nGqzoZNbaw2+/qQuMr+mz4KLq8yVOVM
jzRihQMVvO+q6fcAeB7WVbPnOM2tcEtZV/iPiE/21Xo3lxZ4bZYgq/x8iAT5Zax5Bq77JFGdDNJ5
gZn9si8s4tiYw85WCxg2Cs25Rxy+M3wgao0xgpJPcACATUxATT9ihTOdZvVV16QYHJSj4xWdY0xv
5ciOHPt03GEIbBv6EAdOpEIATE5GsTUfhN3NfKRouooPFEz5mSpTIuvnPCUCUsguka6Jz7geIu1U
kvCH4IUZAW6cPPG5CB4t3BZle/cNIimMztfSDML8ZThjXKIb7lBVkVKwThVyxqd7FRN6rl9fv8+G
B87DDLQqnjfqEjkowRtYxXmwL5S08YWamtP7KukKVuqyGqeIatZ/cPJ+ZYvAG5KJb05bGjLPtWLl
e4IWzroo5PoF0ARbWA5Ugfg+8GMyS5IgONRaWspg7AORdA1XPmn66uovTbdXpT4V9rPInQhqZ+G9
U4J6rVaHQ8akxA5JdhO9b2TBwPcMlQOVnuqjnHU5alJER+9QhWxBF9MwP3zrHvHHIn3DoVp383fN
mJ/HfH+P4qSOHScsg2FFsQSRN7zrA4/AAN0SNeTRd8oIwSUy9szjiI+Ln3wJ7TOi2qbzKkVGu4/L
PyJopQC00qwAf7RLQA==
`protect end_protected
